magic
tech sky130A
magscale 1 2
timestamp 1607544406
<< locali >>
rect 283297 666587 283331 683077
rect 551293 606339 551327 606645
rect 28825 589951 28859 598145
rect 28917 595119 28951 598417
rect 283021 589339 283055 598893
rect 551385 596479 551419 601409
rect 551477 595119 551511 596581
rect 551385 586279 551419 592161
rect 551477 586959 551511 592297
rect 554605 586959 554639 590121
rect 26341 572611 26375 572713
rect 28641 570163 28675 575229
rect 28825 567239 28859 580261
rect 551201 576895 551235 582369
rect 28917 573495 28951 576113
rect 29929 572679 29963 572781
rect 30021 570503 30055 573393
rect 553317 572611 553351 576861
rect 26617 535007 26651 535585
rect 33977 532151 34011 532661
rect 548349 532491 548383 532661
rect 548533 532287 548567 532389
rect 34069 531879 34103 532117
rect 34161 531675 34195 531845
rect 196081 531131 196115 531165
rect 195931 531097 196115 531131
rect 186329 530995 186363 531097
rect 173817 529771 173851 530961
rect 191113 530859 191147 531029
rect 201509 530995 201543 531165
rect 206293 530995 206327 531097
rect 222209 531063 222243 531165
rect 231777 530995 231811 531165
rect 231869 531063 231903 531233
rect 241437 531063 241471 531233
rect 241529 531063 241563 531165
rect 251097 530995 251131 531165
rect 251189 531063 251223 531165
rect 264989 531063 265023 531165
rect 263643 531029 263701 531063
rect 274557 530995 274591 531165
rect 325709 531063 325743 531233
rect 292623 531029 292681 531063
rect 302283 531029 302341 531063
rect 282929 530995 282963 531029
rect 282871 530961 282963 530995
rect 335277 530995 335311 531233
rect 338071 530961 338129 530995
rect 342913 529907 342947 530961
rect 543749 530247 543783 530485
rect 547889 530247 547923 531097
rect 547981 530995 548015 531097
rect 550097 530859 550131 531165
rect 550005 530519 550039 530825
rect 550189 530587 550223 530689
rect 549913 530179 549947 530485
rect 550097 530383 550131 530553
rect 388855 528173 389189 528207
rect 403633 528139 403667 528445
rect 388947 528105 389223 528139
rect 389189 528071 389223 528105
rect 389557 528105 389833 528139
rect 389557 528071 389591 528105
rect 406393 528003 406427 528377
rect 408693 528139 408727 528445
rect 413293 528003 413327 528377
rect 422953 528003 422987 528309
rect 423689 528003 423723 528309
rect 434729 528003 434763 528173
rect 444297 528071 444331 528173
rect 456717 528071 456751 528173
rect 463617 528071 463651 528173
rect 468125 528139 468159 530145
rect 550005 530111 550039 530349
rect 463709 528003 463743 528105
rect 89729 500055 89763 500157
rect 283021 499579 283055 509201
rect 547889 500667 547923 500769
rect 547889 500191 547923 500497
rect 546601 472039 546635 473433
rect 551661 467347 551695 471869
rect 551753 467483 551787 471733
rect 552765 470951 552799 471529
rect 552949 468503 552983 473365
rect 553133 471155 553167 471529
rect 551661 467313 551753 467347
rect 283113 452659 283147 462281
rect 282929 434843 282963 437529
rect 282929 423691 282963 433245
rect 283113 405739 283147 415361
rect 80345 396627 80379 401965
rect 86969 401863 87003 402033
rect 99297 402033 99481 402067
rect 99297 401999 99331 402033
rect 96537 401863 96571 401965
rect 106289 401863 106323 402033
rect 118651 401965 118835 401999
rect 115857 401863 115891 401965
rect 118801 401931 118835 401965
rect 128369 401931 128403 401965
rect 128311 401897 128403 401931
rect 133889 401863 133923 401965
rect 143457 401863 143491 401965
rect 144929 401795 144963 401897
rect 153209 401795 153243 402305
rect 282377 347803 282411 357357
rect 202889 320671 202923 320773
rect 207673 320671 207707 320841
rect 282101 305643 282135 309077
rect 282101 299523 282135 305609
rect 126345 224519 126379 224757
rect 127817 224587 127851 224825
rect 127725 224179 127759 224485
rect 128829 224383 128863 224893
rect 128553 223839 128587 224077
rect 214481 222207 214515 224961
rect 214481 212551 214515 222037
rect 214481 202895 214515 205649
rect 214481 173927 214515 179537
rect 38577 29087 38611 31297
rect 133153 29903 133187 30141
rect 80069 29359 80103 29461
rect 89729 29359 89763 29529
rect 41371 29053 41429 29087
rect 57989 29019 58023 29325
rect 74457 29019 74491 29257
rect 74549 29019 74583 29189
rect 83013 29019 83047 29189
rect 94237 29019 94271 29189
rect 104173 29019 104207 29189
rect 109969 29019 110003 29257
rect 121469 29019 121503 29257
rect 68017 19363 68051 28917
rect 144745 25755 144779 25789
rect 172529 25755 172563 25857
rect 115857 20723 115891 25721
rect 144745 25721 144837 25755
rect 182097 25755 182131 25857
rect 183569 25823 183603 26197
rect 128369 25687 128403 25721
rect 128311 25653 128403 25687
rect 164249 25483 164283 25653
rect 169033 25483 169067 25721
rect 65993 9707 66027 19261
rect 67189 9707 67223 12461
rect 121653 12427 121687 19261
rect 179429 9707 179463 12461
rect 182189 9707 182223 19261
rect 184857 9707 184891 13277
rect 287069 13039 287103 13753
rect 296637 13039 296671 13753
rect 306389 12971 306423 13753
rect 315957 12971 315991 13753
rect 325709 12971 325743 13753
rect 335277 12971 335311 13753
rect 366867 13685 367017 13719
rect 366591 13481 366741 13515
rect 366683 13413 366925 13447
rect 366867 13277 366925 13311
rect 366591 13141 366833 13175
rect 366683 13073 366925 13107
rect 366959 12869 367017 12903
rect 367017 12563 367051 12733
rect 375297 12563 375331 12733
rect 379529 12563 379563 12733
rect 382381 12495 382415 12869
rect 384221 12631 384255 13753
rect 393145 12563 393179 12801
rect 393237 12631 393271 13753
rect 402989 12563 403023 13753
rect 403081 12835 403115 13753
rect 412465 12835 412499 13753
rect 412557 12563 412591 13753
rect 422401 12835 422435 13753
rect 208685 12155 208719 12393
rect 210433 12087 210467 12325
rect 219265 12087 219299 12325
rect 219357 12155 219391 12393
rect 229201 12087 229235 12393
rect 238585 12087 238619 12393
rect 248521 12087 248555 12393
rect 257905 12087 257939 12393
rect 428933 12359 428967 14433
rect 545681 14195 545715 14297
rect 431785 12835 431819 13753
rect 431969 13651 432003 13753
rect 436201 13175 436235 13753
rect 451933 13175 451967 13413
rect 456809 12835 456843 13005
rect 461501 12903 461535 13005
rect 461501 12869 461685 12903
rect 461777 12835 461811 13005
rect 475393 12903 475427 13005
rect 296453 12121 296637 12155
rect 383703 12121 383887 12155
rect 210341 11679 210375 11985
rect 219357 11679 219391 11985
rect 229109 11679 229143 11985
rect 238677 11679 238711 11985
rect 248429 11679 248463 11985
rect 257997 11679 258031 11985
rect 267749 11679 267783 11985
rect 267841 11611 267875 12053
rect 277225 11611 277259 12053
rect 277317 11679 277351 11985
rect 287069 11679 287103 11985
rect 287161 11611 287195 12053
rect 296453 11543 296487 12121
rect 296545 11611 296579 12053
rect 296637 11679 296671 11985
rect 306389 11679 306423 11985
rect 306481 11611 306515 12053
rect 315865 11611 315899 12053
rect 315957 11679 315991 11985
rect 325709 11679 325743 11985
rect 325801 11611 325835 12053
rect 335185 11611 335219 12053
rect 335277 11679 335311 11985
rect 383669 11407 383703 11985
rect 383761 11339 383795 12053
rect 383853 12019 383887 12121
rect 393053 12121 393237 12155
rect 403023 12121 403207 12155
rect 393053 12019 393087 12121
rect 393145 11339 393179 12053
rect 393237 11407 393271 11985
rect 402989 11135 403023 11985
rect 403081 11067 403115 12053
rect 403173 12019 403207 12121
rect 412373 12121 412557 12155
rect 412373 12019 412407 12121
rect 412465 11067 412499 12053
rect 412557 11135 412591 11985
rect 419457 11815 419491 12121
rect 438225 11951 438259 12053
rect 470609 11883 470643 11985
rect 419365 11067 419399 11781
rect 125609 4199 125643 4301
rect 35909 3723 35943 4097
rect 45661 3383 45695 4097
rect 55263 3825 55355 3859
rect 50353 3043 50387 3281
rect 55229 2975 55263 3689
rect 55321 2907 55355 3825
rect 60105 3247 60139 4097
rect 93869 3859 93903 4165
rect 74583 3825 74675 3859
rect 57989 3111 58023 3213
rect 62313 2975 62347 3689
rect 67005 2907 67039 3825
rect 74549 3043 74583 3689
rect 74641 2907 74675 3825
rect 84025 3825 84117 3859
rect 103437 3859 103471 4165
rect 84025 2907 84059 3825
rect 113189 3723 113223 4165
rect 84117 2975 84151 3689
rect 93869 2907 93903 3689
rect 125517 3723 125551 4165
rect 103437 2771 103471 3689
rect 111015 2805 111257 2839
rect 126621 595 126655 9605
rect 130117 3723 130151 3825
rect 130025 3451 130059 3689
rect 133153 3655 133187 3825
rect 139501 3791 139535 4029
rect 147689 3859 147723 4097
rect 162869 3859 162903 3961
rect 166951 3825 167009 3859
rect 138581 3519 138615 3757
rect 142813 3655 142847 3825
rect 162869 3247 162903 3349
rect 168021 1003 168055 3893
rect 183845 3791 183879 4913
rect 182315 3621 182557 3655
rect 182315 3485 182373 3519
rect 171149 3111 171183 3213
rect 180717 3111 180751 3417
rect 182189 3179 182223 3417
rect 186237 3383 186271 7837
rect 195253 3859 195287 4097
rect 186329 3247 186363 3349
rect 186271 3213 186363 3247
rect 193137 3179 193171 3417
rect 195345 3383 195379 3825
rect 201509 3315 201543 3417
rect 202797 595 202831 9605
rect 443193 9095 443227 9469
rect 451933 9231 451967 9605
rect 204085 3383 204119 4029
rect 441629 3791 441663 4029
rect 430807 3621 430991 3655
rect 430957 3587 430991 3621
rect 303629 3383 303663 3553
rect 432613 3519 432647 3553
rect 360209 3247 360243 3349
rect 383393 3043 383427 3281
rect 390569 3043 390603 3213
rect 406025 3043 406059 3485
rect 418077 3043 418111 3485
rect 422711 3485 423689 3519
rect 432613 3485 432889 3519
rect 419641 2839 419675 3009
rect 419733 2839 419767 3417
rect 421481 3043 421515 3485
rect 448989 2499 449023 8925
rect 502475 4029 502625 4063
rect 347363 2261 347605 2295
rect 328135 2193 328193 2227
rect 386095 2193 386153 2227
rect 347455 2125 347605 2159
rect 386003 2125 386245 2159
rect 453957 2091 453991 3825
rect 463525 3655 463559 3961
rect 463709 3655 463743 3961
rect 502567 3961 502717 3995
rect 473277 3655 473311 3961
rect 502383 3893 502625 3927
rect 515505 3859 515539 4097
rect 483063 3825 483213 3859
rect 483155 3757 483305 3791
rect 502475 3757 502625 3791
rect 559849 3723 559883 3961
rect 483063 3689 483213 3723
rect 483155 3621 483305 3655
rect 463835 3553 463893 3587
rect 483247 3553 483397 3587
rect 483063 3485 483305 3519
rect 473403 3417 473553 3451
rect 492689 3315 492723 3621
rect 502383 3621 502625 3655
rect 501153 3383 501187 3485
rect 502257 3315 502291 3621
rect 564633 3043 564667 3349
rect 328043 2057 328285 2091
rect 347363 2057 347697 2091
rect 328135 1921 328377 1955
rect 328043 1853 328193 1887
rect 347455 1853 347697 1887
rect 386187 1853 386245 1887
<< viali >>
rect 283297 683077 283331 683111
rect 283297 666553 283331 666587
rect 551293 606645 551327 606679
rect 551293 606305 551327 606339
rect 551385 601409 551419 601443
rect 283021 598893 283055 598927
rect 28917 598417 28951 598451
rect 28825 598145 28859 598179
rect 28917 595085 28951 595119
rect 28825 589917 28859 589951
rect 551385 596445 551419 596479
rect 551477 596581 551511 596615
rect 551477 595085 551511 595119
rect 551477 592297 551511 592331
rect 283021 589305 283055 589339
rect 551385 592161 551419 592195
rect 551477 586925 551511 586959
rect 554605 590121 554639 590155
rect 554605 586925 554639 586959
rect 551385 586245 551419 586279
rect 551201 582369 551235 582403
rect 28825 580261 28859 580295
rect 28641 575229 28675 575263
rect 26341 572713 26375 572747
rect 26341 572577 26375 572611
rect 28641 570129 28675 570163
rect 551201 576861 551235 576895
rect 553317 576861 553351 576895
rect 28917 576113 28951 576147
rect 28917 573461 28951 573495
rect 30021 573393 30055 573427
rect 29929 572781 29963 572815
rect 29929 572645 29963 572679
rect 553317 572577 553351 572611
rect 30021 570469 30055 570503
rect 28825 567205 28859 567239
rect 26617 535585 26651 535619
rect 26617 534973 26651 535007
rect 33977 532661 34011 532695
rect 548349 532661 548383 532695
rect 548349 532457 548383 532491
rect 548533 532389 548567 532423
rect 548533 532253 548567 532287
rect 33977 532117 34011 532151
rect 34069 532117 34103 532151
rect 34069 531845 34103 531879
rect 34161 531845 34195 531879
rect 34161 531641 34195 531675
rect 231869 531233 231903 531267
rect 196081 531165 196115 531199
rect 186329 531097 186363 531131
rect 195897 531097 195931 531131
rect 201509 531165 201543 531199
rect 173817 530961 173851 530995
rect 186329 530961 186363 530995
rect 191113 531029 191147 531063
rect 222209 531165 222243 531199
rect 201509 530961 201543 530995
rect 206293 531097 206327 531131
rect 222209 531029 222243 531063
rect 231777 531165 231811 531199
rect 206293 530961 206327 530995
rect 231869 531029 231903 531063
rect 241437 531233 241471 531267
rect 325709 531233 325743 531267
rect 241437 531029 241471 531063
rect 241529 531165 241563 531199
rect 241529 531029 241563 531063
rect 251097 531165 251131 531199
rect 231777 530961 231811 530995
rect 251189 531165 251223 531199
rect 264989 531165 265023 531199
rect 251189 531029 251223 531063
rect 263609 531029 263643 531063
rect 263701 531029 263735 531063
rect 264989 531029 265023 531063
rect 274557 531165 274591 531199
rect 251097 530961 251131 530995
rect 282929 531029 282963 531063
rect 292589 531029 292623 531063
rect 292681 531029 292715 531063
rect 302249 531029 302283 531063
rect 302341 531029 302375 531063
rect 325709 531029 325743 531063
rect 335277 531233 335311 531267
rect 274557 530961 274591 530995
rect 282837 530961 282871 530995
rect 550097 531165 550131 531199
rect 547889 531097 547923 531131
rect 335277 530961 335311 530995
rect 338037 530961 338071 530995
rect 338129 530961 338163 530995
rect 342913 530961 342947 530995
rect 191113 530825 191147 530859
rect 543749 530485 543783 530519
rect 543749 530213 543783 530247
rect 547981 531097 548015 531131
rect 547981 530961 548015 530995
rect 550005 530825 550039 530859
rect 550097 530825 550131 530859
rect 550189 530689 550223 530723
rect 547889 530213 547923 530247
rect 549913 530485 549947 530519
rect 550005 530485 550039 530519
rect 550097 530553 550131 530587
rect 550189 530553 550223 530587
rect 342913 529873 342947 529907
rect 468125 530145 468159 530179
rect 549913 530145 549947 530179
rect 550005 530349 550039 530383
rect 550097 530349 550131 530383
rect 173817 529737 173851 529771
rect 403633 528445 403667 528479
rect 388821 528173 388855 528207
rect 389189 528173 389223 528207
rect 408693 528445 408727 528479
rect 388913 528105 388947 528139
rect 389189 528037 389223 528071
rect 389833 528105 389867 528139
rect 403633 528105 403667 528139
rect 406393 528377 406427 528411
rect 389557 528037 389591 528071
rect 408693 528105 408727 528139
rect 413293 528377 413327 528411
rect 406393 527969 406427 528003
rect 413293 527969 413327 528003
rect 422953 528309 422987 528343
rect 422953 527969 422987 528003
rect 423689 528309 423723 528343
rect 423689 527969 423723 528003
rect 434729 528173 434763 528207
rect 444297 528173 444331 528207
rect 444297 528037 444331 528071
rect 456717 528173 456751 528207
rect 456717 528037 456751 528071
rect 463617 528173 463651 528207
rect 550005 530077 550039 530111
rect 463617 528037 463651 528071
rect 463709 528105 463743 528139
rect 468125 528105 468159 528139
rect 434729 527969 434763 528003
rect 463709 527969 463743 528003
rect 283021 509201 283055 509235
rect 89729 500157 89763 500191
rect 89729 500021 89763 500055
rect 547889 500769 547923 500803
rect 547889 500633 547923 500667
rect 547889 500497 547923 500531
rect 547889 500157 547923 500191
rect 283021 499545 283055 499579
rect 546601 473433 546635 473467
rect 546601 472005 546635 472039
rect 552949 473365 552983 473399
rect 551661 471869 551695 471903
rect 551753 471733 551787 471767
rect 552765 471529 552799 471563
rect 552765 470917 552799 470951
rect 553133 471529 553167 471563
rect 553133 471121 553167 471155
rect 552949 468469 552983 468503
rect 551753 467449 551787 467483
rect 551753 467313 551787 467347
rect 283113 462281 283147 462315
rect 283113 452625 283147 452659
rect 282929 437529 282963 437563
rect 282929 434809 282963 434843
rect 282929 433245 282963 433279
rect 282929 423657 282963 423691
rect 283113 415361 283147 415395
rect 283113 405705 283147 405739
rect 153209 402305 153243 402339
rect 86969 402033 87003 402067
rect 80345 401965 80379 401999
rect 99481 402033 99515 402067
rect 106289 402033 106323 402067
rect 86969 401829 87003 401863
rect 96537 401965 96571 401999
rect 99297 401965 99331 401999
rect 96537 401829 96571 401863
rect 106289 401829 106323 401863
rect 115857 401965 115891 401999
rect 118617 401965 118651 401999
rect 128369 401965 128403 401999
rect 118801 401897 118835 401931
rect 128277 401897 128311 401931
rect 133889 401965 133923 401999
rect 115857 401829 115891 401863
rect 133889 401829 133923 401863
rect 143457 401965 143491 401999
rect 143457 401829 143491 401863
rect 144929 401897 144963 401931
rect 144929 401761 144963 401795
rect 153209 401761 153243 401795
rect 80345 396593 80379 396627
rect 282377 357357 282411 357391
rect 282377 347769 282411 347803
rect 207673 320841 207707 320875
rect 202889 320773 202923 320807
rect 202889 320637 202923 320671
rect 207673 320637 207707 320671
rect 282101 309077 282135 309111
rect 282101 305609 282135 305643
rect 282101 299489 282135 299523
rect 214481 224961 214515 224995
rect 128829 224893 128863 224927
rect 127817 224825 127851 224859
rect 126345 224757 126379 224791
rect 127817 224553 127851 224587
rect 126345 224485 126379 224519
rect 127725 224485 127759 224519
rect 128829 224349 128863 224383
rect 127725 224145 127759 224179
rect 128553 224077 128587 224111
rect 128553 223805 128587 223839
rect 214481 222173 214515 222207
rect 214481 222037 214515 222071
rect 214481 212517 214515 212551
rect 214481 205649 214515 205683
rect 214481 202861 214515 202895
rect 214481 179537 214515 179571
rect 214481 173893 214515 173927
rect 38577 31297 38611 31331
rect 133153 30141 133187 30175
rect 133153 29869 133187 29903
rect 89729 29529 89763 29563
rect 80069 29461 80103 29495
rect 57989 29325 58023 29359
rect 80069 29325 80103 29359
rect 89729 29325 89763 29359
rect 38577 29053 38611 29087
rect 41337 29053 41371 29087
rect 41429 29053 41463 29087
rect 57989 28985 58023 29019
rect 74457 29257 74491 29291
rect 109969 29257 110003 29291
rect 74457 28985 74491 29019
rect 74549 29189 74583 29223
rect 74549 28985 74583 29019
rect 83013 29189 83047 29223
rect 83013 28985 83047 29019
rect 94237 29189 94271 29223
rect 94237 28985 94271 29019
rect 104173 29189 104207 29223
rect 104173 28985 104207 29019
rect 109969 28985 110003 29019
rect 121469 29257 121503 29291
rect 121469 28985 121503 29019
rect 68017 28917 68051 28951
rect 183569 26197 183603 26231
rect 172529 25857 172563 25891
rect 144745 25789 144779 25823
rect 115857 25721 115891 25755
rect 128369 25721 128403 25755
rect 144837 25721 144871 25755
rect 169033 25721 169067 25755
rect 172529 25721 172563 25755
rect 182097 25857 182131 25891
rect 183569 25789 183603 25823
rect 182097 25721 182131 25755
rect 128277 25653 128311 25687
rect 164249 25653 164283 25687
rect 164249 25449 164283 25483
rect 169033 25449 169067 25483
rect 115857 20689 115891 20723
rect 68017 19329 68051 19363
rect 65993 19261 66027 19295
rect 121653 19261 121687 19295
rect 65993 9673 66027 9707
rect 67189 12461 67223 12495
rect 182189 19261 182223 19295
rect 121653 12393 121687 12427
rect 179429 12461 179463 12495
rect 67189 9673 67223 9707
rect 179429 9673 179463 9707
rect 428933 14433 428967 14467
rect 287069 13753 287103 13787
rect 182189 9673 182223 9707
rect 184857 13277 184891 13311
rect 287069 13005 287103 13039
rect 296637 13753 296671 13787
rect 296637 13005 296671 13039
rect 306389 13753 306423 13787
rect 306389 12937 306423 12971
rect 315957 13753 315991 13787
rect 315957 12937 315991 12971
rect 325709 13753 325743 13787
rect 325709 12937 325743 12971
rect 335277 13753 335311 13787
rect 384221 13753 384255 13787
rect 366833 13685 366867 13719
rect 367017 13685 367051 13719
rect 366557 13481 366591 13515
rect 366741 13481 366775 13515
rect 366649 13413 366683 13447
rect 366925 13413 366959 13447
rect 366833 13277 366867 13311
rect 366925 13277 366959 13311
rect 366557 13141 366591 13175
rect 366833 13141 366867 13175
rect 366649 13073 366683 13107
rect 366925 13073 366959 13107
rect 335277 12937 335311 12971
rect 366925 12869 366959 12903
rect 367017 12869 367051 12903
rect 382381 12869 382415 12903
rect 367017 12733 367051 12767
rect 367017 12529 367051 12563
rect 375297 12733 375331 12767
rect 375297 12529 375331 12563
rect 379529 12733 379563 12767
rect 379529 12529 379563 12563
rect 393237 13753 393271 13787
rect 384221 12597 384255 12631
rect 393145 12801 393179 12835
rect 393237 12597 393271 12631
rect 402989 13753 403023 13787
rect 393145 12529 393179 12563
rect 403081 13753 403115 13787
rect 403081 12801 403115 12835
rect 412465 13753 412499 13787
rect 412465 12801 412499 12835
rect 412557 13753 412591 13787
rect 402989 12529 403023 12563
rect 422401 13753 422435 13787
rect 422401 12801 422435 12835
rect 412557 12529 412591 12563
rect 382381 12461 382415 12495
rect 208685 12393 208719 12427
rect 219357 12393 219391 12427
rect 208685 12121 208719 12155
rect 210433 12325 210467 12359
rect 210433 12053 210467 12087
rect 219265 12325 219299 12359
rect 219357 12121 219391 12155
rect 229201 12393 229235 12427
rect 219265 12053 219299 12087
rect 229201 12053 229235 12087
rect 238585 12393 238619 12427
rect 238585 12053 238619 12087
rect 248521 12393 248555 12427
rect 248521 12053 248555 12087
rect 257905 12393 257939 12427
rect 545681 14297 545715 14331
rect 545681 14161 545715 14195
rect 431785 13753 431819 13787
rect 431969 13753 432003 13787
rect 431969 13617 432003 13651
rect 436201 13753 436235 13787
rect 436201 13141 436235 13175
rect 451933 13413 451967 13447
rect 451933 13141 451967 13175
rect 431785 12801 431819 12835
rect 456809 13005 456843 13039
rect 461501 13005 461535 13039
rect 461777 13005 461811 13039
rect 461685 12869 461719 12903
rect 456809 12801 456843 12835
rect 475393 13005 475427 13039
rect 475393 12869 475427 12903
rect 461777 12801 461811 12835
rect 428933 12325 428967 12359
rect 296637 12121 296671 12155
rect 383669 12121 383703 12155
rect 257905 12053 257939 12087
rect 267841 12053 267875 12087
rect 210341 11985 210375 12019
rect 210341 11645 210375 11679
rect 219357 11985 219391 12019
rect 219357 11645 219391 11679
rect 229109 11985 229143 12019
rect 229109 11645 229143 11679
rect 238677 11985 238711 12019
rect 238677 11645 238711 11679
rect 248429 11985 248463 12019
rect 248429 11645 248463 11679
rect 257997 11985 258031 12019
rect 257997 11645 258031 11679
rect 267749 11985 267783 12019
rect 267749 11645 267783 11679
rect 267841 11577 267875 11611
rect 277225 12053 277259 12087
rect 287161 12053 287195 12087
rect 277317 11985 277351 12019
rect 277317 11645 277351 11679
rect 287069 11985 287103 12019
rect 287069 11645 287103 11679
rect 277225 11577 277259 11611
rect 287161 11577 287195 11611
rect 296545 12053 296579 12087
rect 306481 12053 306515 12087
rect 296637 11985 296671 12019
rect 296637 11645 296671 11679
rect 306389 11985 306423 12019
rect 306389 11645 306423 11679
rect 296545 11577 296579 11611
rect 306481 11577 306515 11611
rect 315865 12053 315899 12087
rect 325801 12053 325835 12087
rect 315957 11985 315991 12019
rect 315957 11645 315991 11679
rect 325709 11985 325743 12019
rect 325709 11645 325743 11679
rect 315865 11577 315899 11611
rect 325801 11577 325835 11611
rect 335185 12053 335219 12087
rect 383761 12053 383795 12087
rect 335277 11985 335311 12019
rect 335277 11645 335311 11679
rect 383669 11985 383703 12019
rect 335185 11577 335219 11611
rect 296453 11509 296487 11543
rect 383669 11373 383703 11407
rect 383853 11985 383887 12019
rect 393237 12121 393271 12155
rect 402989 12121 403023 12155
rect 393053 11985 393087 12019
rect 393145 12053 393179 12087
rect 383761 11305 383795 11339
rect 403081 12053 403115 12087
rect 393237 11985 393271 12019
rect 393237 11373 393271 11407
rect 402989 11985 403023 12019
rect 393145 11305 393179 11339
rect 402989 11101 403023 11135
rect 403173 11985 403207 12019
rect 412557 12121 412591 12155
rect 419457 12121 419491 12155
rect 412373 11985 412407 12019
rect 412465 12053 412499 12087
rect 403081 11033 403115 11067
rect 412557 11985 412591 12019
rect 438225 12053 438259 12087
rect 438225 11917 438259 11951
rect 470609 11985 470643 12019
rect 470609 11849 470643 11883
rect 412557 11101 412591 11135
rect 419365 11781 419399 11815
rect 419457 11781 419491 11815
rect 412465 11033 412499 11067
rect 419365 11033 419399 11067
rect 184857 9673 184891 9707
rect 126621 9605 126655 9639
rect 125609 4301 125643 4335
rect 93869 4165 93903 4199
rect 35909 4097 35943 4131
rect 35909 3689 35943 3723
rect 45661 4097 45695 4131
rect 60105 4097 60139 4131
rect 55229 3825 55263 3859
rect 45661 3349 45695 3383
rect 55229 3689 55263 3723
rect 50353 3281 50387 3315
rect 50353 3009 50387 3043
rect 55229 2941 55263 2975
rect 67005 3825 67039 3859
rect 74549 3825 74583 3859
rect 57989 3213 58023 3247
rect 60105 3213 60139 3247
rect 62313 3689 62347 3723
rect 57989 3077 58023 3111
rect 62313 2941 62347 2975
rect 55321 2873 55355 2907
rect 74549 3689 74583 3723
rect 74549 3009 74583 3043
rect 67005 2873 67039 2907
rect 74641 2873 74675 2907
rect 84117 3825 84151 3859
rect 93869 3825 93903 3859
rect 103437 4165 103471 4199
rect 103437 3825 103471 3859
rect 113189 4165 113223 4199
rect 84117 3689 84151 3723
rect 84117 2941 84151 2975
rect 93869 3689 93903 3723
rect 84025 2873 84059 2907
rect 93869 2873 93903 2907
rect 103437 3689 103471 3723
rect 113189 3689 113223 3723
rect 125517 4165 125551 4199
rect 125609 4165 125643 4199
rect 125517 3689 125551 3723
rect 110981 2805 111015 2839
rect 111257 2805 111291 2839
rect 103437 2737 103471 2771
rect 202797 9605 202831 9639
rect 186237 7837 186271 7871
rect 183845 4913 183879 4947
rect 147689 4097 147723 4131
rect 139501 4029 139535 4063
rect 130117 3825 130151 3859
rect 130025 3689 130059 3723
rect 130117 3689 130151 3723
rect 133153 3825 133187 3859
rect 133153 3621 133187 3655
rect 138581 3757 138615 3791
rect 139501 3757 139535 3791
rect 142813 3825 142847 3859
rect 147689 3825 147723 3859
rect 162869 3961 162903 3995
rect 168021 3893 168055 3927
rect 162869 3825 162903 3859
rect 166917 3825 166951 3859
rect 167009 3825 167043 3859
rect 142813 3621 142847 3655
rect 138581 3485 138615 3519
rect 130025 3417 130059 3451
rect 162869 3349 162903 3383
rect 162869 3213 162903 3247
rect 183845 3757 183879 3791
rect 182281 3621 182315 3655
rect 182557 3621 182591 3655
rect 182281 3485 182315 3519
rect 182373 3485 182407 3519
rect 180717 3417 180751 3451
rect 171149 3213 171183 3247
rect 171149 3077 171183 3111
rect 182189 3417 182223 3451
rect 195253 4097 195287 4131
rect 195253 3825 195287 3859
rect 195345 3825 195379 3859
rect 193137 3417 193171 3451
rect 186237 3349 186271 3383
rect 186329 3349 186363 3383
rect 186237 3213 186271 3247
rect 182189 3145 182223 3179
rect 195345 3349 195379 3383
rect 201509 3417 201543 3451
rect 201509 3281 201543 3315
rect 193137 3145 193171 3179
rect 180717 3077 180751 3111
rect 168021 969 168055 1003
rect 126621 561 126655 595
rect 451933 9605 451967 9639
rect 443193 9469 443227 9503
rect 451933 9197 451967 9231
rect 443193 9061 443227 9095
rect 448989 8925 449023 8959
rect 204085 4029 204119 4063
rect 441629 4029 441663 4063
rect 441629 3757 441663 3791
rect 430773 3621 430807 3655
rect 204085 3349 204119 3383
rect 303629 3553 303663 3587
rect 430957 3553 430991 3587
rect 432613 3553 432647 3587
rect 406025 3485 406059 3519
rect 303629 3349 303663 3383
rect 360209 3349 360243 3383
rect 360209 3213 360243 3247
rect 383393 3281 383427 3315
rect 383393 3009 383427 3043
rect 390569 3213 390603 3247
rect 390569 3009 390603 3043
rect 406025 3009 406059 3043
rect 418077 3485 418111 3519
rect 421481 3485 421515 3519
rect 422677 3485 422711 3519
rect 423689 3485 423723 3519
rect 432889 3485 432923 3519
rect 419733 3417 419767 3451
rect 418077 3009 418111 3043
rect 419641 3009 419675 3043
rect 419641 2805 419675 2839
rect 421481 3009 421515 3043
rect 419733 2805 419767 2839
rect 515505 4097 515539 4131
rect 502441 4029 502475 4063
rect 502625 4029 502659 4063
rect 463525 3961 463559 3995
rect 448989 2465 449023 2499
rect 453957 3825 453991 3859
rect 347329 2261 347363 2295
rect 347605 2261 347639 2295
rect 328101 2193 328135 2227
rect 328193 2193 328227 2227
rect 386061 2193 386095 2227
rect 386153 2193 386187 2227
rect 347421 2125 347455 2159
rect 347605 2125 347639 2159
rect 385969 2125 386003 2159
rect 386245 2125 386279 2159
rect 463525 3621 463559 3655
rect 463709 3961 463743 3995
rect 463709 3621 463743 3655
rect 473277 3961 473311 3995
rect 502533 3961 502567 3995
rect 502717 3961 502751 3995
rect 502349 3893 502383 3927
rect 502625 3893 502659 3927
rect 483029 3825 483063 3859
rect 483213 3825 483247 3859
rect 515505 3825 515539 3859
rect 559849 3961 559883 3995
rect 483121 3757 483155 3791
rect 483305 3757 483339 3791
rect 502441 3757 502475 3791
rect 502625 3757 502659 3791
rect 483029 3689 483063 3723
rect 483213 3689 483247 3723
rect 559849 3689 559883 3723
rect 473277 3621 473311 3655
rect 483121 3621 483155 3655
rect 483305 3621 483339 3655
rect 492689 3621 492723 3655
rect 463801 3553 463835 3587
rect 463893 3553 463927 3587
rect 483213 3553 483247 3587
rect 483397 3553 483431 3587
rect 483029 3485 483063 3519
rect 483305 3485 483339 3519
rect 473369 3417 473403 3451
rect 473553 3417 473587 3451
rect 502257 3621 502291 3655
rect 502349 3621 502383 3655
rect 502625 3621 502659 3655
rect 501153 3485 501187 3519
rect 501153 3349 501187 3383
rect 492689 3281 492723 3315
rect 502257 3281 502291 3315
rect 564633 3349 564667 3383
rect 564633 3009 564667 3043
rect 328009 2057 328043 2091
rect 328285 2057 328319 2091
rect 347329 2057 347363 2091
rect 347697 2057 347731 2091
rect 453957 2057 453991 2091
rect 328101 1921 328135 1955
rect 328377 1921 328411 1955
rect 328009 1853 328043 1887
rect 328193 1853 328227 1887
rect 347421 1853 347455 1887
rect 347697 1853 347731 1887
rect 386153 1853 386187 1887
rect 386245 1853 386279 1887
rect 202797 561 202831 595
<< metal1 >>
rect 305638 700544 305644 700596
rect 305696 700584 305702 700596
rect 332502 700584 332508 700596
rect 305696 700556 332508 700584
rect 305696 700544 305702 700556
rect 332502 700544 332508 700556
rect 332560 700544 332566 700596
rect 138658 700476 138664 700528
rect 138716 700516 138722 700528
rect 154114 700516 154120 700528
rect 138716 700488 154120 700516
rect 138716 700476 138722 700488
rect 154114 700476 154120 700488
rect 154172 700476 154178 700528
rect 202782 700476 202788 700528
rect 202840 700516 202846 700528
rect 250622 700516 250628 700528
rect 202840 700488 250628 700516
rect 202840 700476 202846 700488
rect 250622 700476 250628 700488
rect 250680 700476 250686 700528
rect 267642 700476 267648 700528
rect 267700 700516 267706 700528
rect 282178 700516 282184 700528
rect 267700 700488 282184 700516
rect 267700 700476 267706 700488
rect 282178 700476 282184 700488
rect 282236 700476 282242 700528
rect 301498 700476 301504 700528
rect 301556 700516 301562 700528
rect 397454 700516 397460 700528
rect 301556 700488 397460 700516
rect 301556 700476 301562 700488
rect 397454 700476 397460 700488
rect 397512 700476 397518 700528
rect 51718 700408 51724 700460
rect 51776 700448 51782 700460
rect 72970 700448 72976 700460
rect 51776 700420 72976 700448
rect 51776 700408 51782 700420
rect 72970 700408 72976 700420
rect 73028 700408 73034 700460
rect 89162 700408 89168 700460
rect 89220 700448 89226 700460
rect 138750 700448 138756 700460
rect 89220 700420 138756 700448
rect 89220 700408 89226 700420
rect 138750 700408 138756 700420
rect 138808 700408 138814 700460
rect 218974 700408 218980 700460
rect 219032 700448 219038 700460
rect 282454 700448 282460 700460
rect 219032 700420 282460 700448
rect 219032 700408 219038 700420
rect 282454 700408 282460 700420
rect 282512 700408 282518 700460
rect 313918 700408 313924 700460
rect 313976 700448 313982 700460
rect 413646 700448 413652 700460
rect 313976 700420 413652 700448
rect 313976 700408 313982 700420
rect 413646 700408 413652 700420
rect 413704 700408 413710 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 282362 700380 282368 700392
rect 40552 700352 282368 700380
rect 40552 700340 40558 700352
rect 282362 700340 282368 700352
rect 282420 700340 282426 700392
rect 312538 700340 312544 700392
rect 312596 700380 312602 700392
rect 462314 700380 462320 700392
rect 312596 700352 462320 700380
rect 312596 700340 312602 700352
rect 462314 700340 462320 700352
rect 462372 700340 462378 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 8938 700312 8944 700324
rect 8168 700284 8944 700312
rect 8168 700272 8174 700284
rect 8938 700272 8944 700284
rect 8996 700272 9002 700324
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 282270 700312 282276 700324
rect 24360 700284 282276 700312
rect 24360 700272 24366 700284
rect 282270 700272 282276 700284
rect 282328 700272 282334 700324
rect 315298 700272 315304 700324
rect 315356 700312 315362 700324
rect 527174 700312 527180 700324
rect 315356 700284 527180 700312
rect 315356 700272 315362 700284
rect 527174 700272 527180 700284
rect 527232 700272 527238 700324
rect 250622 698640 250628 698692
rect 250680 698680 250686 698692
rect 252554 698680 252560 698692
rect 250680 698652 252560 698680
rect 250680 698640 250686 698652
rect 252554 698640 252560 698652
rect 252612 698640 252618 698692
rect 283282 698232 283288 698284
rect 283340 698272 283346 698284
rect 283926 698272 283932 698284
rect 283340 698244 283932 698272
rect 283340 698232 283346 698244
rect 283926 698232 283932 698244
rect 283984 698232 283990 698284
rect 136634 697552 136640 697604
rect 136692 697592 136698 697604
rect 137830 697592 137836 697604
rect 136692 697564 137836 697592
rect 136692 697552 136698 697564
rect 137830 697552 137836 697564
rect 137888 697552 137894 697604
rect 576118 696940 576124 696992
rect 576176 696980 576182 696992
rect 580166 696980 580172 696992
rect 576176 696952 580172 696980
rect 576176 696940 576182 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 252554 696872 252560 696924
rect 252612 696912 252618 696924
rect 260006 696912 260012 696924
rect 252612 696884 260012 696912
rect 252612 696872 252618 696884
rect 260006 696872 260012 696884
rect 260064 696872 260070 696924
rect 260006 694764 260012 694816
rect 260064 694804 260070 694816
rect 266998 694804 267004 694816
rect 260064 694776 267004 694804
rect 260064 694764 260070 694776
rect 266998 694764 267004 694776
rect 267056 694764 267062 694816
rect 283098 694084 283104 694136
rect 283156 694124 283162 694136
rect 283282 694124 283288 694136
rect 283156 694096 283288 694124
rect 283156 694084 283162 694096
rect 283282 694084 283288 694096
rect 283340 694084 283346 694136
rect 283098 692724 283104 692776
rect 283156 692764 283162 692776
rect 283282 692764 283288 692776
rect 283156 692736 283288 692764
rect 283156 692724 283162 692736
rect 283282 692724 283288 692736
rect 283340 692724 283346 692776
rect 48498 691364 48504 691416
rect 48556 691404 48562 691416
rect 51718 691404 51724 691416
rect 48556 691376 51724 691404
rect 48556 691364 48562 691376
rect 51718 691364 51724 691376
rect 51776 691364 51782 691416
rect 46934 685176 46940 685228
rect 46992 685216 46998 685228
rect 48498 685216 48504 685228
rect 46992 685188 48504 685216
rect 46992 685176 46998 685188
rect 48498 685176 48504 685188
rect 48556 685176 48562 685228
rect 282914 683068 282920 683120
rect 282972 683108 282978 683120
rect 283285 683111 283343 683117
rect 283285 683108 283297 683111
rect 282972 683080 283297 683108
rect 282972 683068 282978 683080
rect 283285 683077 283297 683080
rect 283331 683077 283343 683111
rect 283285 683071 283343 683077
rect 3510 681708 3516 681760
rect 3568 681748 3574 681760
rect 453298 681748 453304 681760
rect 3568 681720 453304 681748
rect 3568 681708 3574 681720
rect 453298 681708 453304 681720
rect 453356 681708 453362 681760
rect 46934 680388 46940 680400
rect 44192 680360 46940 680388
rect 42058 680212 42064 680264
rect 42116 680252 42122 680264
rect 44192 680252 44220 680360
rect 46934 680348 46940 680360
rect 46992 680348 46998 680400
rect 42116 680224 44220 680252
rect 42116 680212 42122 680224
rect 133874 674772 133880 674824
rect 133932 674812 133938 674824
rect 136634 674812 136640 674824
rect 133932 674784 136640 674812
rect 133932 674772 133938 674784
rect 136634 674772 136640 674784
rect 136692 674772 136698 674824
rect 40034 672052 40040 672104
rect 40092 672092 40098 672104
rect 42058 672092 42064 672104
rect 40092 672064 42064 672092
rect 40092 672052 40098 672064
rect 42058 672052 42064 672064
rect 42116 672052 42122 672104
rect 131758 670692 131764 670744
rect 131816 670732 131822 670744
rect 133874 670732 133880 670744
rect 131816 670704 133880 670732
rect 131816 670692 131822 670704
rect 133874 670692 133880 670704
rect 133932 670692 133938 670744
rect 266998 670624 267004 670676
rect 267056 670664 267062 670676
rect 269758 670664 269764 670676
rect 267056 670636 269764 670664
rect 267056 670624 267062 670636
rect 269758 670624 269764 670636
rect 269816 670624 269822 670676
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 287698 667944 287704 667956
rect 3476 667916 287704 667944
rect 3476 667904 3482 667916
rect 287698 667904 287704 667916
rect 287756 667904 287762 667956
rect 40034 666584 40040 666596
rect 38672 666556 40040 666584
rect 37918 666476 37924 666528
rect 37976 666516 37982 666528
rect 38672 666516 38700 666556
rect 40034 666544 40040 666556
rect 40092 666544 40098 666596
rect 283285 666587 283343 666593
rect 283285 666553 283297 666587
rect 283331 666584 283343 666587
rect 283374 666584 283380 666596
rect 283331 666556 283380 666584
rect 283331 666553 283343 666556
rect 283285 666547 283343 666553
rect 283374 666544 283380 666556
rect 283432 666544 283438 666596
rect 37976 666488 38700 666516
rect 37976 666476 37982 666488
rect 269758 659404 269764 659456
rect 269816 659444 269822 659456
rect 271138 659444 271144 659456
rect 269816 659416 271144 659444
rect 269816 659404 269822 659416
rect 271138 659404 271144 659416
rect 271196 659404 271202 659456
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 10318 652780 10324 652792
rect 3108 652752 10324 652780
rect 3108 652740 3114 652752
rect 10318 652740 10324 652752
rect 10376 652740 10382 652792
rect 271138 651516 271144 651568
rect 271196 651556 271202 651568
rect 271966 651556 271972 651568
rect 271196 651528 271972 651556
rect 271196 651516 271202 651528
rect 271966 651516 271972 651528
rect 272024 651516 272030 651568
rect 36538 650020 36544 650072
rect 36596 650060 36602 650072
rect 37918 650060 37924 650072
rect 36596 650032 37924 650060
rect 36596 650020 36602 650032
rect 37918 650020 37924 650032
rect 37976 650020 37982 650072
rect 577498 650020 577504 650072
rect 577556 650060 577562 650072
rect 579614 650060 579620 650072
rect 577556 650032 579620 650060
rect 577556 650020 577562 650032
rect 579614 650020 579620 650032
rect 579672 650020 579678 650072
rect 271966 648592 271972 648644
rect 272024 648632 272030 648644
rect 272024 648604 273300 648632
rect 272024 648592 272030 648604
rect 273272 648564 273300 648604
rect 274634 648564 274640 648576
rect 273272 648536 274640 648564
rect 274634 648524 274640 648536
rect 274692 648524 274698 648576
rect 128998 648320 129004 648372
rect 129056 648360 129062 648372
rect 131758 648360 131764 648372
rect 129056 648332 131764 648360
rect 129056 648320 129062 648332
rect 131758 648320 131764 648332
rect 131816 648320 131822 648372
rect 283098 647232 283104 647284
rect 283156 647272 283162 647284
rect 283190 647272 283196 647284
rect 283156 647244 283196 647272
rect 283156 647232 283162 647244
rect 283190 647232 283196 647244
rect 283248 647232 283254 647284
rect 274634 645804 274640 645856
rect 274692 645844 274698 645856
rect 276658 645844 276664 645856
rect 274692 645816 276664 645844
rect 274692 645804 274698 645816
rect 276658 645804 276664 645816
rect 276716 645804 276722 645856
rect 283098 640364 283104 640416
rect 283156 640404 283162 640416
rect 283190 640404 283196 640416
rect 283156 640376 283196 640404
rect 283156 640364 283162 640376
rect 283190 640364 283196 640376
rect 283248 640364 283254 640416
rect 126238 640296 126244 640348
rect 126296 640336 126302 640348
rect 128998 640336 129004 640348
rect 126296 640308 129004 640336
rect 126296 640296 126302 640308
rect 128998 640296 129004 640308
rect 129056 640296 129062 640348
rect 35250 634788 35256 634840
rect 35308 634828 35314 634840
rect 36538 634828 36544 634840
rect 35308 634800 36544 634828
rect 35308 634788 35314 634800
rect 36538 634788 36544 634800
rect 36596 634788 36602 634840
rect 276658 633156 276664 633208
rect 276716 633196 276722 633208
rect 278314 633196 278320 633208
rect 276716 633168 278320 633196
rect 276716 633156 276722 633168
rect 278314 633156 278320 633168
rect 278372 633156 278378 633208
rect 283006 630640 283012 630692
rect 283064 630680 283070 630692
rect 283190 630680 283196 630692
rect 283064 630652 283196 630680
rect 283064 630640 283070 630652
rect 283190 630640 283196 630652
rect 283248 630640 283254 630692
rect 116578 629892 116584 629944
rect 116636 629932 116642 629944
rect 126238 629932 126244 629944
rect 116636 629904 126244 629932
rect 116636 629892 116642 629904
rect 126238 629892 126244 629904
rect 126296 629892 126302 629944
rect 33778 629484 33784 629536
rect 33836 629524 33842 629536
rect 35250 629524 35256 629536
rect 33836 629496 35256 629524
rect 33836 629484 33842 629496
rect 35250 629484 35256 629496
rect 35308 629484 35314 629536
rect 278314 627852 278320 627904
rect 278372 627892 278378 627904
rect 279142 627892 279148 627904
rect 278372 627864 279148 627892
rect 278372 627852 278378 627864
rect 279142 627852 279148 627864
rect 279200 627852 279206 627904
rect 551370 627308 551376 627360
rect 551428 627348 551434 627360
rect 551646 627348 551652 627360
rect 551428 627320 551652 627348
rect 551428 627308 551434 627320
rect 551646 627308 551652 627320
rect 551704 627308 551710 627360
rect 23382 619624 23388 619676
rect 23440 619664 23446 619676
rect 84102 619664 84108 619676
rect 23440 619636 84108 619664
rect 23440 619624 23446 619636
rect 84102 619624 84108 619636
rect 84160 619624 84166 619676
rect 551186 618672 551192 618724
rect 551244 618712 551250 618724
rect 551554 618712 551560 618724
rect 551244 618684 551560 618712
rect 551244 618672 551250 618684
rect 551554 618672 551560 618684
rect 551612 618672 551618 618724
rect 29730 618536 29736 618588
rect 29788 618576 29794 618588
rect 33778 618576 33784 618588
rect 29788 618548 33784 618576
rect 29788 618536 29794 618548
rect 33778 618536 33784 618548
rect 33836 618536 33842 618588
rect 453298 616768 453304 616820
rect 453356 616808 453362 616820
rect 456794 616808 456800 616820
rect 453356 616780 456800 616808
rect 453356 616768 453362 616780
rect 456794 616768 456800 616780
rect 456852 616768 456858 616820
rect 282362 614048 282368 614100
rect 282420 614088 282426 614100
rect 313274 614088 313280 614100
rect 282420 614060 313280 614088
rect 282420 614048 282426 614060
rect 313274 614048 313280 614060
rect 313332 614048 313338 614100
rect 283006 611328 283012 611380
rect 283064 611368 283070 611380
rect 283190 611368 283196 611380
rect 283064 611340 283196 611368
rect 283064 611328 283070 611340
rect 283190 611328 283196 611340
rect 283248 611328 283254 611380
rect 551370 611260 551376 611312
rect 551428 611300 551434 611312
rect 551830 611300 551836 611312
rect 551428 611272 551836 611300
rect 551428 611260 551434 611272
rect 551830 611260 551836 611272
rect 551888 611260 551894 611312
rect 3326 609968 3332 610020
rect 3384 610008 3390 610020
rect 13078 610008 13084 610020
rect 3384 609980 13084 610008
rect 3384 609968 3390 609980
rect 13078 609968 13084 609980
rect 13136 609968 13142 610020
rect 551281 606679 551339 606685
rect 551281 606645 551293 606679
rect 551327 606676 551339 606679
rect 551830 606676 551836 606688
rect 551327 606648 551836 606676
rect 551327 606645 551339 606648
rect 551281 606639 551339 606645
rect 551830 606636 551836 606648
rect 551888 606636 551894 606688
rect 551186 606500 551192 606552
rect 551244 606540 551250 606552
rect 551830 606540 551836 606552
rect 551244 606512 551836 606540
rect 551244 606500 551250 606512
rect 551830 606500 551836 606512
rect 551888 606500 551894 606552
rect 551278 606432 551284 606484
rect 551336 606472 551342 606484
rect 551922 606472 551928 606484
rect 551336 606444 551928 606472
rect 551336 606432 551342 606444
rect 551922 606432 551928 606444
rect 551980 606432 551986 606484
rect 551278 606336 551284 606348
rect 551239 606308 551284 606336
rect 551278 606296 551284 606308
rect 551336 606296 551342 606348
rect 551370 601440 551376 601452
rect 551331 601412 551376 601440
rect 551370 601400 551376 601412
rect 551428 601400 551434 601452
rect 283009 598927 283067 598933
rect 283009 598893 283021 598927
rect 283055 598924 283067 598927
rect 283190 598924 283196 598936
rect 283055 598896 283196 598924
rect 283055 598893 283067 598896
rect 283009 598887 283067 598893
rect 283190 598884 283196 598896
rect 283248 598884 283254 598936
rect 28902 598448 28908 598460
rect 28863 598420 28908 598448
rect 28902 598408 28908 598420
rect 28960 598408 28966 598460
rect 28813 598179 28871 598185
rect 28813 598145 28825 598179
rect 28859 598176 28871 598179
rect 28902 598176 28908 598188
rect 28859 598148 28908 598176
rect 28859 598145 28871 598148
rect 28813 598139 28871 598145
rect 28902 598136 28908 598148
rect 28960 598136 28966 598188
rect 551186 598000 551192 598052
rect 551244 598040 551250 598052
rect 551830 598040 551836 598052
rect 551244 598012 551836 598040
rect 551244 598000 551250 598012
rect 551830 598000 551836 598012
rect 551888 598000 551894 598052
rect 26142 597932 26148 597984
rect 26200 597972 26206 597984
rect 28902 597972 28908 597984
rect 26200 597944 28908 597972
rect 26200 597932 26206 597944
rect 28902 597932 28908 597944
rect 28960 597932 28966 597984
rect 551278 597020 551284 597032
rect 551204 596992 551284 597020
rect 551204 596748 551232 596992
rect 551278 596980 551284 596992
rect 551336 596980 551342 597032
rect 551278 596844 551284 596896
rect 551336 596884 551342 596896
rect 551922 596884 551928 596896
rect 551336 596856 551928 596884
rect 551336 596844 551342 596856
rect 551922 596844 551928 596856
rect 551980 596844 551986 596896
rect 551922 596748 551928 596760
rect 551204 596720 551928 596748
rect 551922 596708 551928 596720
rect 551980 596708 551986 596760
rect 551370 596572 551376 596624
rect 551428 596612 551434 596624
rect 551465 596615 551523 596621
rect 551465 596612 551477 596615
rect 551428 596584 551477 596612
rect 551428 596572 551434 596584
rect 551465 596581 551477 596584
rect 551511 596581 551523 596615
rect 551465 596575 551523 596581
rect 551370 596476 551376 596488
rect 551331 596448 551376 596476
rect 551370 596436 551376 596448
rect 551428 596436 551434 596488
rect 28902 595116 28908 595128
rect 28863 595088 28908 595116
rect 28902 595076 28908 595088
rect 28960 595076 28966 595128
rect 551370 595076 551376 595128
rect 551428 595116 551434 595128
rect 551465 595119 551523 595125
rect 551465 595116 551477 595119
rect 551428 595088 551477 595116
rect 551428 595076 551434 595088
rect 551465 595085 551477 595088
rect 551511 595085 551523 595119
rect 551465 595079 551523 595085
rect 3510 594804 3516 594856
rect 3568 594844 3574 594856
rect 9030 594844 9036 594856
rect 3568 594816 9036 594844
rect 3568 594804 3574 594816
rect 9030 594804 9036 594816
rect 9088 594804 9094 594856
rect 139210 594668 139216 594720
rect 139268 594708 139274 594720
rect 139578 594708 139584 594720
rect 139268 594680 139584 594708
rect 139268 594668 139274 594680
rect 139578 594668 139584 594680
rect 139636 594668 139642 594720
rect 551370 592288 551376 592340
rect 551428 592328 551434 592340
rect 551465 592331 551523 592337
rect 551465 592328 551477 592331
rect 551428 592300 551477 592328
rect 551428 592288 551434 592300
rect 551465 592297 551477 592300
rect 551511 592297 551523 592331
rect 551465 592291 551523 592297
rect 551370 592192 551376 592204
rect 551331 592164 551376 592192
rect 551370 592152 551376 592164
rect 551428 592152 551434 592204
rect 551370 592016 551376 592068
rect 551428 592056 551434 592068
rect 551922 592056 551928 592068
rect 551428 592028 551928 592056
rect 551428 592016 551434 592028
rect 551922 592016 551928 592028
rect 551980 592016 551986 592068
rect 554590 590152 554596 590164
rect 554551 590124 554596 590152
rect 554590 590112 554596 590124
rect 554648 590112 554654 590164
rect 28813 589951 28871 589957
rect 28813 589917 28825 589951
rect 28859 589948 28871 589951
rect 28902 589948 28908 589960
rect 28859 589920 28908 589948
rect 28859 589917 28871 589920
rect 28813 589911 28871 589917
rect 28902 589908 28908 589920
rect 28960 589908 28966 589960
rect 28258 589364 28264 589416
rect 28316 589404 28322 589416
rect 28902 589404 28908 589416
rect 28316 589376 28908 589404
rect 28316 589364 28322 589376
rect 28902 589364 28908 589376
rect 28960 589364 28966 589416
rect 283006 589336 283012 589348
rect 282967 589308 283012 589336
rect 283006 589296 283012 589308
rect 283064 589296 283070 589348
rect 554590 589296 554596 589348
rect 554648 589336 554654 589348
rect 556154 589336 556160 589348
rect 554648 589308 556160 589336
rect 554648 589296 554654 589308
rect 556154 589296 556160 589308
rect 556212 589296 556218 589348
rect 28442 589228 28448 589280
rect 28500 589268 28506 589280
rect 28902 589268 28908 589280
rect 28500 589240 28908 589268
rect 28500 589228 28506 589240
rect 28902 589228 28908 589240
rect 28960 589228 28966 589280
rect 554590 588752 554596 588804
rect 554648 588792 554654 588804
rect 557626 588792 557632 588804
rect 554648 588764 557632 588792
rect 554648 588752 554654 588764
rect 557626 588752 557632 588764
rect 557684 588752 557690 588804
rect 28350 588548 28356 588600
rect 28408 588588 28414 588600
rect 28902 588588 28908 588600
rect 28408 588560 28908 588588
rect 28408 588548 28414 588560
rect 28902 588548 28908 588560
rect 28960 588548 28966 588600
rect 551278 587188 551284 587240
rect 551336 587228 551342 587240
rect 551922 587228 551928 587240
rect 551336 587200 551928 587228
rect 551336 587188 551342 587200
rect 551922 587188 551928 587200
rect 551980 587188 551986 587240
rect 554590 587052 554596 587104
rect 554648 587092 554654 587104
rect 556798 587092 556804 587104
rect 554648 587064 556804 587092
rect 554648 587052 554654 587064
rect 556798 587052 556804 587064
rect 556856 587052 556862 587104
rect 551370 586916 551376 586968
rect 551428 586956 551434 586968
rect 551465 586959 551523 586965
rect 551465 586956 551477 586959
rect 551428 586928 551477 586956
rect 551428 586916 551434 586928
rect 551465 586925 551477 586928
rect 551511 586925 551523 586959
rect 554590 586956 554596 586968
rect 554551 586928 554596 586956
rect 551465 586919 551523 586925
rect 554590 586916 554596 586928
rect 554648 586916 554654 586968
rect 554866 586304 554872 586356
rect 554924 586344 554930 586356
rect 558178 586344 558184 586356
rect 554924 586316 558184 586344
rect 554924 586304 554930 586316
rect 558178 586304 558184 586316
rect 558236 586304 558242 586356
rect 551370 586276 551376 586288
rect 551331 586248 551376 586276
rect 551370 586236 551376 586248
rect 551428 586236 551434 586288
rect 24118 586032 24124 586084
rect 24176 586072 24182 586084
rect 26142 586072 26148 586084
rect 24176 586044 26148 586072
rect 24176 586032 24182 586044
rect 26142 586032 26148 586044
rect 26200 586032 26206 586084
rect 554866 585148 554872 585200
rect 554924 585188 554930 585200
rect 560294 585188 560300 585200
rect 554924 585160 560300 585188
rect 554924 585148 554930 585160
rect 560294 585148 560300 585160
rect 560352 585148 560358 585200
rect 554866 583720 554872 583772
rect 554924 583760 554930 583772
rect 561766 583760 561772 583772
rect 554924 583732 561772 583760
rect 554924 583720 554930 583732
rect 561766 583720 561772 583732
rect 561824 583720 561830 583772
rect 551186 582400 551192 582412
rect 551147 582372 551192 582400
rect 551186 582360 551192 582372
rect 551244 582360 551250 582412
rect 554866 581000 554872 581052
rect 554924 581040 554930 581052
rect 563054 581040 563060 581052
rect 554924 581012 563060 581040
rect 554924 581000 554930 581012
rect 563054 581000 563060 581012
rect 563112 581000 563118 581052
rect 28813 580295 28871 580301
rect 28813 580261 28825 580295
rect 28859 580292 28871 580295
rect 28902 580292 28908 580304
rect 28859 580264 28908 580292
rect 28859 580261 28871 580264
rect 28813 580255 28871 580261
rect 28902 580252 28908 580264
rect 28960 580252 28966 580304
rect 283006 579640 283012 579692
rect 283064 579680 283070 579692
rect 283098 579680 283104 579692
rect 283064 579652 283104 579680
rect 283064 579640 283070 579652
rect 283098 579640 283104 579652
rect 283156 579640 283162 579692
rect 554866 579640 554872 579692
rect 554924 579680 554930 579692
rect 564434 579680 564440 579692
rect 554924 579652 564440 579680
rect 554924 579640 554930 579652
rect 564434 579640 564440 579652
rect 564492 579640 564498 579692
rect 576210 579640 576216 579692
rect 576268 579680 576274 579692
rect 580166 579680 580172 579692
rect 576268 579652 580172 579680
rect 576268 579640 576274 579652
rect 580166 579640 580172 579652
rect 580224 579640 580230 579692
rect 554866 578212 554872 578264
rect 554924 578252 554930 578264
rect 565814 578252 565820 578264
rect 554924 578224 565820 578252
rect 554924 578212 554930 578224
rect 565814 578212 565820 578224
rect 565872 578212 565878 578264
rect 551186 576892 551192 576904
rect 551147 576864 551192 576892
rect 551186 576852 551192 576864
rect 551244 576852 551250 576904
rect 551278 576852 551284 576904
rect 551336 576892 551342 576904
rect 551922 576892 551928 576904
rect 551336 576864 551928 576892
rect 551336 576852 551342 576864
rect 551922 576852 551928 576864
rect 551980 576852 551986 576904
rect 553302 576892 553308 576904
rect 553263 576864 553308 576892
rect 553302 576852 553308 576864
rect 553360 576852 553366 576904
rect 554866 576852 554872 576904
rect 554924 576892 554930 576904
rect 567286 576892 567292 576904
rect 554924 576864 567292 576892
rect 554924 576852 554930 576864
rect 567286 576852 567292 576864
rect 567344 576852 567350 576904
rect 28626 576104 28632 576156
rect 28684 576104 28690 576156
rect 28902 576144 28908 576156
rect 28863 576116 28908 576144
rect 28902 576104 28908 576116
rect 28960 576104 28966 576156
rect 28644 575872 28672 576104
rect 28902 575872 28908 575884
rect 28644 575844 28908 575872
rect 28902 575832 28908 575844
rect 28960 575832 28966 575884
rect 553302 575492 553308 575544
rect 553360 575532 553366 575544
rect 560938 575532 560944 575544
rect 553360 575504 560944 575532
rect 553360 575492 553366 575504
rect 560938 575492 560944 575504
rect 560996 575492 561002 575544
rect 28626 575260 28632 575272
rect 28587 575232 28632 575260
rect 28626 575220 28632 575232
rect 28684 575220 28690 575272
rect 28626 575084 28632 575136
rect 28684 575124 28690 575136
rect 28902 575124 28908 575136
rect 28684 575096 28908 575124
rect 28684 575084 28690 575096
rect 28902 575084 28908 575096
rect 28960 575084 28966 575136
rect 28810 575016 28816 575068
rect 28868 575016 28874 575068
rect 28626 574988 28632 575000
rect 28552 574960 28632 574988
rect 28552 574784 28580 574960
rect 28626 574948 28632 574960
rect 28684 574948 28690 575000
rect 28626 574812 28632 574864
rect 28684 574852 28690 574864
rect 28828 574852 28856 575016
rect 28684 574824 28856 574852
rect 28684 574812 28690 574824
rect 28810 574784 28816 574796
rect 28552 574756 28816 574784
rect 28810 574744 28816 574756
rect 28868 574744 28874 574796
rect 553302 574200 553308 574252
rect 553360 574240 553366 574252
rect 568574 574240 568580 574252
rect 553360 574212 568580 574240
rect 553360 574200 553366 574212
rect 568574 574200 568580 574212
rect 568632 574200 568638 574252
rect 553302 574064 553308 574116
rect 553360 574104 553366 574116
rect 569954 574104 569960 574116
rect 553360 574076 569960 574104
rect 553360 574064 553366 574076
rect 569954 574064 569960 574076
rect 570012 574064 570018 574116
rect 28905 573495 28963 573501
rect 28905 573461 28917 573495
rect 28951 573492 28963 573495
rect 29362 573492 29368 573504
rect 28951 573464 29368 573492
rect 28951 573461 28963 573464
rect 28905 573455 28963 573461
rect 29362 573452 29368 573464
rect 29420 573452 29426 573504
rect 30006 573424 30012 573436
rect 29967 573396 30012 573424
rect 30006 573384 30012 573396
rect 30064 573384 30070 573436
rect 29086 572772 29092 572824
rect 29144 572812 29150 572824
rect 29917 572815 29975 572821
rect 29144 572784 29316 572812
rect 29144 572772 29150 572784
rect 29288 572756 29316 572784
rect 29917 572781 29929 572815
rect 29963 572812 29975 572815
rect 30098 572812 30104 572824
rect 29963 572784 30104 572812
rect 29963 572781 29975 572784
rect 29917 572775 29975 572781
rect 30098 572772 30104 572784
rect 30156 572772 30162 572824
rect 26329 572747 26387 572753
rect 26329 572713 26341 572747
rect 26375 572744 26387 572747
rect 26418 572744 26424 572756
rect 26375 572716 26424 572744
rect 26375 572713 26387 572716
rect 26329 572707 26387 572713
rect 26418 572704 26424 572716
rect 26476 572704 26482 572756
rect 29270 572704 29276 572756
rect 29328 572704 29334 572756
rect 553302 572704 553308 572756
rect 553360 572744 553366 572756
rect 571426 572744 571432 572756
rect 553360 572716 571432 572744
rect 553360 572704 553366 572716
rect 571426 572704 571432 572716
rect 571484 572704 571490 572756
rect 29914 572676 29920 572688
rect 29875 572648 29920 572676
rect 29914 572636 29920 572648
rect 29972 572636 29978 572688
rect 26329 572611 26387 572617
rect 26329 572577 26341 572611
rect 26375 572608 26387 572611
rect 26418 572608 26424 572620
rect 26375 572580 26424 572608
rect 26375 572577 26387 572580
rect 26329 572571 26387 572577
rect 26418 572568 26424 572580
rect 26476 572568 26482 572620
rect 551922 572568 551928 572620
rect 551980 572608 551986 572620
rect 553305 572611 553363 572617
rect 553305 572608 553317 572611
rect 551980 572580 553317 572608
rect 551980 572568 551986 572580
rect 553305 572577 553317 572580
rect 553351 572577 553363 572611
rect 553305 572571 553363 572577
rect 199286 572432 199292 572484
rect 199344 572472 199350 572484
rect 204254 572472 204260 572484
rect 199344 572444 204260 572472
rect 199344 572432 199350 572444
rect 204254 572432 204260 572444
rect 204312 572432 204318 572484
rect 189534 572296 189540 572348
rect 189592 572336 189598 572348
rect 195974 572336 195980 572348
rect 189592 572308 195980 572336
rect 189592 572296 189598 572308
rect 195974 572296 195980 572308
rect 196032 572296 196038 572348
rect 198090 572296 198096 572348
rect 198148 572336 198154 572348
rect 202874 572336 202880 572348
rect 198148 572308 202880 572336
rect 198148 572296 198154 572308
rect 202874 572296 202880 572308
rect 202932 572296 202938 572348
rect 188338 572160 188344 572212
rect 188396 572200 188402 572212
rect 194594 572200 194600 572212
rect 188396 572172 194600 572200
rect 188396 572160 188402 572172
rect 194594 572160 194600 572172
rect 194652 572160 194658 572212
rect 196802 572160 196808 572212
rect 196860 572200 196866 572212
rect 202966 572200 202972 572212
rect 196860 572172 202972 572200
rect 196860 572160 196866 572172
rect 202966 572160 202972 572172
rect 203024 572160 203030 572212
rect 209038 572160 209044 572212
rect 209096 572200 209102 572212
rect 213914 572200 213920 572212
rect 209096 572172 213920 572200
rect 209096 572160 209102 572172
rect 213914 572160 213920 572172
rect 213972 572160 213978 572212
rect 206646 572092 206652 572144
rect 206704 572132 206710 572144
rect 211154 572132 211160 572144
rect 206704 572104 211160 572132
rect 206704 572092 206710 572104
rect 211154 572092 211160 572104
rect 211212 572092 211218 572144
rect 218882 572092 218888 572144
rect 218940 572132 218946 572144
rect 222194 572132 222200 572144
rect 218940 572104 222200 572132
rect 218940 572092 218946 572104
rect 222194 572092 222200 572104
rect 222252 572092 222258 572144
rect 190270 572024 190276 572076
rect 190328 572064 190334 572076
rect 197354 572064 197360 572076
rect 190328 572036 197360 572064
rect 190328 572024 190334 572036
rect 197354 572024 197360 572036
rect 197412 572024 197418 572076
rect 207842 572024 207848 572076
rect 207900 572064 207906 572076
rect 212534 572064 212540 572076
rect 207900 572036 212540 572064
rect 207900 572024 207906 572036
rect 212534 572024 212540 572036
rect 212592 572024 212598 572076
rect 194410 571888 194416 571940
rect 194468 571928 194474 571940
rect 200114 571928 200120 571940
rect 194468 571900 200120 571928
rect 194468 571888 194474 571900
rect 200114 571888 200120 571900
rect 200172 571888 200178 571940
rect 205358 571888 205364 571940
rect 205416 571928 205422 571940
rect 209774 571928 209780 571940
rect 205416 571900 209780 571928
rect 205416 571888 205422 571900
rect 209774 571888 209780 571900
rect 209832 571888 209838 571940
rect 227438 571888 227444 571940
rect 227496 571928 227502 571940
rect 229094 571928 229100 571940
rect 227496 571900 229100 571928
rect 227496 571888 227502 571900
rect 229094 571888 229100 571900
rect 229152 571888 229158 571940
rect 195606 571820 195612 571872
rect 195664 571860 195670 571872
rect 201494 571860 201500 571872
rect 195664 571832 201500 571860
rect 195664 571820 195670 571832
rect 201494 571820 201500 571832
rect 201552 571820 201558 571872
rect 23290 571752 23296 571804
rect 23348 571792 23354 571804
rect 24670 571792 24676 571804
rect 23348 571764 24676 571792
rect 23348 571752 23354 571764
rect 24670 571752 24676 571764
rect 24728 571752 24734 571804
rect 267642 571752 267648 571804
rect 267700 571792 267706 571804
rect 268286 571792 268292 571804
rect 267700 571764 268292 571792
rect 267700 571752 267706 571764
rect 268286 571752 268292 571764
rect 268344 571752 268350 571804
rect 217594 571684 217600 571736
rect 217652 571724 217658 571736
rect 220814 571724 220820 571736
rect 217652 571696 220820 571724
rect 217652 571684 217658 571696
rect 220814 571684 220820 571696
rect 220872 571684 220878 571736
rect 216398 571616 216404 571668
rect 216456 571656 216462 571668
rect 219434 571656 219440 571668
rect 216456 571628 219440 571656
rect 216456 571616 216462 571628
rect 219434 571616 219440 571628
rect 219492 571616 219498 571668
rect 228634 571616 228640 571668
rect 228692 571656 228698 571668
rect 230474 571656 230480 571668
rect 228692 571628 230480 571656
rect 228692 571616 228698 571628
rect 230474 571616 230480 571628
rect 230532 571616 230538 571668
rect 553302 571616 553308 571668
rect 553360 571656 553366 571668
rect 558270 571656 558276 571668
rect 553360 571628 558276 571656
rect 553360 571616 553366 571628
rect 558270 571616 558276 571628
rect 558328 571616 558334 571668
rect 202782 571548 202788 571600
rect 202840 571588 202846 571600
rect 208394 571588 208400 571600
rect 202840 571560 208400 571588
rect 202840 571548 202846 571560
rect 208394 571548 208400 571560
rect 208452 571548 208458 571600
rect 213822 571548 213828 571600
rect 213880 571588 213886 571600
rect 218054 571588 218060 571600
rect 213880 571560 218060 571588
rect 213880 571548 213886 571560
rect 218054 571548 218060 571560
rect 218112 571548 218118 571600
rect 220078 571548 220084 571600
rect 220136 571588 220142 571600
rect 223666 571588 223672 571600
rect 220136 571560 223672 571588
rect 220136 571548 220142 571560
rect 223666 571548 223672 571560
rect 223724 571548 223730 571600
rect 224862 571548 224868 571600
rect 224920 571588 224926 571600
rect 227806 571588 227812 571600
rect 224920 571560 227812 571588
rect 224920 571548 224926 571560
rect 227806 571548 227812 571560
rect 227864 571548 227870 571600
rect 201402 571480 201408 571532
rect 201460 571520 201466 571532
rect 207014 571520 207020 571532
rect 201460 571492 207020 571520
rect 201460 571480 201466 571492
rect 207014 571480 207020 571492
rect 207072 571480 207078 571532
rect 212442 571480 212448 571532
rect 212500 571520 212506 571532
rect 216674 571520 216680 571532
rect 212500 571492 216680 571520
rect 212500 571480 212506 571492
rect 216674 571480 216680 571492
rect 216732 571480 216738 571532
rect 223482 571480 223488 571532
rect 223540 571520 223546 571532
rect 226334 571520 226340 571532
rect 223540 571492 226340 571520
rect 223540 571480 223546 571492
rect 226334 571480 226340 571492
rect 226392 571480 226398 571532
rect 231026 571480 231032 571532
rect 231084 571520 231090 571532
rect 233326 571520 233332 571532
rect 231084 571492 233332 571520
rect 231084 571480 231090 571492
rect 233326 571480 233332 571492
rect 233384 571480 233390 571532
rect 273070 571480 273076 571532
rect 273128 571520 273134 571532
rect 275646 571520 275652 571532
rect 273128 571492 275652 571520
rect 273128 571480 273134 571492
rect 275646 571480 275652 571492
rect 275704 571480 275710 571532
rect 278682 571480 278688 571532
rect 278740 571520 278746 571532
rect 281718 571520 281724 571532
rect 278740 571492 281724 571520
rect 278740 571480 278746 571492
rect 281718 571480 281724 571492
rect 281776 571480 281782 571532
rect 191742 571412 191748 571464
rect 191800 571452 191806 571464
rect 198826 571452 198832 571464
rect 191800 571424 198832 571452
rect 191800 571412 191806 571424
rect 198826 571412 198832 571424
rect 198884 571412 198890 571464
rect 200482 571412 200488 571464
rect 200540 571452 200546 571464
rect 205634 571452 205640 571464
rect 200540 571424 205640 571452
rect 200540 571412 200546 571424
rect 205634 571412 205640 571424
rect 205692 571412 205698 571464
rect 211522 571412 211528 571464
rect 211580 571452 211586 571464
rect 215294 571452 215300 571464
rect 211580 571424 215300 571452
rect 211580 571412 211586 571424
rect 215294 571412 215300 571424
rect 215352 571412 215358 571464
rect 222102 571412 222108 571464
rect 222160 571452 222166 571464
rect 224954 571452 224960 571464
rect 222160 571424 224960 571452
rect 222160 571412 222166 571424
rect 224954 571412 224960 571424
rect 225012 571412 225018 571464
rect 233142 571412 233148 571464
rect 233200 571452 233206 571464
rect 234614 571452 234620 571464
rect 233200 571424 234620 571452
rect 233200 571412 233206 571424
rect 234614 571412 234620 571424
rect 234672 571412 234678 571464
rect 235902 571412 235908 571464
rect 235960 571452 235966 571464
rect 237466 571452 237472 571464
rect 235960 571424 237472 571452
rect 235960 571412 235966 571424
rect 237466 571412 237472 571424
rect 237524 571412 237530 571464
rect 269022 571412 269028 571464
rect 269080 571452 269086 571464
rect 270770 571452 270776 571464
rect 269080 571424 270776 571452
rect 269080 571412 269086 571424
rect 270770 571412 270776 571424
rect 270828 571412 270834 571464
rect 271782 571412 271788 571464
rect 271840 571452 271846 571464
rect 273254 571452 273260 571464
rect 271840 571424 273260 571452
rect 271840 571412 271846 571424
rect 273254 571412 273260 571424
rect 273312 571412 273318 571464
rect 274542 571412 274548 571464
rect 274600 571452 274606 571464
rect 276842 571452 276848 571464
rect 274600 571424 276848 571452
rect 274600 571412 274606 571424
rect 276842 571412 276848 571424
rect 276900 571412 276906 571464
rect 277302 571412 277308 571464
rect 277360 571452 277366 571464
rect 279326 571452 279332 571464
rect 277360 571424 279332 571452
rect 277360 571412 277366 571424
rect 279326 571412 279332 571424
rect 279384 571412 279390 571464
rect 193122 571344 193128 571396
rect 193180 571384 193186 571396
rect 198734 571384 198740 571396
rect 193180 571356 198740 571384
rect 193180 571344 193186 571356
rect 198734 571344 198740 571356
rect 198792 571344 198798 571396
rect 204162 571344 204168 571396
rect 204220 571384 204226 571396
rect 208486 571384 208492 571396
rect 204220 571356 208492 571384
rect 204220 571344 204226 571356
rect 208486 571344 208492 571356
rect 208544 571344 208550 571396
rect 210326 571344 210332 571396
rect 210384 571384 210390 571396
rect 214006 571384 214012 571396
rect 210384 571356 214012 571384
rect 210384 571344 210390 571356
rect 214006 571344 214012 571356
rect 214064 571344 214070 571396
rect 215202 571344 215208 571396
rect 215260 571384 215266 571396
rect 218146 571384 218152 571396
rect 215260 571356 218152 571384
rect 215260 571344 215266 571356
rect 218146 571344 218152 571356
rect 218204 571344 218210 571396
rect 221274 571344 221280 571396
rect 221332 571384 221338 571396
rect 223574 571384 223580 571396
rect 221332 571356 223580 571384
rect 221332 571344 221338 571356
rect 223574 571344 223580 571356
rect 223632 571344 223638 571396
rect 226150 571344 226156 571396
rect 226208 571384 226214 571396
rect 227714 571384 227720 571396
rect 226208 571356 227720 571384
rect 226208 571344 226214 571356
rect 227714 571344 227720 571356
rect 227772 571344 227778 571396
rect 229830 571344 229836 571396
rect 229888 571384 229894 571396
rect 231854 571384 231860 571396
rect 229888 571356 231860 571384
rect 229888 571344 229894 571356
rect 231854 571344 231860 571356
rect 231912 571344 231918 571396
rect 232314 571344 232320 571396
rect 232372 571384 232378 571396
rect 233234 571384 233240 571396
rect 232372 571356 233240 571384
rect 232372 571344 232378 571356
rect 233234 571344 233240 571356
rect 233292 571344 233298 571396
rect 234522 571344 234528 571396
rect 234580 571384 234586 571396
rect 235994 571384 236000 571396
rect 234580 571356 236000 571384
rect 234580 571344 234586 571356
rect 235994 571344 236000 571356
rect 236052 571344 236058 571396
rect 239582 571344 239588 571396
rect 239640 571384 239646 571396
rect 240134 571384 240140 571396
rect 239640 571356 240140 571384
rect 239640 571344 239646 571356
rect 240134 571344 240140 571356
rect 240192 571344 240198 571396
rect 240870 571344 240876 571396
rect 240928 571384 240934 571396
rect 241514 571384 241520 571396
rect 240928 571356 241520 571384
rect 240928 571344 240934 571356
rect 241514 571344 241520 571356
rect 241572 571344 241578 571396
rect 242066 571344 242072 571396
rect 242124 571384 242130 571396
rect 242894 571384 242900 571396
rect 242124 571356 242900 571384
rect 242124 571344 242130 571356
rect 242894 571344 242900 571356
rect 242952 571344 242958 571396
rect 254854 571384 254860 571396
rect 253952 571356 254860 571384
rect 253952 571328 253980 571356
rect 254854 571344 254860 571356
rect 254912 571344 254918 571396
rect 255314 571344 255320 571396
rect 255372 571384 255378 571396
rect 256050 571384 256056 571396
rect 255372 571356 256056 571384
rect 255372 571344 255378 571356
rect 256050 571344 256056 571356
rect 256108 571344 256114 571396
rect 256694 571344 256700 571396
rect 256752 571384 256758 571396
rect 257338 571384 257344 571396
rect 256752 571356 257344 571384
rect 256752 571344 256758 571356
rect 257338 571344 257344 571356
rect 257396 571344 257402 571396
rect 263410 571344 263416 571396
rect 263468 571384 263474 571396
rect 264606 571384 264612 571396
rect 263468 571356 264612 571384
rect 263468 571344 263474 571356
rect 264606 571344 264612 571356
rect 264664 571344 264670 571396
rect 264882 571344 264888 571396
rect 264940 571384 264946 571396
rect 265894 571384 265900 571396
rect 264940 571356 265900 571384
rect 264940 571344 264946 571356
rect 265894 571344 265900 571356
rect 265952 571344 265958 571396
rect 266262 571344 266268 571396
rect 266320 571384 266326 571396
rect 267090 571384 267096 571396
rect 266320 571356 267096 571384
rect 266320 571344 266326 571356
rect 267090 571344 267096 571356
rect 267148 571344 267154 571396
rect 268930 571344 268936 571396
rect 268988 571384 268994 571396
rect 269482 571384 269488 571396
rect 268988 571356 269488 571384
rect 268988 571344 268994 571356
rect 269482 571344 269488 571356
rect 269540 571344 269546 571396
rect 270402 571344 270408 571396
rect 270460 571384 270466 571396
rect 271966 571384 271972 571396
rect 270460 571356 271972 571384
rect 270460 571344 270466 571356
rect 271966 571344 271972 571356
rect 272024 571344 272030 571396
rect 273162 571344 273168 571396
rect 273220 571384 273226 571396
rect 274634 571384 274640 571396
rect 273220 571356 274640 571384
rect 273220 571344 273226 571356
rect 274634 571344 274640 571356
rect 274692 571344 274698 571396
rect 275922 571344 275928 571396
rect 275980 571384 275986 571396
rect 278038 571384 278044 571396
rect 275980 571356 278044 571384
rect 275980 571344 275986 571356
rect 278038 571344 278044 571356
rect 278096 571344 278102 571396
rect 278590 571344 278596 571396
rect 278648 571384 278654 571396
rect 280522 571384 280528 571396
rect 278648 571356 280528 571384
rect 278648 571344 278654 571356
rect 280522 571344 280528 571356
rect 280580 571344 280586 571396
rect 28994 571276 29000 571328
rect 29052 571316 29058 571328
rect 31846 571316 31852 571328
rect 29052 571288 31852 571316
rect 29052 571276 29058 571288
rect 31846 571276 31852 571288
rect 31904 571276 31910 571328
rect 253934 571276 253940 571328
rect 253992 571276 253998 571328
rect 30282 570596 30288 570648
rect 30340 570636 30346 570648
rect 74534 570636 74540 570648
rect 30340 570608 74540 570636
rect 30340 570596 30346 570608
rect 74534 570596 74540 570608
rect 74592 570596 74598 570648
rect 30009 570503 30067 570509
rect 30009 570469 30021 570503
rect 30055 570500 30067 570503
rect 30282 570500 30288 570512
rect 30055 570472 30288 570500
rect 30055 570469 30067 570472
rect 30009 570463 30067 570469
rect 30282 570460 30288 570472
rect 30340 570460 30346 570512
rect 28629 570163 28687 570169
rect 28629 570129 28641 570163
rect 28675 570160 28687 570163
rect 31754 570160 31760 570172
rect 28675 570132 31760 570160
rect 28675 570129 28687 570132
rect 28629 570123 28687 570129
rect 31754 570120 31760 570132
rect 31812 570120 31818 570172
rect 28994 569984 29000 570036
rect 29052 570024 29058 570036
rect 29638 570024 29644 570036
rect 29052 569996 29644 570024
rect 29052 569984 29058 569996
rect 29638 569984 29644 569996
rect 29696 569984 29702 570036
rect 318518 569916 318524 569968
rect 318576 569956 318582 569968
rect 318702 569956 318708 569968
rect 318576 569928 318708 569956
rect 318576 569916 318582 569928
rect 318702 569916 318708 569928
rect 318760 569916 318766 569968
rect 354398 569916 354404 569968
rect 354456 569956 354462 569968
rect 354582 569956 354588 569968
rect 354456 569928 354588 569956
rect 354456 569916 354462 569928
rect 354582 569916 354588 569928
rect 354640 569916 354646 569968
rect 553302 569916 553308 569968
rect 553360 569956 553366 569968
rect 572714 569956 572720 569968
rect 553360 569928 572720 569956
rect 553360 569916 553366 569928
rect 572714 569916 572720 569928
rect 572772 569916 572778 569968
rect 112530 569848 112536 569900
rect 112588 569888 112594 569900
rect 138658 569888 138664 569900
rect 112588 569860 138664 569888
rect 112588 569848 112594 569860
rect 138658 569848 138664 569860
rect 138716 569848 138722 569900
rect 282270 569848 282276 569900
rect 282328 569888 282334 569900
rect 284294 569888 284300 569900
rect 282328 569860 284300 569888
rect 282328 569848 282334 569860
rect 284294 569848 284300 569860
rect 284352 569848 284358 569900
rect 30190 569236 30196 569288
rect 30248 569276 30254 569288
rect 78674 569276 78680 569288
rect 30248 569248 78680 569276
rect 30248 569236 30254 569248
rect 78674 569236 78680 569248
rect 78732 569236 78738 569288
rect 56410 569168 56416 569220
rect 56468 569208 56474 569220
rect 281534 569208 281540 569220
rect 56468 569180 281540 569208
rect 56468 569168 56474 569180
rect 281534 569168 281540 569180
rect 281592 569208 281598 569220
rect 282270 569208 282276 569220
rect 281592 569180 282276 569208
rect 281592 569168 281598 569180
rect 282270 569168 282276 569180
rect 282328 569168 282334 569220
rect 286318 569168 286324 569220
rect 286376 569208 286382 569220
rect 580442 569208 580448 569220
rect 286376 569180 580448 569208
rect 286376 569168 286382 569180
rect 580442 569168 580448 569180
rect 580500 569168 580506 569220
rect 327534 568488 327540 568540
rect 327592 568528 327598 568540
rect 328270 568528 328276 568540
rect 327592 568500 328276 568528
rect 327592 568488 327598 568500
rect 328270 568488 328276 568500
rect 328328 568488 328334 568540
rect 338298 568488 338304 568540
rect 338356 568528 338362 568540
rect 339310 568528 339316 568540
rect 338356 568500 339316 568528
rect 338356 568488 338362 568500
rect 339310 568488 339316 568500
rect 339368 568488 339374 568540
rect 346118 568488 346124 568540
rect 346176 568528 346182 568540
rect 408218 568528 408224 568540
rect 346176 568500 408224 568528
rect 346176 568488 346182 568500
rect 408218 568488 408224 568500
rect 408276 568488 408282 568540
rect 456058 568488 456064 568540
rect 456116 568528 456122 568540
rect 483014 568528 483020 568540
rect 456116 568500 483020 568528
rect 456116 568488 456122 568500
rect 483014 568488 483020 568500
rect 483072 568488 483078 568540
rect 529014 568488 529020 568540
rect 529072 568528 529078 568540
rect 529842 568528 529848 568540
rect 529072 568500 529848 568528
rect 529072 568488 529078 568500
rect 529842 568488 529848 568500
rect 529900 568488 529906 568540
rect 329374 568420 329380 568472
rect 329432 568460 329438 568472
rect 392026 568460 392032 568472
rect 329432 568432 392032 568460
rect 329432 568420 329438 568432
rect 392026 568420 392032 568432
rect 392084 568420 392090 568472
rect 343542 568352 343548 568404
rect 343600 568392 343606 568404
rect 411806 568392 411812 568404
rect 343600 568364 411812 568392
rect 343600 568352 343606 568364
rect 411806 568352 411812 568364
rect 411864 568352 411870 568404
rect 325786 568284 325792 568336
rect 325844 568324 325850 568336
rect 394878 568324 394884 568336
rect 325844 568296 394884 568324
rect 325844 568284 325850 568296
rect 394878 568284 394884 568296
rect 394936 568284 394942 568336
rect 341978 568216 341984 568268
rect 342036 568256 342042 568268
rect 415394 568256 415400 568268
rect 342036 568228 415400 568256
rect 342036 568216 342042 568228
rect 415394 568216 415400 568228
rect 415452 568216 415458 568268
rect 339402 568148 339408 568200
rect 339460 568188 339466 568200
rect 418982 568188 418988 568200
rect 339460 568160 418988 568188
rect 339460 568148 339466 568160
rect 418982 568148 418988 568160
rect 419040 568148 419046 568200
rect 336550 568080 336556 568132
rect 336608 568120 336614 568132
rect 422570 568120 422576 568132
rect 336608 568092 422576 568120
rect 336608 568080 336614 568092
rect 422570 568080 422576 568092
rect 422628 568080 422634 568132
rect 335262 568012 335268 568064
rect 335320 568052 335326 568064
rect 426158 568052 426164 568064
rect 335320 568024 426164 568052
rect 335320 568012 335326 568024
rect 426158 568012 426164 568024
rect 426216 568012 426222 568064
rect 332410 567944 332416 567996
rect 332468 567984 332474 567996
rect 429746 567984 429752 567996
rect 332468 567956 429752 567984
rect 332468 567944 332474 567956
rect 429746 567944 429752 567956
rect 429804 567944 429810 567996
rect 29270 567876 29276 567928
rect 29328 567916 29334 567928
rect 56594 567916 56600 567928
rect 29328 567888 56600 567916
rect 29328 567876 29334 567888
rect 56594 567876 56600 567888
rect 56652 567876 56658 567928
rect 331122 567876 331128 567928
rect 331180 567916 331186 567928
rect 433334 567916 433340 567928
rect 331180 567888 433340 567916
rect 331180 567876 331186 567888
rect 433334 567876 433340 567888
rect 433392 567876 433398 567928
rect 29454 567808 29460 567860
rect 29512 567848 29518 567860
rect 66346 567848 66352 567860
rect 29512 567820 66352 567848
rect 29512 567808 29518 567820
rect 66346 567808 66352 567820
rect 66404 567808 66410 567860
rect 328362 567808 328368 567860
rect 328420 567848 328426 567860
rect 436922 567848 436928 567860
rect 328420 567820 436928 567848
rect 328420 567808 328426 567820
rect 436922 567808 436928 567820
rect 436980 567808 436986 567860
rect 347682 567740 347688 567792
rect 347740 567780 347746 567792
rect 404630 567780 404636 567792
rect 347740 567752 404636 567780
rect 347740 567740 347746 567752
rect 404630 567740 404636 567752
rect 404688 567740 404694 567792
rect 332962 567672 332968 567724
rect 333020 567712 333026 567724
rect 389174 567712 389180 567724
rect 333020 567684 389180 567712
rect 333020 567672 333026 567684
rect 389174 567672 389180 567684
rect 389232 567672 389238 567724
rect 336458 567604 336464 567656
rect 336516 567644 336522 567656
rect 387794 567644 387800 567656
rect 336516 567616 387800 567644
rect 336516 567604 336522 567616
rect 387794 567604 387800 567616
rect 387852 567604 387858 567656
rect 350442 567536 350448 567588
rect 350500 567576 350506 567588
rect 401042 567576 401048 567588
rect 350500 567548 401048 567576
rect 350500 567536 350506 567548
rect 401042 567536 401048 567548
rect 401100 567536 401106 567588
rect 351730 567468 351736 567520
rect 351788 567508 351794 567520
rect 397454 567508 397460 567520
rect 351788 567480 397460 567508
rect 351788 567468 351794 567480
rect 397454 567468 397460 567480
rect 397512 567468 397518 567520
rect 340138 567400 340144 567452
rect 340196 567440 340202 567452
rect 385034 567440 385040 567452
rect 340196 567412 385040 567440
rect 340196 567400 340202 567412
rect 385034 567400 385040 567412
rect 385092 567400 385098 567452
rect 343726 567332 343732 567384
rect 343784 567372 343790 567384
rect 383654 567372 383660 567384
rect 343784 567344 383660 567372
rect 343784 567332 343790 567344
rect 383654 567332 383660 567344
rect 383712 567332 383718 567384
rect 347314 567264 347320 567316
rect 347372 567304 347378 567316
rect 380986 567304 380992 567316
rect 347372 567276 380992 567304
rect 347372 567264 347378 567276
rect 380986 567264 380992 567276
rect 381044 567264 381050 567316
rect 3510 567196 3516 567248
rect 3568 567236 3574 567248
rect 9122 567236 9128 567248
rect 3568 567208 9128 567236
rect 3568 567196 3574 567208
rect 9122 567196 9128 567208
rect 9180 567196 9186 567248
rect 28813 567239 28871 567245
rect 28813 567205 28825 567239
rect 28859 567236 28871 567239
rect 29086 567236 29092 567248
rect 28859 567208 29092 567236
rect 28859 567205 28871 567208
rect 28813 567199 28871 567205
rect 29086 567196 29092 567208
rect 29144 567196 29150 567248
rect 320358 567196 320364 567248
rect 320416 567236 320422 567248
rect 321462 567236 321468 567248
rect 320416 567208 321468 567236
rect 320416 567196 320422 567208
rect 321462 567196 321468 567208
rect 321520 567196 321526 567248
rect 350902 567196 350908 567248
rect 350960 567236 350966 567248
rect 350960 567208 356192 567236
rect 350960 567196 350966 567208
rect 356164 567168 356192 567208
rect 356238 567196 356244 567248
rect 356296 567236 356302 567248
rect 357342 567236 357348 567248
rect 356296 567208 357348 567236
rect 356296 567196 356302 567208
rect 357342 567196 357348 567208
rect 357400 567196 357406 567248
rect 357452 567208 358768 567236
rect 357452 567168 357480 567208
rect 356164 567140 357480 567168
rect 358740 567168 358768 567208
rect 358814 567196 358820 567248
rect 358872 567236 358878 567248
rect 359826 567236 359832 567248
rect 358872 567208 359832 567236
rect 358872 567196 358878 567208
rect 359826 567196 359832 567208
rect 359884 567196 359890 567248
rect 379514 567236 379520 567248
rect 359936 567208 379520 567236
rect 359936 567168 359964 567208
rect 379514 567196 379520 567208
rect 379572 567196 379578 567248
rect 358740 567140 359964 567168
rect 29362 566448 29368 566500
rect 29420 566488 29426 566500
rect 60826 566488 60832 566500
rect 29420 566460 60832 566488
rect 29420 566448 29426 566460
rect 60826 566448 60832 566460
rect 60884 566448 60890 566500
rect 361574 566448 361580 566500
rect 361632 566488 361638 566500
rect 372614 566488 372620 566500
rect 361632 566460 372620 566488
rect 361632 566448 361638 566460
rect 372614 566448 372620 566460
rect 372672 566448 372678 566500
rect 368382 565836 368388 565888
rect 368440 565876 368446 565888
rect 369854 565876 369860 565888
rect 368440 565848 369860 565876
rect 368440 565836 368446 565848
rect 369854 565836 369860 565848
rect 369912 565836 369918 565888
rect 29086 565156 29092 565208
rect 29144 565196 29150 565208
rect 49694 565196 49700 565208
rect 29144 565168 49700 565196
rect 29144 565156 29150 565168
rect 49694 565156 49700 565168
rect 49752 565156 49758 565208
rect 358078 565156 358084 565208
rect 358136 565196 358142 565208
rect 358136 565168 364380 565196
rect 358136 565156 358142 565168
rect 29546 565088 29552 565140
rect 29604 565128 29610 565140
rect 63494 565128 63500 565140
rect 29604 565100 63500 565128
rect 29604 565088 29610 565100
rect 63494 565088 63500 565100
rect 63552 565088 63558 565140
rect 364352 565128 364380 565168
rect 375558 565128 375564 565140
rect 364352 565100 375564 565128
rect 375558 565088 375564 565100
rect 375616 565088 375622 565140
rect 29914 563660 29920 563712
rect 29972 563700 29978 563712
rect 67634 563700 67640 563712
rect 29972 563672 67640 563700
rect 29972 563660 29978 563672
rect 67634 563660 67640 563672
rect 67692 563660 67698 563712
rect 355870 563660 355876 563712
rect 355928 563700 355934 563712
rect 389266 563700 389272 563712
rect 355928 563672 389272 563700
rect 355928 563660 355934 563672
rect 389266 563660 389272 563672
rect 389324 563660 389330 563712
rect 29178 563524 29184 563576
rect 29236 563564 29242 563576
rect 29914 563564 29920 563576
rect 29236 563536 29920 563564
rect 29236 563524 29242 563536
rect 29914 563524 29920 563536
rect 29972 563524 29978 563576
rect 364334 563048 364340 563100
rect 364392 563088 364398 563100
rect 369854 563088 369860 563100
rect 364392 563060 369860 563088
rect 364392 563048 364398 563060
rect 369854 563048 369860 563060
rect 369912 563048 369918 563100
rect 30282 562300 30288 562352
rect 30340 562340 30346 562352
rect 71774 562340 71780 562352
rect 30340 562312 71780 562340
rect 30340 562300 30346 562312
rect 71774 562300 71780 562312
rect 71832 562300 71838 562352
rect 362954 562300 362960 562352
rect 363012 562340 363018 562352
rect 364242 562340 364248 562352
rect 363012 562312 364248 562340
rect 363012 562300 363018 562312
rect 364242 562300 364248 562312
rect 364300 562300 364306 562352
rect 365714 562300 365720 562352
rect 365772 562340 365778 562352
rect 367002 562340 367008 562352
rect 365772 562312 367008 562340
rect 365772 562300 365778 562312
rect 367002 562300 367008 562312
rect 367060 562300 367066 562352
rect 375374 562340 375380 562352
rect 367204 562312 375380 562340
rect 365622 562232 365628 562284
rect 365680 562272 365686 562284
rect 367204 562272 367232 562312
rect 375374 562300 375380 562312
rect 375432 562300 375438 562352
rect 365680 562244 367232 562272
rect 365680 562232 365686 562244
rect 29822 560940 29828 560992
rect 29880 560980 29886 560992
rect 86954 560980 86960 560992
rect 29880 560952 86960 560980
rect 29880 560940 29886 560952
rect 86954 560940 86960 560952
rect 87012 560940 87018 560992
rect 362862 560940 362868 560992
rect 362920 560980 362926 560992
rect 379606 560980 379612 560992
rect 362920 560952 379612 560980
rect 362920 560940 362926 560952
rect 379606 560940 379612 560952
rect 379664 560940 379670 560992
rect 283190 560260 283196 560312
rect 283248 560300 283254 560312
rect 283282 560300 283288 560312
rect 283248 560272 283288 560300
rect 283248 560260 283254 560272
rect 283282 560260 283288 560272
rect 283340 560260 283346 560312
rect 358814 558152 358820 558204
rect 358872 558192 358878 558204
rect 360102 558192 360108 558204
rect 358872 558164 360108 558192
rect 358872 558152 358878 558164
rect 360102 558152 360108 558164
rect 360160 558152 360166 558204
rect 304258 556180 304264 556232
rect 304316 556220 304322 556232
rect 580166 556220 580172 556232
rect 304316 556192 580172 556220
rect 304316 556180 304322 556192
rect 580166 556180 580172 556192
rect 580224 556180 580230 556232
rect 364242 554004 364248 554056
rect 364300 554044 364306 554056
rect 371234 554044 371240 554056
rect 364300 554016 371240 554044
rect 364300 554004 364306 554016
rect 371234 554004 371240 554016
rect 371292 554004 371298 554056
rect 317322 552644 317328 552696
rect 317380 552684 317386 552696
rect 400306 552684 400312 552696
rect 317380 552656 400312 552684
rect 317380 552644 317386 552656
rect 400306 552644 400312 552656
rect 400364 552644 400370 552696
rect 3142 552032 3148 552084
rect 3200 552072 3206 552084
rect 279510 552072 279516 552084
rect 3200 552044 279516 552072
rect 3200 552032 3206 552044
rect 279510 552032 279516 552044
rect 279568 552032 279574 552084
rect 29546 551284 29552 551336
rect 29604 551324 29610 551336
rect 95234 551324 95240 551336
rect 29604 551296 95240 551324
rect 29604 551284 29610 551296
rect 95234 551284 95240 551296
rect 95292 551284 95298 551336
rect 543642 547204 543648 547256
rect 543700 547244 543706 547256
rect 553118 547244 553124 547256
rect 543700 547216 553124 547244
rect 543700 547204 543706 547216
rect 553118 547204 553124 547216
rect 553176 547204 553182 547256
rect 540882 547136 540888 547188
rect 540940 547176 540946 547188
rect 553026 547176 553032 547188
rect 540940 547148 553032 547176
rect 540940 547136 540946 547148
rect 553026 547136 553032 547148
rect 553084 547136 553090 547188
rect 545022 547068 545028 547120
rect 545080 547108 545086 547120
rect 553210 547108 553216 547120
rect 545080 547080 553216 547108
rect 545080 547068 545086 547080
rect 553210 547068 553216 547080
rect 553268 547068 553274 547120
rect 366910 546456 366916 546508
rect 366968 546496 366974 546508
rect 371326 546496 371332 546508
rect 366968 546468 371332 546496
rect 366968 546456 366974 546468
rect 371326 546456 371332 546468
rect 371384 546456 371390 546508
rect 354490 542988 354496 543040
rect 354548 543028 354554 543040
rect 393314 543028 393320 543040
rect 354548 543000 393320 543028
rect 354548 542988 354554 543000
rect 393314 542988 393320 543000
rect 393372 542988 393378 543040
rect 322842 541628 322848 541680
rect 322900 541668 322906 541680
rect 396074 541668 396080 541680
rect 322900 541640 396080 541668
rect 322900 541628 322906 541640
rect 396074 541628 396080 541640
rect 396132 541628 396138 541680
rect 282914 540948 282920 541000
rect 282972 540988 282978 541000
rect 283190 540988 283196 541000
rect 282972 540960 283196 540988
rect 282972 540948 282978 540960
rect 283190 540948 283196 540960
rect 283248 540948 283254 541000
rect 358722 540200 358728 540252
rect 358780 540240 358786 540252
rect 386414 540240 386420 540252
rect 358780 540212 386420 540240
rect 358780 540200 358786 540212
rect 386414 540200 386420 540212
rect 386472 540200 386478 540252
rect 366818 538840 366824 538892
rect 366876 538880 366882 538892
rect 373994 538880 374000 538892
rect 366876 538852 374000 538880
rect 366876 538840 366882 538852
rect 373994 538840 374000 538852
rect 374052 538840 374058 538892
rect 3510 538228 3516 538280
rect 3568 538268 3574 538280
rect 10410 538268 10416 538280
rect 3568 538240 10416 538268
rect 3568 538228 3574 538240
rect 10410 538228 10416 538240
rect 10468 538228 10474 538280
rect 360102 537480 360108 537532
rect 360160 537520 360166 537532
rect 374086 537520 374092 537532
rect 360160 537492 374092 537520
rect 360160 537480 360166 537492
rect 374086 537480 374092 537492
rect 374144 537480 374150 537532
rect 357158 536120 357164 536172
rect 357216 536160 357222 536172
rect 376110 536160 376116 536172
rect 357216 536132 376116 536160
rect 357216 536120 357222 536132
rect 376110 536120 376116 536132
rect 376168 536120 376174 536172
rect 360562 536052 360568 536104
rect 360620 536092 360626 536104
rect 382274 536092 382280 536104
rect 360620 536064 382280 536092
rect 360620 536052 360626 536064
rect 382274 536052 382280 536064
rect 382332 536052 382338 536104
rect 26602 535616 26608 535628
rect 26563 535588 26608 535616
rect 26602 535576 26608 535588
rect 26660 535576 26666 535628
rect 26786 535440 26792 535492
rect 26844 535440 26850 535492
rect 26804 535288 26832 535440
rect 26786 535236 26792 535288
rect 26844 535236 26850 535288
rect 367002 535236 367008 535288
rect 367060 535276 367066 535288
rect 369854 535276 369860 535288
rect 367060 535248 369860 535276
rect 367060 535236 367066 535248
rect 369854 535236 369860 535248
rect 369912 535236 369918 535288
rect 353202 535168 353208 535220
rect 353260 535208 353266 535220
rect 378226 535208 378232 535220
rect 353260 535180 378232 535208
rect 353260 535168 353266 535180
rect 378226 535168 378232 535180
rect 378284 535168 378290 535220
rect 152458 535100 152464 535152
rect 152516 535140 152522 535152
rect 436002 535140 436008 535152
rect 152516 535112 436008 535140
rect 152516 535100 152522 535112
rect 436002 535100 436008 535112
rect 436060 535100 436066 535152
rect 156322 535032 156328 535084
rect 156380 535072 156386 535084
rect 446122 535072 446128 535084
rect 156380 535044 446128 535072
rect 156380 535032 156386 535044
rect 446122 535032 446128 535044
rect 446180 535032 446186 535084
rect 26605 535007 26663 535013
rect 26605 534973 26617 535007
rect 26651 535004 26663 535007
rect 27062 535004 27068 535016
rect 26651 534976 27068 535004
rect 26651 534973 26663 534976
rect 26605 534967 26663 534973
rect 27062 534964 27068 534976
rect 27120 534964 27126 535016
rect 148134 534964 148140 535016
rect 148192 535004 148198 535016
rect 442902 535004 442908 535016
rect 148192 534976 442908 535004
rect 148192 534964 148198 534976
rect 442902 534964 442908 534976
rect 442960 534964 442966 535016
rect 147950 534896 147956 534948
rect 148008 534936 148014 534948
rect 450446 534936 450452 534948
rect 148008 534908 450452 534936
rect 148008 534896 148014 534908
rect 450446 534896 450452 534908
rect 450504 534896 450510 534948
rect 143810 534828 143816 534880
rect 143868 534868 143874 534880
rect 452562 534868 452568 534880
rect 143868 534840 452568 534868
rect 143868 534828 143874 534840
rect 452562 534828 452568 534840
rect 452620 534828 452626 534880
rect 166994 534760 167000 534812
rect 167052 534800 167058 534812
rect 483842 534800 483848 534812
rect 167052 534772 483848 534800
rect 167052 534760 167058 534772
rect 483842 534760 483848 534772
rect 483900 534760 483906 534812
rect 139486 534692 139492 534744
rect 139544 534732 139550 534744
rect 456978 534732 456984 534744
rect 139544 534704 456984 534732
rect 139544 534692 139550 534704
rect 456978 534692 456984 534704
rect 457036 534692 457042 534744
rect 137370 534624 137376 534676
rect 137428 534664 137434 534676
rect 459094 534664 459100 534676
rect 137428 534636 459100 534664
rect 137428 534624 137434 534636
rect 459094 534624 459100 534636
rect 459152 534624 459158 534676
rect 135254 534556 135260 534608
rect 135312 534596 135318 534608
rect 461210 534596 461216 534608
rect 135312 534568 461216 534596
rect 135312 534556 135318 534568
rect 461210 534556 461216 534568
rect 461268 534556 461274 534608
rect 131942 534488 131948 534540
rect 132000 534528 132006 534540
rect 464522 534528 464528 534540
rect 132000 534500 464528 534528
rect 132000 534488 132006 534500
rect 464522 534488 464528 534500
rect 464580 534488 464586 534540
rect 129826 534420 129832 534472
rect 129884 534460 129890 534472
rect 466638 534460 466644 534472
rect 129884 534432 466644 534460
rect 129884 534420 129890 534432
rect 466638 534420 466644 534432
rect 466696 534420 466702 534472
rect 127710 534352 127716 534404
rect 127768 534392 127774 534404
rect 468754 534392 468760 534404
rect 127768 534364 468760 534392
rect 127768 534352 127774 534364
rect 468754 534352 468760 534364
rect 468812 534352 468818 534404
rect 125502 534284 125508 534336
rect 125560 534324 125566 534336
rect 470962 534324 470968 534336
rect 125560 534296 470968 534324
rect 125560 534284 125566 534296
rect 470962 534284 470968 534296
rect 471020 534284 471026 534336
rect 123386 534216 123392 534268
rect 123444 534256 123450 534268
rect 473446 534256 473452 534268
rect 123444 534228 473452 534256
rect 123444 534216 123450 534228
rect 473446 534216 473452 534228
rect 473504 534216 473510 534268
rect 121178 534148 121184 534200
rect 121236 534188 121242 534200
rect 475286 534188 475292 534200
rect 121236 534160 475292 534188
rect 121236 534148 121242 534160
rect 475286 534148 475292 534160
rect 475344 534148 475350 534200
rect 111058 534080 111064 534132
rect 111116 534120 111122 534132
rect 487154 534120 487160 534132
rect 111116 534092 487160 534120
rect 111116 534080 111122 534092
rect 487154 534080 487160 534092
rect 487212 534080 487218 534132
rect 339310 534012 339316 534064
rect 339368 534052 339374 534064
rect 386874 534052 386880 534064
rect 339368 534024 386880 534052
rect 339368 534012 339374 534024
rect 386874 534012 386880 534024
rect 386932 534012 386938 534064
rect 335170 533944 335176 533996
rect 335228 533984 335234 533996
rect 389174 533984 389180 533996
rect 335228 533956 389180 533984
rect 335228 533944 335234 533956
rect 389174 533944 389180 533956
rect 389232 533944 389238 533996
rect 26142 533876 26148 533928
rect 26200 533916 26206 533928
rect 34974 533916 34980 533928
rect 26200 533888 34980 533916
rect 26200 533876 26206 533888
rect 34974 533876 34980 533888
rect 35032 533876 35038 533928
rect 331030 533876 331036 533928
rect 331088 533916 331094 533928
rect 391198 533916 391204 533928
rect 331088 533888 391204 533916
rect 331088 533876 331094 533888
rect 391198 533876 391204 533888
rect 391256 533876 391262 533928
rect 25038 533808 25044 533860
rect 25096 533848 25102 533860
rect 37182 533848 37188 533860
rect 25096 533820 37188 533848
rect 25096 533808 25102 533820
rect 37182 533808 37188 533820
rect 37240 533808 37246 533860
rect 328270 533808 328276 533860
rect 328328 533848 328334 533860
rect 393314 533848 393320 533860
rect 328328 533820 393320 533848
rect 328328 533808 328334 533820
rect 393314 533808 393320 533820
rect 393372 533808 393378 533860
rect 25130 533740 25136 533792
rect 25188 533780 25194 533792
rect 39298 533780 39304 533792
rect 25188 533752 39304 533780
rect 25188 533740 25194 533752
rect 39298 533740 39304 533752
rect 39356 533740 39362 533792
rect 318702 533740 318708 533792
rect 318760 533780 318766 533792
rect 398926 533780 398932 533792
rect 318760 533752 398932 533780
rect 318760 533740 318766 533752
rect 398926 533740 398932 533752
rect 398984 533740 398990 533792
rect 25222 533672 25228 533724
rect 25280 533712 25286 533724
rect 41414 533712 41420 533724
rect 25280 533684 41420 533712
rect 25280 533672 25286 533684
rect 41414 533672 41420 533684
rect 41472 533672 41478 533724
rect 323946 533672 323952 533724
rect 324004 533712 324010 533724
rect 442994 533712 443000 533724
rect 324004 533684 443000 533712
rect 324004 533672 324010 533684
rect 442994 533672 443000 533684
rect 443052 533672 443058 533724
rect 25314 533604 25320 533656
rect 25372 533644 25378 533656
rect 43622 533644 43628 533656
rect 25372 533616 43628 533644
rect 25372 533604 25378 533616
rect 43622 533604 43628 533616
rect 43680 533604 43686 533656
rect 322842 533604 322848 533656
rect 322900 533644 322906 533656
rect 445754 533644 445760 533656
rect 322900 533616 445760 533644
rect 322900 533604 322906 533616
rect 445754 533604 445760 533616
rect 445812 533604 445818 533656
rect 530854 533604 530860 533656
rect 530912 533644 530918 533656
rect 551462 533644 551468 533656
rect 530912 533616 551468 533644
rect 530912 533604 530918 533616
rect 551462 533604 551468 533616
rect 551520 533604 551526 533656
rect 27154 533536 27160 533588
rect 27212 533536 27218 533588
rect 29730 533536 29736 533588
rect 29788 533576 29794 533588
rect 56502 533576 56508 533588
rect 29788 533548 56508 533576
rect 29788 533536 29794 533548
rect 56502 533536 56508 533548
rect 56560 533536 56566 533588
rect 321278 533536 321284 533588
rect 321336 533576 321342 533588
rect 447134 533576 447140 533588
rect 321336 533548 447140 533576
rect 321336 533536 321342 533548
rect 447134 533536 447140 533548
rect 447192 533536 447198 533588
rect 514662 533536 514668 533588
rect 514720 533576 514726 533588
rect 552290 533576 552296 533588
rect 514720 533548 552296 533576
rect 514720 533536 514726 533548
rect 552290 533536 552296 533548
rect 552348 533536 552354 533588
rect 27172 533440 27200 533536
rect 27246 533468 27252 533520
rect 27304 533508 27310 533520
rect 84562 533508 84568 533520
rect 27304 533480 84568 533508
rect 27304 533468 27310 533480
rect 84562 533468 84568 533480
rect 84620 533468 84626 533520
rect 320726 533468 320732 533520
rect 320784 533508 320790 533520
rect 448514 533508 448520 533520
rect 320784 533480 448520 533508
rect 320784 533468 320790 533480
rect 448514 533468 448520 533480
rect 448572 533468 448578 533520
rect 512546 533468 512552 533520
rect 512604 533508 512610 533520
rect 552198 533508 552204 533520
rect 512604 533480 552204 533508
rect 512604 533468 512610 533480
rect 552198 533468 552204 533480
rect 552256 533468 552262 533520
rect 86678 533440 86684 533452
rect 27172 533412 86684 533440
rect 86678 533400 86684 533412
rect 86736 533400 86742 533452
rect 319622 533400 319628 533452
rect 319680 533440 319686 533452
rect 451274 533440 451280 533452
rect 319680 533412 451280 533440
rect 319680 533400 319686 533412
rect 451274 533400 451280 533412
rect 451332 533400 451338 533452
rect 510430 533400 510436 533452
rect 510488 533440 510494 533452
rect 552014 533440 552020 533452
rect 510488 533412 552020 533440
rect 510488 533400 510494 533412
rect 552014 533400 552020 533412
rect 552072 533400 552078 533452
rect 26234 533332 26240 533384
rect 26292 533372 26298 533384
rect 27062 533372 27068 533384
rect 26292 533344 27068 533372
rect 26292 533332 26298 533344
rect 27062 533332 27068 533344
rect 27120 533332 27126 533384
rect 27706 533332 27712 533384
rect 27764 533372 27770 533384
rect 91002 533372 91008 533384
rect 27764 533344 91008 533372
rect 27764 533332 27770 533344
rect 91002 533332 91008 533344
rect 91060 533332 91066 533384
rect 266722 533332 266728 533384
rect 266780 533372 266786 533384
rect 267642 533372 267648 533384
rect 266780 533344 267648 533372
rect 266780 533332 266786 533344
rect 267642 533332 267648 533344
rect 267700 533332 267706 533384
rect 318518 533332 318524 533384
rect 318576 533372 318582 533384
rect 452654 533372 452660 533384
rect 318576 533344 452660 533372
rect 318576 533332 318582 533344
rect 452654 533332 452660 533344
rect 452712 533332 452718 533384
rect 529842 533332 529848 533384
rect 529900 533372 529906 533384
rect 574370 533372 574376 533384
rect 529900 533344 574376 533372
rect 529900 533332 529906 533344
rect 574370 533332 574376 533344
rect 574428 533332 574434 533384
rect 342070 533264 342076 533316
rect 342128 533304 342134 533316
rect 385126 533304 385132 533316
rect 342128 533276 385132 533304
rect 342128 533264 342134 533276
rect 385126 533264 385132 533276
rect 385184 533264 385190 533316
rect 346210 533196 346216 533248
rect 346268 533236 346274 533248
rect 382550 533236 382556 533248
rect 346268 533208 382556 533236
rect 346268 533196 346274 533208
rect 382550 533196 382556 533208
rect 382608 533196 382614 533248
rect 349062 533128 349068 533180
rect 349120 533168 349126 533180
rect 380434 533168 380440 533180
rect 349120 533140 380440 533168
rect 349120 533128 349126 533140
rect 380434 533128 380440 533140
rect 380492 533128 380498 533180
rect 354582 533060 354588 533112
rect 354640 533100 354646 533112
rect 377214 533100 377220 533112
rect 354640 533072 377220 533100
rect 354640 533060 354646 533072
rect 377214 533060 377220 533072
rect 377272 533060 377278 533112
rect 193398 532992 193404 533044
rect 193456 533032 193462 533044
rect 403066 533032 403072 533044
rect 193456 533004 403072 533032
rect 193456 532992 193462 533004
rect 403066 532992 403072 533004
rect 403124 532992 403130 533044
rect 192386 532924 192392 532976
rect 192444 532964 192450 532976
rect 404446 532964 404452 532976
rect 192444 532936 404452 532964
rect 192444 532924 192450 532936
rect 404446 532924 404452 532936
rect 404504 532924 404510 532976
rect 189074 532856 189080 532908
rect 189132 532896 189138 532908
rect 407390 532896 407396 532908
rect 189132 532868 407396 532896
rect 189132 532856 189138 532868
rect 407390 532856 407396 532868
rect 407448 532856 407454 532908
rect 183738 532788 183744 532840
rect 183796 532828 183802 532840
rect 412726 532828 412732 532840
rect 183796 532800 412732 532828
rect 183796 532788 183802 532800
rect 412726 532788 412732 532800
rect 412784 532788 412790 532840
rect 177298 532720 177304 532772
rect 177356 532760 177362 532772
rect 419626 532760 419632 532772
rect 177356 532732 419632 532760
rect 177356 532720 177362 532732
rect 419626 532720 419632 532732
rect 419684 532720 419690 532772
rect 28718 532652 28724 532704
rect 28776 532692 28782 532704
rect 33870 532692 33876 532704
rect 28776 532664 33876 532692
rect 28776 532652 28782 532664
rect 33870 532652 33876 532664
rect 33928 532652 33934 532704
rect 33965 532695 34023 532701
rect 33965 532661 33977 532695
rect 34011 532692 34023 532695
rect 42518 532692 42524 532704
rect 34011 532664 42524 532692
rect 34011 532661 34023 532664
rect 33965 532655 34023 532661
rect 42518 532652 42524 532664
rect 42576 532652 42582 532704
rect 344370 532652 344376 532704
rect 344428 532692 344434 532704
rect 409874 532692 409880 532704
rect 344428 532664 409880 532692
rect 344428 532652 344434 532664
rect 409874 532652 409880 532664
rect 409932 532652 409938 532704
rect 548337 532695 548395 532701
rect 548337 532661 548349 532695
rect 548383 532692 548395 532695
rect 554314 532692 554320 532704
rect 548383 532664 554320 532692
rect 548383 532661 548395 532664
rect 548337 532655 548395 532661
rect 554314 532652 554320 532664
rect 554372 532652 554378 532704
rect 25498 532584 25504 532636
rect 25556 532624 25562 532636
rect 45738 532624 45744 532636
rect 25556 532596 45744 532624
rect 25556 532584 25562 532596
rect 45738 532584 45744 532596
rect 45796 532584 45802 532636
rect 342162 532584 342168 532636
rect 342220 532624 342226 532636
rect 412634 532624 412640 532636
rect 342220 532596 412640 532624
rect 342220 532584 342226 532596
rect 412634 532584 412640 532596
rect 412692 532584 412698 532636
rect 547046 532584 547052 532636
rect 547104 532624 547110 532636
rect 551738 532624 551744 532636
rect 547104 532596 551744 532624
rect 547104 532584 547110 532596
rect 551738 532584 551744 532596
rect 551796 532584 551802 532636
rect 25682 532516 25688 532568
rect 25740 532556 25746 532568
rect 47946 532556 47952 532568
rect 25740 532528 47952 532556
rect 25740 532516 25746 532528
rect 47946 532516 47952 532528
rect 48004 532516 48010 532568
rect 324130 532516 324136 532568
rect 324188 532556 324194 532568
rect 395522 532556 395528 532568
rect 324188 532528 395528 532556
rect 324188 532516 324194 532528
rect 395522 532516 395528 532528
rect 395580 532516 395586 532568
rect 536282 532516 536288 532568
rect 536340 532556 536346 532568
rect 551554 532556 551560 532568
rect 536340 532528 551560 532556
rect 536340 532516 536346 532528
rect 551554 532516 551560 532528
rect 551612 532516 551618 532568
rect 21358 532448 21364 532500
rect 21416 532488 21422 532500
rect 24118 532488 24124 532500
rect 21416 532460 24124 532488
rect 21416 532448 21422 532460
rect 24118 532448 24124 532460
rect 24176 532448 24182 532500
rect 25774 532448 25780 532500
rect 25832 532488 25838 532500
rect 52270 532488 52276 532500
rect 25832 532460 52276 532488
rect 25832 532448 25838 532460
rect 52270 532448 52276 532460
rect 52328 532448 52334 532500
rect 340138 532448 340144 532500
rect 340196 532488 340202 532500
rect 416774 532488 416780 532500
rect 340196 532460 416780 532488
rect 340196 532448 340202 532460
rect 416774 532448 416780 532460
rect 416832 532448 416838 532500
rect 538122 532448 538128 532500
rect 538180 532488 538186 532500
rect 548337 532491 548395 532497
rect 548337 532488 548349 532491
rect 538180 532460 548349 532488
rect 538180 532448 538186 532460
rect 548337 532457 548349 532460
rect 548383 532457 548395 532491
rect 554130 532488 554136 532500
rect 548337 532451 548395 532457
rect 548444 532460 554136 532488
rect 28442 532380 28448 532432
rect 28500 532420 28506 532432
rect 54386 532420 54392 532432
rect 28500 532392 54392 532420
rect 28500 532380 28506 532392
rect 54386 532380 54392 532392
rect 54444 532380 54450 532432
rect 321462 532380 321468 532432
rect 321520 532420 321526 532432
rect 397638 532420 397644 532432
rect 321520 532392 397644 532420
rect 321520 532380 321526 532392
rect 397638 532380 397644 532392
rect 397696 532380 397702 532432
rect 401502 532380 401508 532432
rect 401560 532420 401566 532432
rect 455414 532420 455420 532432
rect 401560 532392 455420 532420
rect 401560 532380 401566 532392
rect 455414 532380 455420 532392
rect 455472 532380 455478 532432
rect 531958 532380 531964 532432
rect 532016 532420 532022 532432
rect 548444 532420 548472 532460
rect 554130 532448 554136 532460
rect 554188 532448 554194 532500
rect 532016 532392 548472 532420
rect 548521 532423 548579 532429
rect 532016 532380 532022 532392
rect 548521 532389 548533 532423
rect 548567 532420 548579 532423
rect 553946 532420 553952 532432
rect 548567 532392 553952 532420
rect 548567 532389 548579 532392
rect 548521 532383 548579 532389
rect 553946 532380 553952 532392
rect 554004 532380 554010 532432
rect 25866 532312 25872 532364
rect 25924 532352 25930 532364
rect 58710 532352 58716 532364
rect 25924 532324 58716 532352
rect 25924 532312 25930 532324
rect 58710 532312 58716 532324
rect 58768 532312 58774 532364
rect 337930 532312 337936 532364
rect 337988 532352 337994 532364
rect 419534 532352 419540 532364
rect 337988 532324 419540 532352
rect 337988 532312 337994 532324
rect 419534 532312 419540 532324
rect 419592 532312 419598 532364
rect 527634 532312 527640 532364
rect 527692 532352 527698 532364
rect 551370 532352 551376 532364
rect 527692 532324 551376 532352
rect 527692 532312 527698 532324
rect 551370 532312 551376 532324
rect 551428 532312 551434 532364
rect 26050 532244 26056 532296
rect 26108 532284 26114 532296
rect 60826 532284 60832 532296
rect 26108 532256 60832 532284
rect 26108 532244 26114 532256
rect 60826 532244 60832 532256
rect 60884 532244 60890 532296
rect 335814 532244 335820 532296
rect 335872 532284 335878 532296
rect 423674 532284 423680 532296
rect 335872 532256 423680 532284
rect 335872 532244 335878 532256
rect 423674 532244 423680 532256
rect 423732 532244 423738 532296
rect 529750 532244 529756 532296
rect 529808 532284 529814 532296
rect 548521 532287 548579 532293
rect 548521 532284 548533 532287
rect 529808 532256 548533 532284
rect 529808 532244 529814 532256
rect 548521 532253 548533 532256
rect 548567 532253 548579 532287
rect 553854 532284 553860 532296
rect 548521 532247 548579 532253
rect 548628 532256 553860 532284
rect 24946 532176 24952 532228
rect 25004 532216 25010 532228
rect 63034 532216 63040 532228
rect 25004 532188 63040 532216
rect 25004 532176 25010 532188
rect 63034 532176 63040 532188
rect 63092 532176 63098 532228
rect 333606 532176 333612 532228
rect 333664 532216 333670 532228
rect 427814 532216 427820 532228
rect 333664 532188 427820 532216
rect 333664 532176 333670 532188
rect 427814 532176 427820 532188
rect 427872 532176 427878 532228
rect 525518 532176 525524 532228
rect 525576 532216 525582 532228
rect 548628 532216 548656 532256
rect 553854 532244 553860 532256
rect 553912 532244 553918 532296
rect 553762 532216 553768 532228
rect 525576 532188 548656 532216
rect 548720 532188 553768 532216
rect 525576 532176 525582 532188
rect 26510 532108 26516 532160
rect 26568 532148 26574 532160
rect 33965 532151 34023 532157
rect 33965 532148 33977 532151
rect 26568 532120 33977 532148
rect 26568 532108 26574 532120
rect 33965 532117 33977 532120
rect 34011 532117 34023 532151
rect 33965 532111 34023 532117
rect 34057 532151 34115 532157
rect 34057 532117 34069 532151
rect 34103 532148 34115 532151
rect 67358 532148 67364 532160
rect 34103 532120 67364 532148
rect 34103 532117 34115 532120
rect 34057 532111 34115 532117
rect 67358 532108 67364 532120
rect 67416 532108 67422 532160
rect 331490 532108 331496 532160
rect 331548 532148 331554 532160
rect 430574 532148 430580 532160
rect 331548 532120 430580 532148
rect 331548 532108 331554 532120
rect 430574 532108 430580 532120
rect 430632 532108 430638 532160
rect 523310 532108 523316 532160
rect 523368 532148 523374 532160
rect 548720 532148 548748 532188
rect 553762 532176 553768 532188
rect 553820 532176 553826 532228
rect 523368 532120 548748 532148
rect 523368 532108 523374 532120
rect 549162 532108 549168 532160
rect 549220 532148 549226 532160
rect 551830 532148 551836 532160
rect 549220 532120 551836 532148
rect 549220 532108 549226 532120
rect 551830 532108 551836 532120
rect 551888 532108 551894 532160
rect 28166 532040 28172 532092
rect 28224 532080 28230 532092
rect 69474 532080 69480 532092
rect 28224 532052 69480 532080
rect 28224 532040 28230 532052
rect 69474 532040 69480 532052
rect 69532 532040 69538 532092
rect 329282 532040 329288 532092
rect 329340 532080 329346 532092
rect 434714 532080 434720 532092
rect 329340 532052 434720 532080
rect 329340 532040 329346 532052
rect 434714 532040 434720 532052
rect 434772 532040 434778 532092
rect 521194 532040 521200 532092
rect 521252 532080 521258 532092
rect 553578 532080 553584 532092
rect 521252 532052 553584 532080
rect 521252 532040 521258 532052
rect 553578 532040 553584 532052
rect 553636 532040 553642 532092
rect 26970 531972 26976 532024
rect 27028 532012 27034 532024
rect 75914 532012 75920 532024
rect 27028 531984 75920 532012
rect 27028 531972 27034 531984
rect 75914 531972 75920 531984
rect 75972 531972 75978 532024
rect 326982 531972 326988 532024
rect 327040 532012 327046 532024
rect 437474 532012 437480 532024
rect 327040 531984 437480 532012
rect 327040 531972 327046 531984
rect 437474 531972 437480 531984
rect 437532 531972 437538 532024
rect 518710 531972 518716 532024
rect 518768 532012 518774 532024
rect 551094 532012 551100 532024
rect 518768 531984 551100 532012
rect 518768 531972 518774 531984
rect 551094 531972 551100 531984
rect 551152 531972 551158 532024
rect 25406 531904 25412 531956
rect 25464 531944 25470 531956
rect 40402 531944 40408 531956
rect 25464 531916 40408 531944
rect 25464 531904 25470 531916
rect 40402 531904 40408 531916
rect 40460 531904 40466 531956
rect 346302 531904 346308 531956
rect 346360 531944 346366 531956
rect 405734 531944 405740 531956
rect 346360 531916 405740 531944
rect 346360 531904 346366 531916
rect 405734 531904 405740 531916
rect 405792 531904 405798 531956
rect 26786 531836 26792 531888
rect 26844 531876 26850 531888
rect 34057 531879 34115 531885
rect 34057 531876 34069 531879
rect 26844 531848 34069 531876
rect 26844 531836 26850 531848
rect 34057 531845 34069 531848
rect 34103 531845 34115 531879
rect 34057 531839 34115 531845
rect 34149 531879 34207 531885
rect 34149 531845 34161 531879
rect 34195 531876 34207 531879
rect 36078 531876 36084 531888
rect 34195 531848 36084 531876
rect 34195 531845 34207 531848
rect 34149 531839 34207 531845
rect 36078 531836 36084 531848
rect 36136 531836 36142 531888
rect 348694 531836 348700 531888
rect 348752 531876 348758 531888
rect 401594 531876 401600 531888
rect 348752 531848 401600 531876
rect 348752 531836 348758 531848
rect 401594 531836 401600 531848
rect 401652 531836 401658 531888
rect 28626 531768 28632 531820
rect 28684 531808 28690 531820
rect 38194 531808 38200 531820
rect 28684 531780 38200 531808
rect 28684 531768 28690 531780
rect 38194 531768 38200 531780
rect 38252 531768 38258 531820
rect 350902 531768 350908 531820
rect 350960 531808 350966 531820
rect 398834 531808 398840 531820
rect 350960 531780 398840 531808
rect 350960 531768 350966 531780
rect 398834 531768 398840 531780
rect 398892 531768 398898 531820
rect 353018 531700 353024 531752
rect 353076 531740 353082 531752
rect 394786 531740 394792 531752
rect 353076 531712 394792 531740
rect 353076 531700 353082 531712
rect 394786 531700 394792 531712
rect 394844 531700 394850 531752
rect 26418 531632 26424 531684
rect 26476 531672 26482 531684
rect 34149 531675 34207 531681
rect 34149 531672 34161 531675
rect 26476 531644 34161 531672
rect 26476 531632 26482 531644
rect 34149 531641 34161 531644
rect 34195 531641 34207 531675
rect 34149 531635 34207 531641
rect 355226 531632 355232 531684
rect 355284 531672 355290 531684
rect 391934 531672 391940 531684
rect 355284 531644 391940 531672
rect 355284 531632 355290 531644
rect 391934 531632 391940 531644
rect 391992 531632 391998 531684
rect 167546 531564 167552 531616
rect 167604 531604 167610 531616
rect 339494 531604 339500 531616
rect 167604 531576 339500 531604
rect 167604 531564 167610 531576
rect 339494 531564 339500 531576
rect 339552 531564 339558 531616
rect 357342 531564 357348 531616
rect 357400 531604 357406 531616
rect 387886 531604 387892 531616
rect 357400 531576 387892 531604
rect 357400 531564 357406 531576
rect 387886 531564 387892 531576
rect 387944 531564 387950 531616
rect 163222 531496 163228 531548
rect 163280 531536 163286 531548
rect 344922 531536 344928 531548
rect 163280 531508 344928 531536
rect 163280 531496 163286 531508
rect 344922 531496 344928 531508
rect 344980 531496 344986 531548
rect 359458 531496 359464 531548
rect 359516 531536 359522 531548
rect 383746 531536 383752 531548
rect 359516 531508 383752 531536
rect 359516 531496 359522 531508
rect 383746 531496 383752 531508
rect 383804 531496 383810 531548
rect 161106 531428 161112 531480
rect 161164 531468 161170 531480
rect 347774 531468 347780 531480
rect 161164 531440 347780 531468
rect 161164 531428 161170 531440
rect 347774 531428 347780 531440
rect 347832 531428 347838 531480
rect 361482 531428 361488 531480
rect 361540 531468 361546 531480
rect 380894 531468 380900 531480
rect 361540 531440 380900 531468
rect 361540 531428 361546 531440
rect 380894 531428 380900 531440
rect 380952 531428 380958 531480
rect 158898 531360 158904 531412
rect 158956 531400 158962 531412
rect 353202 531400 353208 531412
rect 158956 531372 353208 531400
rect 158956 531360 158962 531372
rect 353202 531360 353208 531372
rect 353260 531360 353266 531412
rect 363782 531360 363788 531412
rect 363840 531400 363846 531412
rect 376754 531400 376760 531412
rect 363840 531372 376760 531400
rect 363840 531360 363846 531372
rect 376754 531360 376760 531372
rect 376812 531360 376818 531412
rect 29840 531304 30788 531332
rect 26602 531224 26608 531276
rect 26660 531264 26666 531276
rect 29840 531264 29868 531304
rect 26660 531236 29868 531264
rect 26660 531224 26666 531236
rect 29914 531224 29920 531276
rect 29972 531264 29978 531276
rect 30650 531264 30656 531276
rect 29972 531236 30656 531264
rect 29972 531224 29978 531236
rect 30650 531224 30656 531236
rect 30708 531224 30714 531276
rect 30760 531264 30788 531304
rect 156782 531292 156788 531344
rect 156840 531332 156846 531344
rect 156840 531304 356100 531332
rect 156840 531292 156846 531304
rect 59814 531264 59820 531276
rect 30760 531236 59820 531264
rect 59814 531224 59820 531236
rect 59872 531224 59878 531276
rect 231857 531267 231915 531273
rect 231857 531233 231869 531267
rect 231903 531264 231915 531267
rect 241425 531267 241483 531273
rect 241425 531264 241437 531267
rect 231903 531236 241437 531264
rect 231903 531233 231915 531236
rect 231857 531227 231915 531233
rect 241425 531233 241437 531236
rect 241471 531233 241483 531267
rect 241425 531227 241483 531233
rect 325697 531267 325755 531273
rect 325697 531233 325709 531267
rect 325743 531264 325755 531267
rect 335265 531267 335323 531273
rect 335265 531264 335277 531267
rect 325743 531236 335277 531264
rect 325743 531233 325755 531236
rect 325697 531227 325755 531233
rect 335265 531233 335277 531236
rect 335311 531233 335323 531267
rect 335265 531227 335323 531233
rect 353202 531224 353208 531276
rect 353260 531264 353266 531276
rect 356072 531264 356100 531304
rect 439682 531264 439688 531276
rect 353260 531236 355456 531264
rect 356072 531236 439688 531264
rect 353260 531224 353266 531236
rect 27982 531156 27988 531208
rect 28040 531196 28046 531208
rect 70578 531196 70584 531208
rect 28040 531168 70584 531196
rect 28040 531156 28046 531168
rect 70578 531156 70584 531168
rect 70636 531156 70642 531208
rect 196069 531199 196127 531205
rect 196069 531165 196081 531199
rect 196115 531196 196127 531199
rect 201497 531199 201555 531205
rect 201497 531196 201509 531199
rect 196115 531168 201509 531196
rect 196115 531165 196127 531168
rect 196069 531159 196127 531165
rect 201497 531165 201509 531168
rect 201543 531165 201555 531199
rect 201497 531159 201555 531165
rect 222197 531199 222255 531205
rect 222197 531165 222209 531199
rect 222243 531196 222255 531199
rect 231765 531199 231823 531205
rect 231765 531196 231777 531199
rect 222243 531168 231777 531196
rect 222243 531165 222255 531168
rect 222197 531159 222255 531165
rect 231765 531165 231777 531168
rect 231811 531165 231823 531199
rect 231765 531159 231823 531165
rect 241517 531199 241575 531205
rect 241517 531165 241529 531199
rect 241563 531196 241575 531199
rect 251085 531199 251143 531205
rect 251085 531196 251097 531199
rect 241563 531168 251097 531196
rect 241563 531165 241575 531168
rect 241517 531159 241575 531165
rect 251085 531165 251097 531168
rect 251131 531165 251143 531199
rect 251085 531159 251143 531165
rect 251177 531199 251235 531205
rect 251177 531165 251189 531199
rect 251223 531196 251235 531199
rect 264977 531199 265035 531205
rect 251223 531168 254164 531196
rect 251223 531165 251235 531168
rect 251177 531159 251235 531165
rect 22094 531088 22100 531140
rect 22152 531128 22158 531140
rect 23382 531128 23388 531140
rect 22152 531100 23388 531128
rect 22152 531088 22158 531100
rect 23382 531088 23388 531100
rect 23440 531088 23446 531140
rect 26694 531088 26700 531140
rect 26752 531128 26758 531140
rect 65150 531128 65156 531140
rect 26752 531100 65156 531128
rect 26752 531088 26758 531100
rect 65150 531088 65156 531100
rect 65208 531088 65214 531140
rect 150342 531088 150348 531140
rect 150400 531128 150406 531140
rect 156322 531128 156328 531140
rect 150400 531100 156328 531128
rect 150400 531088 150406 531100
rect 156322 531088 156328 531100
rect 156380 531088 156386 531140
rect 186317 531131 186375 531137
rect 186317 531097 186329 531131
rect 186363 531128 186375 531131
rect 195885 531131 195943 531137
rect 195885 531128 195897 531131
rect 186363 531100 195897 531128
rect 186363 531097 186375 531100
rect 186317 531091 186375 531097
rect 195885 531097 195897 531100
rect 195931 531097 195943 531131
rect 195885 531091 195943 531097
rect 206281 531131 206339 531137
rect 206281 531097 206293 531131
rect 206327 531128 206339 531131
rect 206327 531100 215340 531128
rect 206327 531097 206339 531100
rect 206281 531091 206339 531097
rect 26878 531020 26884 531072
rect 26936 531060 26942 531072
rect 71590 531060 71596 531072
rect 26936 531032 71596 531060
rect 26936 531020 26942 531032
rect 71590 531020 71596 531032
rect 71648 531020 71654 531072
rect 184842 531020 184848 531072
rect 184900 531060 184906 531072
rect 191101 531063 191159 531069
rect 191101 531060 191113 531063
rect 184900 531032 191113 531060
rect 184900 531020 184906 531032
rect 191101 531029 191113 531032
rect 191147 531029 191159 531063
rect 191101 531023 191159 531029
rect 198734 531020 198740 531072
rect 198792 531060 198798 531072
rect 199654 531060 199660 531072
rect 198792 531032 199660 531060
rect 198792 531020 198798 531032
rect 199654 531020 199660 531032
rect 199712 531020 199718 531072
rect 202874 531020 202880 531072
rect 202932 531060 202938 531072
rect 203886 531060 203892 531072
rect 202932 531032 203892 531060
rect 202932 531020 202938 531032
rect 203886 531020 203892 531032
rect 203944 531020 203950 531072
rect 215312 531060 215340 531100
rect 223574 531088 223580 531140
rect 223632 531128 223638 531140
rect 224310 531128 224316 531140
rect 223632 531100 224316 531128
rect 223632 531088 223638 531100
rect 224310 531088 224316 531100
rect 224368 531088 224374 531140
rect 227714 531088 227720 531140
rect 227772 531128 227778 531140
rect 228726 531128 228732 531140
rect 227772 531100 228732 531128
rect 227772 531088 227778 531100
rect 228726 531088 228732 531100
rect 228784 531088 228790 531140
rect 233234 531088 233240 531140
rect 233292 531128 233298 531140
rect 234062 531128 234068 531140
rect 233292 531100 234068 531128
rect 233292 531088 233298 531100
rect 234062 531088 234068 531100
rect 234120 531088 234126 531140
rect 237374 531088 237380 531140
rect 237432 531128 237438 531140
rect 238294 531128 238300 531140
rect 237432 531100 238300 531128
rect 237432 531088 237438 531100
rect 238294 531088 238300 531100
rect 238352 531088 238358 531140
rect 254136 531128 254164 531168
rect 264977 531165 264989 531199
rect 265023 531196 265035 531199
rect 274545 531199 274603 531205
rect 274545 531196 274557 531199
rect 265023 531168 274557 531196
rect 265023 531165 265035 531168
rect 264977 531159 265035 531165
rect 274545 531165 274557 531168
rect 274591 531165 274603 531199
rect 274545 531159 274603 531165
rect 339494 531156 339500 531208
rect 339552 531196 339558 531208
rect 339552 531168 345060 531196
rect 339552 531156 339558 531168
rect 254136 531100 261248 531128
rect 222197 531063 222255 531069
rect 222197 531060 222209 531063
rect 215312 531032 222209 531060
rect 222197 531029 222209 531032
rect 222243 531029 222255 531063
rect 222197 531023 222255 531029
rect 231857 531063 231915 531069
rect 231857 531029 231869 531063
rect 231903 531029 231915 531063
rect 231857 531023 231915 531029
rect 241425 531063 241483 531069
rect 241425 531029 241437 531063
rect 241471 531060 241483 531063
rect 241517 531063 241575 531069
rect 241517 531060 241529 531063
rect 241471 531032 241529 531060
rect 241471 531029 241483 531032
rect 241425 531023 241483 531029
rect 241517 531029 241529 531032
rect 241563 531029 241575 531063
rect 241517 531023 241575 531029
rect 251177 531063 251235 531069
rect 251177 531029 251189 531063
rect 251223 531029 251235 531063
rect 261220 531060 261248 531100
rect 261294 531088 261300 531140
rect 261352 531128 261358 531140
rect 262122 531128 262128 531140
rect 261352 531100 262128 531128
rect 261352 531088 261358 531100
rect 262122 531088 262128 531100
rect 262180 531088 262186 531140
rect 262398 531088 262404 531140
rect 262456 531128 262462 531140
rect 263502 531128 263508 531140
rect 262456 531100 263508 531128
rect 262456 531088 262462 531100
rect 263502 531088 263508 531100
rect 263560 531088 263566 531140
rect 267826 531088 267832 531140
rect 267884 531128 267890 531140
rect 268930 531128 268936 531140
rect 267884 531100 268936 531128
rect 267884 531088 267890 531100
rect 268930 531088 268936 531100
rect 268988 531088 268994 531140
rect 271046 531088 271052 531140
rect 271104 531128 271110 531140
rect 271782 531128 271788 531140
rect 271104 531100 271788 531128
rect 271104 531088 271110 531100
rect 271782 531088 271788 531100
rect 271840 531088 271846 531140
rect 272058 531088 272064 531140
rect 272116 531128 272122 531140
rect 273162 531128 273168 531140
rect 272116 531100 273168 531128
rect 272116 531088 272122 531100
rect 273162 531088 273168 531100
rect 273220 531088 273226 531140
rect 276382 531088 276388 531140
rect 276440 531128 276446 531140
rect 277302 531128 277308 531140
rect 276440 531100 277308 531128
rect 276440 531088 276446 531100
rect 277302 531088 277308 531100
rect 277360 531088 277366 531140
rect 277486 531088 277492 531140
rect 277544 531128 277550 531140
rect 278590 531128 278596 531140
rect 277544 531100 278596 531128
rect 277544 531088 277550 531100
rect 278590 531088 278596 531100
rect 278648 531088 278654 531140
rect 318904 531100 322244 531128
rect 263597 531063 263655 531069
rect 263597 531060 263609 531063
rect 261220 531032 263609 531060
rect 251177 531023 251235 531029
rect 263597 531029 263609 531032
rect 263643 531029 263655 531063
rect 263597 531023 263655 531029
rect 263689 531063 263747 531069
rect 263689 531029 263701 531063
rect 263735 531060 263747 531063
rect 264977 531063 265035 531069
rect 264977 531060 264989 531063
rect 263735 531032 264989 531060
rect 263735 531029 263747 531032
rect 263689 531023 263747 531029
rect 264977 531029 264989 531032
rect 265023 531029 265035 531063
rect 264977 531023 265035 531029
rect 282917 531063 282975 531069
rect 282917 531029 282929 531063
rect 282963 531060 282975 531063
rect 292577 531063 292635 531069
rect 292577 531060 292589 531063
rect 282963 531032 292589 531060
rect 282963 531029 282975 531032
rect 282917 531023 282975 531029
rect 292577 531029 292589 531032
rect 292623 531029 292635 531063
rect 292577 531023 292635 531029
rect 292669 531063 292727 531069
rect 292669 531029 292681 531063
rect 292715 531060 292727 531063
rect 292715 531032 296668 531060
rect 292715 531029 292727 531032
rect 292669 531023 292727 531029
rect 28074 530952 28080 531004
rect 28132 530992 28138 531004
rect 77018 530992 77024 531004
rect 28132 530964 77024 530992
rect 28132 530952 28138 530964
rect 77018 530952 77024 530964
rect 77076 530952 77082 531004
rect 173805 530995 173863 531001
rect 173805 530961 173817 530995
rect 173851 530992 173863 530995
rect 186317 530995 186375 531001
rect 186317 530992 186329 530995
rect 173851 530964 186329 530992
rect 173851 530961 173863 530964
rect 173805 530955 173863 530961
rect 186317 530961 186329 530964
rect 186363 530961 186375 530995
rect 186317 530955 186375 530961
rect 201497 530995 201555 531001
rect 201497 530961 201509 530995
rect 201543 530992 201555 530995
rect 206281 530995 206339 531001
rect 206281 530992 206293 530995
rect 201543 530964 206293 530992
rect 201543 530961 201555 530964
rect 201497 530955 201555 530961
rect 206281 530961 206293 530964
rect 206327 530961 206339 530995
rect 206281 530955 206339 530961
rect 231765 530995 231823 531001
rect 231765 530961 231777 530995
rect 231811 530992 231823 530995
rect 231872 530992 231900 531023
rect 231811 530964 231900 530992
rect 251085 530995 251143 531001
rect 231811 530961 231823 530964
rect 231765 530955 231823 530961
rect 251085 530961 251097 530995
rect 251131 530992 251143 530995
rect 251192 530992 251220 531023
rect 251131 530964 251220 530992
rect 274545 530995 274603 531001
rect 251131 530961 251143 530964
rect 251085 530955 251143 530961
rect 274545 530961 274557 530995
rect 274591 530992 274603 530995
rect 282825 530995 282883 531001
rect 282825 530992 282837 530995
rect 274591 530964 282837 530992
rect 274591 530961 274603 530964
rect 274545 530955 274603 530961
rect 282825 530961 282837 530964
rect 282871 530961 282883 530995
rect 296640 530992 296668 531032
rect 298186 531020 298192 531072
rect 298244 531060 298250 531072
rect 302237 531063 302295 531069
rect 302237 531060 302249 531063
rect 298244 531032 302249 531060
rect 298244 531020 298250 531032
rect 302237 531029 302249 531032
rect 302283 531029 302295 531063
rect 302237 531023 302295 531029
rect 302329 531063 302387 531069
rect 302329 531029 302341 531063
rect 302375 531060 302387 531063
rect 318904 531060 318932 531100
rect 302375 531032 318932 531060
rect 322216 531060 322244 531100
rect 326062 531088 326068 531140
rect 326120 531128 326126 531140
rect 326890 531128 326896 531140
rect 326120 531100 326896 531128
rect 326120 531088 326126 531100
rect 326890 531088 326896 531100
rect 326948 531088 326954 531140
rect 330386 531088 330392 531140
rect 330444 531128 330450 531140
rect 331122 531128 331128 531140
rect 330444 531100 331128 531128
rect 330444 531088 330450 531100
rect 331122 531088 331128 531100
rect 331180 531088 331186 531140
rect 334710 531088 334716 531140
rect 334768 531128 334774 531140
rect 335262 531128 335268 531140
rect 334768 531100 335268 531128
rect 334768 531088 334774 531100
rect 335262 531088 335268 531100
rect 335320 531088 335326 531140
rect 341150 531088 341156 531140
rect 341208 531128 341214 531140
rect 341978 531128 341984 531140
rect 341208 531100 341984 531128
rect 341208 531088 341214 531100
rect 341978 531088 341984 531100
rect 342036 531088 342042 531140
rect 325697 531063 325755 531069
rect 325697 531060 325709 531063
rect 322216 531032 325709 531060
rect 302375 531029 302387 531032
rect 302329 531023 302387 531029
rect 325697 531029 325709 531032
rect 325743 531029 325755 531063
rect 345032 531060 345060 531168
rect 347774 531156 347780 531208
rect 347832 531196 347838 531208
rect 355428 531196 355456 531236
rect 439682 531224 439688 531236
rect 439740 531224 439746 531276
rect 442902 531224 442908 531276
rect 442960 531264 442966 531276
rect 448514 531264 448520 531276
rect 442960 531236 448520 531264
rect 442960 531224 442966 531236
rect 448514 531224 448520 531236
rect 448572 531224 448578 531276
rect 535178 531224 535184 531276
rect 535236 531264 535242 531276
rect 535236 531236 550220 531264
rect 535236 531224 535242 531236
rect 437658 531196 437664 531208
rect 347832 531168 355364 531196
rect 355428 531168 437664 531196
rect 347832 531156 347838 531168
rect 345474 531088 345480 531140
rect 345532 531128 345538 531140
rect 346118 531128 346124 531140
rect 345532 531100 346124 531128
rect 345532 531088 345538 531100
rect 346118 531088 346124 531100
rect 346176 531088 346182 531140
rect 349798 531088 349804 531140
rect 349856 531128 349862 531140
rect 350442 531128 350448 531140
rect 349856 531100 350448 531128
rect 349856 531088 349862 531100
rect 350442 531088 350448 531100
rect 350500 531088 350506 531140
rect 354030 531088 354036 531140
rect 354088 531128 354094 531140
rect 354490 531128 354496 531140
rect 354088 531100 354496 531128
rect 354088 531088 354094 531100
rect 354490 531088 354496 531100
rect 354548 531088 354554 531140
rect 355336 531128 355364 531168
rect 437658 531156 437664 531168
rect 437716 531156 437722 531208
rect 533982 531156 533988 531208
rect 534040 531196 534046 531208
rect 550085 531199 550143 531205
rect 550085 531196 550097 531199
rect 534040 531168 550097 531196
rect 534040 531156 534046 531168
rect 550085 531165 550097 531168
rect 550131 531165 550143 531199
rect 550192 531196 550220 531236
rect 551370 531224 551376 531276
rect 551428 531264 551434 531276
rect 551922 531264 551928 531276
rect 551428 531236 551928 531264
rect 551428 531224 551434 531236
rect 551922 531224 551928 531236
rect 551980 531224 551986 531276
rect 552382 531224 552388 531276
rect 552440 531264 552446 531276
rect 552934 531264 552940 531276
rect 552440 531236 552940 531264
rect 552440 531224 552446 531236
rect 552934 531224 552940 531236
rect 552992 531224 552998 531276
rect 552566 531196 552572 531208
rect 550192 531168 552572 531196
rect 550085 531159 550143 531165
rect 552566 531156 552572 531168
rect 552624 531156 552630 531208
rect 435358 531128 435364 531140
rect 355336 531100 435364 531128
rect 435358 531088 435364 531100
rect 435416 531088 435422 531140
rect 533062 531088 533068 531140
rect 533120 531128 533126 531140
rect 547877 531131 547935 531137
rect 547877 531128 547889 531131
rect 533120 531100 547889 531128
rect 533120 531088 533126 531100
rect 547877 531097 547889 531100
rect 547923 531097 547935 531131
rect 547877 531091 547935 531097
rect 547969 531131 548027 531137
rect 547969 531097 547981 531131
rect 548015 531128 548027 531131
rect 552474 531128 552480 531140
rect 548015 531100 552480 531128
rect 548015 531097 548027 531100
rect 547969 531091 548027 531097
rect 552474 531088 552480 531100
rect 552532 531088 552538 531140
rect 429286 531060 429292 531072
rect 345032 531032 429292 531060
rect 325697 531023 325755 531029
rect 429286 531020 429292 531032
rect 429344 531020 429350 531072
rect 528462 531020 528468 531072
rect 528520 531060 528526 531072
rect 551278 531060 551284 531072
rect 528520 531032 551284 531060
rect 528520 531020 528526 531032
rect 551278 531020 551284 531032
rect 551336 531020 551342 531072
rect 298094 530992 298100 531004
rect 296640 530964 298100 530992
rect 282825 530955 282883 530961
rect 298094 530952 298100 530964
rect 298152 530952 298158 531004
rect 335265 530995 335323 531001
rect 335265 530961 335277 530995
rect 335311 530992 335323 530995
rect 338025 530995 338083 531001
rect 338025 530992 338037 530995
rect 335311 530964 338037 530992
rect 335311 530961 335323 530964
rect 335265 530955 335323 530961
rect 338025 530961 338037 530964
rect 338071 530961 338083 530995
rect 338025 530955 338083 530961
rect 338117 530995 338175 531001
rect 338117 530961 338129 530995
rect 338163 530992 338175 530995
rect 342901 530995 342959 531001
rect 342901 530992 342913 530995
rect 338163 530964 342913 530992
rect 338163 530961 338175 530964
rect 338117 530955 338175 530961
rect 342901 530961 342913 530964
rect 342947 530961 342959 530995
rect 342901 530955 342959 530961
rect 344922 530952 344928 531004
rect 344980 530992 344986 531004
rect 433334 530992 433340 531004
rect 344980 530964 433340 530992
rect 344980 530952 344986 530964
rect 433334 530952 433340 530964
rect 433392 530952 433398 531004
rect 526530 530952 526536 531004
rect 526588 530992 526594 531004
rect 547969 530995 548027 531001
rect 547969 530992 547981 530995
rect 526588 530964 547981 530992
rect 526588 530952 526594 530964
rect 547969 530961 547981 530964
rect 548015 530961 548027 530995
rect 551186 530992 551192 531004
rect 547969 530955 548027 530961
rect 548076 530964 551192 530992
rect 27890 530884 27896 530936
rect 27948 530924 27954 530936
rect 78122 530924 78128 530936
rect 27948 530896 78128 530924
rect 27948 530884 27954 530896
rect 78122 530884 78128 530896
rect 78180 530884 78186 530936
rect 186958 530884 186964 530936
rect 187016 530924 187022 530936
rect 409874 530924 409880 530936
rect 187016 530896 409880 530924
rect 187016 530884 187022 530896
rect 409874 530884 409880 530896
rect 409932 530884 409938 530936
rect 522206 530884 522212 530936
rect 522264 530924 522270 530936
rect 548076 530924 548104 530964
rect 551186 530952 551192 530964
rect 551244 530952 551250 531004
rect 522264 530896 548104 530924
rect 522264 530884 522270 530896
rect 548150 530884 548156 530936
rect 548208 530924 548214 530936
rect 552750 530924 552756 530936
rect 548208 530896 552756 530924
rect 548208 530884 548214 530896
rect 552750 530884 552756 530896
rect 552808 530884 552814 530936
rect 27338 530816 27344 530868
rect 27396 530856 27402 530868
rect 81342 530856 81348 530868
rect 27396 530828 81348 530856
rect 27396 530816 27402 530828
rect 81342 530816 81348 530828
rect 81400 530816 81406 530868
rect 146018 530816 146024 530868
rect 146076 530856 146082 530868
rect 147950 530856 147956 530868
rect 146076 530828 147956 530856
rect 146076 530816 146082 530828
rect 147950 530816 147956 530828
rect 148008 530816 148014 530868
rect 191101 530859 191159 530865
rect 191101 530825 191113 530859
rect 191147 530856 191159 530859
rect 411622 530856 411628 530868
rect 191147 530828 411628 530856
rect 191147 530825 191159 530828
rect 191101 530819 191159 530825
rect 411622 530816 411628 530828
rect 411680 530816 411686 530868
rect 524322 530816 524328 530868
rect 524380 530856 524386 530868
rect 549993 530859 550051 530865
rect 549993 530856 550005 530859
rect 524380 530828 550005 530856
rect 524380 530816 524386 530828
rect 549993 530825 550005 530828
rect 550039 530825 550051 530859
rect 549993 530819 550051 530825
rect 550085 530859 550143 530865
rect 550085 530825 550097 530859
rect 550131 530856 550143 530859
rect 554038 530856 554044 530868
rect 550131 530828 554044 530856
rect 550131 530825 550143 530828
rect 550085 530819 550143 530825
rect 554038 530816 554044 530828
rect 554096 530816 554102 530868
rect 27798 530748 27804 530800
rect 27856 530788 27862 530800
rect 83458 530788 83464 530800
rect 27856 530760 83464 530788
rect 27856 530748 27862 530760
rect 83458 530748 83464 530760
rect 83516 530748 83522 530800
rect 182634 530748 182640 530800
rect 182692 530788 182698 530800
rect 414014 530788 414020 530800
rect 182692 530760 414020 530788
rect 182692 530748 182698 530760
rect 414014 530748 414020 530760
rect 414072 530748 414078 530800
rect 520090 530748 520096 530800
rect 520148 530788 520154 530800
rect 552290 530788 552296 530800
rect 520148 530760 552296 530788
rect 520148 530748 520154 530760
rect 552290 530748 552296 530760
rect 552348 530748 552354 530800
rect 27430 530680 27436 530732
rect 27488 530720 27494 530732
rect 85666 530720 85672 530732
rect 27488 530692 85672 530720
rect 27488 530680 27494 530692
rect 85666 530680 85672 530692
rect 85724 530680 85730 530732
rect 180518 530680 180524 530732
rect 180576 530720 180582 530732
rect 415946 530720 415952 530732
rect 180576 530692 415952 530720
rect 180576 530680 180582 530692
rect 415946 530680 415952 530692
rect 416004 530680 416010 530732
rect 517974 530680 517980 530732
rect 518032 530720 518038 530732
rect 550177 530723 550235 530729
rect 550177 530720 550189 530723
rect 518032 530692 550189 530720
rect 518032 530680 518038 530692
rect 550177 530689 550189 530692
rect 550223 530689 550235 530723
rect 550177 530683 550235 530689
rect 550266 530680 550272 530732
rect 550324 530720 550330 530732
rect 552842 530720 552848 530732
rect 550324 530692 552848 530720
rect 550324 530680 550330 530692
rect 552842 530680 552848 530692
rect 552900 530680 552906 530732
rect 27614 530612 27620 530664
rect 27672 530652 27678 530664
rect 88886 530652 88892 530664
rect 27672 530624 88892 530652
rect 27672 530612 27678 530624
rect 88886 530612 88892 530624
rect 88944 530612 88950 530664
rect 90358 530612 90364 530664
rect 90416 530652 90422 530664
rect 99650 530652 99656 530664
rect 90416 530624 99656 530652
rect 90416 530612 90422 530624
rect 99650 530612 99656 530624
rect 99708 530612 99714 530664
rect 178310 530612 178316 530664
rect 178368 530652 178374 530664
rect 418246 530652 418252 530664
rect 178368 530624 418252 530652
rect 178368 530612 178374 530624
rect 418246 530612 418252 530624
rect 418304 530612 418310 530664
rect 513650 530612 513656 530664
rect 513708 530652 513714 530664
rect 552106 530652 552112 530664
rect 513708 530624 552112 530652
rect 513708 530612 513714 530624
rect 552106 530612 552112 530624
rect 552164 530612 552170 530664
rect 555418 530612 555424 530664
rect 555476 530652 555482 530664
rect 562594 530652 562600 530664
rect 555476 530624 562600 530652
rect 555476 530612 555482 530624
rect 562594 530612 562600 530624
rect 562652 530612 562658 530664
rect 27522 530544 27528 530596
rect 27580 530584 27586 530596
rect 89990 530584 89996 530596
rect 27580 530556 89996 530584
rect 27580 530544 27586 530556
rect 89990 530544 89996 530556
rect 90048 530544 90054 530596
rect 90542 530544 90548 530596
rect 90600 530584 90606 530596
rect 105078 530584 105084 530596
rect 90600 530556 105084 530584
rect 90600 530544 90606 530556
rect 105078 530544 105084 530556
rect 105136 530544 105142 530596
rect 112622 530544 112628 530596
rect 112680 530584 112686 530596
rect 166994 530584 167000 530596
rect 112680 530556 167000 530584
rect 112680 530544 112686 530556
rect 166994 530544 167000 530556
rect 167052 530544 167058 530596
rect 176194 530544 176200 530596
rect 176252 530584 176258 530596
rect 420270 530584 420276 530596
rect 176252 530556 420276 530584
rect 176252 530544 176258 530556
rect 420270 530544 420276 530556
rect 420328 530544 420334 530596
rect 436002 530544 436008 530596
rect 436060 530584 436066 530596
rect 444374 530584 444380 530596
rect 436060 530556 444380 530584
rect 436060 530544 436066 530556
rect 444374 530544 444380 530556
rect 444432 530544 444438 530596
rect 511442 530544 511448 530596
rect 511500 530584 511506 530596
rect 550085 530587 550143 530593
rect 550085 530584 550097 530587
rect 511500 530556 550097 530584
rect 511500 530544 511506 530556
rect 550085 530553 550097 530556
rect 550131 530553 550143 530587
rect 550085 530547 550143 530553
rect 550177 530587 550235 530593
rect 550177 530553 550189 530587
rect 550223 530584 550235 530587
rect 553486 530584 553492 530596
rect 550223 530556 553492 530584
rect 550223 530553 550235 530556
rect 550177 530547 550235 530553
rect 553486 530544 553492 530556
rect 553544 530544 553550 530596
rect 558270 530544 558276 530596
rect 558328 530584 558334 530596
rect 572254 530584 572260 530596
rect 558328 530556 572260 530584
rect 558328 530544 558334 530556
rect 572254 530544 572260 530556
rect 572312 530544 572318 530596
rect 25958 530476 25964 530528
rect 26016 530516 26022 530528
rect 55490 530516 55496 530528
rect 26016 530488 55496 530516
rect 26016 530476 26022 530488
rect 55490 530476 55496 530488
rect 55548 530476 55554 530528
rect 173986 530476 173992 530528
rect 174044 530516 174050 530528
rect 422478 530516 422484 530528
rect 174044 530488 422484 530516
rect 174044 530476 174050 530488
rect 422478 530476 422484 530488
rect 422536 530476 422542 530528
rect 542722 530476 542728 530528
rect 542780 530516 542786 530528
rect 543642 530516 543648 530528
rect 542780 530488 543648 530516
rect 542780 530476 542786 530488
rect 543642 530476 543648 530488
rect 543700 530476 543706 530528
rect 543737 530519 543795 530525
rect 543737 530485 543749 530519
rect 543783 530516 543795 530519
rect 549901 530519 549959 530525
rect 549901 530516 549913 530519
rect 543783 530488 549913 530516
rect 543783 530485 543795 530488
rect 543737 530479 543795 530485
rect 549901 530485 549913 530488
rect 549947 530485 549959 530519
rect 549901 530479 549959 530485
rect 549993 530519 550051 530525
rect 549993 530485 550005 530519
rect 550039 530516 550051 530519
rect 553670 530516 553676 530528
rect 550039 530488 553676 530516
rect 550039 530485 550051 530488
rect 549993 530479 550051 530485
rect 553670 530476 553676 530488
rect 553728 530476 553734 530528
rect 28258 530408 28264 530460
rect 28316 530448 28322 530460
rect 53282 530448 53288 530460
rect 28316 530420 53288 530448
rect 28316 530408 28322 530420
rect 53282 530408 53288 530420
rect 53340 530408 53346 530460
rect 171870 530408 171876 530460
rect 171928 530448 171934 530460
rect 424594 530448 424600 530460
rect 171928 530420 424600 530448
rect 171928 530408 171934 530420
rect 424594 530408 424600 530420
rect 424652 530408 424658 530460
rect 537294 530408 537300 530460
rect 537352 530448 537358 530460
rect 551646 530448 551652 530460
rect 537352 530420 551652 530448
rect 537352 530408 537358 530420
rect 551646 530408 551652 530420
rect 551704 530408 551710 530460
rect 553302 530408 553308 530460
rect 553360 530448 553366 530460
rect 554590 530448 554596 530460
rect 553360 530420 554596 530448
rect 553360 530408 553366 530420
rect 554590 530408 554596 530420
rect 554648 530408 554654 530460
rect 28350 530340 28356 530392
rect 28408 530380 28414 530392
rect 51166 530380 51172 530392
rect 28408 530352 51172 530380
rect 28408 530340 28414 530352
rect 51166 530340 51172 530352
rect 51224 530340 51230 530392
rect 169754 530340 169760 530392
rect 169812 530380 169818 530392
rect 426710 530380 426716 530392
rect 169812 530352 426716 530380
rect 169812 530340 169818 530352
rect 426710 530340 426716 530352
rect 426768 530340 426774 530392
rect 541618 530340 541624 530392
rect 541676 530380 541682 530392
rect 549993 530383 550051 530389
rect 549993 530380 550005 530383
rect 541676 530352 550005 530380
rect 541676 530340 541682 530352
rect 549993 530349 550005 530352
rect 550039 530349 550051 530383
rect 549993 530343 550051 530349
rect 550085 530383 550143 530389
rect 550085 530349 550097 530383
rect 550131 530380 550143 530383
rect 553394 530380 553400 530392
rect 550131 530352 553400 530380
rect 550131 530349 550143 530352
rect 550085 530343 550143 530349
rect 553394 530340 553400 530352
rect 553452 530340 553458 530392
rect 28534 530272 28540 530324
rect 28592 530312 28598 530324
rect 48958 530312 48964 530324
rect 28592 530284 48964 530312
rect 28592 530272 28598 530284
rect 48958 530272 48964 530284
rect 49016 530272 49022 530324
rect 133046 530272 133052 530324
rect 133104 530312 133110 530324
rect 463786 530312 463792 530324
rect 133104 530284 463792 530312
rect 133104 530272 133110 530284
rect 463786 530272 463792 530284
rect 463844 530272 463850 530324
rect 543642 530272 543648 530324
rect 543700 530312 543706 530324
rect 552658 530312 552664 530324
rect 543700 530284 552664 530312
rect 543700 530272 543706 530284
rect 552658 530272 552664 530284
rect 552716 530272 552722 530324
rect 558178 530272 558184 530324
rect 558236 530312 558242 530324
rect 559282 530312 559288 530324
rect 558236 530284 559288 530312
rect 558236 530272 558242 530284
rect 559282 530272 559288 530284
rect 559340 530272 559346 530324
rect 27154 530204 27160 530256
rect 27212 530244 27218 530256
rect 46842 530244 46848 530256
rect 27212 530216 46848 530244
rect 27212 530204 27218 530216
rect 46842 530204 46848 530216
rect 46900 530204 46906 530256
rect 109310 530204 109316 530256
rect 109368 530244 109374 530256
rect 111058 530244 111064 530256
rect 109368 530216 111064 530244
rect 109368 530204 109374 530216
rect 111058 530204 111064 530216
rect 111116 530204 111122 530256
rect 130930 530204 130936 530256
rect 130988 530244 130994 530256
rect 465534 530244 465540 530256
rect 130988 530216 465540 530244
rect 130988 530204 130994 530216
rect 465534 530204 465540 530216
rect 465592 530204 465598 530256
rect 471698 530204 471704 530256
rect 471756 530244 471762 530256
rect 481726 530244 481732 530256
rect 471756 530216 481732 530244
rect 471756 530204 471762 530216
rect 481726 530204 481732 530216
rect 481784 530204 481790 530256
rect 539502 530204 539508 530256
rect 539560 530244 539566 530256
rect 543737 530247 543795 530253
rect 543737 530244 543749 530247
rect 539560 530216 543749 530244
rect 539560 530204 539566 530216
rect 543737 530213 543749 530216
rect 543783 530213 543795 530247
rect 543737 530207 543795 530213
rect 547877 530247 547935 530253
rect 547877 530213 547889 530247
rect 547923 530244 547935 530247
rect 554222 530244 554228 530256
rect 547923 530216 554228 530244
rect 547923 530213 547935 530216
rect 547877 530207 547935 530213
rect 554222 530204 554228 530216
rect 554280 530204 554286 530256
rect 25590 530136 25596 530188
rect 25648 530176 25654 530188
rect 44726 530176 44732 530188
rect 25648 530148 44732 530176
rect 25648 530136 25654 530148
rect 44726 530136 44732 530148
rect 44784 530136 44790 530188
rect 128722 530136 128728 530188
rect 128780 530176 128786 530188
rect 467834 530176 467840 530188
rect 128780 530148 467840 530176
rect 128780 530136 128786 530148
rect 467834 530136 467840 530148
rect 467892 530136 467898 530188
rect 468113 530179 468171 530185
rect 468113 530145 468125 530179
rect 468159 530176 468171 530179
rect 478874 530176 478880 530188
rect 468159 530148 478880 530176
rect 468159 530145 468171 530148
rect 468113 530139 468171 530145
rect 478874 530136 478880 530148
rect 478932 530136 478938 530188
rect 493134 530136 493140 530188
rect 493192 530176 493198 530188
rect 493962 530176 493968 530188
rect 493192 530148 493968 530176
rect 493192 530136 493198 530148
rect 493962 530136 493968 530148
rect 494020 530136 494026 530188
rect 549901 530179 549959 530185
rect 549901 530145 549913 530179
rect 549947 530176 549959 530179
rect 554406 530176 554412 530188
rect 549947 530148 554412 530176
rect 549947 530145 549959 530148
rect 549901 530139 549959 530145
rect 554406 530136 554412 530148
rect 554464 530136 554470 530188
rect 126606 530068 126612 530120
rect 126664 530108 126670 530120
rect 469858 530108 469864 530120
rect 126664 530080 469864 530108
rect 126664 530068 126670 530080
rect 469858 530068 469864 530080
rect 469916 530068 469922 530120
rect 549993 530111 550051 530117
rect 549993 530077 550005 530111
rect 550039 530108 550051 530111
rect 554498 530108 554504 530120
rect 550039 530080 554504 530108
rect 550039 530077 550051 530080
rect 549993 530071 550051 530077
rect 554498 530068 554504 530080
rect 554556 530068 554562 530120
rect 124398 530000 124404 530052
rect 124456 530040 124462 530052
rect 472066 530040 472072 530052
rect 124456 530012 472072 530040
rect 124456 530000 124462 530012
rect 472066 530000 472072 530012
rect 472124 530000 472130 530052
rect 482922 530000 482928 530052
rect 482980 530040 482986 530052
rect 488534 530040 488540 530052
rect 482980 530012 488540 530040
rect 482980 530000 482986 530012
rect 488534 530000 488540 530012
rect 488592 530000 488598 530052
rect 556798 530000 556804 530052
rect 556856 530040 556862 530052
rect 558270 530040 558276 530052
rect 556856 530012 558276 530040
rect 556856 530000 556862 530012
rect 558270 530000 558276 530012
rect 558328 530000 558334 530052
rect 122282 529932 122288 529984
rect 122340 529972 122346 529984
rect 474182 529972 474188 529984
rect 122340 529944 474188 529972
rect 122340 529932 122346 529944
rect 474182 529932 474188 529944
rect 474240 529932 474246 529984
rect 481542 529932 481548 529984
rect 481600 529972 481606 529984
rect 484946 529972 484952 529984
rect 481600 529944 484952 529972
rect 481600 529932 481606 529944
rect 484946 529932 484952 529944
rect 485004 529932 485010 529984
rect 560938 529932 560944 529984
rect 560996 529972 561002 529984
rect 567930 529972 567936 529984
rect 560996 529944 567936 529972
rect 560996 529932 561002 529944
rect 567930 529932 567936 529944
rect 567988 529932 567994 529984
rect 342901 529907 342959 529913
rect 342901 529873 342913 529907
rect 342947 529904 342959 529907
rect 431034 529904 431040 529916
rect 342947 529876 431040 529904
rect 342947 529873 342959 529876
rect 342901 529867 342959 529873
rect 431034 529864 431040 529876
rect 431092 529864 431098 529916
rect 191282 529796 191288 529848
rect 191340 529836 191346 529848
rect 405182 529836 405188 529848
rect 191340 529808 405188 529836
rect 191340 529796 191346 529808
rect 405182 529796 405188 529808
rect 405240 529796 405246 529848
rect 165430 529728 165436 529780
rect 165488 529768 165494 529780
rect 173805 529771 173863 529777
rect 173805 529768 173817 529771
rect 165488 529740 173817 529768
rect 165488 529728 165494 529740
rect 173805 529737 173817 529740
rect 173851 529737 173863 529771
rect 173805 529731 173863 529737
rect 179414 529728 179420 529780
rect 179472 529768 179478 529780
rect 417050 529768 417056 529780
rect 179472 529740 417056 529768
rect 179472 529728 179478 529740
rect 417050 529728 417056 529740
rect 417108 529728 417114 529780
rect 160002 529660 160008 529712
rect 160060 529700 160066 529712
rect 436462 529700 436468 529712
rect 160060 529672 436468 529700
rect 160060 529660 160066 529672
rect 436462 529660 436468 529672
rect 436520 529660 436526 529712
rect 157886 529592 157892 529644
rect 157944 529632 157950 529644
rect 438946 529632 438952 529644
rect 157944 529604 438952 529632
rect 157944 529592 157950 529604
rect 438946 529592 438952 529604
rect 439004 529592 439010 529644
rect 151354 529524 151360 529576
rect 151412 529564 151418 529576
rect 445110 529564 445116 529576
rect 151412 529536 445116 529564
rect 151412 529524 151418 529536
rect 445110 529524 445116 529536
rect 445168 529524 445174 529576
rect 149238 529456 149244 529508
rect 149296 529496 149302 529508
rect 447318 529496 447324 529508
rect 149296 529468 447324 529496
rect 149296 529456 149302 529468
rect 447318 529456 447324 529468
rect 447376 529456 447382 529508
rect 147030 529388 147036 529440
rect 147088 529428 147094 529440
rect 449434 529428 449440 529440
rect 147088 529400 449440 529428
rect 147088 529388 147094 529400
rect 449434 529388 449440 529400
rect 449492 529388 449498 529440
rect 144914 529320 144920 529372
rect 144972 529360 144978 529372
rect 451550 529360 451556 529372
rect 144972 529332 451556 529360
rect 144972 529320 144978 529332
rect 451550 529320 451556 529332
rect 451608 529320 451614 529372
rect 111518 529252 111524 529304
rect 111576 529292 111582 529304
rect 481542 529292 481548 529304
rect 111576 529264 481548 529292
rect 111576 529252 111582 529264
rect 481542 529252 481548 529264
rect 481600 529252 481606 529304
rect 108298 529184 108304 529236
rect 108356 529224 108362 529236
rect 482922 529224 482928 529236
rect 108356 529196 482928 529224
rect 108356 529184 108362 529196
rect 482922 529184 482928 529196
rect 482980 529184 482986 529236
rect 142798 529116 142804 529168
rect 142856 529156 142862 529168
rect 454034 529156 454040 529168
rect 142856 529128 454040 529156
rect 142856 529116 142862 529128
rect 454034 529116 454040 529128
rect 454092 529116 454098 529168
rect 140590 529048 140596 529100
rect 140648 529088 140654 529100
rect 456196 529088 456202 529100
rect 140648 529060 456202 529088
rect 140648 529048 140654 529060
rect 456196 529048 456202 529060
rect 456254 529048 456260 529100
rect 138474 528980 138480 529032
rect 138532 529020 138538 529032
rect 458312 529020 458318 529032
rect 138532 528992 458318 529020
rect 138532 528980 138538 528992
rect 458312 528980 458318 528992
rect 458370 528980 458376 529032
rect 136542 528912 136548 528964
rect 136600 528952 136606 528964
rect 460198 528952 460204 528964
rect 136600 528924 460204 528952
rect 136600 528912 136606 528924
rect 460198 528912 460204 528924
rect 460256 528912 460262 528964
rect 134426 528844 134432 528896
rect 134484 528884 134490 528896
rect 462314 528884 462320 528896
rect 134484 528856 462320 528884
rect 134484 528844 134490 528856
rect 462314 528844 462320 528856
rect 462372 528844 462378 528896
rect 120442 528776 120448 528828
rect 120500 528816 120506 528828
rect 476298 528816 476304 528828
rect 120500 528788 476304 528816
rect 120500 528776 120506 528788
rect 476298 528776 476304 528788
rect 476356 528776 476362 528828
rect 117130 528708 117136 528760
rect 117188 528748 117194 528760
rect 479610 528748 479616 528760
rect 117188 528720 479616 528748
rect 117188 528708 117194 528720
rect 479610 528708 479616 528720
rect 479668 528708 479674 528760
rect 114002 528640 114008 528692
rect 114060 528680 114066 528692
rect 483014 528680 483020 528692
rect 114060 528652 483020 528680
rect 114060 528640 114066 528652
rect 483014 528640 483020 528652
rect 483072 528640 483078 528692
rect 110690 528572 110696 528624
rect 110748 528612 110754 528624
rect 486050 528612 486056 528624
rect 110748 528584 486056 528612
rect 110748 528572 110754 528584
rect 486050 528572 486056 528584
rect 486108 528572 486114 528624
rect 315942 528504 315948 528556
rect 316000 528544 316006 528556
rect 456058 528544 456064 528556
rect 316000 528516 456064 528544
rect 316000 528504 316006 528516
rect 456058 528504 456064 528516
rect 456116 528504 456122 528556
rect 194594 528436 194600 528488
rect 194652 528476 194658 528488
rect 401962 528476 401968 528488
rect 194652 528448 401968 528476
rect 194652 528436 194658 528448
rect 401962 528436 401968 528448
rect 402020 528436 402026 528488
rect 403621 528479 403679 528485
rect 403621 528445 403633 528479
rect 403667 528476 403679 528479
rect 408681 528479 408739 528485
rect 408681 528476 408693 528479
rect 403667 528448 408693 528476
rect 403667 528445 403679 528448
rect 403621 528439 403679 528445
rect 408681 528445 408693 528448
rect 408727 528445 408739 528479
rect 408681 528439 408739 528445
rect 190362 528368 190368 528420
rect 190420 528408 190426 528420
rect 406286 528408 406292 528420
rect 190420 528380 406292 528408
rect 190420 528368 190426 528380
rect 406286 528368 406292 528380
rect 406344 528368 406350 528420
rect 406381 528411 406439 528417
rect 406381 528377 406393 528411
rect 406427 528408 406439 528411
rect 413281 528411 413339 528417
rect 413281 528408 413293 528411
rect 406427 528380 413293 528408
rect 406427 528377 406439 528380
rect 406381 528371 406439 528377
rect 413281 528377 413293 528380
rect 413327 528377 413339 528411
rect 413281 528371 413339 528377
rect 186130 528300 186136 528352
rect 186188 528340 186194 528352
rect 410610 528340 410616 528352
rect 186188 528312 410616 528340
rect 186188 528300 186194 528312
rect 410610 528300 410616 528312
rect 410668 528300 410674 528352
rect 422941 528343 422999 528349
rect 422941 528309 422953 528343
rect 422987 528340 422999 528343
rect 423677 528343 423735 528349
rect 423677 528340 423689 528343
rect 422987 528312 423689 528340
rect 422987 528309 422999 528312
rect 422941 528303 422999 528309
rect 423677 528309 423689 528312
rect 423723 528309 423735 528343
rect 423677 528303 423735 528309
rect 115934 528232 115940 528284
rect 115992 528272 115998 528284
rect 125318 528272 125324 528284
rect 115992 528244 125324 528272
rect 115992 528232 115998 528244
rect 125318 528232 125324 528244
rect 125376 528232 125382 528284
rect 181898 528232 181904 528284
rect 181956 528272 181962 528284
rect 414934 528272 414940 528284
rect 181956 528244 414940 528272
rect 181956 528232 181962 528244
rect 414934 528232 414940 528244
rect 414992 528232 414998 528284
rect 118234 528164 118240 528216
rect 118292 528164 118298 528216
rect 164510 528164 164516 528216
rect 164568 528164 164574 528216
rect 169018 528164 169024 528216
rect 169076 528164 169082 528216
rect 173250 528164 173256 528216
rect 173308 528204 173314 528216
rect 388809 528207 388867 528213
rect 388809 528204 388821 528207
rect 173308 528176 388821 528204
rect 173308 528164 173314 528176
rect 388809 528173 388821 528176
rect 388855 528173 388867 528207
rect 388809 528167 388867 528173
rect 389177 528207 389235 528213
rect 389177 528173 389189 528207
rect 389223 528204 389235 528207
rect 423674 528204 423680 528216
rect 389223 528176 423680 528204
rect 389223 528173 389235 528176
rect 389177 528167 389235 528173
rect 423674 528164 423680 528176
rect 423732 528164 423738 528216
rect 427814 528164 427820 528216
rect 427872 528164 427878 528216
rect 432138 528164 432144 528216
rect 432196 528164 432202 528216
rect 434717 528207 434775 528213
rect 434717 528173 434729 528207
rect 434763 528204 434775 528207
rect 444285 528207 444343 528213
rect 444285 528204 444297 528207
rect 434763 528176 444297 528204
rect 434763 528173 434775 528176
rect 434717 528167 434775 528173
rect 444285 528173 444297 528176
rect 444331 528173 444343 528207
rect 444285 528167 444343 528173
rect 456705 528207 456763 528213
rect 456705 528173 456717 528207
rect 456751 528204 456763 528207
rect 463605 528207 463663 528213
rect 463605 528204 463617 528207
rect 456751 528176 463617 528204
rect 456751 528173 456763 528176
rect 456705 528167 456763 528173
rect 463605 528173 463617 528176
rect 463651 528173 463663 528207
rect 463605 528167 463663 528173
rect 118252 528000 118280 528164
rect 164528 528068 164556 528164
rect 169036 528136 169064 528164
rect 388901 528139 388959 528145
rect 388901 528136 388913 528139
rect 169036 528108 388913 528136
rect 388901 528105 388913 528108
rect 388947 528105 388959 528139
rect 389821 528139 389879 528145
rect 388901 528099 388959 528105
rect 389008 528108 389772 528136
rect 389008 528068 389036 528108
rect 164528 528040 389036 528068
rect 389177 528071 389235 528077
rect 389177 528037 389189 528071
rect 389223 528068 389235 528071
rect 389545 528071 389603 528077
rect 389545 528068 389557 528071
rect 389223 528040 389557 528068
rect 389223 528037 389235 528040
rect 389177 528031 389235 528037
rect 389545 528037 389557 528040
rect 389591 528037 389603 528071
rect 389744 528068 389772 528108
rect 389821 528105 389833 528139
rect 389867 528136 389879 528139
rect 403621 528139 403679 528145
rect 403621 528136 403633 528139
rect 389867 528108 403633 528136
rect 389867 528105 389879 528108
rect 389821 528099 389879 528105
rect 403621 528105 403633 528108
rect 403667 528105 403679 528139
rect 403621 528099 403679 528105
rect 408681 528139 408739 528145
rect 408681 528105 408693 528139
rect 408727 528136 408739 528139
rect 427832 528136 427860 528164
rect 408727 528108 427860 528136
rect 408727 528105 408739 528108
rect 408681 528099 408739 528105
rect 432156 528068 432184 528164
rect 463697 528139 463755 528145
rect 463697 528105 463709 528139
rect 463743 528136 463755 528139
rect 468113 528139 468171 528145
rect 468113 528136 468125 528139
rect 463743 528108 468125 528136
rect 463743 528105 463755 528108
rect 463697 528099 463755 528105
rect 468113 528105 468125 528108
rect 468159 528105 468171 528139
rect 468113 528099 468171 528105
rect 389744 528040 432184 528068
rect 444285 528071 444343 528077
rect 389545 528031 389603 528037
rect 444285 528037 444297 528071
rect 444331 528037 444343 528071
rect 456705 528071 456763 528077
rect 456705 528068 456717 528071
rect 444285 528031 444343 528037
rect 454006 528040 456717 528068
rect 406381 528003 406439 528009
rect 406381 528000 406393 528003
rect 118252 527972 406393 528000
rect 406381 527969 406393 527972
rect 406427 527969 406439 528003
rect 406381 527963 406439 527969
rect 413281 528003 413339 528009
rect 413281 527969 413293 528003
rect 413327 528000 413339 528003
rect 422941 528003 422999 528009
rect 422941 528000 422953 528003
rect 413327 527972 422953 528000
rect 413327 527969 413339 527972
rect 413281 527963 413339 527969
rect 422941 527969 422953 527972
rect 422987 527969 422999 528003
rect 422941 527963 422999 527969
rect 423677 528003 423735 528009
rect 423677 527969 423689 528003
rect 423723 528000 423735 528003
rect 434717 528003 434775 528009
rect 434717 528000 434729 528003
rect 423723 527972 434729 528000
rect 423723 527969 423735 527972
rect 423677 527963 423735 527969
rect 434717 527969 434729 527972
rect 434763 527969 434775 528003
rect 444300 528000 444328 528031
rect 454006 528000 454034 528040
rect 456705 528037 456717 528040
rect 456751 528037 456763 528071
rect 456705 528031 456763 528037
rect 463605 528071 463663 528077
rect 463605 528037 463617 528071
rect 463651 528068 463663 528071
rect 463651 528040 463740 528068
rect 463651 528037 463663 528040
rect 463605 528031 463663 528037
rect 463712 528009 463740 528040
rect 444300 527972 454034 528000
rect 463697 528003 463755 528009
rect 434717 527963 434775 527969
rect 463697 527969 463709 528003
rect 463743 527969 463755 528003
rect 463697 527963 463755 527969
rect 298094 527416 298100 527468
rect 298152 527456 298158 527468
rect 302970 527456 302976 527468
rect 298152 527428 302976 527456
rect 298152 527416 298158 527428
rect 302970 527416 302976 527428
rect 303028 527416 303034 527468
rect 288526 527212 288532 527264
rect 288584 527252 288590 527264
rect 296622 527252 296628 527264
rect 288584 527224 296628 527252
rect 288584 527212 288590 527224
rect 296622 527212 296628 527224
rect 296680 527212 296686 527264
rect 282914 514700 282920 514752
rect 282972 514740 282978 514752
rect 283098 514740 283104 514752
rect 282972 514712 283104 514740
rect 282972 514700 282978 514712
rect 283098 514700 283104 514712
rect 283156 514700 283162 514752
rect 577590 509600 577596 509652
rect 577648 509640 577654 509652
rect 579614 509640 579620 509652
rect 577648 509612 579620 509640
rect 577648 509600 577654 509612
rect 579614 509600 579620 509612
rect 579672 509600 579678 509652
rect 2866 509260 2872 509312
rect 2924 509300 2930 509312
rect 14550 509300 14556 509312
rect 2924 509272 14556 509300
rect 2924 509260 2930 509272
rect 14550 509260 14556 509272
rect 14608 509260 14614 509312
rect 283009 509235 283067 509241
rect 283009 509201 283021 509235
rect 283055 509232 283067 509235
rect 283098 509232 283104 509244
rect 283055 509204 283104 509232
rect 283055 509201 283067 509204
rect 283009 509195 283067 509201
rect 283098 509192 283104 509204
rect 283156 509192 283162 509244
rect 416590 503004 416596 503056
rect 416648 503044 416654 503056
rect 418154 503044 418160 503056
rect 416648 503016 418160 503044
rect 416648 503004 416654 503016
rect 418154 503004 418160 503016
rect 418212 503004 418218 503056
rect 418798 503004 418804 503056
rect 418856 503044 418862 503056
rect 420270 503044 420276 503056
rect 418856 503016 420276 503044
rect 418856 503004 418862 503016
rect 420270 503004 420276 503016
rect 420328 503004 420334 503056
rect 413278 502936 413284 502988
rect 413336 502976 413342 502988
rect 580350 502976 580356 502988
rect 413336 502948 580356 502976
rect 413336 502936 413342 502948
rect 580350 502936 580356 502948
rect 580408 502936 580414 502988
rect 481266 502868 481272 502920
rect 481324 502908 481330 502920
rect 484302 502908 484308 502920
rect 481324 502880 484308 502908
rect 481324 502868 481330 502880
rect 484302 502868 484308 502880
rect 484360 502908 484366 502920
rect 487154 502908 487160 502920
rect 484360 502880 487160 502908
rect 484360 502868 484366 502880
rect 487154 502868 487160 502880
rect 487212 502868 487218 502920
rect 459462 502664 459468 502716
rect 459520 502704 459526 502716
rect 461210 502704 461216 502716
rect 459520 502676 461216 502704
rect 459520 502664 459526 502676
rect 461210 502664 461216 502676
rect 461268 502664 461274 502716
rect 114554 502596 114560 502648
rect 114612 502636 114618 502648
rect 115566 502636 115572 502648
rect 114612 502608 115572 502636
rect 114612 502596 114618 502608
rect 115566 502596 115572 502608
rect 115624 502596 115630 502648
rect 158714 501168 158720 501220
rect 158772 501208 158778 501220
rect 159726 501208 159732 501220
rect 158772 501180 159732 501208
rect 158772 501168 158778 501180
rect 159726 501168 159732 501180
rect 159784 501168 159790 501220
rect 164234 501168 164240 501220
rect 164292 501208 164298 501220
rect 165062 501208 165068 501220
rect 164292 501180 165068 501208
rect 164292 501168 164298 501180
rect 165062 501168 165068 501180
rect 165120 501168 165126 501220
rect 173894 501168 173900 501220
rect 173952 501208 173958 501220
rect 174814 501208 174820 501220
rect 173952 501180 174820 501208
rect 173952 501168 173958 501180
rect 174814 501168 174820 501180
rect 174872 501168 174878 501220
rect 183646 501168 183652 501220
rect 183704 501208 183710 501220
rect 184566 501208 184572 501220
rect 183704 501180 184572 501208
rect 183704 501168 183710 501180
rect 184566 501168 184572 501180
rect 184624 501168 184630 501220
rect 24210 500896 24216 500948
rect 24268 500936 24274 500948
rect 25314 500936 25320 500948
rect 24268 500908 25320 500936
rect 24268 500896 24274 500908
rect 25314 500896 25320 500908
rect 25372 500896 25378 500948
rect 27522 500896 27528 500948
rect 27580 500936 27586 500948
rect 29638 500936 29644 500948
rect 27580 500908 29644 500936
rect 27580 500896 27586 500908
rect 29638 500896 29644 500908
rect 29696 500896 29702 500948
rect 50062 500896 50068 500948
rect 50120 500936 50126 500948
rect 50982 500936 50988 500948
rect 50120 500908 50988 500936
rect 50120 500896 50126 500908
rect 50982 500896 50988 500908
rect 51040 500896 51046 500948
rect 59814 500896 59820 500948
rect 59872 500936 59878 500948
rect 60642 500936 60648 500948
rect 59872 500908 60648 500936
rect 59872 500896 59878 500908
rect 60642 500896 60648 500908
rect 60700 500896 60706 500948
rect 60826 500896 60832 500948
rect 60884 500936 60890 500948
rect 61930 500936 61936 500948
rect 60884 500908 61936 500936
rect 60884 500896 60890 500908
rect 61930 500896 61936 500908
rect 61988 500896 61994 500948
rect 64046 500896 64052 500948
rect 64104 500936 64110 500948
rect 64782 500936 64788 500948
rect 64104 500908 64788 500936
rect 64104 500896 64110 500908
rect 64782 500896 64788 500908
rect 64840 500896 64846 500948
rect 69474 500896 69480 500948
rect 69532 500936 69538 500948
rect 70302 500936 70308 500948
rect 69532 500908 70308 500936
rect 69532 500896 69538 500908
rect 70302 500896 70308 500908
rect 70360 500896 70366 500948
rect 99650 500896 99656 500948
rect 99708 500936 99714 500948
rect 100662 500936 100668 500948
rect 99708 500908 100668 500936
rect 99708 500896 99714 500908
rect 100662 500896 100668 500908
rect 100720 500896 100726 500948
rect 100754 500896 100760 500948
rect 100812 500936 100818 500948
rect 102042 500936 102048 500948
rect 100812 500908 102048 500936
rect 100812 500896 100818 500908
rect 102042 500896 102048 500908
rect 102100 500896 102106 500948
rect 105078 500896 105084 500948
rect 105136 500936 105142 500948
rect 106182 500936 106188 500948
rect 105136 500908 106188 500936
rect 105136 500896 105142 500908
rect 106182 500896 106188 500908
rect 106240 500896 106246 500948
rect 121454 500896 121460 500948
rect 121512 500936 121518 500948
rect 153470 500936 153476 500948
rect 121512 500908 153476 500936
rect 121512 500896 121518 500908
rect 153470 500896 153476 500908
rect 153528 500896 153534 500948
rect 195238 500896 195244 500948
rect 195296 500936 195302 500948
rect 197722 500936 197728 500948
rect 195296 500908 197728 500936
rect 195296 500896 195302 500908
rect 197722 500896 197728 500908
rect 197780 500896 197786 500948
rect 201678 500896 201684 500948
rect 201736 500936 201742 500948
rect 203150 500936 203156 500948
rect 201736 500908 203156 500936
rect 201736 500896 201742 500908
rect 203150 500896 203156 500908
rect 203208 500896 203214 500948
rect 204622 500896 204628 500948
rect 204680 500936 204686 500948
rect 208486 500936 208492 500948
rect 204680 500908 208492 500936
rect 204680 500896 204686 500908
rect 208486 500896 208492 500908
rect 208544 500896 208550 500948
rect 214650 500896 214656 500948
rect 214708 500936 214714 500948
rect 217134 500936 217140 500948
rect 214708 500908 217140 500936
rect 214708 500896 214714 500908
rect 217134 500896 217140 500908
rect 217192 500896 217198 500948
rect 224862 500896 224868 500948
rect 224920 500936 224926 500948
rect 225782 500936 225788 500948
rect 224920 500908 225788 500936
rect 224920 500896 224926 500908
rect 225782 500896 225788 500908
rect 225840 500896 225846 500948
rect 229094 500896 229100 500948
rect 229152 500936 229158 500948
rect 230106 500936 230112 500948
rect 229152 500908 230112 500936
rect 229152 500896 229158 500908
rect 230106 500896 230112 500908
rect 230164 500896 230170 500948
rect 230566 500896 230572 500948
rect 230624 500936 230630 500948
rect 232222 500936 232228 500948
rect 230624 500908 232228 500936
rect 230624 500896 230630 500908
rect 232222 500896 232228 500908
rect 232280 500896 232286 500948
rect 234522 500896 234528 500948
rect 234580 500936 234586 500948
rect 235442 500936 235448 500948
rect 234580 500908 235448 500936
rect 234580 500896 234586 500908
rect 235442 500896 235448 500908
rect 235500 500896 235506 500948
rect 235902 500896 235908 500948
rect 235960 500936 235966 500948
rect 236546 500936 236552 500948
rect 235960 500908 236552 500936
rect 235960 500896 235966 500908
rect 236546 500896 236552 500908
rect 236604 500896 236610 500948
rect 255314 500896 255320 500948
rect 255372 500936 255378 500948
rect 256970 500936 256976 500948
rect 255372 500908 256976 500936
rect 255372 500896 255378 500908
rect 256970 500896 256976 500908
rect 257028 500896 257034 500948
rect 259454 500896 259460 500948
rect 259512 500936 259518 500948
rect 261294 500936 261300 500948
rect 259512 500908 261300 500936
rect 259512 500896 259518 500908
rect 261294 500896 261300 500908
rect 261352 500896 261358 500948
rect 262306 500896 262312 500948
rect 262364 500936 262370 500948
rect 263502 500936 263508 500948
rect 262364 500908 263508 500936
rect 262364 500896 262370 500908
rect 263502 500896 263508 500908
rect 263560 500896 263566 500948
rect 267918 500896 267924 500948
rect 267976 500936 267982 500948
rect 268838 500936 268844 500948
rect 267976 500908 268844 500936
rect 267976 500896 267982 500908
rect 268838 500896 268844 500908
rect 268896 500896 268902 500948
rect 269114 500896 269120 500948
rect 269172 500936 269178 500948
rect 269942 500936 269948 500948
rect 269172 500908 269948 500936
rect 269172 500896 269178 500908
rect 269942 500896 269948 500908
rect 270000 500896 270006 500948
rect 340138 500896 340144 500948
rect 340196 500936 340202 500948
rect 340782 500936 340788 500948
rect 340196 500908 340788 500936
rect 340196 500896 340202 500908
rect 340782 500896 340788 500908
rect 340840 500896 340846 500948
rect 341150 500896 341156 500948
rect 341208 500936 341214 500948
rect 342070 500936 342076 500948
rect 341208 500908 342076 500936
rect 341208 500896 341214 500908
rect 342070 500896 342076 500908
rect 342128 500896 342134 500948
rect 343174 500896 343180 500948
rect 343232 500936 343238 500948
rect 343726 500936 343732 500948
rect 343232 500908 343732 500936
rect 343232 500896 343238 500908
rect 343726 500896 343732 500908
rect 343784 500896 343790 500948
rect 345474 500896 345480 500948
rect 345532 500936 345538 500948
rect 346210 500936 346216 500948
rect 345532 500908 346216 500936
rect 345532 500896 345538 500908
rect 346210 500896 346216 500908
rect 346268 500896 346274 500948
rect 354122 500896 354128 500948
rect 354180 500936 354186 500948
rect 354582 500936 354588 500948
rect 354180 500908 354588 500936
rect 354180 500896 354186 500908
rect 354582 500896 354588 500908
rect 354640 500896 354646 500948
rect 359458 500896 359464 500948
rect 359516 500936 359522 500948
rect 360102 500936 360108 500948
rect 359516 500908 360108 500936
rect 359516 500896 359522 500908
rect 360102 500896 360108 500908
rect 360160 500896 360166 500948
rect 364886 500896 364892 500948
rect 364944 500936 364950 500948
rect 365622 500936 365628 500948
rect 364944 500908 365628 500936
rect 364944 500896 364950 500908
rect 365622 500896 365628 500908
rect 365680 500896 365686 500948
rect 365990 500896 365996 500948
rect 366048 500936 366054 500948
rect 367002 500936 367008 500948
rect 366048 500908 367008 500936
rect 366048 500896 366054 500908
rect 367002 500896 367008 500908
rect 367060 500896 367066 500948
rect 370314 500896 370320 500948
rect 370372 500936 370378 500948
rect 371142 500936 371148 500948
rect 370372 500908 371148 500936
rect 370372 500896 370378 500908
rect 371142 500896 371148 500908
rect 371200 500896 371206 500948
rect 375650 500896 375656 500948
rect 375708 500936 375714 500948
rect 376570 500936 376576 500948
rect 375708 500908 376576 500936
rect 375708 500896 375714 500908
rect 376570 500896 376576 500908
rect 376628 500896 376634 500948
rect 384298 500896 384304 500948
rect 384356 500936 384362 500948
rect 384942 500936 384948 500948
rect 384356 500908 384948 500936
rect 384356 500896 384362 500908
rect 384942 500896 384948 500908
rect 385000 500896 385006 500948
rect 385402 500896 385408 500948
rect 385460 500936 385466 500948
rect 386322 500936 386328 500948
rect 385460 500908 386328 500936
rect 385460 500896 385466 500908
rect 386322 500896 386328 500908
rect 386380 500896 386386 500948
rect 395062 500896 395068 500948
rect 395120 500936 395126 500948
rect 395982 500936 395988 500948
rect 395120 500908 395988 500936
rect 395120 500896 395126 500908
rect 395982 500896 395988 500908
rect 396040 500896 396046 500948
rect 400490 500896 400496 500948
rect 400548 500936 400554 500948
rect 401410 500936 401416 500948
rect 400548 500908 401416 500936
rect 400548 500896 400554 500908
rect 401410 500896 401416 500908
rect 401468 500896 401474 500948
rect 404722 500896 404728 500948
rect 404780 500936 404786 500948
rect 411622 500936 411628 500948
rect 404780 500908 411628 500936
rect 404780 500896 404786 500908
rect 411622 500896 411628 500908
rect 411680 500896 411686 500948
rect 420822 500896 420828 500948
rect 420880 500936 420886 500948
rect 423122 500936 423128 500948
rect 420880 500908 423128 500936
rect 420880 500896 420886 500908
rect 423122 500896 423128 500908
rect 423180 500936 423186 500948
rect 424962 500936 424968 500948
rect 423180 500908 424968 500936
rect 423180 500896 423186 500908
rect 424962 500896 424968 500908
rect 425020 500936 425026 500948
rect 427078 500936 427084 500948
rect 425020 500908 427084 500936
rect 425020 500896 425026 500908
rect 427078 500896 427084 500908
rect 427136 500936 427142 500948
rect 429286 500936 429292 500948
rect 427136 500908 429292 500936
rect 427136 500896 427142 500908
rect 429286 500896 429292 500908
rect 429344 500936 429350 500948
rect 431402 500936 431408 500948
rect 429344 500908 431408 500936
rect 429344 500896 429350 500908
rect 431402 500896 431408 500908
rect 431460 500936 431466 500948
rect 433426 500936 433432 500948
rect 431460 500908 433432 500936
rect 431460 500896 431466 500908
rect 433426 500896 433432 500908
rect 433484 500936 433490 500948
rect 435542 500936 435548 500948
rect 433484 500908 435548 500936
rect 433484 500896 433490 500908
rect 435542 500896 435548 500908
rect 435600 500936 435606 500948
rect 437566 500936 437572 500948
rect 435600 500908 437572 500936
rect 435600 500896 435606 500908
rect 437566 500896 437572 500908
rect 437624 500936 437630 500948
rect 439682 500936 439688 500948
rect 437624 500908 439688 500936
rect 437624 500896 437630 500908
rect 439682 500896 439688 500908
rect 439740 500936 439746 500948
rect 441982 500936 441988 500948
rect 439740 500908 441988 500936
rect 439740 500896 439746 500908
rect 441982 500896 441988 500908
rect 442040 500936 442046 500948
rect 444374 500936 444380 500948
rect 442040 500908 444380 500936
rect 442040 500896 442046 500908
rect 444374 500896 444380 500908
rect 444432 500936 444438 500948
rect 446306 500936 446312 500948
rect 444432 500908 446312 500936
rect 444432 500896 444438 500908
rect 446306 500896 446312 500908
rect 446364 500936 446370 500948
rect 448514 500936 448520 500948
rect 446364 500908 448520 500936
rect 446364 500896 446370 500908
rect 448514 500896 448520 500908
rect 448572 500936 448578 500948
rect 450446 500936 450452 500948
rect 448572 500908 450452 500936
rect 448572 500896 448578 500908
rect 450446 500896 450452 500908
rect 450504 500936 450510 500948
rect 453298 500936 453304 500948
rect 450504 500908 453304 500936
rect 450504 500896 450510 500908
rect 453298 500896 453304 500908
rect 453356 500936 453362 500948
rect 455322 500936 455328 500948
rect 453356 500908 455328 500936
rect 453356 500896 453362 500908
rect 455322 500896 455328 500908
rect 455380 500936 455386 500948
rect 457346 500936 457352 500948
rect 455380 500908 457352 500936
rect 455380 500896 455386 500908
rect 457346 500896 457352 500908
rect 457404 500936 457410 500948
rect 461854 500936 461860 500948
rect 457404 500908 461860 500936
rect 457404 500896 457410 500908
rect 461854 500896 461860 500908
rect 461912 500936 461918 500948
rect 464062 500936 464068 500948
rect 461912 500908 464068 500936
rect 461912 500896 461918 500908
rect 464062 500896 464068 500908
rect 464120 500936 464126 500948
rect 465902 500936 465908 500948
rect 464120 500908 465908 500936
rect 464120 500896 464126 500908
rect 465902 500896 465908 500908
rect 465960 500936 465966 500948
rect 468110 500936 468116 500948
rect 465960 500908 468116 500936
rect 465960 500896 465966 500908
rect 468110 500896 468116 500908
rect 468168 500936 468174 500948
rect 470226 500936 470232 500948
rect 468168 500908 470232 500936
rect 468168 500896 468174 500908
rect 470226 500896 470232 500908
rect 470284 500936 470290 500948
rect 472710 500936 472716 500948
rect 470284 500908 472716 500936
rect 470284 500896 470290 500908
rect 472710 500896 472716 500908
rect 472768 500936 472774 500948
rect 474642 500936 474648 500948
rect 472768 500908 474648 500936
rect 472768 500896 472774 500908
rect 474642 500896 474648 500908
rect 474700 500936 474706 500948
rect 477770 500936 477776 500948
rect 474700 500908 477776 500936
rect 474700 500896 474706 500908
rect 477770 500896 477776 500908
rect 477828 500936 477834 500948
rect 480806 500936 480812 500948
rect 477828 500908 480812 500936
rect 477828 500896 477834 500908
rect 480806 500896 480812 500908
rect 480864 500896 480870 500948
rect 492030 500896 492036 500948
rect 492088 500936 492094 500948
rect 492582 500936 492588 500948
rect 492088 500908 492588 500936
rect 492088 500896 492094 500908
rect 492582 500896 492588 500908
rect 492640 500896 492646 500948
rect 498378 500896 498384 500948
rect 498436 500936 498442 500948
rect 498930 500936 498936 500948
rect 498436 500908 498936 500936
rect 498436 500896 498442 500908
rect 498930 500896 498936 500908
rect 498988 500896 498994 500948
rect 502426 500896 502432 500948
rect 502484 500936 502490 500948
rect 503254 500936 503260 500948
rect 502484 500908 503260 500936
rect 502484 500896 502490 500908
rect 503254 500896 503260 500908
rect 503312 500896 503318 500948
rect 509234 500896 509240 500948
rect 509292 500936 509298 500948
rect 509786 500936 509792 500948
rect 509292 500908 509792 500936
rect 509292 500896 509298 500908
rect 509786 500896 509792 500908
rect 509844 500896 509850 500948
rect 511442 500896 511448 500948
rect 511500 500936 511506 500948
rect 511902 500936 511908 500948
rect 511500 500908 511908 500936
rect 511500 500896 511506 500908
rect 511902 500896 511908 500908
rect 511960 500896 511966 500948
rect 522206 500896 522212 500948
rect 522264 500936 522270 500948
rect 522942 500936 522948 500948
rect 522264 500908 522948 500936
rect 522264 500896 522270 500908
rect 522942 500896 522948 500908
rect 523000 500896 523006 500948
rect 527634 500896 527640 500948
rect 527692 500936 527698 500948
rect 528370 500936 528376 500948
rect 527692 500908 528376 500936
rect 527692 500896 527698 500908
rect 528370 500896 528376 500908
rect 528428 500896 528434 500948
rect 531958 500896 531964 500948
rect 532016 500936 532022 500948
rect 532602 500936 532608 500948
rect 532016 500908 532608 500936
rect 532016 500896 532022 500908
rect 532602 500896 532608 500908
rect 532660 500896 532666 500948
rect 533062 500896 533068 500948
rect 533120 500936 533126 500948
rect 533982 500936 533988 500948
rect 533120 500908 533988 500936
rect 533120 500896 533126 500908
rect 533982 500896 533988 500908
rect 534040 500896 534046 500948
rect 536282 500896 536288 500948
rect 536340 500936 536346 500948
rect 536742 500936 536748 500948
rect 536340 500908 536748 500936
rect 536340 500896 536346 500908
rect 536742 500896 536748 500908
rect 536800 500896 536806 500948
rect 541618 500896 541624 500948
rect 541676 500936 541682 500948
rect 542262 500936 542268 500948
rect 541676 500908 542268 500936
rect 541676 500896 541682 500908
rect 542262 500896 542268 500908
rect 542320 500896 542326 500948
rect 545942 500896 545948 500948
rect 546000 500936 546006 500948
rect 546402 500936 546408 500948
rect 546000 500908 546408 500936
rect 546000 500896 546006 500908
rect 546402 500896 546408 500908
rect 546460 500896 546466 500948
rect 547046 500896 547052 500948
rect 547104 500936 547110 500948
rect 547782 500936 547788 500948
rect 547104 500908 547788 500936
rect 547104 500896 547110 500908
rect 547782 500896 547788 500908
rect 547840 500896 547846 500948
rect 553302 500896 553308 500948
rect 553360 500936 553366 500948
rect 554038 500936 554044 500948
rect 553360 500908 554044 500936
rect 553360 500896 553366 500908
rect 554038 500896 554044 500908
rect 554096 500896 554102 500948
rect 558178 500896 558184 500948
rect 558236 500936 558242 500948
rect 559282 500936 559288 500948
rect 558236 500908 559288 500936
rect 558236 500896 558242 500908
rect 559282 500896 559288 500908
rect 559340 500896 559346 500948
rect 31662 500828 31668 500880
rect 31720 500868 31726 500880
rect 31754 500868 31760 500880
rect 31720 500840 31760 500868
rect 31720 500828 31726 500840
rect 31754 500828 31760 500840
rect 31812 500828 31818 500880
rect 45738 500828 45744 500880
rect 45796 500868 45802 500880
rect 53926 500868 53932 500880
rect 45796 500840 53932 500868
rect 45796 500828 45802 500840
rect 53926 500828 53932 500840
rect 53984 500828 53990 500880
rect 126606 500828 126612 500880
rect 126664 500868 126670 500880
rect 153378 500868 153384 500880
rect 126664 500840 153384 500868
rect 126664 500828 126670 500840
rect 153378 500828 153384 500840
rect 153436 500828 153442 500880
rect 195330 500828 195336 500880
rect 195388 500868 195394 500880
rect 198826 500868 198832 500880
rect 195388 500840 198832 500868
rect 195388 500828 195394 500840
rect 198826 500828 198832 500840
rect 198884 500828 198890 500880
rect 200206 500828 200212 500880
rect 200264 500868 200270 500880
rect 205266 500868 205272 500880
rect 200264 500840 205272 500868
rect 200264 500828 200270 500840
rect 205266 500828 205272 500840
rect 205324 500828 205330 500880
rect 205634 500828 205640 500880
rect 205692 500868 205698 500880
rect 209590 500868 209596 500880
rect 205692 500840 209596 500868
rect 205692 500828 205698 500840
rect 209590 500828 209596 500840
rect 209648 500828 209654 500880
rect 213454 500828 213460 500880
rect 213512 500868 213518 500880
rect 216030 500868 216036 500880
rect 213512 500840 216036 500868
rect 213512 500828 213518 500840
rect 216030 500828 216036 500840
rect 216088 500828 216094 500880
rect 251174 500828 251180 500880
rect 251232 500868 251238 500880
rect 253750 500868 253756 500880
rect 251232 500840 253756 500868
rect 251232 500828 251238 500840
rect 253750 500828 253756 500840
rect 253808 500828 253814 500880
rect 253934 500828 253940 500880
rect 253992 500868 253998 500880
rect 255958 500868 255964 500880
rect 253992 500840 255964 500868
rect 253992 500828 253998 500840
rect 255958 500828 255964 500840
rect 256016 500828 256022 500880
rect 260834 500828 260840 500880
rect 260892 500868 260898 500880
rect 262398 500868 262404 500880
rect 260892 500840 262404 500868
rect 260892 500828 260898 500840
rect 262398 500828 262404 500840
rect 262456 500828 262462 500880
rect 403710 500828 403716 500880
rect 403768 500868 403774 500880
rect 409874 500868 409880 500880
rect 403768 500840 409880 500868
rect 403768 500828 403774 500840
rect 409874 500828 409880 500840
rect 409932 500828 409938 500880
rect 129826 500760 129832 500812
rect 129884 500800 129890 500812
rect 153286 500800 153292 500812
rect 129884 500772 153292 500800
rect 129884 500760 129890 500772
rect 153286 500760 153292 500772
rect 153344 500760 153350 500812
rect 214926 500760 214932 500812
rect 214984 500800 214990 500812
rect 218238 500800 218244 500812
rect 214984 500772 218244 500800
rect 214984 500760 214990 500772
rect 218238 500760 218244 500772
rect 218296 500760 218302 500812
rect 355226 500760 355232 500812
rect 355284 500800 355290 500812
rect 355962 500800 355968 500812
rect 355284 500772 355968 500800
rect 355284 500760 355290 500772
rect 355962 500760 355968 500772
rect 356020 500760 356026 500812
rect 547877 500803 547935 500809
rect 547877 500769 547889 500803
rect 547923 500800 547935 500803
rect 554130 500800 554136 500812
rect 547923 500772 554136 500800
rect 547923 500769 547935 500772
rect 547877 500763 547935 500769
rect 554130 500760 554136 500772
rect 554188 500760 554194 500812
rect 41414 500692 41420 500744
rect 41472 500732 41478 500744
rect 47026 500732 47032 500744
rect 41472 500704 47032 500732
rect 41472 500692 41478 500704
rect 47026 500692 47032 500704
rect 47084 500692 47090 500744
rect 128722 500692 128728 500744
rect 128780 500732 128786 500744
rect 151906 500732 151912 500744
rect 128780 500704 151912 500732
rect 128780 500692 128786 500704
rect 151906 500692 151912 500704
rect 151964 500692 151970 500744
rect 197170 500692 197176 500744
rect 197228 500732 197234 500744
rect 202046 500732 202052 500744
rect 197228 500704 202052 500732
rect 197228 500692 197234 500704
rect 202046 500692 202052 500704
rect 202104 500692 202110 500744
rect 211338 500692 211344 500744
rect 211396 500732 211402 500744
rect 215018 500732 215024 500744
rect 211396 500704 215024 500732
rect 211396 500692 211402 500704
rect 215018 500692 215024 500704
rect 215076 500692 215082 500744
rect 542722 500692 542728 500744
rect 542780 500732 542786 500744
rect 551370 500732 551376 500744
rect 542780 500704 551376 500732
rect 542780 500692 542786 500704
rect 551370 500692 551376 500704
rect 551428 500692 551434 500744
rect 130930 500624 130936 500676
rect 130988 500664 130994 500676
rect 154758 500664 154764 500676
rect 130988 500636 154764 500664
rect 130988 500624 130994 500636
rect 154758 500624 154764 500636
rect 154816 500624 154822 500676
rect 223482 500624 223488 500676
rect 223540 500664 223546 500676
rect 224678 500664 224684 500676
rect 223540 500636 224684 500664
rect 223540 500624 223546 500636
rect 224678 500624 224684 500636
rect 224736 500624 224742 500676
rect 350902 500624 350908 500676
rect 350960 500664 350966 500676
rect 351822 500664 351828 500676
rect 350960 500636 351828 500664
rect 350960 500624 350966 500636
rect 351822 500624 351828 500636
rect 351880 500624 351886 500676
rect 507118 500624 507124 500676
rect 507176 500664 507182 500676
rect 507762 500664 507768 500676
rect 507176 500636 507768 500664
rect 507176 500624 507182 500636
rect 507762 500624 507768 500636
rect 507820 500624 507826 500676
rect 544838 500624 544844 500676
rect 544896 500664 544902 500676
rect 547877 500667 547935 500673
rect 547877 500664 547889 500667
rect 544896 500636 547889 500664
rect 544896 500624 544902 500636
rect 547877 500633 547889 500636
rect 547923 500633 547935 500667
rect 547877 500627 547935 500633
rect 127710 500556 127716 500608
rect 127768 500596 127774 500608
rect 154482 500596 154488 500608
rect 127768 500568 154488 500596
rect 127768 500556 127774 500568
rect 154482 500556 154488 500568
rect 154540 500556 154546 500608
rect 201586 500556 201592 500608
rect 201644 500596 201650 500608
rect 206370 500596 206376 500608
rect 201644 500568 206376 500596
rect 201644 500556 201650 500568
rect 206370 500556 206376 500568
rect 206428 500556 206434 500608
rect 215294 500556 215300 500608
rect 215352 500596 215358 500608
rect 219250 500596 219256 500608
rect 215352 500568 219256 500596
rect 215352 500556 215358 500568
rect 219250 500556 219256 500568
rect 219308 500556 219314 500608
rect 219526 500556 219532 500608
rect 219584 500596 219590 500608
rect 222562 500596 222568 500608
rect 219584 500568 222568 500596
rect 219584 500556 219590 500568
rect 222562 500556 222568 500568
rect 222620 500556 222626 500608
rect 533890 500556 533896 500608
rect 533948 500596 533954 500608
rect 554222 500596 554228 500608
rect 533948 500568 554228 500596
rect 533948 500556 533954 500568
rect 554222 500556 554228 500568
rect 554280 500556 554286 500608
rect 124398 500488 124404 500540
rect 124456 500528 124462 500540
rect 151998 500528 152004 500540
rect 124456 500500 152004 500528
rect 124456 500488 124462 500500
rect 151998 500488 152004 500500
rect 152056 500488 152062 500540
rect 196066 500488 196072 500540
rect 196124 500528 196130 500540
rect 200942 500528 200948 500540
rect 196124 500500 200948 500528
rect 196124 500488 196130 500500
rect 200942 500488 200948 500500
rect 201000 500488 201006 500540
rect 363782 500488 363788 500540
rect 363840 500528 363846 500540
rect 364242 500528 364248 500540
rect 363840 500500 364248 500528
rect 363840 500488 363846 500500
rect 364242 500488 364248 500500
rect 364300 500488 364306 500540
rect 523310 500488 523316 500540
rect 523368 500528 523374 500540
rect 547877 500531 547935 500537
rect 547877 500528 547889 500531
rect 523368 500500 547889 500528
rect 523368 500488 523374 500500
rect 547877 500497 547889 500500
rect 547923 500497 547935 500531
rect 547877 500491 547935 500497
rect 548150 500488 548156 500540
rect 548208 500528 548214 500540
rect 549162 500528 549168 500540
rect 548208 500500 549168 500528
rect 548208 500488 548214 500500
rect 549162 500488 549168 500500
rect 549220 500488 549226 500540
rect 42518 500420 42524 500472
rect 42576 500460 42582 500472
rect 47578 500460 47584 500472
rect 42576 500432 47584 500460
rect 42576 500420 42582 500432
rect 47578 500420 47584 500432
rect 47636 500420 47642 500472
rect 125502 500420 125508 500472
rect 125560 500460 125566 500472
rect 153378 500460 153384 500472
rect 125560 500432 153384 500460
rect 125560 500420 125566 500432
rect 153378 500420 153384 500432
rect 153436 500420 153442 500472
rect 187786 500420 187792 500472
rect 187844 500460 187850 500472
rect 192386 500460 192392 500472
rect 187844 500432 192392 500460
rect 187844 500420 187850 500432
rect 192386 500420 192392 500432
rect 192444 500420 192450 500472
rect 199470 500420 199476 500472
rect 199528 500460 199534 500472
rect 204162 500460 204168 500472
rect 199528 500432 204168 500460
rect 199528 500420 199534 500432
rect 204162 500420 204168 500432
rect 204220 500420 204226 500472
rect 209866 500420 209872 500472
rect 209924 500460 209930 500472
rect 213914 500460 213920 500472
rect 209924 500432 213920 500460
rect 209924 500420 209930 500432
rect 213914 500420 213920 500432
rect 213972 500420 213978 500472
rect 218146 500420 218152 500472
rect 218204 500460 218210 500472
rect 221458 500460 221464 500472
rect 218204 500432 221464 500460
rect 218204 500420 218210 500432
rect 221458 500420 221464 500432
rect 221516 500420 221522 500472
rect 224218 500420 224224 500472
rect 224276 500460 224282 500472
rect 226794 500460 226800 500472
rect 224276 500432 226800 500460
rect 224276 500420 224282 500432
rect 226794 500420 226800 500432
rect 226852 500420 226858 500472
rect 515766 500420 515772 500472
rect 515824 500460 515830 500472
rect 551462 500460 551468 500472
rect 515824 500432 551468 500460
rect 515824 500420 515830 500432
rect 551462 500420 551468 500432
rect 551520 500420 551526 500472
rect 43622 500352 43628 500404
rect 43680 500392 43686 500404
rect 48958 500392 48964 500404
rect 43680 500364 48964 500392
rect 43680 500352 43686 500364
rect 48958 500352 48964 500364
rect 49016 500352 49022 500404
rect 123386 500352 123392 500404
rect 123444 500392 123450 500404
rect 153470 500392 153476 500404
rect 123444 500364 153476 500392
rect 123444 500352 123450 500364
rect 153470 500352 153476 500364
rect 153528 500352 153534 500404
rect 209130 500352 209136 500404
rect 209188 500392 209194 500404
rect 212810 500392 212816 500404
rect 209188 500364 212816 500392
rect 209188 500352 209194 500364
rect 212810 500352 212816 500364
rect 212868 500352 212874 500404
rect 322842 500352 322848 500404
rect 322900 500392 322906 500404
rect 323302 500392 323308 500404
rect 322900 500364 323308 500392
rect 322900 500352 322906 500364
rect 323302 500352 323308 500364
rect 323360 500352 323366 500404
rect 349798 500352 349804 500404
rect 349856 500392 349862 500404
rect 350442 500392 350448 500404
rect 349856 500364 350448 500392
rect 349856 500352 349862 500364
rect 350442 500352 350448 500364
rect 350500 500352 350506 500404
rect 398282 500352 398288 500404
rect 398340 500392 398346 500404
rect 398742 500392 398748 500404
rect 398340 500364 398748 500392
rect 398340 500352 398346 500364
rect 398742 500352 398748 500364
rect 398800 500352 398806 500404
rect 506106 500352 506112 500404
rect 506164 500392 506170 500404
rect 512638 500392 512644 500404
rect 506164 500364 512644 500392
rect 506164 500352 506170 500364
rect 512638 500352 512644 500364
rect 512696 500352 512702 500404
rect 513650 500352 513656 500404
rect 513708 500392 513714 500404
rect 551554 500392 551560 500404
rect 513708 500364 551560 500392
rect 513708 500352 513714 500364
rect 551554 500352 551560 500364
rect 551612 500352 551618 500404
rect 44726 500284 44732 500336
rect 44784 500324 44790 500336
rect 52546 500324 52552 500336
rect 44784 500296 52552 500324
rect 44784 500284 44790 500296
rect 52546 500284 52552 500296
rect 52604 500284 52610 500336
rect 55490 500284 55496 500336
rect 55548 500324 55554 500336
rect 56410 500324 56416 500336
rect 55548 500296 56416 500324
rect 55548 500284 55554 500296
rect 56410 500284 56416 500296
rect 56468 500284 56474 500336
rect 120258 500284 120264 500336
rect 120316 500324 120322 500336
rect 153838 500324 153844 500336
rect 120316 500296 153844 500324
rect 120316 500284 120322 500296
rect 153838 500284 153844 500296
rect 153896 500284 153902 500336
rect 509050 500284 509056 500336
rect 509108 500324 509114 500336
rect 551646 500324 551652 500336
rect 509108 500296 551652 500324
rect 509108 500284 509114 500296
rect 551646 500284 551652 500296
rect 551704 500284 551710 500336
rect 85666 500216 85672 500268
rect 85724 500256 85730 500268
rect 112438 500256 112444 500268
rect 85724 500228 112444 500256
rect 85724 500216 85730 500228
rect 112438 500216 112444 500228
rect 112496 500216 112502 500268
rect 117314 500216 117320 500268
rect 117372 500256 117378 500268
rect 153102 500256 153108 500268
rect 117372 500228 153108 500256
rect 117372 500216 117378 500228
rect 153102 500216 153108 500228
rect 153160 500216 153166 500268
rect 187878 500216 187884 500268
rect 187936 500256 187942 500268
rect 193398 500256 193404 500268
rect 187936 500228 193404 500256
rect 187936 500216 187942 500228
rect 193398 500216 193404 500228
rect 193456 500216 193462 500268
rect 195606 500216 195612 500268
rect 195664 500256 195670 500268
rect 279602 500256 279608 500268
rect 195664 500228 279608 500256
rect 195664 500216 195670 500228
rect 279602 500216 279608 500228
rect 279660 500216 279666 500268
rect 289722 500216 289728 500268
rect 289780 500256 289786 500268
rect 416130 500256 416136 500268
rect 289780 500228 416136 500256
rect 289780 500216 289786 500228
rect 416130 500216 416136 500228
rect 416188 500216 416194 500268
rect 498562 500216 498568 500268
rect 498620 500256 498626 500268
rect 499482 500256 499488 500268
rect 498620 500228 499488 500256
rect 498620 500216 498626 500228
rect 499482 500216 499488 500228
rect 499540 500216 499546 500268
rect 502886 500216 502892 500268
rect 502944 500256 502950 500268
rect 551738 500256 551744 500268
rect 502944 500228 551744 500256
rect 502944 500216 502950 500228
rect 551738 500216 551744 500228
rect 551796 500216 551802 500268
rect 556798 500216 556804 500268
rect 556856 500256 556862 500268
rect 571334 500256 571340 500268
rect 556856 500228 571340 500256
rect 556856 500216 556862 500228
rect 571334 500216 571340 500228
rect 571392 500216 571398 500268
rect 70578 500148 70584 500200
rect 70636 500188 70642 500200
rect 89717 500191 89775 500197
rect 89717 500188 89729 500191
rect 70636 500160 89729 500188
rect 70636 500148 70642 500160
rect 89717 500157 89729 500160
rect 89763 500157 89775 500191
rect 89717 500151 89775 500157
rect 131942 500148 131948 500200
rect 132000 500188 132006 500200
rect 154390 500188 154396 500200
rect 132000 500160 154396 500188
rect 132000 500148 132006 500160
rect 154390 500148 154396 500160
rect 154448 500148 154454 500200
rect 547877 500191 547935 500197
rect 547877 500157 547889 500191
rect 547923 500188 547935 500191
rect 549898 500188 549904 500200
rect 547923 500160 549904 500188
rect 547923 500157 547935 500160
rect 547877 500151 547935 500157
rect 549898 500148 549904 500160
rect 549956 500148 549962 500200
rect 65150 500080 65156 500132
rect 65208 500120 65214 500132
rect 66162 500120 66168 500132
rect 65208 500092 66168 500120
rect 65208 500080 65214 500092
rect 66162 500080 66168 500092
rect 66220 500080 66226 500132
rect 135254 500080 135260 500132
rect 135312 500120 135318 500132
rect 154298 500120 154304 500132
rect 135312 500092 154304 500120
rect 135312 500080 135318 500092
rect 154298 500080 154304 500092
rect 154356 500080 154362 500132
rect 220814 500080 220820 500132
rect 220872 500120 220878 500132
rect 223574 500120 223580 500132
rect 220872 500092 223580 500120
rect 220872 500080 220878 500092
rect 223574 500080 223580 500092
rect 223632 500080 223638 500132
rect 369210 500080 369216 500132
rect 369268 500120 369274 500132
rect 369762 500120 369768 500132
rect 369268 500092 369768 500120
rect 369268 500080 369274 500092
rect 369762 500080 369768 500092
rect 369820 500080 369826 500132
rect 379974 500080 379980 500132
rect 380032 500120 380038 500132
rect 380802 500120 380808 500132
rect 380032 500092 380808 500120
rect 380032 500080 380038 500092
rect 380802 500080 380808 500092
rect 380860 500080 380866 500132
rect 89717 500055 89775 500061
rect 89717 500021 89729 500055
rect 89763 500052 89775 500055
rect 94498 500052 94504 500064
rect 89763 500024 94504 500052
rect 89763 500021 89775 500024
rect 89717 500015 89775 500021
rect 94498 500012 94504 500024
rect 94556 500012 94562 500064
rect 137370 500012 137376 500064
rect 137428 500052 137434 500064
rect 154114 500052 154120 500064
rect 137428 500024 154120 500052
rect 137428 500012 137434 500024
rect 154114 500012 154120 500024
rect 154172 500012 154178 500064
rect 191834 500012 191840 500064
rect 191892 500052 191898 500064
rect 199930 500052 199936 500064
rect 191892 500024 199936 500052
rect 191892 500012 191898 500024
rect 199930 500012 199936 500024
rect 199988 500012 199994 500064
rect 501782 500012 501788 500064
rect 501840 500052 501846 500064
rect 502242 500052 502248 500064
rect 501840 500024 502248 500052
rect 501840 500012 501846 500024
rect 502242 500012 502248 500024
rect 502300 500012 502306 500064
rect 516870 500012 516876 500064
rect 516928 500052 516934 500064
rect 517422 500052 517428 500064
rect 516928 500024 517428 500052
rect 516928 500012 516934 500024
rect 517422 500012 517428 500024
rect 517480 500012 517486 500064
rect 140590 499944 140596 499996
rect 140648 499984 140654 499996
rect 154206 499984 154212 499996
rect 140648 499956 154212 499984
rect 140648 499944 140654 499956
rect 154206 499944 154212 499956
rect 154264 499944 154270 499996
rect 360562 499944 360568 499996
rect 360620 499984 360626 499996
rect 361482 499984 361488 499996
rect 360620 499956 361488 499984
rect 360620 499944 360626 499956
rect 361482 499944 361488 499956
rect 361540 499944 361546 499996
rect 374546 499944 374552 499996
rect 374604 499984 374610 499996
rect 375282 499984 375288 499996
rect 374604 499956 375288 499984
rect 374604 499944 374610 499956
rect 375282 499944 375288 499956
rect 375340 499944 375346 499996
rect 378870 499944 378876 499996
rect 378928 499984 378934 499996
rect 379422 499984 379428 499996
rect 378928 499956 379428 499984
rect 378928 499944 378934 499956
rect 379422 499944 379428 499956
rect 379480 499944 379486 499996
rect 389634 499944 389640 499996
rect 389692 499984 389698 499996
rect 390462 499984 390468 499996
rect 389692 499956 390468 499984
rect 389692 499944 389698 499956
rect 390462 499944 390468 499956
rect 390520 499944 390526 499996
rect 393958 499944 393964 499996
rect 394016 499984 394022 499996
rect 394602 499984 394608 499996
rect 394016 499956 394608 499984
rect 394016 499944 394022 499956
rect 394602 499944 394608 499956
rect 394660 499944 394666 499996
rect 399386 499944 399392 499996
rect 399444 499984 399450 499996
rect 400122 499984 400128 499996
rect 399444 499956 400128 499984
rect 399444 499944 399450 499956
rect 400122 499944 400128 499956
rect 400180 499944 400186 499996
rect 526530 499944 526536 499996
rect 526588 499984 526594 499996
rect 527082 499984 527088 499996
rect 526588 499956 527088 499984
rect 526588 499944 526594 499956
rect 527082 499944 527088 499956
rect 527140 499944 527146 499996
rect 537294 499944 537300 499996
rect 537352 499984 537358 499996
rect 538122 499984 538128 499996
rect 537352 499956 538128 499984
rect 537352 499944 537358 499956
rect 538122 499944 538128 499956
rect 538180 499944 538186 499996
rect 139486 499876 139492 499928
rect 139544 499916 139550 499928
rect 154022 499916 154028 499928
rect 139544 499888 154028 499916
rect 139544 499876 139550 499888
rect 154022 499876 154028 499888
rect 154080 499876 154086 499928
rect 223574 499876 223580 499928
rect 223632 499916 223638 499928
rect 229002 499916 229008 499928
rect 223632 499888 229008 499916
rect 223632 499876 223638 499888
rect 229002 499876 229008 499888
rect 229060 499876 229066 499928
rect 388622 499876 388628 499928
rect 388680 499916 388686 499928
rect 389082 499916 389088 499928
rect 388680 499888 389088 499916
rect 388680 499876 388686 499888
rect 389082 499876 389088 499888
rect 389140 499876 389146 499928
rect 141694 499808 141700 499860
rect 141752 499848 141758 499860
rect 153930 499848 153936 499860
rect 141752 499820 153936 499848
rect 141752 499808 141758 499820
rect 153930 499808 153936 499820
rect 153988 499808 153994 499860
rect 344370 499808 344376 499860
rect 344428 499848 344434 499860
rect 344922 499848 344928 499860
rect 344428 499820 344928 499848
rect 344428 499808 344434 499820
rect 344922 499808 344928 499820
rect 344980 499808 344986 499860
rect 493134 499808 493140 499860
rect 493192 499848 493198 499860
rect 494698 499848 494704 499860
rect 493192 499820 494704 499848
rect 493192 499808 493198 499820
rect 494698 499808 494704 499820
rect 494756 499808 494762 499860
rect 517974 499808 517980 499860
rect 518032 499848 518038 499860
rect 518802 499848 518808 499860
rect 518032 499820 518808 499848
rect 518032 499808 518038 499820
rect 518802 499808 518808 499820
rect 518860 499808 518866 499860
rect 22094 499740 22100 499792
rect 22152 499780 22158 499792
rect 24118 499780 24124 499792
rect 22152 499752 24124 499780
rect 22152 499740 22158 499752
rect 24118 499740 24124 499752
rect 24176 499740 24182 499792
rect 51166 499740 51172 499792
rect 51224 499780 51230 499792
rect 52362 499780 52368 499792
rect 51224 499752 52368 499780
rect 51224 499740 51230 499752
rect 52362 499740 52368 499752
rect 52420 499740 52426 499792
rect 66254 499740 66260 499792
rect 66312 499780 66318 499792
rect 67542 499780 67548 499792
rect 66312 499752 67548 499780
rect 66312 499740 66318 499752
rect 67542 499740 67548 499752
rect 67600 499740 67606 499792
rect 142798 499740 142804 499792
rect 142856 499780 142862 499792
rect 153654 499780 153660 499792
rect 142856 499752 153660 499780
rect 142856 499740 142862 499752
rect 153654 499740 153660 499752
rect 153712 499740 153718 499792
rect 191926 499740 191932 499792
rect 191984 499780 191990 499792
rect 196618 499780 196624 499792
rect 191984 499752 196624 499780
rect 191984 499740 191990 499752
rect 196618 499740 196624 499752
rect 196676 499740 196682 499792
rect 233050 499740 233056 499792
rect 233108 499780 233114 499792
rect 234338 499780 234344 499792
rect 233108 499752 234344 499780
rect 233108 499740 233114 499752
rect 234338 499740 234344 499752
rect 234396 499740 234402 499792
rect 259362 499740 259368 499792
rect 259420 499780 259426 499792
rect 260282 499780 260288 499792
rect 259420 499752 260288 499780
rect 259420 499740 259426 499752
rect 260282 499740 260288 499752
rect 260340 499740 260346 499792
rect 263594 499740 263600 499792
rect 263652 499780 263658 499792
rect 264514 499780 264520 499792
rect 263652 499752 264520 499780
rect 263652 499740 263658 499752
rect 264514 499740 264520 499752
rect 264572 499740 264578 499792
rect 549070 499740 549076 499792
rect 549128 499780 549134 499792
rect 551278 499780 551284 499792
rect 549128 499752 551284 499780
rect 549128 499740 549134 499752
rect 551278 499740 551284 499752
rect 551336 499740 551342 499792
rect 24302 499672 24308 499724
rect 24360 499712 24366 499724
rect 26326 499712 26332 499724
rect 24360 499684 26332 499712
rect 24360 499672 24366 499684
rect 26326 499672 26332 499684
rect 26384 499672 26390 499724
rect 143810 499672 143816 499724
rect 143868 499712 143874 499724
rect 153562 499712 153568 499724
rect 143868 499684 153568 499712
rect 143868 499672 143874 499684
rect 153562 499672 153568 499684
rect 153620 499672 153626 499724
rect 206370 499672 206376 499724
rect 206428 499712 206434 499724
rect 210694 499712 210700 499724
rect 206428 499684 210700 499712
rect 206428 499672 206434 499684
rect 210694 499672 210700 499684
rect 210752 499672 210758 499724
rect 26142 499604 26148 499656
rect 26200 499644 26206 499656
rect 28534 499644 28540 499656
rect 26200 499616 28540 499644
rect 26200 499604 26206 499616
rect 28534 499604 28540 499616
rect 28592 499604 28598 499656
rect 103974 499604 103980 499656
rect 104032 499644 104038 499656
rect 104802 499644 104808 499656
rect 104032 499616 104808 499644
rect 104032 499604 104038 499616
rect 104802 499604 104808 499616
rect 104860 499604 104866 499656
rect 203702 499604 203708 499656
rect 203760 499644 203766 499656
rect 207474 499644 207480 499656
rect 203760 499616 207480 499644
rect 203760 499604 203766 499616
rect 207474 499604 207480 499616
rect 207532 499604 207538 499656
rect 207750 499604 207756 499656
rect 207808 499644 207814 499656
rect 211706 499644 211712 499656
rect 207808 499616 211712 499644
rect 207808 499604 207814 499616
rect 211706 499604 211712 499616
rect 211764 499604 211770 499656
rect 216674 499604 216680 499656
rect 216732 499644 216738 499656
rect 220354 499644 220360 499656
rect 216732 499616 220360 499644
rect 216732 499604 216738 499616
rect 220354 499604 220360 499616
rect 220412 499604 220418 499656
rect 252646 499604 252652 499656
rect 252704 499644 252710 499656
rect 254854 499644 254860 499656
rect 252704 499616 254860 499644
rect 252704 499604 252710 499616
rect 254854 499604 254860 499616
rect 254912 499604 254918 499656
rect 271966 499604 271972 499656
rect 272024 499644 272030 499656
rect 273162 499644 273168 499656
rect 272024 499616 273168 499644
rect 272024 499604 272030 499616
rect 273162 499604 273168 499616
rect 273220 499604 273226 499656
rect 25498 499536 25504 499588
rect 25556 499576 25562 499588
rect 27430 499576 27436 499588
rect 25556 499548 27436 499576
rect 25556 499536 25562 499548
rect 27430 499536 27436 499548
rect 27488 499536 27494 499588
rect 31938 499536 31944 499588
rect 31996 499576 32002 499588
rect 32858 499576 32864 499588
rect 31996 499548 32864 499576
rect 31996 499536 32002 499548
rect 32858 499536 32864 499548
rect 32916 499536 32922 499588
rect 34974 499536 34980 499588
rect 35032 499576 35038 499588
rect 35802 499576 35808 499588
rect 35032 499548 35808 499576
rect 35032 499536 35038 499548
rect 35802 499536 35808 499548
rect 35860 499536 35866 499588
rect 36078 499536 36084 499588
rect 36136 499576 36142 499588
rect 37090 499576 37096 499588
rect 36136 499548 37096 499576
rect 36136 499536 36142 499548
rect 37090 499536 37096 499548
rect 37148 499536 37154 499588
rect 40402 499536 40408 499588
rect 40460 499576 40466 499588
rect 41322 499576 41328 499588
rect 40460 499548 41328 499576
rect 40460 499536 40466 499548
rect 41322 499536 41328 499548
rect 41380 499536 41386 499588
rect 75914 499536 75920 499588
rect 75972 499576 75978 499588
rect 77202 499576 77208 499588
rect 75972 499548 77208 499576
rect 75972 499536 75978 499548
rect 77202 499536 77208 499548
rect 77260 499536 77266 499588
rect 79134 499536 79140 499588
rect 79192 499576 79198 499588
rect 79962 499576 79968 499588
rect 79192 499548 79968 499576
rect 79192 499536 79198 499548
rect 79962 499536 79968 499548
rect 80020 499536 80026 499588
rect 80238 499536 80244 499588
rect 80296 499576 80302 499588
rect 81250 499576 81256 499588
rect 80296 499548 81256 499576
rect 80296 499536 80302 499548
rect 81250 499536 81256 499548
rect 81308 499536 81314 499588
rect 84562 499536 84568 499588
rect 84620 499576 84626 499588
rect 85482 499576 85488 499588
rect 84620 499548 85488 499576
rect 84620 499536 84626 499548
rect 85482 499536 85488 499548
rect 85540 499536 85546 499588
rect 86954 499536 86960 499588
rect 87012 499576 87018 499588
rect 87782 499576 87788 499588
rect 87012 499548 87788 499576
rect 87012 499536 87018 499548
rect 87782 499536 87788 499548
rect 87840 499536 87846 499588
rect 88886 499536 88892 499588
rect 88944 499576 88950 499588
rect 89622 499576 89628 499588
rect 88944 499548 89628 499576
rect 88944 499536 88950 499548
rect 89622 499536 89628 499548
rect 89680 499536 89686 499588
rect 89990 499536 89996 499588
rect 90048 499576 90054 499588
rect 91002 499576 91008 499588
rect 90048 499548 91008 499576
rect 90048 499536 90054 499548
rect 91002 499536 91008 499548
rect 91060 499536 91066 499588
rect 94222 499536 94228 499588
rect 94280 499576 94286 499588
rect 95142 499576 95148 499588
rect 94280 499548 95148 499576
rect 94280 499536 94286 499548
rect 95142 499536 95148 499548
rect 95200 499536 95206 499588
rect 95326 499536 95332 499588
rect 95384 499576 95390 499588
rect 96522 499576 96528 499588
rect 95384 499548 96528 499576
rect 95384 499536 95390 499548
rect 96522 499536 96528 499548
rect 96580 499536 96586 499588
rect 144914 499536 144920 499588
rect 144972 499576 144978 499588
rect 153746 499576 153752 499588
rect 144972 499548 153752 499576
rect 144972 499536 144978 499548
rect 153746 499536 153752 499548
rect 153804 499536 153810 499588
rect 230382 499536 230388 499588
rect 230440 499576 230446 499588
rect 231118 499576 231124 499588
rect 230440 499548 231124 499576
rect 230440 499536 230446 499548
rect 231118 499536 231124 499548
rect 231176 499536 231182 499588
rect 247034 499536 247040 499588
rect 247092 499576 247098 499588
rect 249426 499576 249432 499588
rect 247092 499548 249432 499576
rect 247092 499536 247098 499548
rect 249426 499536 249432 499548
rect 249484 499536 249490 499588
rect 256786 499536 256792 499588
rect 256844 499576 256850 499588
rect 259178 499576 259184 499588
rect 256844 499548 259184 499576
rect 256844 499536 256850 499548
rect 259178 499536 259184 499548
rect 259236 499536 259242 499588
rect 266354 499536 266360 499588
rect 266412 499576 266418 499588
rect 267826 499576 267832 499588
rect 266412 499548 267832 499576
rect 266412 499536 266418 499548
rect 267826 499536 267832 499548
rect 267884 499536 267890 499588
rect 277578 499536 277584 499588
rect 277636 499576 277642 499588
rect 278590 499576 278596 499588
rect 277636 499548 278596 499576
rect 277636 499536 277642 499548
rect 278590 499536 278596 499548
rect 278648 499536 278654 499588
rect 283006 499576 283012 499588
rect 282967 499548 283012 499576
rect 283006 499536 283012 499548
rect 283064 499536 283070 499588
rect 317322 499536 317328 499588
rect 317380 499576 317386 499588
rect 317874 499576 317880 499588
rect 317380 499548 317880 499576
rect 317380 499536 317386 499548
rect 317874 499536 317880 499548
rect 317932 499536 317938 499588
rect 560938 499536 560944 499588
rect 560996 499576 561002 499588
rect 567194 499576 567200 499588
rect 560996 499548 567200 499576
rect 560996 499536 561002 499548
rect 567194 499536 567200 499548
rect 567252 499536 567258 499588
rect 551462 499468 551468 499520
rect 551520 499508 551526 499520
rect 551830 499508 551836 499520
rect 551520 499480 551836 499508
rect 551520 499468 551526 499480
rect 551830 499468 551836 499480
rect 551888 499468 551894 499520
rect 81342 498788 81348 498840
rect 81400 498828 81406 498840
rect 113174 498828 113180 498840
rect 81400 498800 113180 498828
rect 81400 498788 81406 498800
rect 113174 498788 113180 498800
rect 113232 498788 113238 498840
rect 527818 498788 527824 498840
rect 527876 498828 527882 498840
rect 574094 498828 574100 498840
rect 527876 498800 574100 498828
rect 527876 498788 527882 498800
rect 574094 498788 574100 498800
rect 574152 498788 574158 498840
rect 77018 497428 77024 497480
rect 77076 497468 77082 497480
rect 106274 497468 106280 497480
rect 77076 497440 106280 497468
rect 77076 497428 77082 497440
rect 106274 497428 106280 497440
rect 106332 497428 106338 497480
rect 132494 497428 132500 497480
rect 132552 497468 132558 497480
rect 154850 497468 154856 497480
rect 132552 497440 154856 497468
rect 132552 497428 132558 497440
rect 154850 497428 154856 497440
rect 154908 497428 154914 497480
rect 498378 497428 498384 497480
rect 498436 497468 498442 497480
rect 553302 497468 553308 497480
rect 498436 497440 553308 497468
rect 498436 497428 498442 497440
rect 553302 497428 553308 497440
rect 553360 497428 553366 497480
rect 299382 496068 299388 496120
rect 299440 496108 299446 496120
rect 414014 496108 414020 496120
rect 299440 496080 414020 496108
rect 299440 496068 299446 496080
rect 414014 496068 414020 496080
rect 414072 496068 414078 496120
rect 3510 495456 3516 495508
rect 3568 495496 3574 495508
rect 298094 495496 298100 495508
rect 3568 495468 298100 495496
rect 3568 495456 3574 495468
rect 298094 495456 298100 495468
rect 298152 495496 298158 495508
rect 299382 495496 299388 495508
rect 298152 495468 299388 495496
rect 298152 495456 298158 495468
rect 299382 495456 299388 495468
rect 299440 495456 299446 495508
rect 320450 495456 320456 495508
rect 320508 495496 320514 495508
rect 321094 495496 321100 495508
rect 320508 495468 321100 495496
rect 320508 495456 320514 495468
rect 321094 495456 321100 495468
rect 321152 495456 321158 495508
rect 283006 495388 283012 495440
rect 283064 495428 283070 495440
rect 283190 495428 283196 495440
rect 283064 495400 283196 495428
rect 283064 495388 283070 495400
rect 283190 495388 283196 495400
rect 283248 495388 283254 495440
rect 13078 494708 13084 494760
rect 13136 494748 13142 494760
rect 443638 494748 443644 494760
rect 13136 494720 443644 494748
rect 13136 494708 13142 494720
rect 443638 494708 443644 494720
rect 443696 494708 443702 494760
rect 502426 494708 502432 494760
rect 502484 494748 502490 494760
rect 553210 494748 553216 494760
rect 502484 494720 553216 494748
rect 502484 494708 502490 494720
rect 553210 494708 553216 494720
rect 553268 494708 553274 494760
rect 190914 493960 190920 494012
rect 190972 494000 190978 494012
rect 195330 494000 195336 494012
rect 190972 493972 195336 494000
rect 190972 493960 190978 493972
rect 195330 493960 195336 493972
rect 195388 493960 195394 494012
rect 196894 493960 196900 494012
rect 196952 494000 196958 494012
rect 199470 494000 199476 494012
rect 196952 493972 199476 494000
rect 196952 493960 196958 493972
rect 199470 493960 199476 493972
rect 199528 493960 199534 494012
rect 200482 493960 200488 494012
rect 200540 494000 200546 494012
rect 203702 494000 203708 494012
rect 200540 493972 203708 494000
rect 200540 493960 200546 493972
rect 203702 493960 203708 493972
rect 203760 493960 203766 494012
rect 205266 493960 205272 494012
rect 205324 494000 205330 494012
rect 207750 494000 207756 494012
rect 205324 493972 207756 494000
rect 205324 493960 205330 493972
rect 207750 493960 207756 493972
rect 207808 493960 207814 494012
rect 213638 493960 213644 494012
rect 213696 494000 213702 494012
rect 215294 494000 215300 494012
rect 213696 493972 215300 494000
rect 213696 493960 213702 493972
rect 215294 493960 215300 493972
rect 215352 493960 215358 494012
rect 216030 493960 216036 494012
rect 216088 494000 216094 494012
rect 218146 494000 218152 494012
rect 216088 493972 218152 494000
rect 216088 493960 216094 493972
rect 218146 493960 218152 493972
rect 218204 493960 218210 494012
rect 231578 493960 231584 494012
rect 231636 494000 231642 494012
rect 234522 494000 234528 494012
rect 231636 493972 234528 494000
rect 231636 493960 231642 493972
rect 234522 493960 234528 493972
rect 234580 493960 234586 494012
rect 235166 493960 235172 494012
rect 235224 494000 235230 494012
rect 237558 494000 237564 494012
rect 235224 493972 237564 494000
rect 235224 493960 235230 493972
rect 237558 493960 237564 493972
rect 237616 493960 237622 494012
rect 241146 493960 241152 494012
rect 241204 494000 241210 494012
rect 243078 494000 243084 494012
rect 241204 493972 243084 494000
rect 241204 493960 241210 493972
rect 243078 493960 243084 493972
rect 243136 493960 243142 494012
rect 245930 493960 245936 494012
rect 245988 494000 245994 494012
rect 248414 494000 248420 494012
rect 245988 493972 248420 494000
rect 245988 493960 245994 493972
rect 248414 493960 248420 493972
rect 248472 493960 248478 494012
rect 256786 493960 256792 494012
rect 256844 494000 256850 494012
rect 257890 494000 257896 494012
rect 256844 493972 257896 494000
rect 256844 493960 256850 493972
rect 257890 493960 257896 493972
rect 257948 493960 257954 494012
rect 259454 493960 259460 494012
rect 259512 494000 259518 494012
rect 260282 494000 260288 494012
rect 259512 493972 260288 494000
rect 259512 493960 259518 493972
rect 260282 493960 260288 493972
rect 260340 493960 260346 494012
rect 266354 493960 266360 494012
rect 266412 494000 266418 494012
rect 267458 494000 267464 494012
rect 266412 493972 267464 494000
rect 266412 493960 266418 493972
rect 267458 493960 267464 493972
rect 267516 493960 267522 494012
rect 226794 493892 226800 493944
rect 226852 493932 226858 493944
rect 230382 493932 230388 493944
rect 226852 493904 230388 493932
rect 226852 493892 226858 493904
rect 230382 493892 230388 493904
rect 230440 493892 230446 493944
rect 232774 493892 232780 493944
rect 232832 493932 232838 493944
rect 235902 493932 235908 493944
rect 232832 493904 235908 493932
rect 232832 493892 232838 493904
rect 235902 493892 235908 493904
rect 235960 493892 235966 493944
rect 201678 493824 201684 493876
rect 201736 493864 201742 493876
rect 204622 493864 204628 493876
rect 201736 493836 204628 493864
rect 201736 493824 201742 493836
rect 204622 493824 204628 493836
rect 204680 493824 204686 493876
rect 210050 493824 210056 493876
rect 210108 493864 210114 493876
rect 213454 493864 213460 493876
rect 210108 493836 213460 493864
rect 210108 493824 210114 493836
rect 213454 493824 213460 493836
rect 213512 493824 213518 493876
rect 219618 493824 219624 493876
rect 219676 493864 219682 493876
rect 223482 493864 223488 493876
rect 219676 493836 223488 493864
rect 219676 493824 219682 493836
rect 223482 493824 223488 493836
rect 223540 493824 223546 493876
rect 229186 493824 229192 493876
rect 229244 493864 229250 493876
rect 233142 493864 233148 493876
rect 229244 493836 233148 493864
rect 229244 493824 229250 493836
rect 233142 493824 233148 493836
rect 233200 493824 233206 493876
rect 237558 493824 237564 493876
rect 237616 493864 237622 493876
rect 240134 493864 240140 493876
rect 237616 493836 240140 493864
rect 237616 493824 237622 493836
rect 240134 493824 240140 493836
rect 240192 493824 240198 493876
rect 236362 493756 236368 493808
rect 236420 493796 236426 493808
rect 238754 493796 238760 493808
rect 236420 493768 238760 493796
rect 236420 493756 236426 493768
rect 238754 493756 238760 493768
rect 238812 493756 238818 493808
rect 248322 493756 248328 493808
rect 248380 493796 248386 493808
rect 249794 493796 249800 493808
rect 248380 493768 249800 493796
rect 248380 493756 248386 493768
rect 249794 493756 249800 493768
rect 249852 493756 249858 493808
rect 206462 493688 206468 493740
rect 206520 493728 206526 493740
rect 209130 493728 209136 493740
rect 206520 493700 209136 493728
rect 206520 493688 206526 493700
rect 209130 493688 209136 493700
rect 209188 493688 209194 493740
rect 212442 493688 212448 493740
rect 212500 493728 212506 493740
rect 214926 493728 214932 493740
rect 212500 493700 214932 493728
rect 212500 493688 212506 493700
rect 214926 493688 214932 493700
rect 214984 493688 214990 493740
rect 193306 493620 193312 493672
rect 193364 493660 193370 493672
rect 196066 493660 196072 493672
rect 193364 493632 196072 493660
rect 193364 493620 193370 493632
rect 196066 493620 196072 493632
rect 196124 493620 196130 493672
rect 204070 493620 204076 493672
rect 204128 493660 204134 493672
rect 206370 493660 206376 493672
rect 204128 493632 206376 493660
rect 204128 493620 204134 493632
rect 206370 493620 206376 493632
rect 206428 493620 206434 493672
rect 211246 493620 211252 493672
rect 211304 493660 211310 493672
rect 214650 493660 214656 493672
rect 211304 493632 214656 493660
rect 211304 493620 211310 493632
rect 214650 493620 214656 493632
rect 214708 493620 214714 493672
rect 222010 493620 222016 493672
rect 222068 493660 222074 493672
rect 224218 493660 224224 493672
rect 222068 493632 224224 493660
rect 222068 493620 222074 493632
rect 224218 493620 224224 493632
rect 224276 493620 224282 493672
rect 198090 493552 198096 493604
rect 198148 493592 198154 493604
rect 200206 493592 200212 493604
rect 198148 493564 200212 493592
rect 198148 493552 198154 493564
rect 200206 493552 200212 493564
rect 200264 493552 200270 493604
rect 218422 493552 218428 493604
rect 218480 493592 218486 493604
rect 220814 493592 220820 493604
rect 218480 493564 220820 493592
rect 218480 493552 218486 493564
rect 220814 493552 220820 493564
rect 220872 493552 220878 493604
rect 225598 493552 225604 493604
rect 225656 493592 225662 493604
rect 229002 493592 229008 493604
rect 225656 493564 229008 493592
rect 225656 493552 225662 493564
rect 229002 493552 229008 493564
rect 229060 493552 229066 493604
rect 230382 493552 230388 493604
rect 230440 493592 230446 493604
rect 233050 493592 233056 493604
rect 230440 493564 233056 493592
rect 230440 493552 230446 493564
rect 233050 493552 233056 493564
rect 233108 493552 233114 493604
rect 233970 493552 233976 493604
rect 234028 493592 234034 493604
rect 237282 493592 237288 493604
rect 234028 493564 237288 493592
rect 234028 493552 234034 493564
rect 237282 493552 237288 493564
rect 237340 493552 237346 493604
rect 194502 493484 194508 493536
rect 194560 493524 194566 493536
rect 197170 493524 197176 493536
rect 194560 493496 197176 493524
rect 194560 493484 194566 493496
rect 197170 493484 197176 493496
rect 197228 493484 197234 493536
rect 217226 493484 217232 493536
rect 217284 493524 217290 493536
rect 219526 493524 219532 493536
rect 217284 493496 219532 493524
rect 217284 493484 217290 493496
rect 219526 493484 219532 493496
rect 219584 493484 219590 493536
rect 239950 493484 239956 493536
rect 240008 493524 240014 493536
rect 242802 493524 242808 493536
rect 240008 493496 242808 493524
rect 240008 493484 240014 493496
rect 242802 493484 242808 493496
rect 242860 493484 242866 493536
rect 202874 493416 202880 493468
rect 202932 493456 202938 493468
rect 205634 493456 205640 493468
rect 202932 493428 205640 493456
rect 202932 493416 202938 493428
rect 205634 493416 205640 493428
rect 205692 493416 205698 493468
rect 207658 493416 207664 493468
rect 207716 493456 207722 493468
rect 209866 493456 209872 493468
rect 207716 493428 209872 493456
rect 207716 493416 207722 493428
rect 209866 493416 209872 493428
rect 209924 493416 209930 493468
rect 220814 493416 220820 493468
rect 220872 493456 220878 493468
rect 224862 493456 224868 493468
rect 220872 493428 224868 493456
rect 220872 493416 220878 493428
rect 224862 493416 224868 493428
rect 224920 493416 224926 493468
rect 238754 493416 238760 493468
rect 238812 493456 238818 493468
rect 241514 493456 241520 493468
rect 238812 493428 241520 493456
rect 238812 493416 238818 493428
rect 241514 493416 241520 493428
rect 241572 493416 241578 493468
rect 243538 493416 243544 493468
rect 243596 493456 243602 493468
rect 245654 493456 245660 493468
rect 243596 493428 245660 493456
rect 243596 493416 243602 493428
rect 245654 493416 245660 493428
rect 245712 493416 245718 493468
rect 74534 493348 74540 493400
rect 74592 493388 74598 493400
rect 102134 493388 102140 493400
rect 74592 493360 102140 493388
rect 74592 493348 74598 493360
rect 102134 493348 102140 493360
rect 102192 493348 102198 493400
rect 189718 493348 189724 493400
rect 189776 493388 189782 493400
rect 195238 493388 195244 493400
rect 189776 493360 195244 493388
rect 189776 493348 189782 493360
rect 195238 493348 195244 493360
rect 195296 493348 195302 493400
rect 86954 493280 86960 493332
rect 87012 493320 87018 493332
rect 124214 493320 124220 493332
rect 87012 493292 124220 493320
rect 87012 493280 87018 493292
rect 124214 493280 124220 493292
rect 124272 493280 124278 493332
rect 199286 493280 199292 493332
rect 199344 493320 199350 493332
rect 201586 493320 201592 493332
rect 199344 493292 201592 493320
rect 199344 493280 199350 493292
rect 201586 493280 201592 493292
rect 201644 493280 201650 493332
rect 244734 493280 244740 493332
rect 244792 493320 244798 493332
rect 247218 493320 247224 493332
rect 244792 493292 247224 493320
rect 244792 493280 244798 493292
rect 247218 493280 247224 493292
rect 247276 493280 247282 493332
rect 249518 493280 249524 493332
rect 249576 493320 249582 493332
rect 251266 493320 251272 493332
rect 249576 493292 251272 493320
rect 249576 493280 249582 493292
rect 251266 493280 251272 493292
rect 251324 493280 251330 493332
rect 509234 493280 509240 493332
rect 509292 493320 509298 493332
rect 553118 493320 553124 493332
rect 509292 493292 553124 493320
rect 509292 493280 509298 493292
rect 553118 493280 553124 493292
rect 553176 493280 553182 493332
rect 214834 493212 214840 493264
rect 214892 493252 214898 493264
rect 216674 493252 216680 493264
rect 214892 493224 216680 493252
rect 214892 493212 214898 493224
rect 216674 493212 216680 493224
rect 216732 493212 216738 493264
rect 242342 493212 242348 493264
rect 242400 493252 242406 493264
rect 244274 493252 244280 493264
rect 242400 493224 244280 493252
rect 242400 493212 242406 493224
rect 244274 493212 244280 493224
rect 244332 493212 244338 493264
rect 195698 493144 195704 493196
rect 195756 493184 195762 493196
rect 201862 493184 201868 493196
rect 195756 493156 201868 493184
rect 195756 493144 195762 493156
rect 201862 493144 201868 493156
rect 201920 493144 201926 493196
rect 208854 493144 208860 493196
rect 208912 493184 208918 493196
rect 211338 493184 211344 493196
rect 208912 493156 211344 493184
rect 208912 493144 208918 493156
rect 211338 493144 211344 493156
rect 211396 493144 211402 493196
rect 256694 493144 256700 493196
rect 256752 493184 256758 493196
rect 257982 493184 257988 493196
rect 256752 493156 257988 493184
rect 256752 493144 256758 493156
rect 257982 493144 257988 493156
rect 258040 493144 258046 493196
rect 277578 493144 277584 493196
rect 277636 493184 277642 493196
rect 279418 493184 279424 493196
rect 277636 493156 279424 493184
rect 277636 493144 277642 493156
rect 279418 493144 279424 493156
rect 279476 493144 279482 493196
rect 188614 493008 188620 493060
rect 188672 493048 188678 493060
rect 191926 493048 191932 493060
rect 188672 493020 191932 493048
rect 188672 493008 188678 493020
rect 191926 493008 191932 493020
rect 191984 493008 191990 493060
rect 227990 493008 227996 493060
rect 228048 493048 228054 493060
rect 230566 493048 230572 493060
rect 228048 493020 230572 493048
rect 228048 493008 228054 493020
rect 230566 493008 230572 493020
rect 230624 493008 230630 493060
rect 250714 492940 250720 492992
rect 250772 492980 250778 492992
rect 252738 492980 252744 492992
rect 250772 492952 252744 492980
rect 250772 492940 250778 492952
rect 252738 492940 252744 492952
rect 252796 492940 252802 492992
rect 223206 492872 223212 492924
rect 223264 492912 223270 492924
rect 227898 492912 227904 492924
rect 223264 492884 227904 492912
rect 223264 492872 223270 492884
rect 227898 492872 227904 492884
rect 227956 492872 227962 492924
rect 271966 492804 271972 492856
rect 272024 492844 272030 492856
rect 273438 492844 273444 492856
rect 272024 492816 273444 492844
rect 272024 492804 272030 492816
rect 273438 492804 273444 492816
rect 273496 492804 273502 492856
rect 223574 492736 223580 492788
rect 223632 492776 223638 492788
rect 224402 492776 224408 492788
rect 223632 492748 224408 492776
rect 223632 492736 223638 492748
rect 224402 492736 224408 492748
rect 224460 492736 224466 492788
rect 282914 492600 282920 492652
rect 282972 492640 282978 492652
rect 283190 492640 283196 492652
rect 282972 492612 283196 492640
rect 282972 492600 282978 492612
rect 283190 492600 283196 492612
rect 283248 492600 283254 492652
rect 320266 492600 320272 492652
rect 320324 492640 320330 492652
rect 320726 492640 320732 492652
rect 320324 492612 320732 492640
rect 320324 492600 320330 492612
rect 320726 492600 320732 492612
rect 320784 492600 320790 492652
rect 73062 491988 73068 492040
rect 73120 492028 73126 492040
rect 99006 492028 99012 492040
rect 73120 492000 99012 492028
rect 73120 491988 73126 492000
rect 99006 491988 99012 492000
rect 99064 491988 99070 492040
rect 84102 491920 84108 491972
rect 84160 491960 84166 491972
rect 117130 491960 117136 491972
rect 84160 491932 117136 491960
rect 84160 491920 84166 491932
rect 117130 491920 117136 491932
rect 117188 491920 117194 491972
rect 495342 491920 495348 491972
rect 495400 491960 495406 491972
rect 555694 491960 555700 491972
rect 495400 491932 555700 491960
rect 495400 491920 495406 491932
rect 555694 491920 555700 491932
rect 555752 491920 555758 491972
rect 94498 491240 94504 491292
rect 94556 491280 94562 491292
rect 95694 491280 95700 491292
rect 94556 491252 95700 491280
rect 94556 491240 94562 491252
rect 95694 491240 95700 491252
rect 95752 491240 95758 491292
rect 68922 490628 68928 490680
rect 68980 490668 68986 490680
rect 92106 490668 92112 490680
rect 68980 490640 92112 490668
rect 68980 490628 68986 490640
rect 92106 490628 92112 490640
rect 92164 490628 92170 490680
rect 79962 490560 79968 490612
rect 80020 490600 80026 490612
rect 109954 490600 109960 490612
rect 80020 490572 109960 490600
rect 80020 490560 80026 490572
rect 109954 490560 109960 490572
rect 110012 490560 110018 490612
rect 112438 490560 112444 490612
rect 112496 490600 112502 490612
rect 120718 490600 120724 490612
rect 112496 490572 120724 490600
rect 112496 490560 112502 490572
rect 120718 490560 120724 490572
rect 120776 490560 120782 490612
rect 499482 490560 499488 490612
rect 499540 490600 499546 490612
rect 555970 490600 555976 490612
rect 499540 490572 555976 490600
rect 499540 490560 499546 490572
rect 555970 490560 555976 490572
rect 556028 490560 556034 490612
rect 551462 489880 551468 489932
rect 551520 489920 551526 489932
rect 551830 489920 551836 489932
rect 551520 489892 551836 489920
rect 551520 489880 551526 489892
rect 551830 489880 551836 489892
rect 551888 489880 551894 489932
rect 35802 489812 35808 489864
rect 35860 489852 35866 489864
rect 36538 489852 36544 489864
rect 35860 489824 36544 489852
rect 35860 489812 35866 489824
rect 36538 489812 36544 489824
rect 36596 489812 36602 489864
rect 61930 489812 61936 489864
rect 61988 489852 61994 489864
rect 79502 489852 79508 489864
rect 61988 489824 79508 489852
rect 61988 489812 61994 489824
rect 79502 489812 79508 489824
rect 79560 489812 79566 489864
rect 95142 489812 95148 489864
rect 95200 489852 95206 489864
rect 135070 489852 135076 489864
rect 95200 489824 135076 489852
rect 95200 489812 95206 489824
rect 135070 489812 135076 489824
rect 135128 489812 135134 489864
rect 62022 489744 62028 489796
rect 62080 489784 62086 489796
rect 81342 489784 81348 489796
rect 62080 489756 81348 489784
rect 62080 489744 62086 489756
rect 81342 489744 81348 489756
rect 81400 489744 81406 489796
rect 90910 489744 90916 489796
rect 90968 489784 90974 489796
rect 129734 489784 129740 489796
rect 90968 489756 129740 489784
rect 90968 489744 90974 489756
rect 129734 489744 129740 489756
rect 129792 489744 129798 489796
rect 64782 489676 64788 489728
rect 64840 489716 64846 489728
rect 84930 489716 84936 489728
rect 64840 489688 84936 489716
rect 64840 489676 64846 489688
rect 84930 489676 84936 489688
rect 84988 489676 84994 489728
rect 96522 489676 96528 489728
rect 96580 489716 96586 489728
rect 136910 489716 136916 489728
rect 96580 489688 136916 489716
rect 96580 489676 96586 489688
rect 136910 489676 136916 489688
rect 136968 489676 136974 489728
rect 49602 489608 49608 489660
rect 49660 489648 49666 489660
rect 59814 489648 59820 489660
rect 49660 489620 59820 489648
rect 49660 489608 49666 489620
rect 59814 489608 59820 489620
rect 59872 489608 59878 489660
rect 63402 489608 63408 489660
rect 63460 489648 63466 489660
rect 83090 489648 83096 489660
rect 63460 489620 83096 489648
rect 63460 489608 63466 489620
rect 83090 489608 83096 489620
rect 83148 489608 83154 489660
rect 97902 489608 97908 489660
rect 97960 489648 97966 489660
rect 140498 489648 140504 489660
rect 97960 489620 140504 489648
rect 97960 489608 97966 489620
rect 140498 489608 140504 489620
rect 140556 489608 140562 489660
rect 50982 489540 50988 489592
rect 51040 489580 51046 489592
rect 61654 489580 61660 489592
rect 51040 489552 61660 489580
rect 51040 489540 51046 489552
rect 61654 489540 61660 489552
rect 61712 489540 61718 489592
rect 66162 489540 66168 489592
rect 66220 489580 66226 489592
rect 86678 489580 86684 489592
rect 66220 489552 86684 489580
rect 66220 489540 66226 489552
rect 86678 489540 86684 489552
rect 86736 489540 86742 489592
rect 96430 489540 96436 489592
rect 96488 489580 96494 489592
rect 138658 489580 138664 489592
rect 96488 489552 138664 489580
rect 96488 489540 96494 489552
rect 138658 489540 138664 489552
rect 138716 489540 138722 489592
rect 52362 489472 52368 489524
rect 52420 489512 52426 489524
rect 63402 489512 63408 489524
rect 52420 489484 63408 489512
rect 52420 489472 52426 489484
rect 63402 489472 63408 489484
rect 63460 489472 63466 489524
rect 67542 489472 67548 489524
rect 67600 489512 67606 489524
rect 88518 489512 88524 489524
rect 67600 489484 88524 489512
rect 67600 489472 67606 489484
rect 88518 489472 88524 489484
rect 88576 489472 88582 489524
rect 102042 489472 102048 489524
rect 102100 489512 102106 489524
rect 145834 489512 145840 489524
rect 102100 489484 145840 489512
rect 102100 489472 102106 489484
rect 145834 489472 145840 489484
rect 145892 489472 145898 489524
rect 53742 489404 53748 489456
rect 53800 489444 53806 489456
rect 66990 489444 66996 489456
rect 53800 489416 66996 489444
rect 53800 489404 53806 489416
rect 66990 489404 66996 489416
rect 67048 489404 67054 489456
rect 67450 489404 67456 489456
rect 67508 489444 67514 489456
rect 90266 489444 90272 489456
rect 67508 489416 90272 489444
rect 67508 489404 67514 489416
rect 90266 489404 90272 489416
rect 90324 489404 90330 489456
rect 100662 489404 100668 489456
rect 100720 489444 100726 489456
rect 144086 489444 144092 489456
rect 100720 489416 144092 489444
rect 100720 489404 100726 489416
rect 144086 489404 144092 489416
rect 144144 489404 144150 489456
rect 52270 489336 52276 489388
rect 52328 489376 52334 489388
rect 65150 489376 65156 489388
rect 52328 489348 65156 489376
rect 52328 489336 52334 489348
rect 65150 489336 65156 489348
rect 65208 489336 65214 489388
rect 70302 489336 70308 489388
rect 70360 489376 70366 489388
rect 93854 489376 93860 489388
rect 70360 489348 93860 489376
rect 70360 489336 70366 489348
rect 93854 489336 93860 489348
rect 93912 489336 93918 489388
rect 99282 489336 99288 489388
rect 99340 489376 99346 489388
rect 142246 489376 142252 489388
rect 99340 489348 142252 489376
rect 99340 489336 99346 489348
rect 142246 489336 142252 489348
rect 142304 489336 142310 489388
rect 56410 489268 56416 489320
rect 56468 489308 56474 489320
rect 70578 489308 70584 489320
rect 56468 489280 70584 489308
rect 56468 489268 56474 489280
rect 70578 489268 70584 489280
rect 70636 489268 70642 489320
rect 71682 489268 71688 489320
rect 71740 489308 71746 489320
rect 97442 489308 97448 489320
rect 71740 489280 97448 489308
rect 71740 489268 71746 489280
rect 97442 489268 97448 489280
rect 97500 489268 97506 489320
rect 103422 489268 103428 489320
rect 103480 489308 103486 489320
rect 149422 489308 149428 489320
rect 103480 489280 149428 489308
rect 103480 489268 103486 489280
rect 149422 489268 149428 489280
rect 149480 489268 149486 489320
rect 37090 489200 37096 489252
rect 37148 489240 37154 489252
rect 38286 489240 38292 489252
rect 37148 489212 38292 489240
rect 37148 489200 37154 489212
rect 38286 489200 38292 489212
rect 38344 489200 38350 489252
rect 48222 489200 48228 489252
rect 48280 489240 48286 489252
rect 58066 489240 58072 489252
rect 48280 489212 58072 489240
rect 48280 489200 48286 489212
rect 58066 489200 58072 489212
rect 58124 489200 58130 489252
rect 59262 489200 59268 489252
rect 59320 489240 59326 489252
rect 75914 489240 75920 489252
rect 59320 489212 75920 489240
rect 59320 489200 59326 489212
rect 75914 489200 75920 489212
rect 75972 489200 75978 489252
rect 77202 489200 77208 489252
rect 77260 489240 77266 489252
rect 104618 489240 104624 489252
rect 77260 489212 104624 489240
rect 77260 489200 77266 489212
rect 104618 489200 104624 489212
rect 104676 489200 104682 489252
rect 104802 489200 104808 489252
rect 104860 489240 104866 489252
rect 151262 489240 151268 489252
rect 104860 489212 151268 489240
rect 104860 489200 104866 489212
rect 151262 489200 151268 489212
rect 151320 489200 151326 489252
rect 37182 489132 37188 489184
rect 37240 489172 37246 489184
rect 40126 489172 40132 489184
rect 37240 489144 40132 489172
rect 37240 489132 37246 489144
rect 40126 489132 40132 489144
rect 40184 489132 40190 489184
rect 46842 489132 46848 489184
rect 46900 489172 46906 489184
rect 56226 489172 56232 489184
rect 46900 489144 56232 489172
rect 46900 489132 46906 489144
rect 56226 489132 56232 489144
rect 56284 489132 56290 489184
rect 56502 489132 56508 489184
rect 56560 489172 56566 489184
rect 72326 489172 72332 489184
rect 56560 489144 72332 489172
rect 56560 489132 56566 489144
rect 72326 489132 72332 489144
rect 72384 489132 72390 489184
rect 74442 489132 74448 489184
rect 74500 489172 74506 489184
rect 101030 489172 101036 489184
rect 74500 489144 101036 489172
rect 74500 489132 74506 489144
rect 101030 489132 101036 489144
rect 101088 489132 101094 489184
rect 101950 489132 101956 489184
rect 102008 489172 102014 489184
rect 147674 489172 147680 489184
rect 102008 489144 147680 489172
rect 102008 489132 102014 489144
rect 147674 489132 147680 489144
rect 147732 489132 147738 489184
rect 60642 489064 60648 489116
rect 60700 489104 60706 489116
rect 77754 489104 77760 489116
rect 60700 489076 77760 489104
rect 60700 489064 60706 489076
rect 77754 489064 77760 489076
rect 77812 489064 77818 489116
rect 93762 489064 93768 489116
rect 93820 489104 93826 489116
rect 133322 489104 133328 489116
rect 93820 489076 133328 489104
rect 93820 489064 93826 489076
rect 133322 489064 133328 489076
rect 133380 489064 133386 489116
rect 57882 488996 57888 489048
rect 57940 489036 57946 489048
rect 74166 489036 74172 489048
rect 57940 489008 74172 489036
rect 57940 488996 57946 489008
rect 74166 488996 74172 489008
rect 74224 488996 74230 489048
rect 92382 488996 92388 489048
rect 92440 489036 92446 489048
rect 131482 489036 131488 489048
rect 92440 489008 131488 489036
rect 92440 488996 92446 489008
rect 131482 488996 131488 489008
rect 131540 488996 131546 489048
rect 55122 488928 55128 488980
rect 55180 488968 55186 488980
rect 68738 488968 68744 488980
rect 55180 488940 68744 488968
rect 55180 488928 55186 488940
rect 68738 488928 68744 488940
rect 68796 488928 68802 488980
rect 89622 488928 89628 488980
rect 89680 488968 89686 488980
rect 126146 488968 126152 488980
rect 89680 488940 126152 488968
rect 89680 488928 89686 488940
rect 126146 488928 126152 488940
rect 126204 488928 126210 488980
rect 91002 488860 91008 488912
rect 91060 488900 91066 488912
rect 127894 488900 127900 488912
rect 91060 488872 127900 488900
rect 91060 488860 91066 488872
rect 127894 488860 127900 488872
rect 127952 488860 127958 488912
rect 86862 488792 86868 488844
rect 86920 488832 86926 488844
rect 122558 488832 122564 488844
rect 86920 488804 122564 488832
rect 86920 488792 86926 488804
rect 122558 488792 122564 488804
rect 122616 488792 122622 488844
rect 20346 488724 20352 488776
rect 20404 488764 20410 488776
rect 24210 488764 24216 488776
rect 20404 488736 24216 488764
rect 20404 488724 20410 488736
rect 24210 488724 24216 488736
rect 24268 488724 24274 488776
rect 39942 488724 39948 488776
rect 40000 488764 40006 488776
rect 43714 488764 43720 488776
rect 40000 488736 43720 488764
rect 40000 488724 40006 488736
rect 43714 488724 43720 488736
rect 43772 488724 43778 488776
rect 85482 488724 85488 488776
rect 85540 488764 85546 488776
rect 118970 488764 118976 488776
rect 85540 488736 118976 488764
rect 85540 488724 85546 488736
rect 118970 488724 118976 488736
rect 119028 488724 119034 488776
rect 16850 488656 16856 488708
rect 16908 488696 16914 488708
rect 22278 488696 22284 488708
rect 16908 488668 22284 488696
rect 16908 488656 16914 488668
rect 22278 488656 22284 488668
rect 22336 488656 22342 488708
rect 38562 488656 38568 488708
rect 38620 488696 38626 488708
rect 41874 488696 41880 488708
rect 38620 488668 41880 488696
rect 38620 488656 38626 488668
rect 41874 488656 41880 488668
rect 41932 488656 41938 488708
rect 82722 488656 82728 488708
rect 82780 488696 82786 488708
rect 115382 488696 115388 488708
rect 82780 488668 115388 488696
rect 82780 488656 82786 488668
rect 115382 488656 115388 488668
rect 115440 488656 115446 488708
rect 22186 488588 22192 488640
rect 22244 488628 22250 488640
rect 24302 488628 24308 488640
rect 22244 488600 24308 488628
rect 22244 488588 22250 488600
rect 24302 488588 24308 488600
rect 24360 488588 24366 488640
rect 48958 488588 48964 488640
rect 49016 488628 49022 488640
rect 50890 488628 50896 488640
rect 49016 488600 50896 488628
rect 49016 488588 49022 488600
rect 50890 488588 50896 488600
rect 50948 488588 50954 488640
rect 81250 488588 81256 488640
rect 81308 488628 81314 488640
rect 111794 488628 111800 488640
rect 81308 488600 111800 488628
rect 81308 488588 81314 488600
rect 111794 488588 111800 488600
rect 111852 488588 111858 488640
rect 18598 488520 18604 488572
rect 18656 488560 18662 488572
rect 23474 488560 23480 488572
rect 18656 488532 23480 488560
rect 18656 488520 18662 488532
rect 23474 488520 23480 488532
rect 23532 488520 23538 488572
rect 23934 488520 23940 488572
rect 23992 488560 23998 488572
rect 25498 488560 25504 488572
rect 23992 488532 25504 488560
rect 23992 488520 23998 488532
rect 25498 488520 25504 488532
rect 25556 488520 25562 488572
rect 29362 488520 29368 488572
rect 29420 488560 29426 488572
rect 30282 488560 30288 488572
rect 29420 488532 30288 488560
rect 29420 488520 29426 488532
rect 30282 488520 30288 488532
rect 30340 488520 30346 488572
rect 41322 488520 41328 488572
rect 41380 488560 41386 488572
rect 45462 488560 45468 488572
rect 41380 488532 45468 488560
rect 41380 488520 41386 488532
rect 45462 488520 45468 488532
rect 45520 488520 45526 488572
rect 47578 488520 47584 488572
rect 47636 488560 47642 488572
rect 49050 488560 49056 488572
rect 47636 488532 49056 488560
rect 47636 488520 47642 488532
rect 49050 488520 49056 488532
rect 49108 488520 49114 488572
rect 78582 488520 78588 488572
rect 78640 488560 78646 488572
rect 108206 488560 108212 488572
rect 78640 488532 108212 488560
rect 78640 488520 78646 488532
rect 108206 488520 108212 488532
rect 108264 488520 108270 488572
rect 24118 486412 24124 486464
rect 24176 486452 24182 486464
rect 156046 486452 156052 486464
rect 24176 486424 156052 486452
rect 24176 486412 24182 486424
rect 156046 486412 156052 486424
rect 156104 486412 156110 486464
rect 505002 486412 505008 486464
rect 505060 486452 505066 486464
rect 555234 486452 555240 486464
rect 505060 486424 555240 486452
rect 505060 486412 505066 486424
rect 555234 486412 555240 486424
rect 555292 486412 555298 486464
rect 3418 485052 3424 485104
rect 3476 485092 3482 485104
rect 185578 485092 185584 485104
rect 3476 485064 185584 485092
rect 3476 485052 3482 485064
rect 185578 485052 185584 485064
rect 185636 485052 185642 485104
rect 521562 483692 521568 483744
rect 521620 483732 521626 483744
rect 552658 483732 552664 483744
rect 521620 483704 552664 483732
rect 521620 483692 521626 483704
rect 552658 483692 552664 483704
rect 552716 483692 552722 483744
rect 511902 483624 511908 483676
rect 511960 483664 511966 483676
rect 555142 483664 555148 483676
rect 511960 483636 555148 483664
rect 511960 483624 511966 483636
rect 555142 483624 555148 483636
rect 555200 483624 555206 483676
rect 528370 482264 528376 482316
rect 528428 482304 528434 482316
rect 552382 482304 552388 482316
rect 528428 482276 552388 482304
rect 528428 482264 528434 482276
rect 552382 482264 552388 482276
rect 552440 482264 552446 482316
rect 529842 481040 529848 481092
rect 529900 481080 529906 481092
rect 555786 481080 555792 481092
rect 529900 481052 555792 481080
rect 529900 481040 529906 481052
rect 555786 481040 555792 481052
rect 555844 481040 555850 481092
rect 520182 480972 520188 481024
rect 520240 481012 520246 481024
rect 554590 481012 554596 481024
rect 520240 480984 554596 481012
rect 520240 480972 520246 480984
rect 554590 480972 554596 480984
rect 554648 480972 554654 481024
rect 517422 480904 517428 480956
rect 517480 480944 517486 480956
rect 517480 480916 548380 480944
rect 517480 480904 517486 480916
rect 548352 480808 548380 480916
rect 551002 480904 551008 480956
rect 551060 480944 551066 480956
rect 551462 480944 551468 480956
rect 551060 480916 551468 480944
rect 551060 480904 551066 480916
rect 551462 480904 551468 480916
rect 551520 480904 551526 480956
rect 553026 480808 553032 480820
rect 548352 480780 553032 480808
rect 553026 480768 553032 480780
rect 553084 480768 553090 480820
rect 3142 480224 3148 480276
rect 3200 480264 3206 480276
rect 14458 480264 14464 480276
rect 3200 480236 14464 480264
rect 3200 480224 3206 480236
rect 14458 480224 14464 480236
rect 14516 480224 14522 480276
rect 183646 480224 183652 480276
rect 183704 480264 183710 480276
rect 183830 480264 183836 480276
rect 183704 480236 183836 480264
rect 183704 480224 183710 480236
rect 183830 480224 183836 480236
rect 183888 480224 183894 480276
rect 525702 479612 525708 479664
rect 525760 479652 525766 479664
rect 552474 479652 552480 479664
rect 525760 479624 552480 479652
rect 525760 479612 525766 479624
rect 552474 479612 552480 479624
rect 552532 479612 552538 479664
rect 527082 479544 527088 479596
rect 527140 479584 527146 479596
rect 554498 479584 554504 479596
rect 527140 479556 554504 479584
rect 527140 479544 527146 479556
rect 554498 479544 554504 479556
rect 554556 479544 554562 479596
rect 494698 479476 494704 479528
rect 494756 479516 494762 479528
rect 554774 479516 554780 479528
rect 494756 479488 554780 479516
rect 494756 479476 494762 479488
rect 554774 479476 554780 479488
rect 554832 479476 554838 479528
rect 542262 478388 542268 478440
rect 542320 478428 542326 478440
rect 553670 478428 553676 478440
rect 542320 478400 553676 478428
rect 542320 478388 542326 478400
rect 553670 478388 553676 478400
rect 553728 478388 553734 478440
rect 540882 478320 540888 478372
rect 540940 478360 540946 478372
rect 555602 478360 555608 478372
rect 540940 478332 555608 478360
rect 540940 478320 540946 478332
rect 555602 478320 555608 478332
rect 555660 478320 555666 478372
rect 532602 478252 532608 478304
rect 532660 478292 532666 478304
rect 552842 478292 552848 478304
rect 532660 478264 552848 478292
rect 532660 478252 532666 478264
rect 552842 478252 552848 478264
rect 552900 478252 552906 478304
rect 522942 478184 522948 478236
rect 523000 478224 523006 478236
rect 551186 478224 551192 478236
rect 523000 478196 551192 478224
rect 523000 478184 523006 478196
rect 551186 478184 551192 478196
rect 551244 478184 551250 478236
rect 496722 478116 496728 478168
rect 496780 478156 496786 478168
rect 555878 478156 555884 478168
rect 496780 478128 555884 478156
rect 496780 478116 496786 478128
rect 555878 478116 555884 478128
rect 555936 478116 555942 478168
rect 344922 477436 344928 477488
rect 344980 477476 344986 477488
rect 346026 477476 346032 477488
rect 344980 477448 346032 477476
rect 344980 477436 344986 477448
rect 346026 477436 346032 477448
rect 346084 477436 346090 477488
rect 353202 477436 353208 477488
rect 353260 477476 353266 477488
rect 355778 477476 355784 477488
rect 353260 477448 355784 477476
rect 353260 477436 353266 477448
rect 355778 477436 355784 477448
rect 355836 477436 355842 477488
rect 369762 477436 369768 477488
rect 369820 477476 369826 477488
rect 374086 477476 374092 477488
rect 369820 477448 374092 477476
rect 369820 477436 369826 477448
rect 374086 477436 374092 477448
rect 374144 477436 374150 477488
rect 354582 477368 354588 477420
rect 354640 477408 354646 477420
rect 356974 477408 356980 477420
rect 354640 477380 356980 477408
rect 354640 477368 354646 477380
rect 356974 477368 356980 477380
rect 357032 477368 357038 477420
rect 378042 477368 378048 477420
rect 378100 477408 378106 477420
rect 383838 477408 383844 477420
rect 378100 477380 383844 477408
rect 378100 477368 378106 477380
rect 383838 477368 383844 477380
rect 383896 477368 383902 477420
rect 390462 477300 390468 477352
rect 390520 477340 390526 477352
rect 397270 477340 397276 477352
rect 390520 477312 397276 477340
rect 390520 477300 390526 477312
rect 397270 477300 397276 477312
rect 397328 477300 397334 477352
rect 395982 477232 395988 477284
rect 396040 477272 396046 477284
rect 403434 477272 403440 477284
rect 396040 477244 403440 477272
rect 396040 477232 396046 477244
rect 403434 477232 403440 477244
rect 403492 477232 403498 477284
rect 362862 477164 362868 477216
rect 362920 477204 362926 477216
rect 366726 477204 366732 477216
rect 362920 477176 366732 477204
rect 362920 477164 362926 477176
rect 366726 477164 366732 477176
rect 366784 477164 366790 477216
rect 383562 477164 383568 477216
rect 383620 477204 383626 477216
rect 390002 477204 390008 477216
rect 383620 477176 390008 477204
rect 383620 477164 383626 477176
rect 390002 477164 390008 477176
rect 390060 477164 390066 477216
rect 391842 477164 391848 477216
rect 391900 477204 391906 477216
rect 399754 477204 399760 477216
rect 391900 477176 399760 477204
rect 391900 477164 391906 477176
rect 399754 477164 399760 477176
rect 399812 477164 399818 477216
rect 400122 477164 400128 477216
rect 400180 477204 400186 477216
rect 408310 477204 408316 477216
rect 400180 477176 408316 477204
rect 400180 477164 400186 477176
rect 408310 477164 408316 477176
rect 408368 477164 408374 477216
rect 375282 477096 375288 477148
rect 375340 477136 375346 477148
rect 380158 477136 380164 477148
rect 375340 477108 380164 477136
rect 375340 477096 375346 477108
rect 380158 477096 380164 477108
rect 380216 477096 380222 477148
rect 386322 477028 386328 477080
rect 386380 477068 386386 477080
rect 392394 477068 392400 477080
rect 386380 477040 392400 477068
rect 386380 477028 386386 477040
rect 392394 477028 392400 477040
rect 392452 477028 392458 477080
rect 393222 477028 393228 477080
rect 393280 477068 393286 477080
rect 400950 477068 400956 477080
rect 393280 477040 400956 477068
rect 393280 477028 393286 477040
rect 400950 477028 400956 477040
rect 401008 477028 401014 477080
rect 401410 477028 401416 477080
rect 401468 477068 401474 477080
rect 409506 477068 409512 477080
rect 401468 477040 409512 477068
rect 401468 477028 401474 477040
rect 409506 477028 409512 477040
rect 409564 477028 409570 477080
rect 546402 477028 546408 477080
rect 546460 477068 546466 477080
rect 553578 477068 553584 477080
rect 546460 477040 553584 477068
rect 546460 477028 546466 477040
rect 553578 477028 553584 477040
rect 553636 477028 553642 477080
rect 317874 476960 317880 477012
rect 317932 477000 317938 477012
rect 318702 477000 318708 477012
rect 317932 476972 318708 477000
rect 317932 476960 317938 476972
rect 318702 476960 318708 476972
rect 318760 476960 318766 477012
rect 319070 476960 319076 477012
rect 319128 477000 319134 477012
rect 320082 477000 320088 477012
rect 319128 476972 320088 477000
rect 319128 476960 319134 476972
rect 320082 476960 320088 476972
rect 320140 476960 320146 477012
rect 364242 476960 364248 477012
rect 364300 477000 364306 477012
rect 368014 477000 368020 477012
rect 364300 476972 368020 477000
rect 364300 476960 364306 476972
rect 368014 476960 368020 476972
rect 368072 476960 368078 477012
rect 371142 476960 371148 477012
rect 371200 477000 371206 477012
rect 375282 477000 375288 477012
rect 371200 476972 375288 477000
rect 371200 476960 371206 476972
rect 375282 476960 375288 476972
rect 375340 476960 375346 477012
rect 376570 476960 376576 477012
rect 376628 477000 376634 477012
rect 381446 477000 381452 477012
rect 376628 476972 381452 477000
rect 376628 476960 376634 476972
rect 381446 476960 381452 476972
rect 381504 476960 381510 477012
rect 382182 476960 382188 477012
rect 382240 477000 382246 477012
rect 388714 477000 388720 477012
rect 382240 476972 388720 477000
rect 382240 476960 382246 476972
rect 388714 476960 388720 476972
rect 388772 476960 388778 477012
rect 389082 476960 389088 477012
rect 389140 477000 389146 477012
rect 396074 477000 396080 477012
rect 389140 476972 396080 477000
rect 389140 476960 389146 476972
rect 396074 476960 396080 476972
rect 396132 476960 396138 477012
rect 397362 476960 397368 477012
rect 397420 477000 397426 477012
rect 405826 477000 405832 477012
rect 397420 476972 405832 477000
rect 397420 476960 397426 476972
rect 405826 476960 405832 476972
rect 405884 476960 405890 477012
rect 536742 476960 536748 477012
rect 536800 477000 536806 477012
rect 552566 477000 552572 477012
rect 536800 476972 552572 477000
rect 536800 476960 536806 476972
rect 552566 476960 552572 476972
rect 552624 476960 552630 477012
rect 351822 476892 351828 476944
rect 351880 476932 351886 476944
rect 353294 476932 353300 476944
rect 351880 476904 353300 476932
rect 351880 476892 351886 476904
rect 353294 476892 353300 476904
rect 353352 476892 353358 476944
rect 355870 476892 355876 476944
rect 355928 476932 355934 476944
rect 359458 476932 359464 476944
rect 355928 476904 359464 476932
rect 355928 476892 355934 476904
rect 359458 476892 359464 476904
rect 359516 476892 359522 476944
rect 361390 476892 361396 476944
rect 361448 476932 361454 476944
rect 365530 476932 365536 476944
rect 361448 476904 365536 476932
rect 361448 476892 361454 476904
rect 365530 476892 365536 476904
rect 365588 476892 365594 476944
rect 372522 476892 372528 476944
rect 372580 476932 372586 476944
rect 377766 476932 377772 476944
rect 372580 476904 377772 476932
rect 372580 476892 372586 476904
rect 377766 476892 377772 476904
rect 377824 476892 377830 476944
rect 380802 476892 380808 476944
rect 380860 476932 380866 476944
rect 386322 476932 386328 476944
rect 380860 476904 386328 476932
rect 380860 476892 380866 476904
rect 386322 476892 386328 476904
rect 386380 476892 386386 476944
rect 398742 476892 398748 476944
rect 398800 476932 398806 476944
rect 407114 476932 407120 476944
rect 398800 476904 407120 476932
rect 398800 476892 398806 476904
rect 407114 476892 407120 476904
rect 407172 476892 407178 476944
rect 535362 476892 535368 476944
rect 535420 476932 535426 476944
rect 554314 476932 554320 476944
rect 535420 476904 554320 476932
rect 535420 476892 535426 476904
rect 554314 476892 554320 476904
rect 554372 476892 554378 476944
rect 332594 476824 332600 476876
rect 332652 476864 332658 476876
rect 333790 476864 333796 476876
rect 332652 476836 333796 476864
rect 332652 476824 332658 476836
rect 333790 476824 333796 476836
rect 333848 476824 333854 476876
rect 335354 476824 335360 476876
rect 335412 476864 335418 476876
rect 336182 476864 336188 476876
rect 335412 476836 336188 476864
rect 335412 476824 335418 476836
rect 336182 476824 336188 476836
rect 336240 476824 336246 476876
rect 336642 476824 336648 476876
rect 336700 476864 336706 476876
rect 337470 476864 337476 476876
rect 336700 476836 337476 476864
rect 336700 476824 336706 476836
rect 337470 476824 337476 476836
rect 337528 476824 337534 476876
rect 342162 476824 342168 476876
rect 342220 476864 342226 476876
rect 343542 476864 343548 476876
rect 342220 476836 343548 476864
rect 342220 476824 342226 476836
rect 343542 476824 343548 476836
rect 343600 476824 343606 476876
rect 346210 476824 346216 476876
rect 346268 476864 346274 476876
rect 347222 476864 347228 476876
rect 346268 476836 347228 476864
rect 346268 476824 346274 476836
rect 347222 476824 347228 476836
rect 347280 476824 347286 476876
rect 350442 476824 350448 476876
rect 350500 476864 350506 476876
rect 352098 476864 352104 476876
rect 350500 476836 352104 476864
rect 350500 476824 350506 476836
rect 352098 476824 352104 476836
rect 352156 476824 352162 476876
rect 355962 476824 355968 476876
rect 356020 476864 356026 476876
rect 358170 476864 358176 476876
rect 356020 476836 358176 476864
rect 356020 476824 356026 476836
rect 358170 476824 358176 476836
rect 358228 476824 358234 476876
rect 358722 476824 358728 476876
rect 358780 476864 358786 476876
rect 361850 476864 361856 476876
rect 358780 476836 361856 476864
rect 358780 476824 358786 476836
rect 361850 476824 361856 476836
rect 361908 476824 361914 476876
rect 365622 476824 365628 476876
rect 365680 476864 365686 476876
rect 369210 476864 369216 476876
rect 365680 476836 369216 476864
rect 365680 476824 365686 476836
rect 369210 476824 369216 476836
rect 369268 476824 369274 476876
rect 373902 476824 373908 476876
rect 373960 476864 373966 476876
rect 378962 476864 378968 476876
rect 373960 476836 378968 476864
rect 373960 476824 373966 476836
rect 378962 476824 378968 476836
rect 379020 476824 379026 476876
rect 380710 476824 380716 476876
rect 380768 476864 380774 476876
rect 387518 476864 387524 476876
rect 380768 476836 387524 476864
rect 380768 476824 380774 476836
rect 387518 476824 387524 476836
rect 387576 476824 387582 476876
rect 390370 476824 390376 476876
rect 390428 476864 390434 476876
rect 398558 476864 398564 476876
rect 390428 476836 398564 476864
rect 390428 476824 390434 476836
rect 398558 476824 398564 476836
rect 398616 476824 398622 476876
rect 401502 476824 401508 476876
rect 401560 476864 401566 476876
rect 410702 476864 410708 476876
rect 401560 476836 410708 476864
rect 401560 476824 401566 476836
rect 410702 476824 410708 476836
rect 410760 476824 410766 476876
rect 524322 476824 524328 476876
rect 524380 476864 524386 476876
rect 551830 476864 551836 476876
rect 524380 476836 551836 476864
rect 524380 476824 524386 476836
rect 551830 476824 551836 476836
rect 551888 476824 551894 476876
rect 351730 476756 351736 476808
rect 351788 476796 351794 476808
rect 354582 476796 354588 476808
rect 351788 476768 354588 476796
rect 351788 476756 351794 476768
rect 354582 476756 354588 476768
rect 354640 476756 354646 476808
rect 371050 476756 371056 476808
rect 371108 476796 371114 476808
rect 376570 476796 376576 476808
rect 371108 476768 376576 476796
rect 371108 476756 371114 476768
rect 376570 476756 376576 476768
rect 376628 476756 376634 476808
rect 386230 476756 386236 476808
rect 386288 476796 386294 476808
rect 393682 476796 393688 476808
rect 386288 476768 393688 476796
rect 386288 476756 386294 476768
rect 393682 476756 393688 476768
rect 393740 476756 393746 476808
rect 395890 476756 395896 476808
rect 395948 476796 395954 476808
rect 404630 476796 404636 476808
rect 395948 476768 404636 476796
rect 395948 476756 395954 476768
rect 404630 476756 404636 476768
rect 404688 476756 404694 476808
rect 492582 476756 492588 476808
rect 492640 476796 492646 476808
rect 552106 476796 552112 476808
rect 492640 476768 552112 476796
rect 492640 476756 492646 476768
rect 552106 476756 552112 476768
rect 552164 476756 552170 476808
rect 361482 476688 361488 476740
rect 361540 476728 361546 476740
rect 364334 476728 364340 476740
rect 361540 476700 364340 476728
rect 361540 476688 361546 476700
rect 364334 476688 364340 476700
rect 364392 476688 364398 476740
rect 368382 476688 368388 476740
rect 368440 476728 368446 476740
rect 372890 476728 372896 476740
rect 368440 476700 372896 476728
rect 368440 476688 368446 476700
rect 372890 476688 372896 476700
rect 372948 476688 372954 476740
rect 394602 476688 394608 476740
rect 394660 476728 394666 476740
rect 402238 476728 402244 476740
rect 394660 476700 402244 476728
rect 394660 476688 394666 476700
rect 402238 476688 402244 476700
rect 402296 476688 402302 476740
rect 367002 476620 367008 476672
rect 367060 476660 367066 476672
rect 370406 476660 370412 476672
rect 367060 476632 370412 476660
rect 367060 476620 367066 476632
rect 370406 476620 370412 476632
rect 370464 476620 370470 476672
rect 316678 476552 316684 476604
rect 316736 476592 316742 476604
rect 317322 476592 317328 476604
rect 316736 476564 317328 476592
rect 316736 476552 316742 476564
rect 317322 476552 317328 476564
rect 317380 476552 317386 476604
rect 333974 476552 333980 476604
rect 334032 476592 334038 476604
rect 334986 476592 334992 476604
rect 334032 476564 334992 476592
rect 334032 476552 334038 476564
rect 334986 476552 334992 476564
rect 335044 476552 335050 476604
rect 349062 476552 349068 476604
rect 349120 476592 349126 476604
rect 350902 476592 350908 476604
rect 349120 476564 350908 476592
rect 349120 476552 349126 476564
rect 350902 476552 350908 476564
rect 350960 476552 350966 476604
rect 357342 476552 357348 476604
rect 357400 476592 357406 476604
rect 360654 476592 360660 476604
rect 357400 476564 360660 476592
rect 357400 476552 357406 476564
rect 360654 476552 360660 476564
rect 360712 476552 360718 476604
rect 366910 476552 366916 476604
rect 366968 476592 366974 476604
rect 371602 476592 371608 476604
rect 366968 476564 371608 476592
rect 366968 476552 366974 476564
rect 371602 476552 371608 476564
rect 371660 476552 371666 476604
rect 360102 476484 360108 476536
rect 360160 476524 360166 476536
rect 363046 476524 363052 476536
rect 360160 476496 363052 476524
rect 360160 476484 360166 476496
rect 363046 476484 363052 476496
rect 363104 476484 363110 476536
rect 331398 476416 331404 476468
rect 331456 476456 331462 476468
rect 332502 476456 332508 476468
rect 331456 476428 332508 476456
rect 331456 476416 331462 476428
rect 332502 476416 332508 476428
rect 332560 476416 332566 476468
rect 387702 476416 387708 476468
rect 387760 476456 387766 476468
rect 394878 476456 394884 476468
rect 387760 476428 394884 476456
rect 387760 476416 387766 476428
rect 394878 476416 394884 476428
rect 394936 476416 394942 476468
rect 347682 476348 347688 476400
rect 347740 476388 347746 476400
rect 349614 476388 349620 476400
rect 347740 476360 349620 476388
rect 347740 476348 347746 476360
rect 349614 476348 349620 476360
rect 349672 476348 349678 476400
rect 346302 476280 346308 476332
rect 346360 476320 346366 476332
rect 348418 476320 348424 476332
rect 346360 476292 348424 476320
rect 346360 476280 346366 476292
rect 348418 476280 348424 476292
rect 348476 476280 348482 476332
rect 379422 476280 379428 476332
rect 379480 476320 379486 476332
rect 385126 476320 385132 476332
rect 379480 476292 385132 476320
rect 379480 476280 379486 476292
rect 385126 476280 385132 476292
rect 385184 476280 385190 476332
rect 376662 476212 376668 476264
rect 376720 476252 376726 476264
rect 382642 476252 382648 476264
rect 376720 476224 382648 476252
rect 376720 476212 376726 476224
rect 382642 476212 382648 476224
rect 382700 476212 382706 476264
rect 384942 476212 384948 476264
rect 385000 476252 385006 476264
rect 391198 476252 391204 476264
rect 385000 476224 391204 476252
rect 385000 476212 385006 476224
rect 391198 476212 391204 476224
rect 391256 476212 391262 476264
rect 550542 475804 550548 475856
rect 550600 475844 550606 475856
rect 553394 475844 553400 475856
rect 550600 475816 553400 475844
rect 550600 475804 550606 475816
rect 553394 475804 553400 475816
rect 553452 475804 553458 475856
rect 549162 475668 549168 475720
rect 549220 475708 549226 475720
rect 553762 475708 553768 475720
rect 549220 475680 553768 475708
rect 549220 475668 549226 475680
rect 553762 475668 553768 475680
rect 553820 475668 553826 475720
rect 543642 475600 543648 475652
rect 543700 475640 543706 475652
rect 553854 475640 553860 475652
rect 543700 475612 553860 475640
rect 543700 475600 543706 475612
rect 553854 475600 553860 475612
rect 553912 475600 553918 475652
rect 538030 475532 538036 475584
rect 538088 475572 538094 475584
rect 555050 475572 555056 475584
rect 538088 475544 555056 475572
rect 538088 475532 538094 475544
rect 555050 475532 555056 475544
rect 555108 475532 555114 475584
rect 531222 475464 531228 475516
rect 531280 475504 531286 475516
rect 554406 475504 554412 475516
rect 531280 475476 554412 475504
rect 531280 475464 531286 475476
rect 554406 475464 554412 475476
rect 554464 475464 554470 475516
rect 499298 475396 499304 475448
rect 499356 475436 499362 475448
rect 527818 475436 527824 475448
rect 499356 475408 527824 475436
rect 499356 475396 499362 475408
rect 527818 475396 527824 475408
rect 527876 475396 527882 475448
rect 528462 475396 528468 475448
rect 528520 475436 528526 475448
rect 552934 475436 552940 475448
rect 528520 475408 552940 475436
rect 528520 475396 528526 475408
rect 552934 475396 552940 475408
rect 552992 475396 552998 475448
rect 518710 475328 518716 475380
rect 518768 475368 518774 475380
rect 555418 475368 555424 475380
rect 518768 475340 555424 475368
rect 518768 475328 518774 475340
rect 555418 475328 555424 475340
rect 555476 475328 555482 475380
rect 287698 474648 287704 474700
rect 287756 474688 287762 474700
rect 551922 474688 551928 474700
rect 287756 474660 551928 474688
rect 287756 474648 287762 474660
rect 551922 474648 551928 474660
rect 551980 474648 551986 474700
rect 550910 474580 550916 474632
rect 550968 474620 550974 474632
rect 553486 474620 553492 474632
rect 550968 474592 553492 474620
rect 550968 474580 550974 474592
rect 553486 474580 553492 474592
rect 553544 474580 553550 474632
rect 549898 474512 549904 474564
rect 549956 474552 549962 474564
rect 555326 474552 555332 474564
rect 549956 474524 555332 474552
rect 549956 474512 549962 474524
rect 555326 474512 555332 474524
rect 555384 474512 555390 474564
rect 538122 474308 538128 474360
rect 538180 474348 538186 474360
rect 552290 474348 552296 474360
rect 538180 474320 552296 474348
rect 538180 474308 538186 474320
rect 552290 474308 552296 474320
rect 552348 474308 552354 474360
rect 539502 474240 539508 474292
rect 539560 474280 539566 474292
rect 553946 474280 553952 474292
rect 539560 474252 553952 474280
rect 539560 474240 539566 474252
rect 553946 474240 553952 474252
rect 554004 474240 554010 474292
rect 533982 474172 533988 474224
rect 534040 474212 534046 474224
rect 552750 474212 552756 474224
rect 534040 474184 552756 474212
rect 534040 474172 534046 474184
rect 552750 474172 552756 474184
rect 552808 474172 552814 474224
rect 518802 474104 518808 474156
rect 518860 474144 518866 474156
rect 552198 474144 552204 474156
rect 518860 474116 552204 474144
rect 518860 474104 518866 474116
rect 552198 474104 552204 474116
rect 552256 474104 552262 474156
rect 512638 474036 512644 474088
rect 512696 474076 512702 474088
rect 556062 474076 556068 474088
rect 512696 474048 556068 474076
rect 512696 474036 512702 474048
rect 556062 474036 556068 474048
rect 556120 474036 556126 474088
rect 502242 473968 502248 474020
rect 502300 474008 502306 474020
rect 554958 474008 554964 474020
rect 502300 473980 554964 474008
rect 502300 473968 502306 473980
rect 554958 473968 554964 473980
rect 555016 473968 555022 474020
rect 551186 473492 551192 473544
rect 551244 473532 551250 473544
rect 551922 473532 551928 473544
rect 551244 473504 551928 473532
rect 551244 473492 551250 473504
rect 551922 473492 551928 473504
rect 551980 473492 551986 473544
rect 546586 473464 546592 473476
rect 546547 473436 546592 473464
rect 546586 473424 546592 473436
rect 546644 473424 546650 473476
rect 547782 473424 547788 473476
rect 547840 473424 547846 473476
rect 551002 473424 551008 473476
rect 551060 473464 551066 473476
rect 551462 473464 551468 473476
rect 551060 473436 551468 473464
rect 551060 473424 551066 473436
rect 551462 473424 551468 473436
rect 551520 473424 551526 473476
rect 547800 473396 547828 473424
rect 552937 473399 552995 473405
rect 552937 473396 552949 473399
rect 547800 473368 552949 473396
rect 552937 473365 552949 473368
rect 552983 473365 552995 473399
rect 552937 473359 552995 473365
rect 546589 472039 546647 472045
rect 546589 472005 546601 472039
rect 546635 472036 546647 472039
rect 554774 472036 554780 472048
rect 546635 472008 554780 472036
rect 546635 472005 546647 472008
rect 546589 471999 546647 472005
rect 554774 471996 554780 472008
rect 554832 471996 554838 472048
rect 283098 471928 283104 471980
rect 283156 471968 283162 471980
rect 283282 471968 283288 471980
rect 283156 471940 283288 471968
rect 283156 471928 283162 471940
rect 283282 471928 283288 471940
rect 283340 471928 283346 471980
rect 551646 471900 551652 471912
rect 551607 471872 551652 471900
rect 551646 471860 551652 471872
rect 551704 471860 551710 471912
rect 551462 471724 551468 471776
rect 551520 471764 551526 471776
rect 551741 471767 551799 471773
rect 551741 471764 551753 471767
rect 551520 471736 551753 471764
rect 551520 471724 551526 471736
rect 551741 471733 551753 471736
rect 551787 471733 551799 471767
rect 551741 471727 551799 471733
rect 552750 471560 552756 471572
rect 552711 471532 552756 471560
rect 552750 471520 552756 471532
rect 552808 471520 552814 471572
rect 552934 471520 552940 471572
rect 552992 471560 552998 471572
rect 553121 471563 553179 471569
rect 553121 471560 553133 471563
rect 552992 471532 553133 471560
rect 552992 471520 552998 471532
rect 553121 471529 553133 471532
rect 553167 471529 553179 471563
rect 553121 471523 553179 471529
rect 551738 471384 551744 471436
rect 551796 471424 551802 471436
rect 552106 471424 552112 471436
rect 551796 471396 552112 471424
rect 551796 471384 551802 471396
rect 552106 471384 552112 471396
rect 552164 471384 552170 471436
rect 552290 471384 552296 471436
rect 552348 471384 552354 471436
rect 552474 471384 552480 471436
rect 552532 471424 552538 471436
rect 552750 471424 552756 471436
rect 552532 471396 552756 471424
rect 552532 471384 552538 471396
rect 552750 471384 552756 471396
rect 552808 471384 552814 471436
rect 552934 471384 552940 471436
rect 552992 471424 552998 471436
rect 553302 471424 553308 471436
rect 552992 471396 553308 471424
rect 552992 471384 552998 471396
rect 553302 471384 553308 471396
rect 553360 471384 553366 471436
rect 552308 471356 552336 471384
rect 552308 471328 552520 471356
rect 552492 471232 552520 471328
rect 553118 471248 553124 471300
rect 553176 471288 553182 471300
rect 553302 471288 553308 471300
rect 553176 471260 553308 471288
rect 553176 471248 553182 471260
rect 553302 471248 553308 471260
rect 553360 471248 553366 471300
rect 552474 471180 552480 471232
rect 552532 471180 552538 471232
rect 552566 471180 552572 471232
rect 552624 471220 552630 471232
rect 552842 471220 552848 471232
rect 552624 471192 552848 471220
rect 552624 471180 552630 471192
rect 552842 471180 552848 471192
rect 552900 471180 552906 471232
rect 553118 471152 553124 471164
rect 553079 471124 553124 471152
rect 553118 471112 553124 471124
rect 553176 471112 553182 471164
rect 552750 470948 552756 470960
rect 552711 470920 552756 470948
rect 552750 470908 552756 470920
rect 552808 470908 552814 470960
rect 554222 470364 554228 470416
rect 554280 470404 554286 470416
rect 555694 470404 555700 470416
rect 554280 470376 555700 470404
rect 554280 470364 554286 470376
rect 555694 470364 555700 470376
rect 555752 470364 555758 470416
rect 552934 468500 552940 468512
rect 552895 468472 552940 468500
rect 552934 468460 552940 468472
rect 552992 468460 552998 468512
rect 554130 467576 554136 467628
rect 554188 467616 554194 467628
rect 555970 467616 555976 467628
rect 554188 467588 555976 467616
rect 554188 467576 554194 467588
rect 555970 467576 555976 467588
rect 556028 467576 556034 467628
rect 551646 467440 551652 467492
rect 551704 467480 551710 467492
rect 551741 467483 551799 467489
rect 551741 467480 551753 467483
rect 551704 467452 551753 467480
rect 551704 467440 551710 467452
rect 551741 467449 551753 467452
rect 551787 467449 551799 467483
rect 551741 467443 551799 467449
rect 551738 467344 551744 467356
rect 551699 467316 551744 467344
rect 551738 467304 551744 467316
rect 551796 467304 551802 467356
rect 552198 466964 552204 467016
rect 552256 467004 552262 467016
rect 552474 467004 552480 467016
rect 552256 466976 552480 467004
rect 552256 466964 552262 466976
rect 552474 466964 552480 466976
rect 552532 466964 552538 467016
rect 552474 466828 552480 466880
rect 552532 466868 552538 466880
rect 552750 466868 552756 466880
rect 552532 466840 552756 466868
rect 552532 466828 552538 466840
rect 552750 466828 552756 466840
rect 552808 466828 552814 466880
rect 552750 466692 552756 466744
rect 552808 466732 552814 466744
rect 553118 466732 553124 466744
rect 552808 466704 553124 466732
rect 552808 466692 552814 466704
rect 553118 466692 553124 466704
rect 553176 466692 553182 466744
rect 554682 464992 554688 465044
rect 554740 465032 554746 465044
rect 555878 465032 555884 465044
rect 554740 465004 555884 465032
rect 554740 464992 554746 465004
rect 555878 464992 555884 465004
rect 555936 464992 555942 465044
rect 279694 463632 279700 463684
rect 279752 463672 279758 463684
rect 313274 463672 313280 463684
rect 279752 463644 313280 463672
rect 279752 463632 279758 463644
rect 313274 463632 313280 463644
rect 313332 463632 313338 463684
rect 551738 463564 551744 463616
rect 551796 463604 551802 463616
rect 553026 463604 553032 463616
rect 551796 463576 553032 463604
rect 551796 463564 551802 463576
rect 553026 463564 553032 463576
rect 553084 463564 553090 463616
rect 551738 463360 551744 463412
rect 551796 463400 551802 463412
rect 553026 463400 553032 463412
rect 551796 463372 553032 463400
rect 551796 463360 551802 463372
rect 553026 463360 553032 463372
rect 553084 463360 553090 463412
rect 563698 462340 563704 462392
rect 563756 462380 563762 462392
rect 580166 462380 580172 462392
rect 563756 462352 580172 462380
rect 563756 462340 563762 462352
rect 580166 462340 580172 462352
rect 580224 462340 580230 462392
rect 283098 462312 283104 462324
rect 283059 462284 283104 462312
rect 283098 462272 283104 462284
rect 283156 462272 283162 462324
rect 552842 461796 552848 461848
rect 552900 461836 552906 461848
rect 553210 461836 553216 461848
rect 552900 461808 553216 461836
rect 552900 461796 552906 461808
rect 553210 461796 553216 461808
rect 553268 461796 553274 461848
rect 552934 461728 552940 461780
rect 552992 461728 552998 461780
rect 552952 461440 552980 461728
rect 551738 461388 551744 461440
rect 551796 461428 551802 461440
rect 552842 461428 552848 461440
rect 551796 461400 552848 461428
rect 551796 461388 551802 461400
rect 552842 461388 552848 461400
rect 552900 461388 552906 461440
rect 552934 461388 552940 461440
rect 552992 461388 552998 461440
rect 183646 460912 183652 460964
rect 183704 460952 183710 460964
rect 183830 460952 183836 460964
rect 183704 460924 183836 460952
rect 183704 460912 183710 460924
rect 183830 460912 183836 460924
rect 183888 460912 183894 460964
rect 552750 459688 552756 459740
rect 552808 459688 552814 459740
rect 552768 459536 552796 459688
rect 554038 459552 554044 459604
rect 554096 459592 554102 459604
rect 554958 459592 554964 459604
rect 554096 459564 554964 459592
rect 554096 459552 554102 459564
rect 554958 459552 554964 459564
rect 555016 459552 555022 459604
rect 552750 459484 552756 459536
rect 552808 459484 552814 459536
rect 551922 456492 551928 456544
rect 551980 456532 551986 456544
rect 552106 456532 552112 456544
rect 551980 456504 552112 456532
rect 551980 456492 551986 456504
rect 552106 456492 552112 456504
rect 552164 456492 552170 456544
rect 551830 455268 551836 455320
rect 551888 455308 551894 455320
rect 552106 455308 552112 455320
rect 551888 455280 552112 455308
rect 551888 455268 551894 455280
rect 552106 455268 552112 455280
rect 552164 455268 552170 455320
rect 283101 452659 283159 452665
rect 283101 452625 283113 452659
rect 283147 452656 283159 452659
rect 283190 452656 283196 452668
rect 283147 452628 283196 452656
rect 283147 452625 283159 452628
rect 283101 452619 283159 452625
rect 283190 452616 283196 452628
rect 283248 452616 283254 452668
rect 3418 451256 3424 451308
rect 3476 451296 3482 451308
rect 11698 451296 11704 451308
rect 3476 451268 11704 451296
rect 3476 451256 3482 451268
rect 11698 451256 11704 451268
rect 11756 451256 11762 451308
rect 283006 447108 283012 447160
rect 283064 447148 283070 447160
rect 283190 447148 283196 447160
rect 283064 447120 283196 447148
rect 283064 447108 283070 447120
rect 283190 447108 283196 447120
rect 283248 447108 283254 447160
rect 9122 444320 9128 444372
rect 9180 444360 9186 444372
rect 12526 444360 12532 444372
rect 9180 444332 12532 444360
rect 9180 444320 9186 444332
rect 12526 444320 12532 444332
rect 12584 444320 12590 444372
rect 183646 441600 183652 441652
rect 183704 441640 183710 441652
rect 183830 441640 183836 441652
rect 183704 441612 183836 441640
rect 183704 441600 183710 441612
rect 183830 441600 183836 441612
rect 183888 441600 183894 441652
rect 282917 437563 282975 437569
rect 282917 437529 282929 437563
rect 282963 437560 282975 437563
rect 283006 437560 283012 437572
rect 282963 437532 283012 437560
rect 282963 437529 282975 437532
rect 282917 437523 282975 437529
rect 283006 437520 283012 437532
rect 283064 437520 283070 437572
rect 554958 437316 554964 437368
rect 555016 437356 555022 437368
rect 557718 437356 557724 437368
rect 555016 437328 557724 437356
rect 555016 437316 555022 437328
rect 557718 437316 557724 437328
rect 557776 437316 557782 437368
rect 554774 437112 554780 437164
rect 554832 437152 554838 437164
rect 557626 437152 557632 437164
rect 554832 437124 557632 437152
rect 554832 437112 554838 437124
rect 557626 437112 557632 437124
rect 557684 437112 557690 437164
rect 554866 436024 554872 436076
rect 554924 436064 554930 436076
rect 560294 436064 560300 436076
rect 554924 436036 560300 436064
rect 554924 436024 554930 436036
rect 560294 436024 560300 436036
rect 560352 436024 560358 436076
rect 554774 435956 554780 436008
rect 554832 435996 554838 436008
rect 558178 435996 558184 436008
rect 554832 435968 558184 435996
rect 554832 435956 554838 435968
rect 558178 435956 558184 435968
rect 558236 435956 558242 436008
rect 282914 434840 282920 434852
rect 282875 434812 282920 434840
rect 282914 434800 282920 434812
rect 282972 434800 282978 434852
rect 554774 434664 554780 434716
rect 554832 434704 554838 434716
rect 561674 434704 561680 434716
rect 554832 434676 561680 434704
rect 554832 434664 554838 434676
rect 561674 434664 561680 434676
rect 561732 434664 561738 434716
rect 554866 434596 554872 434648
rect 554924 434636 554930 434648
rect 561950 434636 561956 434648
rect 554924 434608 561956 434636
rect 554924 434596 554930 434608
rect 561950 434596 561956 434608
rect 562008 434596 562014 434648
rect 282914 433276 282920 433288
rect 282875 433248 282920 433276
rect 282914 433236 282920 433248
rect 282972 433236 282978 433288
rect 554866 433236 554872 433288
rect 554924 433276 554930 433288
rect 564434 433276 564440 433288
rect 554924 433248 564440 433276
rect 554924 433236 554930 433248
rect 564434 433236 564440 433248
rect 564492 433236 564498 433288
rect 554774 433168 554780 433220
rect 554832 433208 554838 433220
rect 563054 433208 563060 433220
rect 554832 433180 563060 433208
rect 554832 433168 554838 433180
rect 563054 433168 563060 433180
rect 563112 433168 563118 433220
rect 554958 431876 554964 431928
rect 555016 431916 555022 431928
rect 567286 431916 567292 431928
rect 555016 431888 567292 431916
rect 555016 431876 555022 431888
rect 567286 431876 567292 431888
rect 567344 431876 567350 431928
rect 554774 431808 554780 431860
rect 554832 431848 554838 431860
rect 565814 431848 565820 431860
rect 554832 431820 565820 431848
rect 554832 431808 554838 431820
rect 565814 431808 565820 431820
rect 565872 431808 565878 431860
rect 554866 431740 554872 431792
rect 554924 431780 554930 431792
rect 560938 431780 560944 431792
rect 554924 431752 560944 431780
rect 554924 431740 554930 431752
rect 560938 431740 560944 431752
rect 560996 431740 561002 431792
rect 554866 430516 554872 430568
rect 554924 430556 554930 430568
rect 569954 430556 569960 430568
rect 554924 430528 569960 430556
rect 554924 430516 554930 430528
rect 569954 430516 569960 430528
rect 570012 430516 570018 430568
rect 554774 430448 554780 430500
rect 554832 430488 554838 430500
rect 568574 430488 568580 430500
rect 554832 430460 568580 430488
rect 554832 430448 554838 430460
rect 568574 430448 568580 430460
rect 568632 430448 568638 430500
rect 554774 429088 554780 429140
rect 554832 429128 554838 429140
rect 571610 429128 571616 429140
rect 554832 429100 571616 429128
rect 554832 429088 554838 429100
rect 571610 429088 571616 429100
rect 571668 429088 571674 429140
rect 554866 428884 554872 428936
rect 554924 428924 554930 428936
rect 556798 428924 556804 428936
rect 554924 428896 556804 428924
rect 554924 428884 554930 428896
rect 556798 428884 556804 428896
rect 556856 428884 556862 428936
rect 554774 427728 554780 427780
rect 554832 427768 554838 427780
rect 572714 427768 572720 427780
rect 554832 427740 572720 427768
rect 554832 427728 554838 427740
rect 572714 427728 572720 427740
rect 572772 427728 572778 427780
rect 314654 426368 314660 426420
rect 314712 426408 314718 426420
rect 499298 426408 499304 426420
rect 314712 426380 499304 426408
rect 314712 426368 314718 426380
rect 499298 426368 499304 426380
rect 499356 426368 499362 426420
rect 289630 425688 289636 425740
rect 289688 425728 289694 425740
rect 314654 425728 314660 425740
rect 289688 425700 314660 425728
rect 289688 425688 289694 425700
rect 314654 425688 314660 425700
rect 314712 425688 314718 425740
rect 3510 423648 3516 423700
rect 3568 423688 3574 423700
rect 13078 423688 13084 423700
rect 3568 423660 13084 423688
rect 3568 423648 3574 423660
rect 13078 423648 13084 423660
rect 13136 423648 13142 423700
rect 282917 423691 282975 423697
rect 282917 423657 282929 423691
rect 282963 423688 282975 423691
rect 283006 423688 283012 423700
rect 282963 423660 283012 423688
rect 282963 423657 282975 423660
rect 282917 423651 282975 423657
rect 283006 423648 283012 423660
rect 283064 423648 283070 423700
rect 183646 422288 183652 422340
rect 183704 422328 183710 422340
rect 183830 422328 183836 422340
rect 183704 422300 183836 422328
rect 183704 422288 183710 422300
rect 183830 422288 183836 422300
rect 183888 422288 183894 422340
rect 281626 421540 281632 421592
rect 281684 421580 281690 421592
rect 282270 421580 282276 421592
rect 281684 421552 282276 421580
rect 281684 421540 281690 421552
rect 282270 421540 282276 421552
rect 282328 421580 282334 421592
rect 292574 421580 292580 421592
rect 282328 421552 292580 421580
rect 282328 421540 282334 421552
rect 292574 421540 292580 421552
rect 292632 421540 292638 421592
rect 304350 415420 304356 415472
rect 304408 415460 304414 415472
rect 580166 415460 580172 415472
rect 304408 415432 580172 415460
rect 304408 415420 304414 415432
rect 580166 415420 580172 415432
rect 580224 415420 580230 415472
rect 283098 415392 283104 415404
rect 283059 415364 283104 415392
rect 283098 415352 283104 415364
rect 283156 415352 283162 415404
rect 283101 405739 283159 405745
rect 283101 405705 283113 405739
rect 283147 405736 283159 405739
rect 283190 405736 283196 405748
rect 283147 405708 283196 405736
rect 283147 405705 283159 405708
rect 283101 405699 283159 405705
rect 283190 405696 283196 405708
rect 283248 405696 283254 405748
rect 183646 402976 183652 403028
rect 183704 403016 183710 403028
rect 183830 403016 183836 403028
rect 183704 402988 183836 403016
rect 183704 402976 183710 402988
rect 183830 402976 183836 402988
rect 183888 402976 183894 403028
rect 153197 402339 153255 402345
rect 153197 402305 153209 402339
rect 153243 402336 153255 402339
rect 283190 402336 283196 402348
rect 153243 402308 283196 402336
rect 153243 402305 153255 402308
rect 153197 402299 153255 402305
rect 283190 402296 283196 402308
rect 283248 402296 283254 402348
rect 86957 402067 87015 402073
rect 86957 402064 86969 402067
rect 80348 402036 86969 402064
rect 80348 402005 80376 402036
rect 86957 402033 86969 402036
rect 87003 402033 87015 402067
rect 86957 402027 87015 402033
rect 99469 402067 99527 402073
rect 99469 402033 99481 402067
rect 99515 402064 99527 402067
rect 106277 402067 106335 402073
rect 106277 402064 106289 402067
rect 99515 402036 106289 402064
rect 99515 402033 99527 402036
rect 99469 402027 99527 402033
rect 106277 402033 106289 402036
rect 106323 402033 106335 402067
rect 106277 402027 106335 402033
rect 80333 401999 80391 402005
rect 80333 401965 80345 401999
rect 80379 401965 80391 401999
rect 80333 401959 80391 401965
rect 96525 401999 96583 402005
rect 96525 401965 96537 401999
rect 96571 401996 96583 401999
rect 99285 401999 99343 402005
rect 99285 401996 99297 401999
rect 96571 401968 99297 401996
rect 96571 401965 96583 401968
rect 96525 401959 96583 401965
rect 99285 401965 99297 401968
rect 99331 401965 99343 401999
rect 99285 401959 99343 401965
rect 115845 401999 115903 402005
rect 115845 401965 115857 401999
rect 115891 401996 115903 401999
rect 118605 401999 118663 402005
rect 118605 401996 118617 401999
rect 115891 401968 118617 401996
rect 115891 401965 115903 401968
rect 115845 401959 115903 401965
rect 118605 401965 118617 401968
rect 118651 401965 118663 401999
rect 118605 401959 118663 401965
rect 128357 401999 128415 402005
rect 128357 401965 128369 401999
rect 128403 401996 128415 401999
rect 133877 401999 133935 402005
rect 133877 401996 133889 401999
rect 128403 401968 133889 401996
rect 128403 401965 128415 401968
rect 128357 401959 128415 401965
rect 133877 401965 133889 401968
rect 133923 401965 133935 401999
rect 133877 401959 133935 401965
rect 143445 401999 143503 402005
rect 143445 401965 143457 401999
rect 143491 401996 143503 401999
rect 143491 401968 144960 401996
rect 143491 401965 143503 401968
rect 143445 401959 143503 401965
rect 144932 401937 144960 401968
rect 118789 401931 118847 401937
rect 118789 401897 118801 401931
rect 118835 401928 118847 401931
rect 128265 401931 128323 401937
rect 128265 401928 128277 401931
rect 118835 401900 128277 401928
rect 118835 401897 118847 401900
rect 118789 401891 118847 401897
rect 128265 401897 128277 401900
rect 128311 401897 128323 401931
rect 128265 401891 128323 401897
rect 144917 401931 144975 401937
rect 144917 401897 144929 401931
rect 144963 401897 144975 401931
rect 144917 401891 144975 401897
rect 86957 401863 87015 401869
rect 86957 401829 86969 401863
rect 87003 401860 87015 401863
rect 96525 401863 96583 401869
rect 96525 401860 96537 401863
rect 87003 401832 96537 401860
rect 87003 401829 87015 401832
rect 86957 401823 87015 401829
rect 96525 401829 96537 401832
rect 96571 401829 96583 401863
rect 96525 401823 96583 401829
rect 106277 401863 106335 401869
rect 106277 401829 106289 401863
rect 106323 401860 106335 401863
rect 115845 401863 115903 401869
rect 115845 401860 115857 401863
rect 106323 401832 115857 401860
rect 106323 401829 106335 401832
rect 106277 401823 106335 401829
rect 115845 401829 115857 401832
rect 115891 401829 115903 401863
rect 115845 401823 115903 401829
rect 133877 401863 133935 401869
rect 133877 401829 133889 401863
rect 133923 401860 133935 401863
rect 143445 401863 143503 401869
rect 143445 401860 143457 401863
rect 133923 401832 143457 401860
rect 133923 401829 133935 401832
rect 133877 401823 133935 401829
rect 143445 401829 143457 401832
rect 143491 401829 143503 401863
rect 143445 401823 143503 401829
rect 144917 401795 144975 401801
rect 144917 401761 144929 401795
rect 144963 401792 144975 401795
rect 153197 401795 153255 401801
rect 153197 401792 153209 401795
rect 144963 401764 153209 401792
rect 144963 401761 144975 401764
rect 144917 401755 144975 401761
rect 153197 401761 153209 401764
rect 153243 401761 153255 401795
rect 153197 401755 153255 401761
rect 143442 401548 143448 401600
rect 143500 401588 143506 401600
rect 153654 401588 153660 401600
rect 143500 401560 153660 401588
rect 143500 401548 143506 401560
rect 153654 401548 153660 401560
rect 153712 401548 153718 401600
rect 142062 401480 142068 401532
rect 142120 401520 142126 401532
rect 153930 401520 153936 401532
rect 142120 401492 153936 401520
rect 142120 401480 142126 401492
rect 153930 401480 153936 401492
rect 153988 401480 153994 401532
rect 140682 401412 140688 401464
rect 140740 401452 140746 401464
rect 154022 401452 154028 401464
rect 140740 401424 154028 401452
rect 140740 401412 140746 401424
rect 154022 401412 154028 401424
rect 154080 401412 154086 401464
rect 140590 401344 140596 401396
rect 140648 401384 140654 401396
rect 154206 401384 154212 401396
rect 140648 401356 154212 401384
rect 140648 401344 140654 401356
rect 154206 401344 154212 401356
rect 154264 401344 154270 401396
rect 137922 401276 137928 401328
rect 137980 401316 137986 401328
rect 154114 401316 154120 401328
rect 137980 401288 154120 401316
rect 137980 401276 137986 401288
rect 154114 401276 154120 401288
rect 154172 401276 154178 401328
rect 136450 401208 136456 401260
rect 136508 401248 136514 401260
rect 154298 401248 154304 401260
rect 136508 401220 154304 401248
rect 136508 401208 136514 401220
rect 154298 401208 154304 401220
rect 154356 401208 154362 401260
rect 133782 401140 133788 401192
rect 133840 401180 133846 401192
rect 154850 401180 154856 401192
rect 133840 401152 154856 401180
rect 133840 401140 133846 401152
rect 154850 401140 154856 401152
rect 154908 401140 154914 401192
rect 132402 401072 132408 401124
rect 132460 401112 132466 401124
rect 154390 401112 154396 401124
rect 132460 401084 154396 401112
rect 132460 401072 132466 401084
rect 154390 401072 154396 401084
rect 154448 401072 154454 401124
rect 128262 401004 128268 401056
rect 128320 401044 128326 401056
rect 154482 401044 154488 401056
rect 128320 401016 154488 401044
rect 128320 401004 128326 401016
rect 154482 401004 154488 401016
rect 154540 401004 154546 401056
rect 121270 400936 121276 400988
rect 121328 400976 121334 400988
rect 153838 400976 153844 400988
rect 121328 400948 153844 400976
rect 121328 400936 121334 400948
rect 153838 400936 153844 400948
rect 153896 400936 153902 400988
rect 118602 400868 118608 400920
rect 118660 400908 118666 400920
rect 153102 400908 153108 400920
rect 118660 400880 153108 400908
rect 118660 400868 118666 400880
rect 153102 400868 153108 400880
rect 153160 400868 153166 400920
rect 144822 400800 144828 400852
rect 144880 400840 144886 400852
rect 153562 400840 153568 400852
rect 144880 400812 153568 400840
rect 144880 400800 144886 400812
rect 153562 400800 153568 400812
rect 153620 400800 153626 400852
rect 146110 400460 146116 400512
rect 146168 400500 146174 400512
rect 153746 400500 153752 400512
rect 146168 400472 153752 400500
rect 146168 400460 146174 400472
rect 153746 400460 153752 400472
rect 153804 400460 153810 400512
rect 77938 396584 77944 396636
rect 77996 396624 78002 396636
rect 80333 396627 80391 396633
rect 80333 396624 80345 396627
rect 77996 396596 80345 396624
rect 77996 396584 78002 396596
rect 80333 396593 80345 396596
rect 80379 396593 80391 396627
rect 80333 396587 80391 396593
rect 183646 383664 183652 383716
rect 183704 383704 183710 383716
rect 183830 383704 183836 383716
rect 183704 383676 183836 383704
rect 183704 383664 183710 383676
rect 183830 383664 183836 383676
rect 183888 383664 183894 383716
rect 282270 377000 282276 377052
rect 282328 377040 282334 377052
rect 284294 377040 284300 377052
rect 282328 377012 284300 377040
rect 282328 377000 282334 377012
rect 284294 377000 284300 377012
rect 284352 377000 284358 377052
rect 304442 368500 304448 368552
rect 304500 368540 304506 368552
rect 580166 368540 580172 368552
rect 304500 368512 580172 368540
rect 304500 368500 304506 368512
rect 580166 368500 580172 368512
rect 580224 368500 580230 368552
rect 183646 364352 183652 364404
rect 183704 364392 183710 364404
rect 183830 364392 183836 364404
rect 183704 364364 183836 364392
rect 183704 364352 183710 364364
rect 183830 364352 183836 364364
rect 183888 364352 183894 364404
rect 282270 360136 282276 360188
rect 282328 360176 282334 360188
rect 282546 360176 282552 360188
rect 282328 360148 282552 360176
rect 282328 360136 282334 360148
rect 282546 360136 282552 360148
rect 282604 360136 282610 360188
rect 187786 358300 187792 358352
rect 187844 358340 187850 358352
rect 191926 358340 191932 358352
rect 187844 358312 191932 358340
rect 187844 358300 187850 358312
rect 191926 358300 191932 358312
rect 191984 358300 191990 358352
rect 187878 358096 187884 358148
rect 187936 358136 187942 358148
rect 193306 358136 193312 358148
rect 187936 358108 193312 358136
rect 187936 358096 187942 358108
rect 193306 358096 193312 358108
rect 193364 358096 193370 358148
rect 282365 357391 282423 357397
rect 282365 357357 282377 357391
rect 282411 357388 282423 357391
rect 282546 357388 282552 357400
rect 282411 357360 282552 357388
rect 282411 357357 282423 357360
rect 282365 357351 282423 357357
rect 282546 357348 282552 357360
rect 282604 357348 282610 357400
rect 194410 355988 194416 356040
rect 194468 356028 194474 356040
rect 198918 356028 198924 356040
rect 194468 356000 198924 356028
rect 194468 355988 194474 356000
rect 198918 355988 198924 356000
rect 198976 355988 198982 356040
rect 201402 355988 201408 356040
rect 201460 356028 201466 356040
rect 206922 356028 206928 356040
rect 201460 356000 206928 356028
rect 201460 355988 201466 356000
rect 206922 355988 206928 356000
rect 206980 355988 206986 356040
rect 210326 355988 210332 356040
rect 210384 356028 210390 356040
rect 214742 356028 214748 356040
rect 210384 356000 214748 356028
rect 210384 355988 210390 356000
rect 214742 355988 214748 356000
rect 214800 355988 214806 356040
rect 215202 355988 215208 356040
rect 215260 356028 215266 356040
rect 218974 356028 218980 356040
rect 215260 356000 218980 356028
rect 215260 355988 215266 356000
rect 218974 355988 218980 356000
rect 219032 355988 219038 356040
rect 221274 355988 221280 356040
rect 221332 356028 221338 356040
rect 223206 356028 223212 356040
rect 221332 356000 223212 356028
rect 221332 355988 221338 356000
rect 223206 355988 223212 356000
rect 223264 355988 223270 356040
rect 226150 355988 226156 356040
rect 226208 356028 226214 356040
rect 226978 356028 226984 356040
rect 226208 356000 226984 356028
rect 226208 355988 226214 356000
rect 226978 355988 226984 356000
rect 227036 355988 227042 356040
rect 233142 355988 233148 356040
rect 233200 356028 233206 356040
rect 233694 356028 233700 356040
rect 233200 356000 233700 356028
rect 233200 355988 233206 356000
rect 233694 355988 233700 356000
rect 233752 355988 233758 356040
rect 234522 355988 234528 356040
rect 234580 356028 234586 356040
rect 235902 356028 235908 356040
rect 234580 356000 235908 356028
rect 234580 355988 234586 356000
rect 235902 355988 235908 356000
rect 235960 355988 235966 356040
rect 239582 355988 239588 356040
rect 239640 356028 239646 356040
rect 240502 356028 240508 356040
rect 239640 356000 240508 356028
rect 239640 355988 239646 356000
rect 240502 355988 240508 356000
rect 240560 355988 240566 356040
rect 242066 355988 242072 356040
rect 242124 356028 242130 356040
rect 242894 356028 242900 356040
rect 242124 356000 242900 356028
rect 242124 355988 242130 356000
rect 242894 355988 242900 356000
rect 242952 355988 242958 356040
rect 258074 355988 258080 356040
rect 258132 356028 258138 356040
rect 258534 356028 258540 356040
rect 258132 356000 258540 356028
rect 258132 355988 258138 356000
rect 258534 355988 258540 356000
rect 258592 355988 258598 356040
rect 261570 355988 261576 356040
rect 261628 356028 261634 356040
rect 262214 356028 262220 356040
rect 261628 356000 262220 356028
rect 261628 355988 261634 356000
rect 262214 355988 262220 356000
rect 262272 355988 262278 356040
rect 262674 355988 262680 356040
rect 262732 356028 262738 356040
rect 263594 356028 263600 356040
rect 262732 356000 263600 356028
rect 262732 355988 262738 356000
rect 263594 355988 263600 356000
rect 263652 355988 263658 356040
rect 191742 355920 191748 355972
rect 191800 355960 191806 355972
rect 198642 355960 198648 355972
rect 191800 355932 198648 355960
rect 191800 355920 191806 355932
rect 198642 355920 198648 355932
rect 198700 355920 198706 355972
rect 200482 355920 200488 355972
rect 200540 355960 200546 355972
rect 206094 355960 206100 355972
rect 200540 355932 206100 355960
rect 200540 355920 200546 355932
rect 206094 355920 206100 355932
rect 206152 355920 206158 355972
rect 222102 355920 222108 355972
rect 222160 355960 222166 355972
rect 225414 355960 225420 355972
rect 222160 355932 225420 355960
rect 222160 355920 222166 355932
rect 225414 355920 225420 355932
rect 225472 355920 225478 355972
rect 232314 355920 232320 355972
rect 232372 355960 232378 355972
rect 234062 355960 234068 355972
rect 232372 355932 234068 355960
rect 232372 355920 232378 355932
rect 234062 355920 234068 355932
rect 234120 355920 234126 355972
rect 193122 355852 193128 355904
rect 193180 355892 193186 355904
rect 199654 355892 199660 355904
rect 193180 355864 199660 355892
rect 193180 355852 193186 355864
rect 199654 355852 199660 355864
rect 199712 355852 199718 355904
rect 204162 355852 204168 355904
rect 204220 355892 204226 355904
rect 209222 355892 209228 355904
rect 204220 355864 209228 355892
rect 204220 355852 204226 355864
rect 209222 355852 209228 355864
rect 209280 355852 209286 355904
rect 213822 355852 213828 355904
rect 213880 355892 213886 355904
rect 218054 355892 218060 355904
rect 213880 355864 218060 355892
rect 213880 355852 213886 355864
rect 218054 355852 218060 355864
rect 218112 355852 218118 355904
rect 220078 355852 220084 355904
rect 220136 355892 220142 355904
rect 223666 355892 223672 355904
rect 220136 355864 223672 355892
rect 220136 355852 220142 355864
rect 223666 355852 223672 355864
rect 223724 355852 223730 355904
rect 231026 355852 231032 355904
rect 231084 355892 231090 355904
rect 233142 355892 233148 355904
rect 231084 355864 233148 355892
rect 231084 355852 231090 355864
rect 233142 355852 233148 355864
rect 233200 355852 233206 355904
rect 211522 355784 211528 355836
rect 211580 355824 211586 355836
rect 215662 355824 215668 355836
rect 211580 355796 215668 355824
rect 211580 355784 211586 355796
rect 215662 355784 215668 355796
rect 215720 355784 215726 355836
rect 229830 355784 229836 355836
rect 229888 355824 229894 355836
rect 230474 355824 230480 355836
rect 229888 355796 230480 355824
rect 229888 355784 229894 355796
rect 230474 355784 230480 355796
rect 230532 355784 230538 355836
rect 235810 355784 235816 355836
rect 235868 355824 235874 355836
rect 237282 355824 237288 355836
rect 235868 355796 237288 355824
rect 235868 355784 235874 355796
rect 237282 355784 237288 355796
rect 237340 355784 237346 355836
rect 240870 355784 240876 355836
rect 240928 355824 240934 355836
rect 241698 355824 241704 355836
rect 240928 355796 241704 355824
rect 240928 355784 240934 355796
rect 241698 355784 241704 355796
rect 241756 355784 241762 355836
rect 199286 355716 199292 355768
rect 199344 355756 199350 355768
rect 204990 355756 204996 355768
rect 199344 355728 204996 355756
rect 199344 355716 199350 355728
rect 204990 355716 204996 355728
rect 205048 355716 205054 355768
rect 209038 355716 209044 355768
rect 209096 355756 209102 355768
rect 214006 355756 214012 355768
rect 209096 355728 214012 355756
rect 209096 355716 209102 355728
rect 214006 355716 214012 355728
rect 214064 355716 214070 355768
rect 198090 355648 198096 355700
rect 198148 355688 198154 355700
rect 203886 355688 203892 355700
rect 198148 355660 203892 355688
rect 198148 355648 198154 355660
rect 203886 355648 203892 355660
rect 203944 355648 203950 355700
rect 217594 355648 217600 355700
rect 217652 355688 217658 355700
rect 221182 355688 221188 355700
rect 217652 355660 221188 355688
rect 217652 355648 217658 355660
rect 221182 355648 221188 355660
rect 221240 355648 221246 355700
rect 255314 355648 255320 355700
rect 255372 355688 255378 355700
rect 256050 355688 256056 355700
rect 255372 355660 256056 355688
rect 255372 355648 255378 355660
rect 256050 355648 256056 355660
rect 256108 355648 256114 355700
rect 196802 355580 196808 355632
rect 196860 355620 196866 355632
rect 201494 355620 201500 355632
rect 196860 355592 201500 355620
rect 196860 355580 196866 355592
rect 201494 355580 201500 355592
rect 201552 355580 201558 355632
rect 218882 355512 218888 355564
rect 218940 355552 218946 355564
rect 222378 355552 222384 355564
rect 218940 355524 222384 355552
rect 218940 355512 218946 355524
rect 222378 355512 222384 355524
rect 222436 355512 222442 355564
rect 224862 355512 224868 355564
rect 224920 355552 224926 355564
rect 227714 355552 227720 355564
rect 224920 355524 227720 355552
rect 224920 355512 224926 355524
rect 227714 355512 227720 355524
rect 227772 355512 227778 355564
rect 263410 355512 263416 355564
rect 263468 355552 263474 355564
rect 264606 355552 264612 355564
rect 263468 355524 264612 355552
rect 263468 355512 263474 355524
rect 264606 355512 264612 355524
rect 264664 355512 264670 355564
rect 207842 355376 207848 355428
rect 207900 355416 207906 355428
rect 212626 355416 212632 355428
rect 207900 355388 212632 355416
rect 207900 355376 207906 355388
rect 212626 355376 212632 355388
rect 212684 355376 212690 355428
rect 227438 355376 227444 355428
rect 227496 355416 227502 355428
rect 228818 355416 228824 355428
rect 227496 355388 228824 355416
rect 227496 355376 227502 355388
rect 228818 355376 228824 355388
rect 228876 355376 228882 355428
rect 256694 355376 256700 355428
rect 256752 355416 256758 355428
rect 257338 355416 257344 355428
rect 256752 355388 257344 355416
rect 256752 355376 256758 355388
rect 257338 355376 257344 355388
rect 257396 355376 257402 355428
rect 266078 355376 266084 355428
rect 266136 355416 266142 355428
rect 267090 355416 267096 355428
rect 266136 355388 267096 355416
rect 266136 355376 266142 355388
rect 267090 355376 267096 355388
rect 267148 355376 267154 355428
rect 243262 355308 243268 355360
rect 243320 355348 243326 355360
rect 243814 355348 243820 355360
rect 243320 355320 243820 355348
rect 243320 355308 243326 355320
rect 243814 355308 243820 355320
rect 243872 355308 243878 355360
rect 244090 355308 244096 355360
rect 244148 355348 244154 355360
rect 244918 355348 244924 355360
rect 244148 355320 244924 355348
rect 244148 355308 244154 355320
rect 244918 355308 244924 355320
rect 244976 355308 244982 355360
rect 264882 355240 264888 355292
rect 264940 355280 264946 355292
rect 265894 355280 265900 355292
rect 264940 355252 265900 355280
rect 264940 355240 264946 355252
rect 265894 355240 265900 355252
rect 265952 355240 265958 355292
rect 202782 355172 202788 355224
rect 202840 355212 202846 355224
rect 208302 355212 208308 355224
rect 202840 355184 208308 355212
rect 202840 355172 202846 355184
rect 208302 355172 208308 355184
rect 208360 355172 208366 355224
rect 254118 355104 254124 355156
rect 254176 355144 254182 355156
rect 254854 355144 254860 355156
rect 254176 355116 254860 355144
rect 254176 355104 254182 355116
rect 254854 355104 254860 355116
rect 254912 355104 254918 355156
rect 268194 355104 268200 355156
rect 268252 355144 268258 355156
rect 269482 355144 269488 355156
rect 268252 355116 269488 355144
rect 268252 355104 268258 355116
rect 269482 355104 269488 355116
rect 269540 355104 269546 355156
rect 212350 354968 212356 355020
rect 212408 355008 212414 355020
rect 216766 355008 216772 355020
rect 212408 354980 216772 355008
rect 212408 354968 212414 354980
rect 216766 354968 216772 354980
rect 216824 354968 216830 355020
rect 237190 354968 237196 355020
rect 237248 355008 237254 355020
rect 238294 355008 238300 355020
rect 237248 354980 238300 355008
rect 237248 354968 237254 354980
rect 238294 354968 238300 354980
rect 238352 354968 238358 355020
rect 189534 354832 189540 354884
rect 189592 354872 189598 354884
rect 193674 354872 193680 354884
rect 189592 354844 193680 354872
rect 189592 354832 189598 354844
rect 193674 354832 193680 354844
rect 193732 354832 193738 354884
rect 190362 354764 190368 354816
rect 190420 354804 190426 354816
rect 193858 354804 193864 354816
rect 190420 354776 193864 354804
rect 190420 354764 190426 354776
rect 193858 354764 193864 354776
rect 193916 354764 193922 354816
rect 206646 354764 206652 354816
rect 206704 354804 206710 354816
rect 211430 354804 211436 354816
rect 206704 354776 211436 354804
rect 206704 354764 206710 354776
rect 211430 354764 211436 354776
rect 211488 354764 211494 354816
rect 223390 354764 223396 354816
rect 223448 354804 223454 354816
rect 226518 354804 226524 354816
rect 223448 354776 226524 354804
rect 223448 354764 223454 354776
rect 226518 354764 226524 354776
rect 226576 354764 226582 354816
rect 238386 354764 238392 354816
rect 238444 354804 238450 354816
rect 239398 354804 239404 354816
rect 238444 354776 239404 354804
rect 238444 354764 238450 354776
rect 239398 354764 239404 354776
rect 239456 354764 239462 354816
rect 248046 354764 248052 354816
rect 248104 354804 248110 354816
rect 248598 354804 248604 354816
rect 248104 354776 248604 354804
rect 248104 354764 248110 354776
rect 248598 354764 248604 354776
rect 248656 354764 248662 354816
rect 188338 354696 188344 354748
rect 188396 354736 188402 354748
rect 195238 354736 195244 354748
rect 188396 354708 195244 354736
rect 188396 354696 188402 354708
rect 195238 354696 195244 354708
rect 195296 354696 195302 354748
rect 195606 354696 195612 354748
rect 195664 354736 195670 354748
rect 201402 354736 201408 354748
rect 195664 354708 201408 354736
rect 195664 354696 195670 354708
rect 201402 354696 201408 354708
rect 201460 354696 201466 354748
rect 205358 354696 205364 354748
rect 205416 354736 205422 354748
rect 210326 354736 210332 354748
rect 205416 354708 210332 354736
rect 205416 354696 205422 354708
rect 210326 354696 210332 354708
rect 210384 354696 210390 354748
rect 216398 354696 216404 354748
rect 216456 354736 216462 354748
rect 220078 354736 220084 354748
rect 216456 354708 220084 354736
rect 216456 354696 216462 354708
rect 220078 354696 220084 354708
rect 220136 354696 220142 354748
rect 228634 354696 228640 354748
rect 228692 354736 228698 354748
rect 230382 354736 230388 354748
rect 228692 354708 230388 354736
rect 228692 354696 228698 354708
rect 230382 354696 230388 354708
rect 230440 354696 230446 354748
rect 260558 354696 260564 354748
rect 260616 354736 260622 354748
rect 261018 354736 261024 354748
rect 260616 354708 261024 354736
rect 260616 354696 260622 354708
rect 261018 354696 261024 354708
rect 261076 354696 261082 354748
rect 267090 354696 267096 354748
rect 267148 354736 267154 354748
rect 268286 354736 268292 354748
rect 267148 354708 268292 354736
rect 267148 354696 267154 354708
rect 268286 354696 268292 354708
rect 268344 354696 268350 354748
rect 278774 354696 278780 354748
rect 278832 354736 278838 354748
rect 280522 354736 280528 354748
rect 278832 354708 280528 354736
rect 278832 354696 278838 354708
rect 280522 354696 280528 354708
rect 280580 354696 280586 354748
rect 46842 354628 46848 354680
rect 46900 354668 46906 354680
rect 58526 354668 58532 354680
rect 46900 354640 58532 354668
rect 46900 354628 46906 354640
rect 58526 354628 58532 354640
rect 58584 354628 58590 354680
rect 48314 354560 48320 354612
rect 48372 354600 48378 354612
rect 59630 354600 59636 354612
rect 48372 354572 59636 354600
rect 48372 354560 48378 354572
rect 59630 354560 59636 354572
rect 59688 354560 59694 354612
rect 29914 354492 29920 354544
rect 29972 354532 29978 354544
rect 35802 354532 35808 354544
rect 29972 354504 35808 354532
rect 29972 354492 29978 354504
rect 35802 354492 35808 354504
rect 35860 354492 35866 354544
rect 45462 354492 45468 354544
rect 45520 354532 45526 354544
rect 57514 354532 57520 354544
rect 45520 354504 57520 354532
rect 45520 354492 45526 354504
rect 57514 354492 57520 354504
rect 57572 354492 57578 354544
rect 34974 354424 34980 354476
rect 35032 354464 35038 354476
rect 40034 354464 40040 354476
rect 35032 354436 40040 354464
rect 35032 354424 35038 354436
rect 40034 354424 40040 354436
rect 40092 354424 40098 354476
rect 47854 354424 47860 354476
rect 47912 354464 47918 354476
rect 59354 354464 59360 354476
rect 47912 354436 59360 354464
rect 47912 354424 47918 354436
rect 59354 354424 59360 354436
rect 59412 354424 59418 354476
rect 35618 354356 35624 354408
rect 35676 354396 35682 354408
rect 40218 354396 40224 354408
rect 35676 354368 40224 354396
rect 35676 354356 35682 354368
rect 40218 354356 40224 354368
rect 40276 354356 40282 354408
rect 46474 354356 46480 354408
rect 46532 354396 46538 354408
rect 58066 354396 58072 354408
rect 46532 354368 58072 354396
rect 46532 354356 46538 354368
rect 58066 354356 58072 354368
rect 58124 354356 58130 354408
rect 38378 354288 38384 354340
rect 38436 354328 38442 354340
rect 48590 354328 48596 354340
rect 38436 354300 48596 354328
rect 38436 354288 38442 354300
rect 48590 354288 48596 354300
rect 48648 354288 48654 354340
rect 49326 354288 49332 354340
rect 49384 354328 49390 354340
rect 64966 354328 64972 354340
rect 49384 354300 64972 354328
rect 49384 354288 49390 354300
rect 64966 354288 64972 354300
rect 65024 354288 65030 354340
rect 39942 354220 39948 354272
rect 40000 354260 40006 354272
rect 50982 354260 50988 354272
rect 40000 354232 50988 354260
rect 40000 354220 40006 354232
rect 50982 354220 50988 354232
rect 51040 354220 51046 354272
rect 52914 354220 52920 354272
rect 52972 354260 52978 354272
rect 70394 354260 70400 354272
rect 52972 354232 70400 354260
rect 52972 354220 52978 354232
rect 70394 354220 70400 354232
rect 70452 354220 70458 354272
rect 41230 354152 41236 354204
rect 41288 354192 41294 354204
rect 53006 354192 53012 354204
rect 41288 354164 53012 354192
rect 41288 354152 41294 354164
rect 53006 354152 53012 354164
rect 53064 354152 53070 354204
rect 55766 354152 55772 354204
rect 55824 354192 55830 354204
rect 74718 354192 74724 354204
rect 55824 354164 74724 354192
rect 55824 354152 55830 354164
rect 74718 354152 74724 354164
rect 74776 354152 74782 354204
rect 25590 354084 25596 354136
rect 25648 354124 25654 354136
rect 29270 354124 29276 354136
rect 25648 354096 29276 354124
rect 25648 354084 25654 354096
rect 29270 354084 29276 354096
rect 29328 354084 29334 354136
rect 32766 354084 32772 354136
rect 32824 354124 32830 354136
rect 38194 354124 38200 354136
rect 32824 354096 38200 354124
rect 32824 354084 32830 354096
rect 38194 354084 38200 354096
rect 38252 354084 38258 354136
rect 42702 354084 42708 354136
rect 42760 354124 42766 354136
rect 55122 354124 55128 354136
rect 42760 354096 55128 354124
rect 42760 354084 42766 354096
rect 55122 354084 55128 354096
rect 55180 354084 55186 354136
rect 58618 354084 58624 354136
rect 58676 354124 58682 354136
rect 78766 354124 78772 354136
rect 58676 354096 78772 354124
rect 58676 354084 58682 354096
rect 78766 354084 78772 354096
rect 78824 354084 78830 354136
rect 26142 354016 26148 354068
rect 26200 354056 26206 354068
rect 30374 354056 30380 354068
rect 26200 354028 30380 354056
rect 26200 354016 26206 354028
rect 30374 354016 30380 354028
rect 30432 354016 30438 354068
rect 34238 354016 34244 354068
rect 34296 354056 34302 354068
rect 39206 354056 39212 354068
rect 34296 354028 39212 354056
rect 34296 354016 34302 354028
rect 39206 354016 39212 354028
rect 39264 354016 39270 354068
rect 45002 354016 45008 354068
rect 45060 354056 45066 354068
rect 56778 354056 56784 354068
rect 45060 354028 56784 354056
rect 45060 354016 45066 354028
rect 56778 354016 56784 354028
rect 56836 354016 56842 354068
rect 61562 354016 61568 354068
rect 61620 354056 61626 354068
rect 83182 354056 83188 354068
rect 61620 354028 83188 354056
rect 61620 354016 61626 354028
rect 83182 354016 83188 354028
rect 83240 354016 83246 354068
rect 44082 353948 44088 354000
rect 44140 353988 44146 354000
rect 57238 353988 57244 354000
rect 44140 353960 57244 353988
rect 44140 353948 44146 353960
rect 57238 353948 57244 353960
rect 57296 353948 57302 354000
rect 64414 353948 64420 354000
rect 64472 353988 64478 354000
rect 87414 353988 87420 354000
rect 64472 353960 87420 353988
rect 64472 353948 64478 353960
rect 87414 353948 87420 353960
rect 87472 353948 87478 354000
rect 39298 353880 39304 353932
rect 39356 353920 39362 353932
rect 49694 353920 49700 353932
rect 39356 353892 49700 353920
rect 39356 353880 39362 353892
rect 49694 353880 49700 353892
rect 49752 353880 49758 353932
rect 50706 353880 50712 353932
rect 50764 353920 50770 353932
rect 62206 353920 62212 353932
rect 50764 353892 62212 353920
rect 50764 353880 50770 353892
rect 62206 353880 62212 353892
rect 62264 353880 62270 353932
rect 33410 353812 33416 353864
rect 33468 353852 33474 353864
rect 38654 353852 38660 353864
rect 33468 353824 38660 353852
rect 33468 353812 33474 353824
rect 38654 353812 38660 353824
rect 38712 353812 38718 353864
rect 51442 353812 51448 353864
rect 51500 353852 51506 353864
rect 63494 353852 63500 353864
rect 51500 353824 63500 353852
rect 51500 353812 51506 353824
rect 63494 353812 63500 353824
rect 63552 353812 63558 353864
rect 30282 353676 30288 353728
rect 30340 353716 30346 353728
rect 34514 353716 34520 353728
rect 30340 353688 34520 353716
rect 30340 353676 30346 353688
rect 34514 353676 34520 353688
rect 34572 353676 34578 353728
rect 37090 353676 37096 353728
rect 37148 353716 37154 353728
rect 42242 353716 42248 353728
rect 37148 353688 42248 353716
rect 37148 353676 37154 353688
rect 42242 353676 42248 353688
rect 42300 353676 42306 353728
rect 43530 353676 43536 353728
rect 43588 353716 43594 353728
rect 56134 353716 56140 353728
rect 43588 353688 56140 353716
rect 43588 353676 43594 353688
rect 56134 353676 56140 353688
rect 56192 353676 56198 353728
rect 28902 353608 28908 353660
rect 28960 353648 28966 353660
rect 34422 353648 34428 353660
rect 28960 353620 34428 353648
rect 28960 353608 28966 353620
rect 34422 353608 34428 353620
rect 34480 353608 34486 353660
rect 42150 353608 42156 353660
rect 42208 353648 42214 353660
rect 54110 353648 54116 353660
rect 42208 353620 54116 353648
rect 42208 353608 42214 353620
rect 54110 353608 54116 353620
rect 54168 353608 54174 353660
rect 27062 353540 27068 353592
rect 27120 353580 27126 353592
rect 31846 353580 31852 353592
rect 27120 353552 31852 353580
rect 27120 353540 27126 353552
rect 31846 353540 31852 353552
rect 31904 353540 31910 353592
rect 40678 353540 40684 353592
rect 40736 353580 40742 353592
rect 51902 353580 51908 353592
rect 40736 353552 51908 353580
rect 40736 353540 40742 353552
rect 51902 353540 51908 353552
rect 51960 353540 51966 353592
rect 24762 353472 24768 353524
rect 24820 353512 24826 353524
rect 28166 353512 28172 353524
rect 24820 353484 28172 353512
rect 24820 353472 24826 353484
rect 28166 353472 28172 353484
rect 28224 353472 28230 353524
rect 31662 353472 31668 353524
rect 31720 353512 31726 353524
rect 37182 353512 37188 353524
rect 31720 353484 37188 353512
rect 31720 353472 31726 353484
rect 37182 353472 37188 353484
rect 37240 353472 37246 353524
rect 50062 353472 50068 353524
rect 50120 353512 50126 353524
rect 62114 353512 62120 353524
rect 50120 353484 62120 353512
rect 50120 353472 50126 353484
rect 62114 353472 62120 353484
rect 62172 353472 62178 353524
rect 22002 353404 22008 353456
rect 22060 353444 22066 353456
rect 23934 353444 23940 353456
rect 22060 353416 23940 353444
rect 22060 353404 22066 353416
rect 23934 353404 23940 353416
rect 23992 353404 23998 353456
rect 24210 353404 24216 353456
rect 24268 353444 24274 353456
rect 27062 353444 27068 353456
rect 24268 353416 27068 353444
rect 24268 353404 24274 353416
rect 27062 353404 27068 353416
rect 27120 353404 27126 353456
rect 31386 353404 31392 353456
rect 31444 353444 31450 353456
rect 37090 353444 37096 353456
rect 31444 353416 37096 353444
rect 31444 353404 31450 353416
rect 37090 353404 37096 353416
rect 37148 353404 37154 353456
rect 21266 353336 21272 353388
rect 21324 353376 21330 353388
rect 22830 353376 22836 353388
rect 21324 353348 22836 353376
rect 21324 353336 21330 353348
rect 22830 353336 22836 353348
rect 22888 353336 22894 353388
rect 23382 353336 23388 353388
rect 23440 353376 23446 353388
rect 26234 353376 26240 353388
rect 23440 353348 26240 353376
rect 23440 353336 23446 353348
rect 26234 353336 26240 353348
rect 26292 353336 26298 353388
rect 28442 353336 28448 353388
rect 28500 353376 28506 353388
rect 33502 353376 33508 353388
rect 28500 353348 33508 353376
rect 28500 353336 28506 353348
rect 33502 353336 33508 353348
rect 33560 353336 33566 353388
rect 36354 353336 36360 353388
rect 36412 353376 36418 353388
rect 41598 353376 41604 353388
rect 36412 353348 41604 353376
rect 36412 353336 36418 353348
rect 41598 353336 41604 353348
rect 41656 353336 41662 353388
rect 20622 353268 20628 353320
rect 20680 353308 20686 353320
rect 22186 353308 22192 353320
rect 20680 353280 22192 353308
rect 20680 353268 20686 353280
rect 22186 353268 22192 353280
rect 22244 353268 22250 353320
rect 22738 353268 22744 353320
rect 22796 353308 22802 353320
rect 25038 353308 25044 353320
rect 22796 353280 25044 353308
rect 22796 353268 22802 353280
rect 25038 353268 25044 353280
rect 25096 353268 25102 353320
rect 27522 353268 27528 353320
rect 27580 353308 27586 353320
rect 32582 353308 32588 353320
rect 27580 353280 32588 353308
rect 27580 353268 27586 353280
rect 32582 353268 32588 353280
rect 32640 353268 32646 353320
rect 37826 353268 37832 353320
rect 37884 353308 37890 353320
rect 42794 353308 42800 353320
rect 37884 353280 42800 353308
rect 37884 353268 37890 353280
rect 42794 353268 42800 353280
rect 42852 353268 42858 353320
rect 54294 353268 54300 353320
rect 54352 353308 54358 353320
rect 57882 353308 57888 353320
rect 54352 353280 57888 353308
rect 54352 353268 54358 353280
rect 57882 353268 57888 353280
rect 57940 353268 57946 353320
rect 57882 352792 57888 352844
rect 57940 352832 57946 352844
rect 72418 352832 72424 352844
rect 57940 352804 72424 352832
rect 57940 352792 57946 352804
rect 72418 352792 72424 352804
rect 72476 352792 72482 352844
rect 57330 352724 57336 352776
rect 57388 352764 57394 352776
rect 76742 352764 76748 352776
rect 57388 352736 76748 352764
rect 57388 352724 57394 352736
rect 76742 352724 76748 352736
rect 76800 352724 76806 352776
rect 60090 352656 60096 352708
rect 60148 352696 60154 352708
rect 80974 352696 80980 352708
rect 60148 352668 80980 352696
rect 60148 352656 60154 352668
rect 80974 352656 80980 352668
rect 81032 352656 81038 352708
rect 62942 352588 62948 352640
rect 63000 352628 63006 352640
rect 85574 352628 85580 352640
rect 63000 352600 85580 352628
rect 63000 352588 63006 352600
rect 85574 352588 85580 352600
rect 85632 352588 85638 352640
rect 65794 352520 65800 352572
rect 65852 352560 65858 352572
rect 89714 352560 89720 352572
rect 65852 352532 89720 352560
rect 65852 352520 65858 352532
rect 89714 352520 89720 352532
rect 89772 352520 89778 352572
rect 37182 351840 37188 351892
rect 37240 351880 37246 351892
rect 39022 351880 39028 351892
rect 37240 351852 39028 351880
rect 37240 351840 37246 351852
rect 39022 351840 39028 351852
rect 39080 351840 39086 351892
rect 56778 351840 56784 351892
rect 56836 351880 56842 351892
rect 58342 351880 58348 351892
rect 56836 351852 58348 351880
rect 56836 351840 56842 351852
rect 58342 351840 58348 351852
rect 58400 351840 58406 351892
rect 62114 351840 62120 351892
rect 62172 351880 62178 351892
rect 66346 351880 66352 351892
rect 62172 351852 66352 351880
rect 62172 351840 62178 351852
rect 66346 351840 66352 351852
rect 66404 351840 66410 351892
rect 68002 351840 68008 351892
rect 68060 351880 68066 351892
rect 92934 351880 92940 351892
rect 68060 351852 92940 351880
rect 68060 351840 68066 351852
rect 92934 351840 92940 351852
rect 92992 351840 92998 351892
rect 198918 351840 198924 351892
rect 198976 351880 198982 351892
rect 200574 351880 200580 351892
rect 198976 351852 200580 351880
rect 198976 351840 198982 351852
rect 200574 351840 200580 351852
rect 200632 351840 200638 351892
rect 274542 351840 274548 351892
rect 274600 351880 274606 351892
rect 276842 351880 276848 351892
rect 274600 351852 276848 351880
rect 274600 351840 274606 351852
rect 276842 351840 276848 351852
rect 276900 351840 276906 351892
rect 58066 351772 58072 351824
rect 58124 351812 58130 351824
rect 60734 351812 60740 351824
rect 58124 351784 60740 351812
rect 58124 351772 58130 351784
rect 60734 351772 60740 351784
rect 60792 351772 60798 351824
rect 68738 351772 68744 351824
rect 68796 351812 68802 351824
rect 94038 351812 94044 351824
rect 68796 351784 94044 351812
rect 68796 351772 68802 351784
rect 94038 351772 94044 351784
rect 94096 351772 94102 351824
rect 275738 351772 275744 351824
rect 275796 351812 275802 351824
rect 278038 351812 278044 351824
rect 275796 351784 278044 351812
rect 275796 351772 275802 351784
rect 278038 351772 278044 351784
rect 278096 351772 278102 351824
rect 59354 351704 59360 351756
rect 59412 351744 59418 351756
rect 62758 351744 62764 351756
rect 59412 351716 62764 351744
rect 59412 351704 59418 351716
rect 62758 351704 62764 351716
rect 62816 351704 62822 351756
rect 70118 351704 70124 351756
rect 70176 351744 70182 351756
rect 96062 351744 96068 351756
rect 70176 351716 96068 351744
rect 70176 351704 70182 351716
rect 96062 351704 96068 351716
rect 96120 351704 96126 351756
rect 276658 351704 276664 351756
rect 276716 351744 276722 351756
rect 279326 351744 279332 351756
rect 276716 351716 279332 351744
rect 276716 351704 276722 351716
rect 279326 351704 279332 351716
rect 279384 351704 279390 351756
rect 42794 351636 42800 351688
rect 42852 351676 42858 351688
rect 47670 351676 47676 351688
rect 42852 351648 47676 351676
rect 42852 351636 42858 351648
rect 47670 351636 47676 351648
rect 47728 351636 47734 351688
rect 62206 351636 62212 351688
rect 62264 351676 62270 351688
rect 66990 351676 66996 351688
rect 62264 351648 66996 351676
rect 62264 351636 62270 351648
rect 66990 351636 66996 351648
rect 67048 351636 67054 351688
rect 70854 351636 70860 351688
rect 70912 351676 70918 351688
rect 97166 351676 97172 351688
rect 70912 351648 97172 351676
rect 70912 351636 70918 351648
rect 97166 351636 97172 351648
rect 97224 351636 97230 351688
rect 277762 351636 277768 351688
rect 277820 351676 277826 351688
rect 278774 351676 278780 351688
rect 277820 351648 278780 351676
rect 277820 351636 277826 351648
rect 278774 351636 278780 351648
rect 278832 351636 278838 351688
rect 58526 351568 58532 351620
rect 58584 351608 58590 351620
rect 61654 351608 61660 351620
rect 58584 351580 61660 351608
rect 58584 351568 58590 351580
rect 61654 351568 61660 351580
rect 61712 351568 61718 351620
rect 69382 351568 69388 351620
rect 69440 351608 69446 351620
rect 95234 351608 95240 351620
rect 69440 351580 95240 351608
rect 69440 351568 69446 351580
rect 95234 351568 95240 351580
rect 95292 351568 95298 351620
rect 278682 351568 278688 351620
rect 278740 351608 278746 351620
rect 281718 351608 281724 351620
rect 278740 351580 281724 351608
rect 278740 351568 278746 351580
rect 281718 351568 281724 351580
rect 281776 351568 281782 351620
rect 59630 351500 59636 351552
rect 59688 351540 59694 351552
rect 63678 351540 63684 351552
rect 59688 351512 63684 351540
rect 59688 351500 59694 351512
rect 63678 351500 63684 351512
rect 63736 351500 63742 351552
rect 73706 351500 73712 351552
rect 73764 351540 73770 351552
rect 101398 351540 101404 351552
rect 73764 351512 101404 351540
rect 73764 351500 73770 351512
rect 101398 351500 101404 351512
rect 101456 351500 101462 351552
rect 271322 351500 271328 351552
rect 271380 351540 271386 351552
rect 273346 351540 273352 351552
rect 271380 351512 273352 351540
rect 271380 351500 271386 351512
rect 273346 351500 273352 351512
rect 273404 351500 273410 351552
rect 57514 351432 57520 351484
rect 57572 351472 57578 351484
rect 59446 351472 59452 351484
rect 57572 351444 59452 351472
rect 57572 351432 57578 351444
rect 59446 351432 59452 351444
rect 59504 351432 59510 351484
rect 71590 351432 71596 351484
rect 71648 351472 71654 351484
rect 98270 351472 98276 351484
rect 71648 351444 98276 351472
rect 71648 351432 71654 351444
rect 98270 351432 98276 351444
rect 98328 351432 98334 351484
rect 114002 351432 114008 351484
rect 114060 351472 114066 351484
rect 114462 351472 114468 351484
rect 114060 351444 114468 351472
rect 114060 351432 114066 351444
rect 114462 351432 114468 351444
rect 114520 351432 114526 351484
rect 115106 351432 115112 351484
rect 115164 351472 115170 351484
rect 115750 351472 115756 351484
rect 115164 351444 115756 351472
rect 115164 351432 115170 351444
rect 115750 351432 115756 351444
rect 115808 351432 115814 351484
rect 118142 351432 118148 351484
rect 118200 351472 118206 351484
rect 118602 351472 118608 351484
rect 118200 351444 118608 351472
rect 118200 351432 118206 351444
rect 118602 351432 118608 351444
rect 118660 351432 118666 351484
rect 133322 351432 133328 351484
rect 133380 351472 133386 351484
rect 133782 351472 133788 351484
rect 133380 351444 133788 351472
rect 133380 351432 133386 351444
rect 133782 351432 133788 351444
rect 133840 351432 133846 351484
rect 138842 351432 138848 351484
rect 138900 351472 138906 351484
rect 139302 351472 139308 351484
rect 138900 351444 139308 351472
rect 138900 351432 138906 351444
rect 139302 351432 139308 351444
rect 139360 351432 139366 351484
rect 143074 351432 143080 351484
rect 143132 351472 143138 351484
rect 143442 351472 143448 351484
rect 143132 351444 143448 351472
rect 143132 351432 143138 351444
rect 143442 351432 143448 351444
rect 143500 351432 143506 351484
rect 145282 351432 145288 351484
rect 145340 351472 145346 351484
rect 146110 351472 146116 351484
rect 145340 351444 146116 351472
rect 145340 351432 145346 351444
rect 146110 351432 146116 351444
rect 146168 351432 146174 351484
rect 155954 351432 155960 351484
rect 156012 351472 156018 351484
rect 156414 351472 156420 351484
rect 156012 351444 156420 351472
rect 156012 351432 156018 351444
rect 156414 351432 156420 351444
rect 156472 351432 156478 351484
rect 160094 351432 160100 351484
rect 160152 351472 160158 351484
rect 160830 351472 160836 351484
rect 160152 351444 160836 351472
rect 160152 351432 160158 351444
rect 160830 351432 160836 351444
rect 160888 351432 160894 351484
rect 161474 351432 161480 351484
rect 161532 351472 161538 351484
rect 161934 351472 161940 351484
rect 161532 351444 161940 351472
rect 161532 351432 161538 351444
rect 161934 351432 161940 351444
rect 161992 351432 161998 351484
rect 165614 351432 165620 351484
rect 165672 351472 165678 351484
rect 166166 351472 166172 351484
rect 165672 351444 166172 351472
rect 165672 351432 165678 351444
rect 166166 351432 166172 351444
rect 166224 351432 166230 351484
rect 169846 351432 169852 351484
rect 169904 351472 169910 351484
rect 170398 351472 170404 351484
rect 169904 351444 170404 351472
rect 169904 351432 169910 351444
rect 170398 351432 170404 351444
rect 170456 351432 170462 351484
rect 171134 351432 171140 351484
rect 171192 351472 171198 351484
rect 171594 351472 171600 351484
rect 171192 351444 171600 351472
rect 171192 351432 171198 351444
rect 171594 351432 171600 351444
rect 171652 351432 171658 351484
rect 175274 351432 175280 351484
rect 175332 351472 175338 351484
rect 175918 351472 175924 351484
rect 175332 351444 175924 351472
rect 175332 351432 175338 351444
rect 175918 351432 175924 351444
rect 175976 351432 175982 351484
rect 176654 351432 176660 351484
rect 176712 351472 176718 351484
rect 177114 351472 177120 351484
rect 176712 351444 177120 351472
rect 176712 351432 176718 351444
rect 177114 351432 177120 351444
rect 177172 351432 177178 351484
rect 179598 351432 179604 351484
rect 179656 351472 179662 351484
rect 180150 351472 180156 351484
rect 179656 351444 180156 351472
rect 179656 351432 179662 351444
rect 180150 351432 180156 351444
rect 180208 351432 180214 351484
rect 180794 351432 180800 351484
rect 180852 351472 180858 351484
rect 181254 351472 181260 351484
rect 180852 351444 181260 351472
rect 180852 351432 180858 351444
rect 181254 351432 181260 351444
rect 181312 351432 181318 351484
rect 184934 351432 184940 351484
rect 184992 351472 184998 351484
rect 185486 351472 185492 351484
rect 184992 351444 185492 351472
rect 184992 351432 184998 351444
rect 185486 351432 185492 351444
rect 185544 351432 185550 351484
rect 193674 351432 193680 351484
rect 193732 351472 193738 351484
rect 196342 351472 196348 351484
rect 193732 351444 196348 351472
rect 193732 351432 193738 351444
rect 196342 351432 196348 351444
rect 196400 351432 196406 351484
rect 269022 351432 269028 351484
rect 269080 351472 269086 351484
rect 270494 351472 270500 351484
rect 269080 351444 270500 351472
rect 269080 351432 269086 351444
rect 270494 351432 270500 351444
rect 270552 351432 270558 351484
rect 273070 351432 273076 351484
rect 273128 351472 273134 351484
rect 275646 351472 275652 351484
rect 273128 351444 275652 351472
rect 273128 351432 273134 351444
rect 275646 351432 275652 351444
rect 275704 351432 275710 351484
rect 40034 351364 40040 351416
rect 40092 351404 40098 351416
rect 43254 351404 43260 351416
rect 40092 351376 43260 351404
rect 40092 351364 40098 351376
rect 43254 351364 43260 351376
rect 43312 351364 43318 351416
rect 63494 351364 63500 351416
rect 63552 351404 63558 351416
rect 68094 351404 68100 351416
rect 63552 351376 68100 351404
rect 63552 351364 63558 351376
rect 68094 351364 68100 351376
rect 68152 351364 68158 351416
rect 72326 351364 72332 351416
rect 72384 351404 72390 351416
rect 99374 351404 99380 351416
rect 72384 351376 99380 351404
rect 72384 351364 72390 351376
rect 99374 351364 99380 351376
rect 99432 351364 99438 351416
rect 130194 351364 130200 351416
rect 130252 351404 130258 351416
rect 153286 351404 153292 351416
rect 130252 351376 153292 351404
rect 130252 351364 130258 351376
rect 153286 351364 153292 351376
rect 153344 351364 153350 351416
rect 193858 351364 193864 351416
rect 193916 351404 193922 351416
rect 197446 351404 197452 351416
rect 193916 351376 197452 351404
rect 193916 351364 193922 351376
rect 197446 351364 197452 351376
rect 197504 351364 197510 351416
rect 270218 351364 270224 351416
rect 270276 351404 270282 351416
rect 271874 351404 271880 351416
rect 270276 351376 271880 351404
rect 270276 351364 270282 351376
rect 271874 351364 271880 351376
rect 271932 351364 271938 351416
rect 39206 351296 39212 351348
rect 39264 351336 39270 351348
rect 42150 351336 42156 351348
rect 39264 351308 42156 351336
rect 39264 351296 39270 351308
rect 42150 351296 42156 351308
rect 42208 351296 42214 351348
rect 42242 351296 42248 351348
rect 42300 351336 42306 351348
rect 46566 351336 46572 351348
rect 42300 351308 46572 351336
rect 42300 351296 42306 351308
rect 46566 351296 46572 351308
rect 46624 351296 46630 351348
rect 52178 351296 52184 351348
rect 52236 351336 52242 351348
rect 69198 351336 69204 351348
rect 52236 351308 69204 351336
rect 52236 351296 52242 351308
rect 69198 351296 69204 351308
rect 69256 351296 69262 351348
rect 72970 351296 72976 351348
rect 73028 351336 73034 351348
rect 100846 351336 100852 351348
rect 73028 351308 100852 351336
rect 73028 351296 73034 351308
rect 100846 351296 100852 351308
rect 100904 351296 100910 351348
rect 131022 351296 131028 351348
rect 131080 351336 131086 351348
rect 154758 351336 154764 351348
rect 131080 351308 154764 351336
rect 131080 351296 131086 351308
rect 154758 351296 154764 351308
rect 154816 351296 154822 351348
rect 40218 351228 40224 351280
rect 40276 351268 40282 351280
rect 44358 351268 44364 351280
rect 40276 351240 44364 351268
rect 40276 351228 40282 351240
rect 44358 351228 44364 351240
rect 44416 351228 44422 351280
rect 53650 351228 53656 351280
rect 53708 351268 53714 351280
rect 71222 351268 71228 351280
rect 53708 351240 71228 351268
rect 53708 351228 53714 351240
rect 71222 351228 71228 351240
rect 71280 351228 71286 351280
rect 75178 351228 75184 351280
rect 75236 351268 75242 351280
rect 103698 351268 103704 351280
rect 75236 351240 103704 351268
rect 75236 351228 75242 351240
rect 103698 351228 103704 351240
rect 103756 351228 103762 351280
rect 125410 351228 125416 351280
rect 125468 351268 125474 351280
rect 153378 351268 153384 351280
rect 125468 351240 153384 351268
rect 125468 351228 125474 351240
rect 153378 351228 153384 351240
rect 153436 351228 153442 351280
rect 226978 351228 226984 351280
rect 227036 351268 227042 351280
rect 228726 351268 228732 351280
rect 227036 351240 228732 351268
rect 227036 351228 227042 351240
rect 228726 351228 228732 351240
rect 228784 351228 228790 351280
rect 38654 351160 38660 351212
rect 38712 351200 38718 351212
rect 41506 351200 41512 351212
rect 38712 351172 41512 351200
rect 38712 351160 38718 351172
rect 41506 351160 41512 351172
rect 41564 351160 41570 351212
rect 41598 351160 41604 351212
rect 41656 351200 41662 351212
rect 45646 351200 45652 351212
rect 41656 351172 45652 351200
rect 41656 351160 41662 351172
rect 45646 351160 45652 351172
rect 45704 351160 45710 351212
rect 55030 351160 55036 351212
rect 55088 351200 55094 351212
rect 73430 351200 73436 351212
rect 55088 351172 73436 351200
rect 55088 351160 55094 351172
rect 73430 351160 73436 351172
rect 73488 351160 73494 351212
rect 74442 351160 74448 351212
rect 74500 351200 74506 351212
rect 102502 351200 102508 351212
rect 74500 351172 102508 351200
rect 74500 351160 74506 351172
rect 102502 351160 102508 351172
rect 102560 351160 102566 351212
rect 123754 351160 123760 351212
rect 123812 351200 123818 351212
rect 153470 351200 153476 351212
rect 123812 351172 153476 351200
rect 123812 351160 123818 351172
rect 153470 351160 153476 351172
rect 153528 351160 153534 351212
rect 228818 351160 228824 351212
rect 228876 351200 228882 351212
rect 229830 351200 229836 351212
rect 228876 351172 229836 351200
rect 228876 351160 228882 351172
rect 229830 351160 229836 351172
rect 229888 351160 229894 351212
rect 38194 351092 38200 351144
rect 38252 351132 38258 351144
rect 40126 351132 40132 351144
rect 38252 351104 40132 351132
rect 38252 351092 38258 351104
rect 40126 351092 40132 351104
rect 40184 351092 40190 351144
rect 64782 351092 64788 351144
rect 64840 351132 64846 351144
rect 88518 351132 88524 351144
rect 64840 351104 88524 351132
rect 64840 351092 64846 351104
rect 88518 351092 88524 351104
rect 88576 351092 88582 351144
rect 66162 351024 66168 351076
rect 66220 351064 66226 351076
rect 90726 351064 90732 351076
rect 66220 351036 90732 351064
rect 66220 351024 66226 351036
rect 90726 351024 90732 351036
rect 90784 351024 90790 351076
rect 183830 351024 183836 351076
rect 183888 351064 183894 351076
rect 184566 351064 184572 351076
rect 183888 351036 184572 351064
rect 183888 351024 183894 351036
rect 184566 351024 184572 351036
rect 184624 351024 184630 351076
rect 67266 350956 67272 351008
rect 67324 350996 67330 351008
rect 91830 350996 91836 351008
rect 67324 350968 91836 350996
rect 67324 350956 67330 350968
rect 91830 350956 91836 350968
rect 91888 350956 91894 351008
rect 110690 350956 110696 351008
rect 110748 350996 110754 351008
rect 111702 350996 111708 351008
rect 110748 350968 111708 350996
rect 110748 350956 110754 350968
rect 111702 350956 111708 350968
rect 111760 350956 111766 351008
rect 173894 350956 173900 351008
rect 173952 350996 173958 351008
rect 174814 350996 174820 351008
rect 173952 350968 174820 350996
rect 173952 350956 173958 350968
rect 174814 350956 174820 350968
rect 174872 350956 174878 351008
rect 230474 350956 230480 351008
rect 230532 350996 230538 351008
rect 231854 350996 231860 351008
rect 230532 350968 231860 350996
rect 230532 350956 230538 350968
rect 231854 350956 231860 350968
rect 231912 350956 231918 351008
rect 62022 350888 62028 350940
rect 62080 350928 62086 350940
rect 84378 350928 84384 350940
rect 62080 350900 84384 350928
rect 62080 350888 62086 350900
rect 84378 350888 84384 350900
rect 84436 350888 84442 350940
rect 135530 350888 135536 350940
rect 135588 350928 135594 350940
rect 136450 350928 136456 350940
rect 135588 350900 136456 350928
rect 135588 350888 135594 350900
rect 136450 350888 136456 350900
rect 136508 350888 136514 350940
rect 201494 350888 201500 350940
rect 201552 350928 201558 350940
rect 202874 350928 202880 350940
rect 201552 350900 202880 350928
rect 201552 350888 201558 350900
rect 202874 350888 202880 350900
rect 202932 350888 202938 350940
rect 233694 350888 233700 350940
rect 233752 350928 233758 350940
rect 235166 350928 235172 350940
rect 233752 350900 235172 350928
rect 233752 350888 233758 350900
rect 235166 350888 235172 350900
rect 235224 350888 235230 350940
rect 272426 350888 272432 350940
rect 272484 350928 272490 350940
rect 274634 350928 274640 350940
rect 272484 350900 274640 350928
rect 272484 350888 272490 350900
rect 274634 350888 274640 350900
rect 274692 350888 274698 350940
rect 63402 350820 63408 350872
rect 63460 350860 63466 350872
rect 86310 350860 86316 350872
rect 63460 350832 86316 350860
rect 63460 350820 63466 350832
rect 86310 350820 86316 350832
rect 86368 350820 86374 350872
rect 120442 350820 120448 350872
rect 120500 350860 120506 350872
rect 121362 350860 121368 350872
rect 120500 350832 121368 350860
rect 120500 350820 120506 350832
rect 121362 350820 121368 350832
rect 121420 350820 121426 350872
rect 158714 350820 158720 350872
rect 158772 350860 158778 350872
rect 159726 350860 159732 350872
rect 158772 350832 159732 350860
rect 158772 350820 158778 350832
rect 159726 350820 159732 350832
rect 159784 350820 159790 350872
rect 34514 350752 34520 350804
rect 34572 350792 34578 350804
rect 36814 350792 36820 350804
rect 34572 350764 36820 350792
rect 34572 350752 34578 350764
rect 36814 350752 36820 350764
rect 36872 350752 36878 350804
rect 37090 350752 37096 350804
rect 37148 350792 37154 350804
rect 37918 350792 37924 350804
rect 37148 350764 37924 350792
rect 37148 350752 37154 350764
rect 37918 350752 37924 350764
rect 37976 350752 37982 350804
rect 60642 350752 60648 350804
rect 60700 350792 60706 350804
rect 82078 350792 82084 350804
rect 60700 350764 82084 350792
rect 60700 350752 60706 350764
rect 82078 350752 82084 350764
rect 82136 350752 82142 350804
rect 134426 350752 134432 350804
rect 134484 350792 134490 350804
rect 135162 350792 135168 350804
rect 134484 350764 135168 350792
rect 134484 350752 134490 350764
rect 135162 350752 135168 350764
rect 135220 350752 135226 350804
rect 139762 350752 139768 350804
rect 139820 350792 139826 350804
rect 140682 350792 140688 350804
rect 139820 350764 140688 350792
rect 139820 350752 139826 350764
rect 140682 350752 140688 350764
rect 140740 350752 140746 350804
rect 223206 350752 223212 350804
rect 223264 350792 223270 350804
rect 224310 350792 224316 350804
rect 223264 350764 224316 350792
rect 223264 350752 223270 350764
rect 224310 350752 224316 350764
rect 224368 350752 224374 350804
rect 59262 350684 59268 350736
rect 59320 350724 59326 350736
rect 80054 350724 80060 350736
rect 59320 350696 80060 350724
rect 59320 350684 59326 350696
rect 80054 350684 80060 350696
rect 80112 350684 80118 350736
rect 57790 350616 57796 350668
rect 57848 350656 57854 350668
rect 77846 350656 77852 350668
rect 57848 350628 77852 350656
rect 57848 350616 57854 350628
rect 77846 350616 77852 350628
rect 77904 350616 77910 350668
rect 144178 350616 144184 350668
rect 144236 350656 144242 350668
rect 144822 350656 144828 350668
rect 144236 350628 144828 350656
rect 144236 350616 144242 350628
rect 144822 350616 144828 350628
rect 144880 350616 144886 350668
rect 164234 350616 164240 350668
rect 164292 350656 164298 350668
rect 165062 350656 165068 350668
rect 164292 350628 165068 350656
rect 164292 350616 164298 350628
rect 165062 350616 165068 350628
rect 165120 350616 165126 350668
rect 56502 350548 56508 350600
rect 56560 350588 56566 350600
rect 76006 350588 76012 350600
rect 56560 350560 76012 350588
rect 56560 350548 56566 350560
rect 76006 350548 76012 350560
rect 76064 350548 76070 350600
rect 282362 347800 282368 347812
rect 282323 347772 282368 347800
rect 282362 347760 282368 347772
rect 282420 347760 282426 347812
rect 3142 336744 3148 336796
rect 3200 336784 3206 336796
rect 6178 336784 6184 336796
rect 3200 336756 6184 336784
rect 3200 336744 3206 336756
rect 6178 336744 6184 336756
rect 6236 336744 6242 336796
rect 303614 327020 303620 327072
rect 303672 327060 303678 327072
rect 577590 327060 577596 327072
rect 303672 327032 577596 327060
rect 303672 327020 303678 327032
rect 577590 327020 577596 327032
rect 577648 327020 577654 327072
rect 303614 325592 303620 325644
rect 303672 325632 303678 325644
rect 563698 325632 563704 325644
rect 303672 325604 563704 325632
rect 303672 325592 303678 325604
rect 563698 325592 563704 325604
rect 563756 325592 563762 325644
rect 21358 322736 21364 322788
rect 21416 322776 21422 322788
rect 22186 322776 22192 322788
rect 21416 322748 22192 322776
rect 21416 322736 21422 322748
rect 22186 322736 22192 322748
rect 22244 322736 22250 322788
rect 303614 321580 303620 321632
rect 303672 321620 303678 321632
rect 580166 321620 580172 321632
rect 303672 321592 580172 321620
rect 303672 321580 303678 321592
rect 580166 321580 580172 321592
rect 580224 321580 580230 321632
rect 100754 321240 100760 321292
rect 100812 321280 100818 321292
rect 106274 321280 106280 321292
rect 100812 321252 106280 321280
rect 100812 321240 100818 321252
rect 106274 321240 106280 321252
rect 106332 321240 106338 321292
rect 231762 321172 231768 321224
rect 231820 321212 231826 321224
rect 235442 321212 235448 321224
rect 231820 321184 235448 321212
rect 231820 321172 231826 321184
rect 235442 321172 235448 321184
rect 235500 321172 235506 321224
rect 108298 321104 108304 321156
rect 108356 321144 108362 321156
rect 115198 321144 115204 321156
rect 108356 321116 115204 321144
rect 108356 321104 108362 321116
rect 115198 321104 115204 321116
rect 115256 321104 115262 321156
rect 92106 321036 92112 321088
rect 92164 321076 92170 321088
rect 96614 321076 96620 321088
rect 92164 321048 96620 321076
rect 92164 321036 92170 321048
rect 96614 321036 96620 321048
rect 96672 321036 96678 321088
rect 111518 321036 111524 321088
rect 111576 321076 111582 321088
rect 117958 321076 117964 321088
rect 111576 321048 117964 321076
rect 111576 321036 111582 321048
rect 117958 321036 117964 321048
rect 118016 321036 118022 321088
rect 101766 320968 101772 321020
rect 101824 321008 101830 321020
rect 106366 321008 106372 321020
rect 101824 320980 106372 321008
rect 101824 320968 101830 320980
rect 106366 320968 106372 320980
rect 106424 320968 106430 321020
rect 109310 320968 109316 321020
rect 109368 321008 109374 321020
rect 119338 321008 119344 321020
rect 109368 320980 119344 321008
rect 109368 320968 109374 320980
rect 119338 320968 119344 320980
rect 119396 320968 119402 321020
rect 228266 320968 228272 321020
rect 228324 321008 228330 321020
rect 232222 321008 232228 321020
rect 228324 320980 232228 321008
rect 228324 320968 228330 320980
rect 232222 320968 232228 320980
rect 232280 320968 232286 321020
rect 22094 320900 22100 320952
rect 22152 320940 22158 320952
rect 22152 320912 31064 320940
rect 22152 320900 22158 320912
rect 24762 320832 24768 320884
rect 24820 320872 24826 320884
rect 26326 320872 26332 320884
rect 24820 320844 26332 320872
rect 24820 320832 24826 320844
rect 26326 320832 26332 320844
rect 26384 320832 26390 320884
rect 31036 320872 31064 320912
rect 75914 320900 75920 320952
rect 75972 320940 75978 320952
rect 78674 320940 78680 320952
rect 75972 320912 78680 320940
rect 75972 320900 75978 320912
rect 78674 320900 78680 320912
rect 78732 320900 78738 320952
rect 102870 320900 102876 320952
rect 102928 320940 102934 320952
rect 108942 320940 108948 320952
rect 102928 320912 108948 320940
rect 102928 320900 102934 320912
rect 108942 320900 108948 320912
rect 109000 320900 109006 320952
rect 42886 320872 42892 320884
rect 31036 320844 42892 320872
rect 42886 320832 42892 320844
rect 42944 320832 42950 320884
rect 64046 320832 64052 320884
rect 64104 320872 64110 320884
rect 64874 320872 64880 320884
rect 64104 320844 64880 320872
rect 64104 320832 64110 320844
rect 64874 320832 64880 320844
rect 64932 320832 64938 320884
rect 72694 320832 72700 320884
rect 72752 320872 72758 320884
rect 74534 320872 74540 320884
rect 72752 320844 74540 320872
rect 72752 320832 72758 320844
rect 74534 320832 74540 320844
rect 74592 320832 74598 320884
rect 82446 320832 82452 320884
rect 82504 320872 82510 320884
rect 85114 320872 85120 320884
rect 82504 320844 85120 320872
rect 82504 320832 82510 320844
rect 85114 320832 85120 320844
rect 85172 320832 85178 320884
rect 93210 320832 93216 320884
rect 93268 320872 93274 320884
rect 97994 320872 98000 320884
rect 93268 320844 98000 320872
rect 93268 320832 93274 320844
rect 97994 320832 98000 320844
rect 98052 320832 98058 320884
rect 106090 320832 106096 320884
rect 106148 320872 106154 320884
rect 121546 320872 121552 320884
rect 106148 320844 121552 320872
rect 106148 320832 106154 320844
rect 121546 320832 121552 320844
rect 121604 320832 121610 320884
rect 207661 320875 207719 320881
rect 207661 320841 207673 320875
rect 207707 320872 207719 320875
rect 279510 320872 279516 320884
rect 207707 320844 279516 320872
rect 207707 320841 207719 320844
rect 207661 320835 207719 320841
rect 279510 320832 279516 320844
rect 279568 320832 279574 320884
rect 73798 320764 73804 320816
rect 73856 320804 73862 320816
rect 75914 320804 75920 320816
rect 73856 320776 75920 320804
rect 73856 320764 73862 320776
rect 75914 320764 75920 320776
rect 75972 320764 75978 320816
rect 83458 320764 83464 320816
rect 83516 320804 83522 320816
rect 85758 320804 85764 320816
rect 83516 320776 85764 320804
rect 83516 320764 83522 320776
rect 85758 320764 85764 320776
rect 85816 320764 85822 320816
rect 91002 320764 91008 320816
rect 91060 320804 91066 320816
rect 95234 320804 95240 320816
rect 91060 320776 95240 320804
rect 91060 320764 91066 320776
rect 95234 320764 95240 320776
rect 95292 320764 95298 320816
rect 195606 320764 195612 320816
rect 195664 320804 195670 320816
rect 202877 320807 202935 320813
rect 202877 320804 202889 320807
rect 195664 320776 202889 320804
rect 195664 320764 195670 320776
rect 202877 320773 202889 320776
rect 202923 320773 202935 320807
rect 202877 320767 202935 320773
rect 227070 320764 227076 320816
rect 227128 320804 227134 320816
rect 231118 320804 231124 320816
rect 227128 320776 231124 320804
rect 227128 320764 227134 320776
rect 231118 320764 231124 320776
rect 231176 320764 231182 320816
rect 248230 320764 248236 320816
rect 248288 320804 248294 320816
rect 250530 320804 250536 320816
rect 248288 320776 250536 320804
rect 248288 320764 248294 320776
rect 250530 320764 250536 320776
rect 250588 320764 250594 320816
rect 256602 320764 256608 320816
rect 256660 320804 256666 320816
rect 258074 320804 258080 320816
rect 256660 320776 258080 320804
rect 256660 320764 256666 320776
rect 258074 320764 258080 320776
rect 258132 320764 258138 320816
rect 202877 320671 202935 320677
rect 202877 320637 202889 320671
rect 202923 320668 202935 320671
rect 207661 320671 207719 320677
rect 207661 320668 207673 320671
rect 202923 320640 207673 320668
rect 202923 320637 202935 320640
rect 202877 320631 202935 320637
rect 207661 320637 207673 320640
rect 207707 320637 207719 320671
rect 207661 320631 207719 320637
rect 226242 320628 226248 320680
rect 226300 320668 226306 320680
rect 230106 320668 230112 320680
rect 226300 320640 230112 320668
rect 226300 320628 226306 320640
rect 230106 320628 230112 320640
rect 230164 320628 230170 320680
rect 204254 320560 204260 320612
rect 204312 320600 204318 320612
rect 206370 320600 206376 320612
rect 204312 320572 206376 320600
rect 204312 320560 204318 320572
rect 206370 320560 206376 320572
rect 206428 320560 206434 320612
rect 208394 320560 208400 320612
rect 208452 320600 208458 320612
rect 210694 320600 210700 320612
rect 208452 320572 210700 320600
rect 208452 320560 208458 320572
rect 210694 320560 210700 320572
rect 210752 320560 210758 320612
rect 110414 320492 110420 320544
rect 110472 320532 110478 320544
rect 113818 320532 113824 320544
rect 110472 320504 113824 320532
rect 110472 320492 110478 320504
rect 113818 320492 113824 320504
rect 113876 320492 113882 320544
rect 23382 320424 23388 320476
rect 23440 320464 23446 320476
rect 25314 320464 25320 320476
rect 23440 320436 25320 320464
rect 23440 320424 23446 320436
rect 25314 320424 25320 320436
rect 25372 320424 25378 320476
rect 88886 320424 88892 320476
rect 88944 320464 88950 320476
rect 91278 320464 91284 320476
rect 88944 320436 91284 320464
rect 88944 320424 88950 320436
rect 91278 320424 91284 320436
rect 91336 320424 91342 320476
rect 94222 320424 94228 320476
rect 94280 320464 94286 320476
rect 99466 320464 99472 320476
rect 94280 320436 99472 320464
rect 94280 320424 94286 320436
rect 99466 320424 99472 320436
rect 99524 320424 99530 320476
rect 99650 320424 99656 320476
rect 99708 320464 99714 320476
rect 104894 320464 104900 320476
rect 99708 320436 104900 320464
rect 99708 320424 99714 320436
rect 104894 320424 104900 320436
rect 104952 320424 104958 320476
rect 235442 320424 235448 320476
rect 235500 320464 235506 320476
rect 238662 320464 238668 320476
rect 235500 320436 238668 320464
rect 235500 320424 235506 320436
rect 238662 320424 238668 320436
rect 238720 320424 238726 320476
rect 246114 320424 246120 320476
rect 246172 320464 246178 320476
rect 248414 320464 248420 320476
rect 246172 320436 248420 320464
rect 246172 320424 246178 320436
rect 248414 320424 248420 320436
rect 248472 320424 248478 320476
rect 78122 320356 78128 320408
rect 78180 320396 78186 320408
rect 81250 320396 81256 320408
rect 78180 320368 81256 320396
rect 78180 320356 78186 320368
rect 81250 320356 81256 320368
rect 81308 320356 81314 320408
rect 87782 320356 87788 320408
rect 87840 320396 87846 320408
rect 90082 320396 90088 320408
rect 87840 320368 90088 320396
rect 87840 320356 87846 320368
rect 90082 320356 90088 320368
rect 90140 320356 90146 320408
rect 97534 320356 97540 320408
rect 97592 320396 97598 320408
rect 102134 320396 102140 320408
rect 97592 320368 102140 320396
rect 97592 320356 97598 320368
rect 102134 320356 102140 320368
rect 102192 320356 102198 320408
rect 200114 320356 200120 320408
rect 200172 320396 200178 320408
rect 203150 320396 203156 320408
rect 200172 320368 203156 320396
rect 200172 320356 200178 320368
rect 203150 320356 203156 320368
rect 203208 320356 203214 320408
rect 236638 320356 236644 320408
rect 236696 320396 236702 320408
rect 239766 320396 239772 320408
rect 236696 320368 239772 320396
rect 236696 320356 236702 320368
rect 239766 320356 239772 320368
rect 239824 320356 239830 320408
rect 25314 320288 25320 320340
rect 25372 320328 25378 320340
rect 27430 320328 27436 320340
rect 25372 320300 27436 320328
rect 25372 320288 25378 320300
rect 27430 320288 27436 320300
rect 27488 320288 27494 320340
rect 54386 320288 54392 320340
rect 54444 320328 54450 320340
rect 55214 320328 55220 320340
rect 54444 320300 55220 320328
rect 54444 320288 54450 320300
rect 55214 320288 55220 320300
rect 55272 320288 55278 320340
rect 66254 320288 66260 320340
rect 66312 320328 66318 320340
rect 67634 320328 67640 320340
rect 66312 320300 67640 320328
rect 66312 320288 66318 320300
rect 67634 320288 67640 320300
rect 67692 320288 67698 320340
rect 69474 320288 69480 320340
rect 69532 320328 69538 320340
rect 71774 320328 71780 320340
rect 69532 320300 71780 320328
rect 69532 320288 69538 320300
rect 71774 320288 71780 320300
rect 71832 320288 71838 320340
rect 80238 320288 80244 320340
rect 80296 320328 80302 320340
rect 82814 320328 82820 320340
rect 80296 320300 82820 320328
rect 80296 320288 80302 320300
rect 82814 320288 82820 320300
rect 82872 320288 82878 320340
rect 86678 320288 86684 320340
rect 86736 320328 86742 320340
rect 91094 320328 91100 320340
rect 86736 320300 91100 320328
rect 86736 320288 86742 320300
rect 91094 320288 91100 320300
rect 91152 320288 91158 320340
rect 98546 320288 98552 320340
rect 98604 320328 98610 320340
rect 103514 320328 103520 320340
rect 98604 320300 103520 320328
rect 98604 320288 98610 320300
rect 103514 320288 103520 320300
rect 103572 320288 103578 320340
rect 103974 320288 103980 320340
rect 104032 320328 104038 320340
rect 109770 320328 109776 320340
rect 104032 320300 109776 320328
rect 104032 320288 104038 320300
rect 109770 320288 109776 320300
rect 109828 320288 109834 320340
rect 198734 320288 198740 320340
rect 198792 320328 198798 320340
rect 200942 320328 200948 320340
rect 198792 320300 200948 320328
rect 198792 320288 198798 320300
rect 200942 320288 200948 320300
rect 201000 320288 201006 320340
rect 229462 320288 229468 320340
rect 229520 320328 229526 320340
rect 233326 320328 233332 320340
rect 229520 320300 233332 320328
rect 229520 320288 229526 320300
rect 233326 320288 233332 320300
rect 233384 320288 233390 320340
rect 238662 320288 238668 320340
rect 238720 320328 238726 320340
rect 241882 320328 241888 320340
rect 238720 320300 241888 320328
rect 238720 320288 238726 320300
rect 241882 320288 241888 320300
rect 241940 320288 241946 320340
rect 242618 320288 242624 320340
rect 242676 320328 242682 320340
rect 245194 320328 245200 320340
rect 242676 320300 245200 320328
rect 242676 320288 242682 320300
rect 245194 320288 245200 320300
rect 245252 320288 245258 320340
rect 253382 320288 253388 320340
rect 253440 320328 253446 320340
rect 254854 320328 254860 320340
rect 253440 320300 254860 320328
rect 253440 320288 253446 320300
rect 254854 320288 254860 320300
rect 254912 320288 254918 320340
rect 27706 320220 27712 320272
rect 27764 320260 27770 320272
rect 29638 320260 29644 320272
rect 27764 320232 29644 320260
rect 27764 320220 27770 320232
rect 29638 320220 29644 320232
rect 29696 320220 29702 320272
rect 30282 320220 30288 320272
rect 30340 320260 30346 320272
rect 31754 320260 31760 320272
rect 30340 320232 31760 320260
rect 30340 320220 30346 320232
rect 31754 320220 31760 320232
rect 31812 320220 31818 320272
rect 33686 320220 33692 320272
rect 33744 320260 33750 320272
rect 34974 320260 34980 320272
rect 33744 320232 34980 320260
rect 33744 320220 33750 320232
rect 34974 320220 34980 320232
rect 35032 320220 35038 320272
rect 61930 320220 61936 320272
rect 61988 320260 61994 320272
rect 63494 320260 63500 320272
rect 61988 320232 63500 320260
rect 61988 320220 61994 320232
rect 63494 320220 63500 320232
rect 63552 320220 63558 320272
rect 68370 320220 68376 320272
rect 68428 320260 68434 320272
rect 70394 320260 70400 320272
rect 68428 320232 70400 320260
rect 68428 320220 68434 320232
rect 70394 320220 70400 320232
rect 70452 320220 70458 320272
rect 70578 320220 70584 320272
rect 70636 320260 70642 320272
rect 73154 320260 73160 320272
rect 70636 320232 73160 320260
rect 70636 320220 70642 320232
rect 73154 320220 73160 320232
rect 73212 320220 73218 320272
rect 77018 320220 77024 320272
rect 77076 320260 77082 320272
rect 79962 320260 79968 320272
rect 77076 320232 79968 320260
rect 77076 320220 77082 320232
rect 79962 320220 79968 320232
rect 80020 320220 80026 320272
rect 81342 320220 81348 320272
rect 81400 320260 81406 320272
rect 83090 320260 83096 320272
rect 81400 320232 83096 320260
rect 81400 320220 81406 320232
rect 83090 320220 83096 320232
rect 83148 320220 83154 320272
rect 85666 320220 85672 320272
rect 85724 320260 85730 320272
rect 89622 320260 89628 320272
rect 85724 320232 89628 320260
rect 85724 320220 85730 320232
rect 89622 320220 89628 320232
rect 89680 320220 89686 320272
rect 96430 320220 96436 320272
rect 96488 320260 96494 320272
rect 100754 320260 100760 320272
rect 96488 320232 100760 320260
rect 96488 320220 96494 320232
rect 100754 320220 100760 320232
rect 100812 320220 100818 320272
rect 105078 320220 105084 320272
rect 105136 320260 105142 320272
rect 110414 320260 110420 320272
rect 105136 320232 110420 320260
rect 105136 320220 105142 320232
rect 110414 320220 110420 320232
rect 110472 320220 110478 320272
rect 163222 320220 163228 320272
rect 163280 320260 163286 320272
rect 167638 320260 167644 320272
rect 163280 320232 167644 320260
rect 163280 320220 163286 320232
rect 167638 320220 167644 320232
rect 167696 320220 167702 320272
rect 197538 320220 197544 320272
rect 197596 320260 197602 320272
rect 199930 320260 199936 320272
rect 197596 320232 199936 320260
rect 197596 320220 197602 320232
rect 199930 320220 199936 320232
rect 199988 320220 199994 320272
rect 201494 320220 201500 320272
rect 201552 320260 201558 320272
rect 204162 320260 204168 320272
rect 201552 320232 204168 320260
rect 201552 320220 201558 320232
rect 204162 320220 204168 320232
rect 204220 320220 204226 320272
rect 233142 320220 233148 320272
rect 233200 320260 233206 320272
rect 236546 320260 236552 320272
rect 233200 320232 236552 320260
rect 233200 320220 233206 320232
rect 236546 320220 236552 320232
rect 236604 320220 236610 320272
rect 237834 320220 237840 320272
rect 237892 320260 237898 320272
rect 240870 320260 240876 320272
rect 237892 320232 240876 320260
rect 237892 320220 237898 320232
rect 240870 320220 240876 320232
rect 240928 320220 240934 320272
rect 241422 320220 241428 320272
rect 241480 320260 241486 320272
rect 244090 320260 244096 320272
rect 241480 320232 244096 320260
rect 241480 320220 241486 320232
rect 244090 320220 244096 320232
rect 244148 320220 244154 320272
rect 245010 320220 245016 320272
rect 245068 320260 245074 320272
rect 247310 320260 247316 320272
rect 245068 320232 247316 320260
rect 245068 320220 245074 320232
rect 247310 320220 247316 320232
rect 247368 320220 247374 320272
rect 247402 320220 247408 320272
rect 247460 320260 247466 320272
rect 249426 320260 249432 320272
rect 247460 320232 249432 320260
rect 247460 320220 247466 320232
rect 249426 320220 249432 320232
rect 249484 320220 249490 320272
rect 251082 320220 251088 320272
rect 251140 320260 251146 320272
rect 252738 320260 252744 320272
rect 251140 320232 252744 320260
rect 251140 320220 251146 320232
rect 252738 320220 252744 320232
rect 252796 320220 252802 320272
rect 254578 320220 254584 320272
rect 254636 320260 254642 320272
rect 255958 320260 255964 320272
rect 254636 320232 255964 320260
rect 254636 320220 254642 320232
rect 255958 320220 255964 320232
rect 256016 320220 256022 320272
rect 257982 320220 257988 320272
rect 258040 320260 258046 320272
rect 259178 320260 259184 320272
rect 258040 320232 259184 320260
rect 258040 320220 258046 320232
rect 259178 320220 259184 320232
rect 259236 320220 259242 320272
rect 22002 320152 22008 320204
rect 22060 320192 22066 320204
rect 24210 320192 24216 320204
rect 22060 320164 24216 320192
rect 22060 320152 22066 320164
rect 24210 320152 24216 320164
rect 24268 320152 24274 320204
rect 26510 320152 26516 320204
rect 26568 320192 26574 320204
rect 28534 320192 28540 320204
rect 26568 320164 28540 320192
rect 26568 320152 26574 320164
rect 28534 320152 28540 320164
rect 28592 320152 28598 320204
rect 28902 320152 28908 320204
rect 28960 320192 28966 320204
rect 30650 320192 30656 320204
rect 28960 320164 30656 320192
rect 28960 320152 28966 320164
rect 30650 320152 30656 320164
rect 30708 320152 30714 320204
rect 31662 320152 31668 320204
rect 31720 320192 31726 320204
rect 32858 320192 32864 320204
rect 31720 320164 32864 320192
rect 31720 320152 31726 320164
rect 32858 320152 32864 320164
rect 32916 320152 32922 320204
rect 33042 320152 33048 320204
rect 33100 320192 33106 320204
rect 33870 320192 33876 320204
rect 33100 320164 33876 320192
rect 33100 320152 33106 320164
rect 33870 320152 33876 320164
rect 33928 320152 33934 320204
rect 35894 320152 35900 320204
rect 35952 320192 35958 320204
rect 37182 320192 37188 320204
rect 35952 320164 37188 320192
rect 35952 320152 35958 320164
rect 37182 320152 37188 320164
rect 37240 320152 37246 320204
rect 37274 320152 37280 320204
rect 37332 320192 37338 320204
rect 38194 320192 38200 320204
rect 37332 320164 38200 320192
rect 37332 320152 37338 320164
rect 38194 320152 38200 320164
rect 38252 320152 38258 320204
rect 38562 320152 38568 320204
rect 38620 320192 38626 320204
rect 39298 320192 39304 320204
rect 38620 320164 39304 320192
rect 38620 320152 38626 320164
rect 39298 320152 39304 320164
rect 39356 320152 39362 320204
rect 42518 320192 42524 320204
rect 41432 320164 42524 320192
rect 41432 320136 41460 320164
rect 42518 320152 42524 320164
rect 42576 320152 42582 320204
rect 42794 320152 42800 320204
rect 42852 320192 42858 320204
rect 43622 320192 43628 320204
rect 42852 320164 43628 320192
rect 42852 320152 42858 320164
rect 43622 320152 43628 320164
rect 43680 320152 43686 320204
rect 46934 320152 46940 320204
rect 46992 320192 46998 320204
rect 47946 320192 47952 320204
rect 46992 320164 47952 320192
rect 46992 320152 46998 320164
rect 47946 320152 47952 320164
rect 48004 320152 48010 320204
rect 59814 320152 59820 320204
rect 59872 320192 59878 320204
rect 60734 320192 60740 320204
rect 59872 320164 60740 320192
rect 59872 320152 59878 320164
rect 60734 320152 60740 320164
rect 60792 320152 60798 320204
rect 60826 320152 60832 320204
rect 60884 320192 60890 320204
rect 62114 320192 62120 320204
rect 60884 320164 62120 320192
rect 60884 320152 60890 320164
rect 62114 320152 62120 320164
rect 62172 320152 62178 320204
rect 63034 320152 63040 320204
rect 63092 320192 63098 320204
rect 64322 320192 64328 320204
rect 63092 320164 64328 320192
rect 63092 320152 63098 320164
rect 64322 320152 64328 320164
rect 64380 320152 64386 320204
rect 65150 320152 65156 320204
rect 65208 320192 65214 320204
rect 66254 320192 66260 320204
rect 65208 320164 66260 320192
rect 65208 320152 65214 320164
rect 66254 320152 66260 320164
rect 66312 320152 66318 320204
rect 67358 320152 67364 320204
rect 67416 320192 67422 320204
rect 69014 320192 69020 320204
rect 67416 320164 69020 320192
rect 67416 320152 67422 320164
rect 69014 320152 69020 320164
rect 69072 320152 69078 320204
rect 71590 320152 71596 320204
rect 71648 320192 71654 320204
rect 73246 320192 73252 320204
rect 71648 320164 73252 320192
rect 71648 320152 71654 320164
rect 73246 320152 73252 320164
rect 73304 320152 73310 320204
rect 74902 320152 74908 320204
rect 74960 320192 74966 320204
rect 77294 320192 77300 320204
rect 74960 320164 77300 320192
rect 74960 320152 74966 320164
rect 77294 320152 77300 320164
rect 77352 320152 77358 320204
rect 79134 320152 79140 320204
rect 79192 320192 79198 320204
rect 81618 320192 81624 320204
rect 79192 320164 81624 320192
rect 79192 320152 79198 320164
rect 81618 320152 81624 320164
rect 81676 320152 81682 320204
rect 84562 320152 84568 320204
rect 84620 320192 84626 320204
rect 88058 320192 88064 320204
rect 84620 320164 88064 320192
rect 84620 320152 84626 320164
rect 88058 320152 88064 320164
rect 88116 320152 88122 320204
rect 89990 320152 89996 320204
rect 90048 320192 90054 320204
rect 92658 320192 92664 320204
rect 90048 320164 92664 320192
rect 90048 320152 90054 320164
rect 92658 320152 92664 320164
rect 92716 320152 92722 320204
rect 95326 320152 95332 320204
rect 95384 320192 95390 320204
rect 99098 320192 99104 320204
rect 95384 320164 99104 320192
rect 95384 320152 95390 320164
rect 99098 320152 99104 320164
rect 99156 320152 99162 320204
rect 107194 320152 107200 320204
rect 107252 320192 107258 320204
rect 112438 320192 112444 320204
rect 107252 320164 112444 320192
rect 107252 320152 107258 320164
rect 112438 320152 112444 320164
rect 112496 320152 112502 320204
rect 113634 320152 113640 320204
rect 113692 320192 113698 320204
rect 114462 320192 114468 320204
rect 113692 320164 114468 320192
rect 113692 320152 113698 320164
rect 114462 320152 114468 320164
rect 114520 320152 114526 320204
rect 114738 320152 114744 320204
rect 114796 320192 114802 320204
rect 115842 320192 115848 320204
rect 114796 320164 115848 320192
rect 114796 320152 114802 320164
rect 115842 320152 115848 320164
rect 115900 320152 115906 320204
rect 119062 320152 119068 320204
rect 119120 320192 119126 320204
rect 119982 320192 119988 320204
rect 119120 320164 119988 320192
rect 119120 320152 119126 320164
rect 119982 320152 119988 320164
rect 120040 320152 120046 320204
rect 120166 320152 120172 320204
rect 120224 320192 120230 320204
rect 121362 320192 121368 320204
rect 120224 320164 121368 320192
rect 120224 320152 120230 320164
rect 121362 320152 121368 320164
rect 121420 320152 121426 320204
rect 124398 320152 124404 320204
rect 124456 320192 124462 320204
rect 125410 320192 125416 320204
rect 124456 320164 125416 320192
rect 124456 320152 124462 320164
rect 125410 320152 125416 320164
rect 125468 320152 125474 320204
rect 128722 320152 128728 320204
rect 128780 320192 128786 320204
rect 129642 320192 129648 320204
rect 128780 320164 129648 320192
rect 128780 320152 128786 320164
rect 129642 320152 129648 320164
rect 129700 320152 129706 320204
rect 129826 320152 129832 320204
rect 129884 320192 129890 320204
rect 130930 320192 130936 320204
rect 129884 320164 130936 320192
rect 129884 320152 129890 320164
rect 130930 320152 130936 320164
rect 130988 320152 130994 320204
rect 133046 320152 133052 320204
rect 133104 320192 133110 320204
rect 133782 320192 133788 320204
rect 133104 320164 133788 320192
rect 133104 320152 133110 320164
rect 133782 320152 133788 320164
rect 133840 320152 133846 320204
rect 134150 320152 134156 320204
rect 134208 320192 134214 320204
rect 135162 320192 135168 320204
rect 134208 320164 135168 320192
rect 134208 320152 134214 320164
rect 135162 320152 135168 320164
rect 135220 320152 135226 320204
rect 135254 320152 135260 320204
rect 135312 320192 135318 320204
rect 136542 320192 136548 320204
rect 135312 320164 136548 320192
rect 135312 320152 135318 320164
rect 136542 320152 136548 320164
rect 136600 320152 136606 320204
rect 138474 320152 138480 320204
rect 138532 320192 138538 320204
rect 139302 320192 139308 320204
rect 138532 320164 139308 320192
rect 138532 320152 138538 320164
rect 139302 320152 139308 320164
rect 139360 320152 139366 320204
rect 139486 320152 139492 320204
rect 139544 320192 139550 320204
rect 140682 320192 140688 320204
rect 139544 320164 140688 320192
rect 139544 320152 139550 320164
rect 140682 320152 140688 320164
rect 140740 320152 140746 320204
rect 143810 320152 143816 320204
rect 143868 320192 143874 320204
rect 144822 320192 144828 320204
rect 143868 320164 144828 320192
rect 143868 320152 143874 320164
rect 144822 320152 144828 320164
rect 144880 320152 144886 320204
rect 144914 320152 144920 320204
rect 144972 320192 144978 320204
rect 146110 320192 146116 320204
rect 144972 320164 146116 320192
rect 144972 320152 144978 320164
rect 146110 320152 146116 320164
rect 146168 320152 146174 320204
rect 148134 320152 148140 320204
rect 148192 320192 148198 320204
rect 148962 320192 148968 320204
rect 148192 320164 148968 320192
rect 148192 320152 148198 320164
rect 148962 320152 148968 320164
rect 149020 320152 149026 320204
rect 149238 320152 149244 320204
rect 149296 320192 149302 320204
rect 150250 320192 150256 320204
rect 149296 320164 150256 320192
rect 149296 320152 149302 320164
rect 150250 320152 150256 320164
rect 150308 320152 150314 320204
rect 153562 320152 153568 320204
rect 153620 320192 153626 320204
rect 154482 320192 154488 320204
rect 153620 320164 154488 320192
rect 153620 320152 153626 320164
rect 154482 320152 154488 320164
rect 154540 320152 154546 320204
rect 154666 320152 154672 320204
rect 154724 320192 154730 320204
rect 155770 320192 155776 320204
rect 154724 320164 155776 320192
rect 154724 320152 154730 320164
rect 155770 320152 155776 320164
rect 155828 320152 155834 320204
rect 157886 320152 157892 320204
rect 157944 320192 157950 320204
rect 158622 320192 158628 320204
rect 157944 320164 158628 320192
rect 157944 320152 157950 320164
rect 158622 320152 158628 320164
rect 158680 320152 158686 320204
rect 158898 320152 158904 320204
rect 158956 320192 158962 320204
rect 159910 320192 159916 320204
rect 158956 320164 159916 320192
rect 158956 320152 158962 320164
rect 159910 320152 159916 320164
rect 159968 320152 159974 320204
rect 164326 320152 164332 320204
rect 164384 320192 164390 320204
rect 165430 320192 165436 320204
rect 164384 320164 165436 320192
rect 164384 320152 164390 320164
rect 165430 320152 165436 320164
rect 165488 320152 165494 320204
rect 168650 320152 168656 320204
rect 168708 320192 168714 320204
rect 169662 320192 169668 320204
rect 168708 320164 169668 320192
rect 168708 320152 168714 320164
rect 169662 320152 169668 320164
rect 169720 320152 169726 320204
rect 169754 320152 169760 320204
rect 169812 320192 169818 320204
rect 170950 320192 170956 320204
rect 169812 320164 170956 320192
rect 169812 320152 169818 320164
rect 170950 320152 170956 320164
rect 171008 320152 171014 320204
rect 172974 320152 172980 320204
rect 173032 320192 173038 320204
rect 173802 320192 173808 320204
rect 173032 320164 173808 320192
rect 173032 320152 173038 320164
rect 173802 320152 173808 320164
rect 173860 320152 173866 320204
rect 173986 320152 173992 320204
rect 174044 320192 174050 320204
rect 175090 320192 175096 320204
rect 174044 320164 175096 320192
rect 174044 320152 174050 320164
rect 175090 320152 175096 320164
rect 175148 320152 175154 320204
rect 178310 320152 178316 320204
rect 178368 320192 178374 320204
rect 179322 320192 179328 320204
rect 178368 320164 179328 320192
rect 178368 320152 178374 320164
rect 179322 320152 179328 320164
rect 179380 320152 179386 320204
rect 179414 320152 179420 320204
rect 179472 320192 179478 320204
rect 180702 320192 180708 320204
rect 179472 320164 180708 320192
rect 179472 320152 179478 320164
rect 180702 320152 180708 320164
rect 180760 320152 180766 320204
rect 182634 320152 182640 320204
rect 182692 320192 182698 320204
rect 183462 320192 183468 320204
rect 182692 320164 183468 320192
rect 182692 320152 182698 320164
rect 183462 320152 183468 320164
rect 183520 320152 183526 320204
rect 183738 320152 183744 320204
rect 183796 320192 183802 320204
rect 184750 320192 184756 320204
rect 183796 320164 184756 320192
rect 183796 320152 183802 320164
rect 184750 320152 184756 320164
rect 184808 320152 184814 320204
rect 191834 320152 191840 320204
rect 191892 320192 191898 320204
rect 196618 320192 196624 320204
rect 191892 320164 196624 320192
rect 191892 320152 191898 320164
rect 196618 320152 196624 320164
rect 196676 320152 196682 320204
rect 197262 320152 197268 320204
rect 197320 320192 197326 320204
rect 198826 320192 198832 320204
rect 197320 320164 198832 320192
rect 197320 320152 197326 320164
rect 198826 320152 198832 320164
rect 198884 320152 198890 320204
rect 199010 320152 199016 320204
rect 199068 320192 199074 320204
rect 202046 320192 202052 320204
rect 199068 320164 202052 320192
rect 199068 320152 199074 320164
rect 202046 320152 202052 320164
rect 202104 320152 202110 320204
rect 202874 320152 202880 320204
rect 202932 320192 202938 320204
rect 205266 320192 205272 320204
rect 202932 320164 205272 320192
rect 202932 320152 202938 320164
rect 205266 320152 205272 320164
rect 205324 320152 205330 320204
rect 207106 320152 207112 320204
rect 207164 320192 207170 320204
rect 209590 320192 209596 320204
rect 207164 320164 209596 320192
rect 207164 320152 207170 320164
rect 209590 320152 209596 320164
rect 209648 320152 209654 320204
rect 219894 320152 219900 320204
rect 219952 320192 219958 320204
rect 224678 320192 224684 320204
rect 219952 320164 224684 320192
rect 219952 320152 219958 320164
rect 224678 320152 224684 320164
rect 224736 320152 224742 320204
rect 224862 320152 224868 320204
rect 224920 320192 224926 320204
rect 229002 320192 229008 320204
rect 224920 320164 229008 320192
rect 224920 320152 224926 320164
rect 229002 320152 229008 320164
rect 229060 320152 229066 320204
rect 230290 320152 230296 320204
rect 230348 320192 230354 320204
rect 234338 320192 234344 320204
rect 230348 320164 234344 320192
rect 230348 320152 230354 320164
rect 234338 320152 234344 320164
rect 234396 320152 234402 320204
rect 234522 320152 234528 320204
rect 234580 320192 234586 320204
rect 237650 320192 237656 320204
rect 234580 320164 237656 320192
rect 234580 320152 234586 320164
rect 237650 320152 237656 320164
rect 237708 320152 237714 320204
rect 240042 320152 240048 320204
rect 240100 320192 240106 320204
rect 242986 320192 242992 320204
rect 240100 320164 242992 320192
rect 240100 320152 240106 320164
rect 242986 320152 242992 320164
rect 243044 320152 243050 320204
rect 243814 320152 243820 320204
rect 243872 320192 243878 320204
rect 246206 320192 246212 320204
rect 243872 320164 246212 320192
rect 243872 320152 243878 320164
rect 246206 320152 246212 320164
rect 246264 320152 246270 320204
rect 249702 320152 249708 320204
rect 249760 320192 249766 320204
rect 251634 320192 251640 320204
rect 249760 320164 251640 320192
rect 249760 320152 249766 320164
rect 251634 320152 251640 320164
rect 251692 320152 251698 320204
rect 252462 320152 252468 320204
rect 252520 320192 252526 320204
rect 253750 320192 253756 320204
rect 252520 320164 253756 320192
rect 252520 320152 252526 320164
rect 253750 320152 253756 320164
rect 253808 320152 253814 320204
rect 255774 320152 255780 320204
rect 255832 320192 255838 320204
rect 256970 320192 256976 320204
rect 255832 320164 256976 320192
rect 255832 320152 255838 320164
rect 256970 320152 256976 320164
rect 257028 320152 257034 320204
rect 259362 320152 259368 320204
rect 259420 320192 259426 320204
rect 260282 320192 260288 320204
rect 259420 320164 260288 320192
rect 259420 320152 259426 320164
rect 260282 320152 260288 320164
rect 260340 320152 260346 320204
rect 263502 320192 263508 320204
rect 262232 320164 263508 320192
rect 41414 320084 41420 320136
rect 41472 320084 41478 320136
rect 262232 320068 262260 320164
rect 263502 320152 263508 320164
rect 263560 320152 263566 320204
rect 263594 320152 263600 320204
rect 263652 320192 263658 320204
rect 264514 320192 264520 320204
rect 263652 320164 264520 320192
rect 263652 320152 263658 320164
rect 264514 320152 264520 320164
rect 264572 320152 264578 320204
rect 267734 320152 267740 320204
rect 267792 320192 267798 320204
rect 268838 320192 268844 320204
rect 267792 320164 268844 320192
rect 267792 320152 267798 320164
rect 268838 320152 268844 320164
rect 268896 320152 268902 320204
rect 269114 320152 269120 320204
rect 269172 320192 269178 320204
rect 269942 320192 269948 320204
rect 269172 320164 269948 320192
rect 269172 320152 269178 320164
rect 269942 320152 269948 320164
rect 270000 320152 270006 320204
rect 276014 320152 276020 320204
rect 276072 320192 276078 320204
rect 276658 320192 276664 320204
rect 276072 320164 276664 320192
rect 276072 320152 276078 320164
rect 276658 320152 276664 320164
rect 276716 320152 276722 320204
rect 277394 320152 277400 320204
rect 277452 320192 277458 320204
rect 277854 320192 277860 320204
rect 277452 320164 277860 320192
rect 277452 320152 277458 320164
rect 277854 320152 277860 320164
rect 277912 320152 277918 320204
rect 278682 320152 278688 320204
rect 278740 320192 278746 320204
rect 279050 320192 279056 320204
rect 278740 320164 279056 320192
rect 278740 320152 278746 320164
rect 279050 320152 279056 320164
rect 279108 320152 279114 320204
rect 262214 320016 262220 320068
rect 262272 320016 262278 320068
rect 22186 319404 22192 319456
rect 22244 319444 22250 319456
rect 36538 319444 36544 319456
rect 22244 319416 36544 319444
rect 22244 319404 22250 319416
rect 36538 319404 36544 319416
rect 36596 319404 36602 319456
rect 20622 318724 20628 318776
rect 20680 318764 20686 318776
rect 23106 318764 23112 318776
rect 20680 318736 23112 318764
rect 20680 318724 20686 318736
rect 23106 318724 23112 318736
rect 23164 318724 23170 318776
rect 91278 318724 91284 318776
rect 91336 318764 91342 318776
rect 93486 318764 93492 318776
rect 91336 318736 93492 318764
rect 91336 318724 91342 318736
rect 93486 318724 93492 318736
rect 93544 318724 93550 318776
rect 99098 318724 99104 318776
rect 99156 318764 99162 318776
rect 100662 318764 100668 318776
rect 99156 318736 100668 318764
rect 99156 318724 99162 318736
rect 100662 318724 100668 318736
rect 100720 318724 100726 318776
rect 191190 318724 191196 318776
rect 191248 318764 191254 318776
rect 197262 318764 197268 318776
rect 191248 318736 197268 318764
rect 191248 318724 191254 318736
rect 197262 318724 197268 318736
rect 197320 318724 197326 318776
rect 200758 318724 200764 318776
rect 200816 318764 200822 318776
rect 206922 318764 206928 318776
rect 200816 318736 206928 318764
rect 200816 318724 200822 318736
rect 206922 318724 206928 318736
rect 206980 318724 206986 318776
rect 211522 318724 211528 318776
rect 211580 318764 211586 318776
rect 217134 318764 217140 318776
rect 211580 318736 217140 318764
rect 211580 318724 211586 318736
rect 217134 318724 217140 318736
rect 217192 318724 217198 318776
rect 223482 318724 223488 318776
rect 223540 318764 223546 318776
rect 227898 318764 227904 318776
rect 223540 318736 227904 318764
rect 223540 318724 223546 318736
rect 227898 318724 227904 318736
rect 227956 318724 227962 318776
rect 201954 318656 201960 318708
rect 202012 318696 202018 318708
rect 208302 318696 208308 318708
rect 202012 318668 208308 318696
rect 202012 318656 202018 318668
rect 208302 318656 208308 318668
rect 208360 318656 208366 318708
rect 220630 318656 220636 318708
rect 220688 318696 220694 318708
rect 225782 318696 225788 318708
rect 220688 318668 225788 318696
rect 220688 318656 220694 318668
rect 225782 318656 225788 318668
rect 225840 318656 225846 318708
rect 106366 318520 106372 318572
rect 106424 318560 106430 318572
rect 107838 318560 107844 318572
rect 106424 318532 107844 318560
rect 106424 318520 106430 318532
rect 107838 318520 107844 318532
rect 107896 318520 107902 318572
rect 192386 318520 192392 318572
rect 192444 318560 192450 318572
rect 197538 318560 197544 318572
rect 192444 318532 197544 318560
rect 192444 318520 192450 318532
rect 197538 318520 197544 318532
rect 197596 318520 197602 318572
rect 193582 318452 193588 318504
rect 193640 318492 193646 318504
rect 198734 318492 198740 318504
rect 193640 318464 198740 318492
rect 193640 318452 193646 318464
rect 198734 318452 198740 318464
rect 198792 318452 198798 318504
rect 34882 318384 34888 318436
rect 34940 318424 34946 318436
rect 35802 318424 35808 318436
rect 34940 318396 35808 318424
rect 34940 318384 34946 318396
rect 35802 318384 35808 318396
rect 35860 318384 35866 318436
rect 85114 318384 85120 318436
rect 85172 318424 85178 318436
rect 86310 318424 86316 318436
rect 85172 318396 86316 318424
rect 85172 318384 85178 318396
rect 86310 318384 86316 318396
rect 86368 318384 86374 318436
rect 88058 318384 88064 318436
rect 88116 318424 88122 318436
rect 88702 318424 88708 318436
rect 88116 318396 88708 318424
rect 88116 318384 88122 318396
rect 88702 318384 88708 318396
rect 88760 318384 88766 318436
rect 194502 318384 194508 318436
rect 194560 318424 194566 318436
rect 199010 318424 199016 318436
rect 194560 318396 199016 318424
rect 194560 318384 194566 318396
rect 199010 318384 199016 318396
rect 199068 318384 199074 318436
rect 209130 318384 209136 318436
rect 209188 318424 209194 318436
rect 215018 318424 215024 318436
rect 209188 318396 215024 318424
rect 209188 318384 209194 318396
rect 215018 318384 215024 318396
rect 215076 318384 215082 318436
rect 85758 318316 85764 318368
rect 85816 318356 85822 318368
rect 87506 318356 87512 318368
rect 85816 318328 87512 318356
rect 85816 318316 85822 318328
rect 87506 318316 87512 318328
rect 87564 318316 87570 318368
rect 195790 318248 195796 318300
rect 195848 318288 195854 318300
rect 200114 318288 200120 318300
rect 195848 318260 200120 318288
rect 195848 318248 195854 318260
rect 200114 318248 200120 318260
rect 200172 318248 200178 318300
rect 204162 318248 204168 318300
rect 204220 318288 204226 318300
rect 208394 318288 208400 318300
rect 204220 318260 208400 318288
rect 204220 318248 204226 318260
rect 208394 318248 208400 318260
rect 208452 318248 208458 318300
rect 217502 318248 217508 318300
rect 217560 318288 217566 318300
rect 222562 318288 222568 318300
rect 217560 318260 222568 318288
rect 217560 318248 217566 318260
rect 222562 318248 222568 318260
rect 222620 318248 222626 318300
rect 198366 318180 198372 318232
rect 198424 318220 198430 318232
rect 202874 318220 202880 318232
rect 198424 318192 202880 318220
rect 198424 318180 198430 318192
rect 202874 318180 202880 318192
rect 202932 318180 202938 318232
rect 218698 318180 218704 318232
rect 218756 318220 218762 318232
rect 223574 318220 223580 318232
rect 218756 318192 223580 318220
rect 218756 318180 218762 318192
rect 223574 318180 223580 318192
rect 223632 318180 223638 318232
rect 202782 318112 202788 318164
rect 202840 318152 202846 318164
rect 207106 318152 207112 318164
rect 202840 318124 207112 318152
rect 202840 318112 202846 318124
rect 207106 318112 207112 318124
rect 207164 318112 207170 318164
rect 207934 318112 207940 318164
rect 207992 318152 207998 318164
rect 213822 318152 213828 318164
rect 207992 318124 213828 318152
rect 207992 318112 207998 318124
rect 213822 318112 213828 318124
rect 213880 318112 213886 318164
rect 42886 318044 42892 318096
rect 42944 318084 42950 318096
rect 113358 318084 113364 318096
rect 42944 318056 113364 318084
rect 42944 318044 42950 318056
rect 113358 318044 113364 318056
rect 113416 318044 113422 318096
rect 189994 318044 190000 318096
rect 190052 318084 190058 318096
rect 197170 318084 197176 318096
rect 190052 318056 197176 318084
rect 190052 318044 190058 318056
rect 197170 318044 197176 318056
rect 197228 318044 197234 318096
rect 90082 317976 90088 318028
rect 90140 318016 90146 318028
rect 92290 318016 92296 318028
rect 90140 317988 92296 318016
rect 90140 317976 90146 317988
rect 92290 317976 92296 317988
rect 92348 317976 92354 318028
rect 197170 317908 197176 317960
rect 197228 317948 197234 317960
rect 201494 317948 201500 317960
rect 197228 317920 201500 317948
rect 197228 317908 197234 317920
rect 201494 317908 201500 317920
rect 201552 317908 201558 317960
rect 213822 317908 213828 317960
rect 213880 317948 213886 317960
rect 219250 317948 219256 317960
rect 213880 317920 219256 317948
rect 213880 317908 213886 317920
rect 219250 317908 219256 317920
rect 219308 317908 219314 317960
rect 222010 317908 222016 317960
rect 222068 317948 222074 317960
rect 226794 317948 226800 317960
rect 222068 317920 226800 317948
rect 222068 317908 222074 317920
rect 226794 317908 226800 317920
rect 226852 317908 226858 317960
rect 199562 317704 199568 317756
rect 199620 317744 199626 317756
rect 204254 317744 204260 317756
rect 199620 317716 204260 317744
rect 199620 317704 199626 317716
rect 204254 317704 204260 317716
rect 204312 317704 204318 317756
rect 210326 317704 210332 317756
rect 210384 317744 210390 317756
rect 216030 317744 216036 317756
rect 210384 317716 216036 317744
rect 210384 317704 210390 317716
rect 216030 317704 216036 317716
rect 216088 317704 216094 317756
rect 206738 317568 206744 317620
rect 206796 317608 206802 317620
rect 212442 317608 212448 317620
rect 206796 317580 212448 317608
rect 206796 317568 206802 317580
rect 212442 317568 212448 317580
rect 212500 317568 212506 317620
rect 216306 317568 216312 317620
rect 216364 317608 216370 317620
rect 221458 317608 221464 317620
rect 216364 317580 221464 317608
rect 216364 317568 216370 317580
rect 221458 317568 221464 317580
rect 221516 317568 221522 317620
rect 83090 317500 83096 317552
rect 83148 317540 83154 317552
rect 85114 317540 85120 317552
rect 83148 317512 85120 317540
rect 83148 317500 83154 317512
rect 85114 317500 85120 317512
rect 85172 317500 85178 317552
rect 188890 317500 188896 317552
rect 188948 317540 188954 317552
rect 191834 317540 191840 317552
rect 188948 317512 191840 317540
rect 188948 317500 188954 317512
rect 191834 317500 191840 317512
rect 191892 317500 191898 317552
rect 205358 317500 205364 317552
rect 205416 317540 205422 317552
rect 211062 317540 211068 317552
rect 205416 317512 211068 317540
rect 205416 317500 205422 317512
rect 211062 317500 211068 317512
rect 211120 317500 211126 317552
rect 217962 317540 217968 317552
rect 212460 317512 217968 317540
rect 212460 317484 212488 317512
rect 217962 317500 217968 317512
rect 218020 317500 218026 317552
rect 92658 317432 92664 317484
rect 92716 317472 92722 317484
rect 94682 317472 94688 317484
rect 92716 317444 94688 317472
rect 92716 317432 92722 317444
rect 94682 317432 94688 317444
rect 94740 317432 94746 317484
rect 212442 317432 212448 317484
rect 212500 317432 212506 317484
rect 215110 317432 215116 317484
rect 215168 317472 215174 317484
rect 220354 317472 220360 317484
rect 215168 317444 220360 317472
rect 215168 317432 215174 317444
rect 220354 317432 220360 317444
rect 220412 317432 220418 317484
rect 2774 316684 2780 316736
rect 2832 316724 2838 316736
rect 3510 316724 3516 316736
rect 2832 316696 3516 316724
rect 2832 316684 2838 316696
rect 3510 316684 3516 316696
rect 3568 316724 3574 316736
rect 288894 316724 288900 316736
rect 3568 316696 288900 316724
rect 3568 316684 3574 316696
rect 288894 316684 288900 316696
rect 288952 316684 288958 316736
rect 36538 315324 36544 315376
rect 36596 315364 36602 315376
rect 111794 315364 111800 315376
rect 36596 315336 111800 315364
rect 36596 315324 36602 315336
rect 111794 315324 111800 315336
rect 111852 315324 111858 315376
rect 14550 315256 14556 315308
rect 14608 315296 14614 315308
rect 185578 315296 185584 315308
rect 14608 315268 185584 315296
rect 14608 315256 14614 315268
rect 185578 315256 185584 315268
rect 185636 315256 185642 315308
rect 111794 313216 111800 313268
rect 111852 313256 111858 313268
rect 114370 313256 114376 313268
rect 111852 313228 114376 313256
rect 111852 313216 111858 313228
rect 114370 313216 114376 313228
rect 114428 313216 114434 313268
rect 303614 311856 303620 311908
rect 303672 311896 303678 311908
rect 335998 311896 336004 311908
rect 303672 311868 336004 311896
rect 303672 311856 303678 311868
rect 335998 311856 336004 311868
rect 336056 311856 336062 311908
rect 114370 310768 114376 310820
rect 114428 310808 114434 310820
rect 116578 310808 116584 310820
rect 114428 310780 116584 310808
rect 114428 310768 114434 310780
rect 116578 310768 116584 310780
rect 116636 310768 116642 310820
rect 303614 310496 303620 310548
rect 303672 310536 303678 310548
rect 341518 310536 341524 310548
rect 303672 310508 341524 310536
rect 303672 310496 303678 310508
rect 341518 310496 341524 310508
rect 341576 310496 341582 310548
rect 303614 309136 303620 309188
rect 303672 309176 303678 309188
rect 340138 309176 340144 309188
rect 303672 309148 340144 309176
rect 303672 309136 303678 309148
rect 340138 309136 340144 309148
rect 340196 309136 340202 309188
rect 282086 309108 282092 309120
rect 282047 309080 282092 309108
rect 282086 309068 282092 309080
rect 282144 309068 282150 309120
rect 113174 306348 113180 306400
rect 113232 306388 113238 306400
rect 113358 306388 113364 306400
rect 113232 306360 113364 306388
rect 113232 306348 113238 306360
rect 113358 306348 113364 306360
rect 113416 306348 113422 306400
rect 303614 306348 303620 306400
rect 303672 306388 303678 306400
rect 560938 306388 560944 306400
rect 303672 306360 560944 306388
rect 303672 306348 303678 306360
rect 560938 306348 560944 306360
rect 560996 306348 561002 306400
rect 282089 305643 282147 305649
rect 282089 305609 282101 305643
rect 282135 305640 282147 305643
rect 300854 305640 300860 305652
rect 282135 305612 300860 305640
rect 282135 305609 282147 305612
rect 282089 305603 282147 305609
rect 300854 305600 300860 305612
rect 300912 305600 300918 305652
rect 296162 303560 296168 303612
rect 296220 303600 296226 303612
rect 580350 303600 580356 303612
rect 296220 303572 580356 303600
rect 296220 303560 296226 303572
rect 580350 303560 580356 303572
rect 580408 303560 580414 303612
rect 282089 299523 282147 299529
rect 282089 299489 282101 299523
rect 282135 299520 282147 299523
rect 282546 299520 282552 299532
rect 282135 299492 282552 299520
rect 282135 299489 282147 299492
rect 282089 299483 282147 299489
rect 282546 299480 282552 299492
rect 282604 299480 282610 299532
rect 282362 292544 282368 292596
rect 282420 292584 282426 292596
rect 282546 292584 282552 292596
rect 282420 292556 282552 292584
rect 282420 292544 282426 292556
rect 282546 292544 282552 292556
rect 282604 292544 282610 292596
rect 282270 278740 282276 278792
rect 282328 278780 282334 278792
rect 282362 278780 282368 278792
rect 282328 278752 282368 278780
rect 282328 278740 282334 278752
rect 282362 278740 282368 278752
rect 282420 278740 282426 278792
rect 11698 275952 11704 276004
rect 11756 275992 11762 276004
rect 17126 275992 17132 276004
rect 11756 275964 17132 275992
rect 11756 275952 11762 275964
rect 17126 275952 17132 275964
rect 17184 275952 17190 276004
rect 304350 275952 304356 276004
rect 304408 275992 304414 276004
rect 580166 275992 580172 276004
rect 304408 275964 580172 275992
rect 304408 275952 304414 275964
rect 580166 275952 580172 275964
rect 580224 275952 580230 276004
rect 282178 263576 282184 263628
rect 282236 263616 282242 263628
rect 282362 263616 282368 263628
rect 282236 263588 282368 263616
rect 282236 263576 282242 263588
rect 282362 263576 282368 263588
rect 282420 263576 282426 263628
rect 146018 254124 146024 254176
rect 146076 254164 146082 254176
rect 149514 254164 149520 254176
rect 146076 254136 149520 254164
rect 146076 254124 146082 254136
rect 149514 254124 149520 254136
rect 149572 254124 149578 254176
rect 214558 233860 214564 233912
rect 214616 233900 214622 233912
rect 315298 233900 315304 233912
rect 214616 233872 315304 233900
rect 214616 233860 214622 233872
rect 315298 233860 315304 233872
rect 315356 233860 315362 233912
rect 67174 230392 67180 230444
rect 67232 230432 67238 230444
rect 72418 230432 72424 230444
rect 67232 230404 72424 230432
rect 67232 230392 67238 230404
rect 72418 230392 72424 230404
rect 72476 230392 72482 230444
rect 214742 229712 214748 229764
rect 214800 229752 214806 229764
rect 305638 229752 305644 229764
rect 214800 229724 305644 229752
rect 214800 229712 214806 229724
rect 305638 229712 305644 229724
rect 305696 229712 305702 229764
rect 245562 229100 245568 229152
rect 245620 229140 245626 229152
rect 250438 229140 250444 229152
rect 245620 229112 250444 229140
rect 245620 229100 245626 229112
rect 250438 229100 250444 229112
rect 250496 229100 250502 229152
rect 304258 229032 304264 229084
rect 304316 229072 304322 229084
rect 579982 229072 579988 229084
rect 304316 229044 579988 229072
rect 304316 229032 304322 229044
rect 579982 229032 579988 229044
rect 580040 229032 580046 229084
rect 214926 228352 214932 228404
rect 214984 228392 214990 228404
rect 301498 228392 301504 228404
rect 214984 228364 301504 228392
rect 214984 228352 214990 228364
rect 301498 228352 301504 228364
rect 301556 228352 301562 228404
rect 72418 227060 72424 227112
rect 72476 227100 72482 227112
rect 79318 227100 79324 227112
rect 72476 227072 79324 227100
rect 72476 227060 72482 227072
rect 79318 227060 79324 227072
rect 79376 227060 79382 227112
rect 13078 226992 13084 227044
rect 13136 227032 13142 227044
rect 411898 227032 411904 227044
rect 13136 227004 411904 227032
rect 13136 226992 13142 227004
rect 411898 226992 411904 227004
rect 411956 226992 411962 227044
rect 214650 225632 214656 225684
rect 214708 225672 214714 225684
rect 312538 225672 312544 225684
rect 214708 225644 312544 225672
rect 214708 225632 214714 225644
rect 312538 225632 312544 225644
rect 312596 225632 312602 225684
rect 9122 225564 9128 225616
rect 9180 225604 9186 225616
rect 299474 225604 299480 225616
rect 9180 225576 299480 225604
rect 9180 225564 9186 225576
rect 299474 225564 299480 225576
rect 299532 225564 299538 225616
rect 125502 224952 125508 225004
rect 125560 224992 125566 225004
rect 214466 224992 214472 225004
rect 125560 224964 125640 224992
rect 214427 224964 214472 224992
rect 125560 224952 125566 224964
rect 114462 224884 114468 224936
rect 114520 224924 114526 224936
rect 125612 224924 125640 224964
rect 214466 224952 214472 224964
rect 214524 224952 214530 225004
rect 128817 224927 128875 224933
rect 128817 224924 128829 224927
rect 114520 224896 125548 224924
rect 125612 224896 128829 224924
rect 114520 224884 114526 224896
rect 119338 224816 119344 224868
rect 119396 224856 119402 224868
rect 125410 224856 125416 224868
rect 119396 224828 125416 224856
rect 119396 224816 119402 224828
rect 125410 224816 125416 224828
rect 125468 224816 125474 224868
rect 125520 224856 125548 224896
rect 128817 224893 128829 224896
rect 128863 224893 128875 224927
rect 128817 224887 128875 224893
rect 130930 224884 130936 224936
rect 130988 224924 130994 224936
rect 145742 224924 145748 224936
rect 130988 224896 145748 224924
rect 130988 224884 130994 224896
rect 145742 224884 145748 224896
rect 145800 224884 145806 224936
rect 155770 224884 155776 224936
rect 155828 224924 155834 224936
rect 170306 224924 170312 224936
rect 155828 224896 170312 224924
rect 155828 224884 155834 224896
rect 170306 224884 170312 224896
rect 170364 224884 170370 224936
rect 179322 224884 179328 224936
rect 179380 224924 179386 224936
rect 193858 224924 193864 224936
rect 179380 224896 193864 224924
rect 179380 224884 179386 224896
rect 193858 224884 193864 224896
rect 193916 224884 193922 224936
rect 127805 224859 127863 224865
rect 127805 224856 127817 224859
rect 125520 224828 127817 224856
rect 127805 224825 127817 224828
rect 127851 224825 127863 224859
rect 127805 224819 127863 224825
rect 128262 224816 128268 224868
rect 128320 224856 128326 224868
rect 143534 224856 143540 224868
rect 128320 224828 143540 224856
rect 128320 224816 128326 224828
rect 143534 224816 143540 224828
rect 143592 224816 143598 224868
rect 150250 224816 150256 224868
rect 150308 224856 150314 224868
rect 164970 224856 164976 224868
rect 150308 224828 164976 224856
rect 150308 224816 150314 224828
rect 164970 224816 164976 224828
rect 165028 224816 165034 224868
rect 167638 224816 167644 224868
rect 167696 224856 167702 224868
rect 178862 224856 178868 224868
rect 167696 224828 178868 224856
rect 167696 224816 167702 224828
rect 178862 224816 178868 224828
rect 178920 224816 178926 224868
rect 180702 224816 180708 224868
rect 180760 224856 180766 224868
rect 194870 224856 194876 224868
rect 180760 224828 194876 224856
rect 180760 224816 180766 224828
rect 194870 224816 194876 224828
rect 194928 224816 194934 224868
rect 115198 224748 115204 224800
rect 115256 224788 115262 224800
rect 124306 224788 124312 224800
rect 115256 224760 124312 224788
rect 115256 224748 115262 224760
rect 124306 224748 124312 224760
rect 124364 224748 124370 224800
rect 126333 224791 126391 224797
rect 126333 224757 126345 224791
rect 126379 224788 126391 224791
rect 132862 224788 132868 224800
rect 126379 224760 132868 224788
rect 126379 224757 126391 224760
rect 126333 224751 126391 224757
rect 132862 224748 132868 224760
rect 132920 224748 132926 224800
rect 146110 224748 146116 224800
rect 146168 224788 146174 224800
rect 160646 224788 160652 224800
rect 146168 224760 160652 224788
rect 146168 224748 146174 224760
rect 160646 224748 160652 224760
rect 160704 224748 160710 224800
rect 161382 224748 161388 224800
rect 161440 224788 161446 224800
rect 176746 224788 176752 224800
rect 161440 224760 176752 224788
rect 161440 224748 161446 224760
rect 176746 224748 176752 224760
rect 176804 224748 176810 224800
rect 183462 224748 183468 224800
rect 183520 224788 183526 224800
rect 198090 224788 198096 224800
rect 183520 224760 198096 224788
rect 183520 224748 183526 224760
rect 198090 224748 198096 224760
rect 198148 224748 198154 224800
rect 122742 224680 122748 224732
rect 122800 224720 122806 224732
rect 138198 224720 138204 224732
rect 122800 224692 138204 224720
rect 122800 224680 122806 224692
rect 138198 224680 138204 224692
rect 138256 224680 138262 224732
rect 151722 224680 151728 224732
rect 151780 224720 151786 224732
rect 167086 224720 167092 224732
rect 151780 224692 167092 224720
rect 151780 224680 151786 224692
rect 167086 224680 167092 224692
rect 167144 224680 167150 224732
rect 170950 224680 170956 224732
rect 171008 224720 171014 224732
rect 185302 224720 185308 224732
rect 171008 224692 185308 224720
rect 171008 224680 171014 224692
rect 185302 224680 185308 224692
rect 185360 224680 185366 224732
rect 187602 224680 187608 224732
rect 187660 224720 187666 224732
rect 202414 224720 202420 224732
rect 187660 224692 202420 224720
rect 187660 224680 187666 224692
rect 202414 224680 202420 224692
rect 202472 224680 202478 224732
rect 115842 224612 115848 224664
rect 115900 224652 115906 224664
rect 130746 224652 130752 224664
rect 115900 224624 126836 224652
rect 115900 224612 115906 224624
rect 113082 224544 113088 224596
rect 113140 224584 113146 224596
rect 126808 224584 126836 224624
rect 127728 224624 130752 224652
rect 127728 224584 127756 224624
rect 130746 224612 130752 224624
rect 130804 224612 130810 224664
rect 131022 224612 131028 224664
rect 131080 224652 131086 224664
rect 146754 224652 146760 224664
rect 131080 224624 146760 224652
rect 131080 224612 131086 224624
rect 146754 224612 146760 224624
rect 146812 224612 146818 224664
rect 147582 224612 147588 224664
rect 147640 224652 147646 224664
rect 162854 224652 162860 224664
rect 147640 224624 162860 224652
rect 147640 224612 147646 224624
rect 162854 224612 162860 224624
rect 162912 224612 162918 224664
rect 165430 224612 165436 224664
rect 165488 224652 165494 224664
rect 179966 224652 179972 224664
rect 165488 224624 179972 224652
rect 165488 224612 165494 224624
rect 179966 224612 179972 224624
rect 180024 224612 180030 224664
rect 186222 224612 186228 224664
rect 186280 224652 186286 224664
rect 201310 224652 201316 224664
rect 186280 224624 201316 224652
rect 186280 224612 186286 224624
rect 201310 224612 201316 224624
rect 201368 224612 201374 224664
rect 113140 224556 126652 224584
rect 126808 224556 127756 224584
rect 127805 224587 127863 224593
rect 113140 224544 113146 224556
rect 117222 224476 117228 224528
rect 117280 224516 117286 224528
rect 126333 224519 126391 224525
rect 126333 224516 126345 224519
rect 117280 224488 126345 224516
rect 117280 224476 117286 224488
rect 126333 224485 126345 224488
rect 126379 224485 126391 224519
rect 126333 224479 126391 224485
rect 113818 224408 113824 224460
rect 113876 224448 113882 224460
rect 126422 224448 126428 224460
rect 113876 224420 126428 224448
rect 113876 224408 113882 224420
rect 126422 224408 126428 224420
rect 126480 224408 126486 224460
rect 126624 224448 126652 224556
rect 127805 224553 127817 224587
rect 127851 224584 127863 224587
rect 129366 224584 129372 224596
rect 127851 224556 129372 224584
rect 127851 224553 127863 224556
rect 127805 224547 127863 224553
rect 129366 224544 129372 224556
rect 129424 224544 129430 224596
rect 132402 224544 132408 224596
rect 132460 224584 132466 224596
rect 147858 224584 147864 224596
rect 132460 224556 147864 224584
rect 132460 224544 132466 224556
rect 147858 224544 147864 224556
rect 147916 224544 147922 224596
rect 150342 224544 150348 224596
rect 150400 224584 150406 224596
rect 166074 224584 166080 224596
rect 150400 224556 166080 224584
rect 150400 224544 150406 224556
rect 166074 224544 166080 224556
rect 166132 224544 166138 224596
rect 175090 224544 175096 224596
rect 175148 224584 175154 224596
rect 189534 224584 189540 224596
rect 175148 224556 189540 224584
rect 175148 224544 175154 224556
rect 189534 224544 189540 224556
rect 189592 224544 189598 224596
rect 127713 224519 127771 224525
rect 127713 224485 127725 224519
rect 127759 224516 127771 224519
rect 133966 224516 133972 224528
rect 127759 224488 133972 224516
rect 127759 224485 127771 224488
rect 127713 224479 127771 224485
rect 133966 224476 133972 224488
rect 134024 224476 134030 224528
rect 137922 224476 137928 224528
rect 137980 224516 137986 224528
rect 153194 224516 153200 224528
rect 137980 224488 153200 224516
rect 137980 224476 137986 224488
rect 153194 224476 153200 224488
rect 153252 224476 153258 224528
rect 155862 224476 155868 224528
rect 155920 224516 155926 224528
rect 171410 224516 171416 224528
rect 155920 224488 171416 224516
rect 155920 224476 155926 224488
rect 171410 224476 171416 224488
rect 171468 224476 171474 224528
rect 184750 224476 184756 224528
rect 184808 224516 184814 224528
rect 199194 224516 199200 224528
rect 184808 224488 199200 224516
rect 184808 224476 184814 224488
rect 199194 224476 199200 224488
rect 199252 224476 199258 224528
rect 128630 224448 128636 224460
rect 126624 224420 128636 224448
rect 128630 224408 128636 224420
rect 128688 224408 128694 224460
rect 142522 224448 142528 224460
rect 128740 224420 142528 224448
rect 112438 224340 112444 224392
rect 112496 224380 112502 224392
rect 123202 224380 123208 224392
rect 112496 224352 123208 224380
rect 112496 224340 112502 224352
rect 123202 224340 123208 224352
rect 123260 224340 123266 224392
rect 126882 224340 126888 224392
rect 126940 224380 126946 224392
rect 128740 224380 128768 224420
rect 142522 224408 142528 224420
rect 142580 224408 142586 224460
rect 146202 224408 146208 224460
rect 146260 224448 146266 224460
rect 161750 224448 161756 224460
rect 146260 224420 161756 224448
rect 146260 224408 146266 224420
rect 161750 224408 161756 224420
rect 161808 224408 161814 224460
rect 175182 224408 175188 224460
rect 175240 224448 175246 224460
rect 190638 224448 190644 224460
rect 175240 224420 190644 224448
rect 175240 224408 175246 224420
rect 190638 224408 190644 224420
rect 190696 224408 190702 224460
rect 126940 224352 128768 224380
rect 128817 224383 128875 224389
rect 126940 224340 126946 224352
rect 128817 224349 128829 224383
rect 128863 224380 128875 224383
rect 141418 224380 141424 224392
rect 128863 224352 141424 224380
rect 128863 224349 128875 224352
rect 128817 224343 128875 224349
rect 141418 224340 141424 224352
rect 141476 224340 141482 224392
rect 142062 224340 142068 224392
rect 142120 224380 142126 224392
rect 157426 224380 157432 224392
rect 142120 224352 157432 224380
rect 142120 224340 142126 224352
rect 157426 224340 157432 224352
rect 157484 224340 157490 224392
rect 171042 224340 171048 224392
rect 171100 224380 171106 224392
rect 186314 224380 186320 224392
rect 171100 224352 186320 224380
rect 171100 224340 171106 224352
rect 186314 224340 186320 224352
rect 186372 224340 186378 224392
rect 188430 224340 188436 224392
rect 188488 224380 188494 224392
rect 203426 224380 203432 224392
rect 188488 224352 203432 224380
rect 188488 224340 188494 224352
rect 203426 224340 203432 224352
rect 203484 224340 203490 224392
rect 79318 224272 79324 224324
rect 79376 224312 79382 224324
rect 100294 224312 100300 224324
rect 79376 224284 100300 224312
rect 79376 224272 79382 224284
rect 100294 224272 100300 224284
rect 100352 224272 100358 224324
rect 115750 224272 115756 224324
rect 115808 224312 115814 224324
rect 131758 224312 131764 224324
rect 115808 224284 131764 224312
rect 115808 224272 115814 224284
rect 131758 224272 131764 224284
rect 131816 224272 131822 224324
rect 136450 224272 136456 224324
rect 136508 224312 136514 224324
rect 152090 224312 152096 224324
rect 136508 224284 152096 224312
rect 136508 224272 136514 224284
rect 152090 224272 152096 224284
rect 152148 224272 152154 224324
rect 165522 224272 165528 224324
rect 165580 224312 165586 224324
rect 180978 224312 180984 224324
rect 165580 224284 180984 224312
rect 165580 224272 165586 224284
rect 180978 224272 180984 224284
rect 181036 224272 181042 224324
rect 184842 224272 184848 224324
rect 184900 224312 184906 224324
rect 200298 224312 200304 224324
rect 184900 224284 200304 224312
rect 184900 224272 184906 224284
rect 200298 224272 200304 224284
rect 200356 224272 200362 224324
rect 3602 224204 3608 224256
rect 3660 224244 3666 224256
rect 120074 224244 120080 224256
rect 3660 224216 120080 224244
rect 3660 224204 3666 224216
rect 120074 224204 120080 224216
rect 120132 224204 120138 224256
rect 121270 224204 121276 224256
rect 121328 224244 121334 224256
rect 137186 224244 137192 224256
rect 121328 224216 137192 224244
rect 121328 224204 121334 224216
rect 137186 224204 137192 224216
rect 137244 224204 137250 224256
rect 140590 224204 140596 224256
rect 140648 224244 140654 224256
rect 156414 224244 156420 224256
rect 140648 224216 156420 224244
rect 140648 224204 140654 224216
rect 156414 224204 156420 224216
rect 156472 224204 156478 224256
rect 160002 224204 160008 224256
rect 160060 224244 160066 224256
rect 175642 224244 175648 224256
rect 160060 224216 175648 224244
rect 160060 224204 160066 224216
rect 175642 224204 175648 224216
rect 175700 224204 175706 224256
rect 180610 224204 180616 224256
rect 180668 224244 180674 224256
rect 195974 224244 195980 224256
rect 180668 224216 195980 224244
rect 180668 224204 180674 224216
rect 195974 224204 195980 224216
rect 196032 224204 196038 224256
rect 210970 224204 210976 224256
rect 211028 224244 211034 224256
rect 286318 224244 286324 224256
rect 211028 224216 286324 224244
rect 211028 224204 211034 224216
rect 286318 224204 286324 224216
rect 286376 224204 286382 224256
rect 118602 224136 118608 224188
rect 118660 224176 118666 224188
rect 127713 224179 127771 224185
rect 127713 224176 127725 224179
rect 118660 224148 127725 224176
rect 118660 224136 118666 224148
rect 127713 224145 127725 224148
rect 127759 224145 127771 224179
rect 140314 224176 140320 224188
rect 127713 224139 127771 224145
rect 127820 224148 140320 224176
rect 125226 224068 125232 224120
rect 125284 224108 125290 224120
rect 127820 224108 127848 224148
rect 140314 224136 140320 224148
rect 140372 224136 140378 224188
rect 144822 224136 144828 224188
rect 144880 224176 144886 224188
rect 159634 224176 159640 224188
rect 144880 224148 159640 224176
rect 144880 224136 144886 224148
rect 159634 224136 159640 224148
rect 159692 224136 159698 224188
rect 159910 224136 159916 224188
rect 159968 224176 159974 224188
rect 174630 224176 174636 224188
rect 159968 224148 174636 224176
rect 159968 224136 159974 224148
rect 174630 224136 174636 224148
rect 174688 224136 174694 224188
rect 177942 224136 177948 224188
rect 178000 224176 178006 224188
rect 192754 224176 192760 224188
rect 178000 224148 192760 224176
rect 178000 224136 178006 224148
rect 192754 224136 192760 224148
rect 192812 224136 192818 224188
rect 125284 224080 127848 224108
rect 128541 224111 128599 224117
rect 125284 224068 125290 224080
rect 128541 224077 128553 224111
rect 128587 224108 128599 224111
rect 139302 224108 139308 224120
rect 128587 224080 139308 224108
rect 128587 224077 128599 224080
rect 128541 224071 128599 224077
rect 139302 224068 139308 224080
rect 139360 224068 139366 224120
rect 140682 224068 140688 224120
rect 140740 224108 140746 224120
rect 155310 224108 155316 224120
rect 140740 224080 155316 224108
rect 140740 224068 140746 224080
rect 155310 224068 155316 224080
rect 155368 224068 155374 224120
rect 166902 224068 166908 224120
rect 166960 224108 166966 224120
rect 182082 224108 182088 224120
rect 166960 224080 182088 224108
rect 166960 224068 166966 224080
rect 182082 224068 182088 224080
rect 182140 224068 182146 224120
rect 182174 224068 182180 224120
rect 182232 224108 182238 224120
rect 197078 224108 197084 224120
rect 182232 224080 197084 224108
rect 182232 224068 182238 224080
rect 197078 224068 197084 224080
rect 197136 224068 197142 224120
rect 119982 224000 119988 224052
rect 120040 224040 120046 224052
rect 134978 224040 134984 224052
rect 120040 224012 134984 224040
rect 120040 224000 120046 224012
rect 134978 224000 134984 224012
rect 135036 224000 135042 224052
rect 136542 224000 136548 224052
rect 136600 224040 136606 224052
rect 151078 224040 151084 224052
rect 136600 224012 151084 224040
rect 136600 224000 136606 224012
rect 151078 224000 151084 224012
rect 151136 224000 151142 224052
rect 153102 224000 153108 224052
rect 153160 224040 153166 224052
rect 168190 224040 168196 224052
rect 153160 224012 168196 224040
rect 153160 224000 153166 224012
rect 168190 224000 168196 224012
rect 168248 224000 168254 224052
rect 169662 224000 169668 224052
rect 169720 224040 169726 224052
rect 184198 224040 184204 224052
rect 169720 224012 184204 224040
rect 169720 224000 169726 224012
rect 184198 224000 184204 224012
rect 184256 224000 184262 224052
rect 121362 223932 121368 223984
rect 121420 223972 121426 223984
rect 136082 223972 136088 223984
rect 121420 223944 136088 223972
rect 121420 223932 121426 223944
rect 136082 223932 136088 223944
rect 136140 223932 136146 223984
rect 143442 223932 143448 223984
rect 143500 223972 143506 223984
rect 158530 223972 158536 223984
rect 143500 223944 158536 223972
rect 143500 223932 143506 223944
rect 158530 223932 158536 223944
rect 158588 223932 158594 223984
rect 158622 223932 158628 223984
rect 158680 223972 158686 223984
rect 173526 223972 173532 223984
rect 158680 223944 173532 223972
rect 158680 223932 158686 223944
rect 173526 223932 173532 223944
rect 173584 223932 173590 223984
rect 173802 223932 173808 223984
rect 173860 223972 173866 223984
rect 188522 223972 188528 223984
rect 173860 223944 188528 223972
rect 173860 223932 173866 223944
rect 188522 223932 188528 223944
rect 188580 223932 188586 223984
rect 117958 223864 117964 223916
rect 118016 223904 118022 223916
rect 127526 223904 127532 223916
rect 118016 223876 127532 223904
rect 118016 223864 118022 223876
rect 127526 223864 127532 223876
rect 127584 223864 127590 223916
rect 139394 223864 139400 223916
rect 139452 223904 139458 223916
rect 154298 223904 154304 223916
rect 139452 223876 154304 223904
rect 139452 223864 139458 223876
rect 154298 223864 154304 223876
rect 154356 223864 154362 223916
rect 162762 223864 162768 223916
rect 162820 223904 162826 223916
rect 177758 223904 177764 223916
rect 162820 223876 177764 223904
rect 162820 223864 162826 223876
rect 177758 223864 177764 223876
rect 177816 223864 177822 223916
rect 124122 223796 124128 223848
rect 124180 223836 124186 223848
rect 128541 223839 128599 223845
rect 128541 223836 128553 223839
rect 124180 223808 128553 223836
rect 124180 223796 124186 223808
rect 128541 223805 128553 223808
rect 128587 223805 128599 223839
rect 128541 223799 128599 223805
rect 135162 223796 135168 223848
rect 135220 223836 135226 223848
rect 149974 223836 149980 223848
rect 135220 223808 149980 223836
rect 135220 223796 135226 223808
rect 149974 223796 149980 223808
rect 150032 223796 150038 223848
rect 154482 223796 154488 223848
rect 154540 223836 154546 223848
rect 169202 223836 169208 223848
rect 154540 223808 169208 223836
rect 154540 223796 154546 223808
rect 169202 223796 169208 223808
rect 169260 223796 169266 223848
rect 176562 223796 176568 223848
rect 176620 223836 176626 223848
rect 191742 223836 191748 223848
rect 176620 223808 191748 223836
rect 176620 223796 176626 223808
rect 191742 223796 191748 223808
rect 191800 223796 191806 223848
rect 133782 223728 133788 223780
rect 133840 223768 133846 223780
rect 148870 223768 148876 223780
rect 133840 223740 148876 223768
rect 133840 223728 133846 223740
rect 148870 223728 148876 223740
rect 148928 223728 148934 223780
rect 148962 223728 148968 223780
rect 149020 223768 149026 223780
rect 163866 223768 163872 223780
rect 149020 223740 163872 223768
rect 149020 223728 149026 223740
rect 163866 223728 163872 223740
rect 163924 223728 163930 223780
rect 168282 223728 168288 223780
rect 168340 223768 168346 223780
rect 183186 223768 183192 223780
rect 168340 223740 183192 223768
rect 168340 223728 168346 223740
rect 183186 223728 183192 223740
rect 183244 223728 183250 223780
rect 129642 223660 129648 223712
rect 129700 223700 129706 223712
rect 144638 223700 144644 223712
rect 129700 223672 144644 223700
rect 129700 223660 129706 223672
rect 144638 223660 144644 223672
rect 144696 223660 144702 223712
rect 157242 223660 157248 223712
rect 157300 223700 157306 223712
rect 172422 223700 172428 223712
rect 157300 223672 172428 223700
rect 157300 223660 157306 223672
rect 172422 223660 172428 223672
rect 172480 223660 172486 223712
rect 172514 223660 172520 223712
rect 172572 223700 172578 223712
rect 187418 223700 187424 223712
rect 172572 223672 187424 223700
rect 172572 223660 172578 223672
rect 187418 223660 187424 223672
rect 187476 223660 187482 223712
rect 3510 223592 3516 223644
rect 3568 223632 3574 223644
rect 121086 223632 121092 223644
rect 3568 223604 121092 223632
rect 3568 223592 3574 223604
rect 121086 223592 121092 223604
rect 121144 223592 121150 223644
rect 229738 223592 229744 223644
rect 229796 223632 229802 223644
rect 283374 223632 283380 223644
rect 229796 223604 283380 223632
rect 229796 223592 229802 223604
rect 283374 223592 283380 223604
rect 283432 223592 283438 223644
rect 231118 222912 231124 222964
rect 231176 222952 231182 222964
rect 245562 222952 245568 222964
rect 231176 222924 245568 222952
rect 231176 222912 231182 222924
rect 245562 222912 245568 222924
rect 245620 222912 245626 222964
rect 229002 222844 229008 222896
rect 229060 222884 229066 222896
rect 313918 222884 313924 222896
rect 229060 222856 313924 222884
rect 229060 222844 229066 222856
rect 313918 222844 313924 222856
rect 313976 222844 313982 222896
rect 214466 222204 214472 222216
rect 214427 222176 214472 222204
rect 214466 222164 214472 222176
rect 214524 222164 214530 222216
rect 214466 222068 214472 222080
rect 214427 222040 214472 222068
rect 214466 222028 214472 222040
rect 214524 222028 214530 222080
rect 55214 220804 55220 220856
rect 55272 220844 55278 220856
rect 116394 220844 116400 220856
rect 55272 220816 116400 220844
rect 55272 220804 55278 220816
rect 116394 220804 116400 220816
rect 116452 220804 116458 220856
rect 213914 220804 213920 220856
rect 213972 220844 213978 220856
rect 226334 220844 226340 220856
rect 213972 220816 226340 220844
rect 213972 220804 213978 220816
rect 226334 220804 226340 220816
rect 226392 220804 226398 220856
rect 214006 220124 214012 220176
rect 214064 220164 214070 220176
rect 226334 220164 226340 220176
rect 214064 220136 226340 220164
rect 214064 220124 214070 220136
rect 226334 220124 226340 220136
rect 226392 220124 226398 220176
rect 14458 220056 14464 220108
rect 14516 220096 14522 220108
rect 116670 220096 116676 220108
rect 14516 220068 116676 220096
rect 14516 220056 14522 220068
rect 116670 220056 116676 220068
rect 116728 220056 116734 220108
rect 213914 220056 213920 220108
rect 213972 220096 213978 220108
rect 226426 220096 226432 220108
rect 213972 220068 226432 220096
rect 213972 220056 213978 220068
rect 226426 220056 226432 220068
rect 226484 220056 226490 220108
rect 116118 219484 116124 219496
rect 114572 219456 116124 219484
rect 104802 219376 104808 219428
rect 104860 219416 104866 219428
rect 114572 219416 114600 219456
rect 116118 219444 116124 219456
rect 116176 219444 116182 219496
rect 104860 219388 114600 219416
rect 104860 219376 104866 219388
rect 213914 218764 213920 218816
rect 213972 218804 213978 218816
rect 226334 218804 226340 218816
rect 213972 218776 226340 218804
rect 213972 218764 213978 218776
rect 226334 218764 226340 218776
rect 226392 218764 226398 218816
rect 214006 218696 214012 218748
rect 214064 218736 214070 218748
rect 226426 218736 226432 218748
rect 214064 218708 226432 218736
rect 214064 218696 214070 218708
rect 226426 218696 226432 218708
rect 226484 218696 226490 218748
rect 116394 218056 116400 218068
rect 114480 218028 116400 218056
rect 104802 217948 104808 218000
rect 104860 217988 104866 218000
rect 114480 217988 114508 218028
rect 116394 218016 116400 218028
rect 116452 218016 116458 218068
rect 104860 217960 114508 217988
rect 104860 217948 104866 217960
rect 213914 217268 213920 217320
rect 213972 217308 213978 217320
rect 226334 217308 226340 217320
rect 213972 217280 226340 217308
rect 213972 217268 213978 217280
rect 226334 217268 226340 217280
rect 226392 217268 226398 217320
rect 104802 216588 104808 216640
rect 104860 216628 104866 216640
rect 116394 216628 116400 216640
rect 104860 216600 116400 216628
rect 104860 216588 104866 216600
rect 116394 216588 116400 216600
rect 116452 216588 116458 216640
rect 213914 216588 213920 216640
rect 213972 216628 213978 216640
rect 226426 216628 226432 216640
rect 213972 216600 226432 216628
rect 213972 216588 213978 216600
rect 226426 216588 226432 216600
rect 226484 216588 226490 216640
rect 104802 215908 104808 215960
rect 104860 215948 104866 215960
rect 115934 215948 115940 215960
rect 104860 215920 115940 215948
rect 104860 215908 104866 215920
rect 115934 215908 115940 215920
rect 115992 215908 115998 215960
rect 213914 215908 213920 215960
rect 213972 215948 213978 215960
rect 226334 215948 226340 215960
rect 213972 215920 226340 215948
rect 213972 215908 213978 215920
rect 226334 215908 226340 215920
rect 226392 215908 226398 215960
rect 116394 215336 116400 215348
rect 114480 215308 116400 215336
rect 104802 215228 104808 215280
rect 104860 215268 104866 215280
rect 114480 215268 114508 215308
rect 116394 215296 116400 215308
rect 116452 215296 116458 215348
rect 104860 215240 114508 215268
rect 104860 215228 104866 215240
rect 213914 215228 213920 215280
rect 213972 215268 213978 215280
rect 226426 215268 226432 215280
rect 213972 215240 226432 215268
rect 213972 215228 213978 215240
rect 226426 215228 226432 215240
rect 226484 215228 226490 215280
rect 214006 215160 214012 215212
rect 214064 215200 214070 215212
rect 226334 215200 226340 215212
rect 214064 215172 226340 215200
rect 214064 215160 214070 215172
rect 226334 215160 226340 215172
rect 226392 215160 226398 215212
rect 116394 213976 116400 213988
rect 113928 213948 116400 213976
rect 104802 213868 104808 213920
rect 104860 213908 104866 213920
rect 113928 213908 113956 213948
rect 116394 213936 116400 213948
rect 116452 213936 116458 213988
rect 104860 213880 113956 213908
rect 104860 213868 104866 213880
rect 213914 213868 213920 213920
rect 213972 213908 213978 213920
rect 226426 213908 226432 213920
rect 213972 213880 226432 213908
rect 213972 213868 213978 213880
rect 226426 213868 226432 213880
rect 226484 213868 226490 213920
rect 214006 213800 214012 213852
rect 214064 213840 214070 213852
rect 226334 213840 226340 213852
rect 214064 213812 226340 213840
rect 214064 213800 214070 213812
rect 226334 213800 226340 213812
rect 226392 213800 226398 213852
rect 115934 212548 115940 212560
rect 114480 212520 115940 212548
rect 104434 212440 104440 212492
rect 104492 212480 104498 212492
rect 114480 212480 114508 212520
rect 115934 212508 115940 212520
rect 115992 212508 115998 212560
rect 214469 212551 214527 212557
rect 214469 212517 214481 212551
rect 214515 212548 214527 212551
rect 214558 212548 214564 212560
rect 214515 212520 214564 212548
rect 214515 212517 214527 212520
rect 214469 212511 214527 212517
rect 214558 212508 214564 212520
rect 214616 212508 214622 212560
rect 104492 212452 114508 212480
rect 104492 212440 104498 212452
rect 213914 212440 213920 212492
rect 213972 212480 213978 212492
rect 226426 212480 226432 212492
rect 213972 212452 226432 212480
rect 213972 212440 213978 212452
rect 226426 212440 226432 212452
rect 226484 212440 226490 212492
rect 214006 212372 214012 212424
rect 214064 212412 214070 212424
rect 226334 212412 226340 212424
rect 214064 212384 226340 212412
rect 214064 212372 214070 212384
rect 226334 212372 226340 212384
rect 226392 212372 226398 212424
rect 116302 211188 116308 211200
rect 114480 211160 116308 211188
rect 104802 211080 104808 211132
rect 104860 211120 104866 211132
rect 114480 211120 114508 211160
rect 116302 211148 116308 211160
rect 116360 211148 116366 211200
rect 104860 211092 114508 211120
rect 104860 211080 104866 211092
rect 213914 211080 213920 211132
rect 213972 211120 213978 211132
rect 226518 211120 226524 211132
rect 213972 211092 226524 211120
rect 213972 211080 213978 211092
rect 226518 211080 226524 211092
rect 226576 211080 226582 211132
rect 116302 209828 116308 209840
rect 113192 209800 116308 209828
rect 104802 209720 104808 209772
rect 104860 209760 104866 209772
rect 113192 209760 113220 209800
rect 116302 209788 116308 209800
rect 116360 209788 116366 209840
rect 104860 209732 113220 209760
rect 104860 209720 104866 209732
rect 214006 209720 214012 209772
rect 214064 209760 214070 209772
rect 226242 209760 226248 209772
rect 214064 209732 226248 209760
rect 214064 209720 214070 209732
rect 226242 209720 226248 209732
rect 226300 209720 226306 209772
rect 213914 209652 213920 209704
rect 213972 209692 213978 209704
rect 226058 209692 226064 209704
rect 213972 209664 226064 209692
rect 213972 209652 213978 209664
rect 226058 209652 226064 209664
rect 226116 209652 226122 209704
rect 116026 208400 116032 208412
rect 114480 208372 116032 208400
rect 104802 208292 104808 208344
rect 104860 208332 104866 208344
rect 114480 208332 114508 208372
rect 116026 208360 116032 208372
rect 116084 208360 116090 208412
rect 104860 208304 114508 208332
rect 104860 208292 104866 208304
rect 214006 208292 214012 208344
rect 214064 208332 214070 208344
rect 226150 208332 226156 208344
rect 214064 208304 226156 208332
rect 214064 208292 214070 208304
rect 226150 208292 226156 208304
rect 226208 208292 226214 208344
rect 213914 208224 213920 208276
rect 213972 208264 213978 208276
rect 225966 208264 225972 208276
rect 213972 208236 225972 208264
rect 213972 208224 213978 208236
rect 225966 208224 225972 208236
rect 226024 208224 226030 208276
rect 113818 207068 113824 207120
rect 113876 207108 113882 207120
rect 116394 207108 116400 207120
rect 113876 207080 116400 207108
rect 113876 207068 113882 207080
rect 116394 207068 116400 207080
rect 116452 207068 116458 207120
rect 116302 207040 116308 207052
rect 114480 207012 116308 207040
rect 104710 206932 104716 206984
rect 104768 206972 104774 206984
rect 114480 206972 114508 207012
rect 116302 207000 116308 207012
rect 116360 207000 116366 207052
rect 104768 206944 114508 206972
rect 104768 206932 104774 206944
rect 213914 206932 213920 206984
rect 213972 206972 213978 206984
rect 226058 206972 226064 206984
rect 213972 206944 226064 206972
rect 213972 206932 213978 206944
rect 226058 206932 226064 206944
rect 226116 206932 226122 206984
rect 104802 206864 104808 206916
rect 104860 206904 104866 206916
rect 113818 206904 113824 206916
rect 104860 206876 113824 206904
rect 104860 206864 104866 206876
rect 113818 206864 113824 206876
rect 113876 206864 113882 206916
rect 214006 206864 214012 206916
rect 214064 206904 214070 206916
rect 226242 206904 226248 206916
rect 214064 206876 226248 206904
rect 214064 206864 214070 206876
rect 226242 206864 226248 206876
rect 226300 206864 226306 206916
rect 115934 205680 115940 205692
rect 114480 205652 115940 205680
rect 104802 205572 104808 205624
rect 104860 205612 104866 205624
rect 114480 205612 114508 205652
rect 115934 205640 115940 205652
rect 115992 205640 115998 205692
rect 214466 205680 214472 205692
rect 214427 205652 214472 205680
rect 214466 205640 214472 205652
rect 214524 205640 214530 205692
rect 104860 205584 114508 205612
rect 104860 205572 104866 205584
rect 213914 205572 213920 205624
rect 213972 205612 213978 205624
rect 226150 205612 226156 205624
rect 213972 205584 226156 205612
rect 213972 205572 213978 205584
rect 226150 205572 226156 205584
rect 226208 205572 226214 205624
rect 116394 204320 116400 204332
rect 114480 204292 116400 204320
rect 104802 204212 104808 204264
rect 104860 204252 104866 204264
rect 114480 204252 114508 204292
rect 116394 204280 116400 204292
rect 116452 204280 116458 204332
rect 104860 204224 114508 204252
rect 104860 204212 104866 204224
rect 214006 204212 214012 204264
rect 214064 204252 214070 204264
rect 225966 204252 225972 204264
rect 214064 204224 225972 204252
rect 214064 204212 214070 204224
rect 225966 204212 225972 204224
rect 226024 204212 226030 204264
rect 213914 204144 213920 204196
rect 213972 204184 213978 204196
rect 225782 204184 225788 204196
rect 213972 204156 225788 204184
rect 213972 204144 213978 204156
rect 225782 204144 225788 204156
rect 225840 204144 225846 204196
rect 116302 202892 116308 202904
rect 114480 202864 116308 202892
rect 104802 202784 104808 202836
rect 104860 202824 104866 202836
rect 114480 202824 114508 202864
rect 116302 202852 116308 202864
rect 116360 202852 116366 202904
rect 214466 202892 214472 202904
rect 214427 202864 214472 202892
rect 214466 202852 214472 202864
rect 214524 202852 214530 202904
rect 104860 202796 114508 202824
rect 104860 202784 104866 202796
rect 213914 202784 213920 202836
rect 213972 202824 213978 202836
rect 225874 202824 225880 202836
rect 213972 202796 225880 202824
rect 213972 202784 213978 202796
rect 225874 202784 225880 202796
rect 225932 202784 225938 202836
rect 214006 202716 214012 202768
rect 214064 202756 214070 202768
rect 226150 202756 226156 202768
rect 214064 202728 226156 202756
rect 214064 202716 214070 202728
rect 226150 202716 226156 202728
rect 226208 202716 226214 202768
rect 116118 201532 116124 201544
rect 114480 201504 116124 201532
rect 104802 201424 104808 201476
rect 104860 201464 104866 201476
rect 114480 201464 114508 201504
rect 116118 201492 116124 201504
rect 116176 201492 116182 201544
rect 104860 201436 114508 201464
rect 104860 201424 104866 201436
rect 213914 201424 213920 201476
rect 213972 201464 213978 201476
rect 225598 201464 225604 201476
rect 213972 201436 225604 201464
rect 213972 201424 213978 201436
rect 225598 201424 225604 201436
rect 225656 201424 225662 201476
rect 214006 201356 214012 201408
rect 214064 201396 214070 201408
rect 225690 201396 225696 201408
rect 214064 201368 225696 201396
rect 214064 201356 214070 201368
rect 225690 201356 225696 201368
rect 225748 201356 225754 201408
rect 214466 200540 214472 200592
rect 214524 200580 214530 200592
rect 214834 200580 214840 200592
rect 214524 200552 214840 200580
rect 214524 200540 214530 200552
rect 214834 200540 214840 200552
rect 214892 200540 214898 200592
rect 116118 200240 116124 200252
rect 113192 200212 116124 200240
rect 104802 200064 104808 200116
rect 104860 200104 104866 200116
rect 113192 200104 113220 200212
rect 116118 200200 116124 200212
rect 116176 200200 116182 200252
rect 113266 200132 113272 200184
rect 113324 200172 113330 200184
rect 115934 200172 115940 200184
rect 113324 200144 115940 200172
rect 113324 200132 113330 200144
rect 115934 200132 115940 200144
rect 115992 200132 115998 200184
rect 104860 200076 113220 200104
rect 104860 200064 104866 200076
rect 213914 200064 213920 200116
rect 213972 200104 213978 200116
rect 226242 200104 226248 200116
rect 213972 200076 226248 200104
rect 213972 200064 213978 200076
rect 226242 200064 226248 200076
rect 226300 200064 226306 200116
rect 224126 198772 224132 198824
rect 224184 198812 224190 198824
rect 226426 198812 226432 198824
rect 224184 198784 226432 198812
rect 224184 198772 224190 198784
rect 226426 198772 226432 198784
rect 226484 198772 226490 198824
rect 114462 198704 114468 198756
rect 114520 198744 114526 198756
rect 115934 198744 115940 198756
rect 114520 198716 115940 198744
rect 114520 198704 114526 198716
rect 115934 198704 115940 198716
rect 115992 198704 115998 198756
rect 223942 198704 223948 198756
rect 224000 198744 224006 198756
rect 226334 198744 226340 198756
rect 224000 198716 226340 198744
rect 224000 198704 224006 198716
rect 226334 198704 226340 198716
rect 226392 198704 226398 198756
rect 104802 198636 104808 198688
rect 104860 198676 104866 198688
rect 113266 198676 113272 198688
rect 104860 198648 113272 198676
rect 104860 198636 104866 198648
rect 113266 198636 113272 198648
rect 113324 198636 113330 198688
rect 214006 198636 214012 198688
rect 214064 198676 214070 198688
rect 225966 198676 225972 198688
rect 214064 198648 225972 198676
rect 214064 198636 214070 198648
rect 225966 198636 225972 198648
rect 226024 198636 226030 198688
rect 213914 198568 213920 198620
rect 213972 198608 213978 198620
rect 226058 198608 226064 198620
rect 213972 198580 226064 198608
rect 213972 198568 213978 198580
rect 226058 198568 226064 198580
rect 226116 198568 226122 198620
rect 224494 197412 224500 197464
rect 224552 197452 224558 197464
rect 226426 197452 226432 197464
rect 224552 197424 226432 197452
rect 224552 197412 224558 197424
rect 226426 197412 226432 197424
rect 226484 197412 226490 197464
rect 116118 197384 116124 197396
rect 114480 197356 116124 197384
rect 104710 197276 104716 197328
rect 104768 197316 104774 197328
rect 114480 197316 114508 197356
rect 116118 197344 116124 197356
rect 116176 197344 116182 197396
rect 224034 197344 224040 197396
rect 224092 197384 224098 197396
rect 226334 197384 226340 197396
rect 224092 197356 226340 197384
rect 224092 197344 224098 197356
rect 226334 197344 226340 197356
rect 226392 197344 226398 197396
rect 104768 197288 114508 197316
rect 104768 197276 104774 197288
rect 214006 197276 214012 197328
rect 214064 197316 214070 197328
rect 226150 197316 226156 197328
rect 214064 197288 226156 197316
rect 214064 197276 214070 197288
rect 226150 197276 226156 197288
rect 226208 197276 226214 197328
rect 104802 197208 104808 197260
rect 104860 197248 104866 197260
rect 114462 197248 114468 197260
rect 104860 197220 114468 197248
rect 104860 197208 104866 197220
rect 114462 197208 114468 197220
rect 114520 197208 114526 197260
rect 213914 197208 213920 197260
rect 213972 197248 213978 197260
rect 225782 197248 225788 197260
rect 213972 197220 225788 197248
rect 213972 197208 213978 197220
rect 225782 197208 225788 197220
rect 225840 197208 225846 197260
rect 224310 196052 224316 196104
rect 224368 196092 224374 196104
rect 226334 196092 226340 196104
rect 224368 196064 226340 196092
rect 224368 196052 224374 196064
rect 226334 196052 226340 196064
rect 226392 196052 226398 196104
rect 116394 196024 116400 196036
rect 114296 195996 116400 196024
rect 104802 195916 104808 195968
rect 104860 195956 104866 195968
rect 114296 195956 114324 195996
rect 116394 195984 116400 195996
rect 116452 195984 116458 196036
rect 224402 195984 224408 196036
rect 224460 196024 224466 196036
rect 226702 196024 226708 196036
rect 224460 195996 226708 196024
rect 224460 195984 224466 195996
rect 226702 195984 226708 195996
rect 226760 195984 226766 196036
rect 104860 195928 114324 195956
rect 104860 195916 104866 195928
rect 213914 195916 213920 195968
rect 213972 195956 213978 195968
rect 226242 195956 226248 195968
rect 213972 195928 226248 195956
rect 213972 195916 213978 195928
rect 226242 195916 226248 195928
rect 226300 195916 226306 195968
rect 214006 195848 214012 195900
rect 214064 195888 214070 195900
rect 225874 195888 225880 195900
rect 214064 195860 225880 195888
rect 214064 195848 214070 195860
rect 225874 195848 225880 195860
rect 225932 195848 225938 195900
rect 224218 194692 224224 194744
rect 224276 194732 224282 194744
rect 226518 194732 226524 194744
rect 224276 194704 226524 194732
rect 224276 194692 224282 194704
rect 226518 194692 226524 194704
rect 226576 194692 226582 194744
rect 221458 194624 221464 194676
rect 221516 194664 221522 194676
rect 226426 194664 226432 194676
rect 221516 194636 226432 194664
rect 221516 194624 221522 194636
rect 226426 194624 226432 194636
rect 226484 194624 226490 194676
rect 115934 194596 115940 194608
rect 114480 194568 115940 194596
rect 104802 194488 104808 194540
rect 104860 194528 104866 194540
rect 114480 194528 114508 194568
rect 115934 194556 115940 194568
rect 115992 194556 115998 194608
rect 214190 194556 214196 194608
rect 214248 194596 214254 194608
rect 226334 194596 226340 194608
rect 214248 194568 226340 194596
rect 214248 194556 214254 194568
rect 226334 194556 226340 194568
rect 226392 194556 226398 194608
rect 104860 194500 114508 194528
rect 104860 194488 104866 194500
rect 213914 194488 213920 194540
rect 213972 194528 213978 194540
rect 225690 194528 225696 194540
rect 213972 194500 225696 194528
rect 213972 194488 213978 194500
rect 225690 194488 225696 194500
rect 225748 194488 225754 194540
rect 220078 193264 220084 193316
rect 220136 193304 220142 193316
rect 226426 193304 226432 193316
rect 220136 193276 226432 193304
rect 220136 193264 220142 193276
rect 226426 193264 226432 193276
rect 226484 193264 226490 193316
rect 116118 193236 116124 193248
rect 114480 193208 116124 193236
rect 104434 193128 104440 193180
rect 104492 193168 104498 193180
rect 114480 193168 114508 193208
rect 116118 193196 116124 193208
rect 116176 193196 116182 193248
rect 214466 193196 214472 193248
rect 214524 193236 214530 193248
rect 226334 193236 226340 193248
rect 214524 193208 226340 193236
rect 214524 193196 214530 193208
rect 226334 193196 226340 193208
rect 226392 193196 226398 193248
rect 104492 193140 114508 193168
rect 104492 193128 104498 193140
rect 213914 193128 213920 193180
rect 213972 193168 213978 193180
rect 224126 193168 224132 193180
rect 213972 193140 224132 193168
rect 213972 193128 213978 193140
rect 224126 193128 224132 193140
rect 224184 193128 224190 193180
rect 214006 193060 214012 193112
rect 214064 193100 214070 193112
rect 223942 193100 223948 193112
rect 214064 193072 223948 193100
rect 214064 193060 214070 193072
rect 223942 193060 223948 193072
rect 224000 193060 224006 193112
rect 113910 191972 113916 192024
rect 113968 192012 113974 192024
rect 116394 192012 116400 192024
rect 113968 191984 116400 192012
rect 113968 191972 113974 191984
rect 116394 191972 116400 191984
rect 116452 191972 116458 192024
rect 113174 191904 113180 191956
rect 113232 191944 113238 191956
rect 116026 191944 116032 191956
rect 113232 191916 116032 191944
rect 113232 191904 113238 191916
rect 116026 191904 116032 191916
rect 116084 191904 116090 191956
rect 215294 191904 215300 191956
rect 215352 191944 215358 191956
rect 226334 191944 226340 191956
rect 215352 191916 226340 191944
rect 215352 191904 215358 191916
rect 226334 191904 226340 191916
rect 226392 191904 226398 191956
rect 214098 191836 214104 191888
rect 214156 191876 214162 191888
rect 226426 191876 226432 191888
rect 214156 191848 226432 191876
rect 214156 191836 214162 191848
rect 226426 191836 226432 191848
rect 226484 191836 226490 191888
rect 104434 191768 104440 191820
rect 104492 191808 104498 191820
rect 113910 191808 113916 191820
rect 104492 191780 113916 191808
rect 104492 191768 104498 191780
rect 113910 191768 113916 191780
rect 113968 191768 113974 191820
rect 214006 191768 214012 191820
rect 214064 191808 214070 191820
rect 224034 191808 224040 191820
rect 214064 191780 224040 191808
rect 214064 191768 214070 191780
rect 224034 191768 224040 191780
rect 224092 191768 224098 191820
rect 213914 191700 213920 191752
rect 213972 191740 213978 191752
rect 224494 191740 224500 191752
rect 213972 191712 224500 191740
rect 213972 191700 213978 191712
rect 224494 191700 224500 191712
rect 224552 191700 224558 191752
rect 113266 190612 113272 190664
rect 113324 190652 113330 190664
rect 116486 190652 116492 190664
rect 113324 190624 116492 190652
rect 113324 190612 113330 190624
rect 116486 190612 116492 190624
rect 116544 190612 116550 190664
rect 214282 190544 214288 190596
rect 214340 190584 214346 190596
rect 226334 190584 226340 190596
rect 214340 190556 226340 190584
rect 214340 190544 214346 190556
rect 226334 190544 226340 190556
rect 226392 190544 226398 190596
rect 215018 190476 215024 190528
rect 215076 190516 215082 190528
rect 226426 190516 226432 190528
rect 215076 190488 226432 190516
rect 215076 190476 215082 190488
rect 226426 190476 226432 190488
rect 226484 190476 226490 190528
rect 104710 190408 104716 190460
rect 104768 190448 104774 190460
rect 113174 190448 113180 190460
rect 104768 190420 113180 190448
rect 104768 190408 104774 190420
rect 113174 190408 113180 190420
rect 113232 190408 113238 190460
rect 214006 190408 214012 190460
rect 214064 190448 214070 190460
rect 224402 190448 224408 190460
rect 214064 190420 224408 190448
rect 214064 190408 214070 190420
rect 224402 190408 224408 190420
rect 224460 190408 224466 190460
rect 213914 190340 213920 190392
rect 213972 190380 213978 190392
rect 224310 190380 224316 190392
rect 213972 190352 224316 190380
rect 213972 190340 213978 190352
rect 224310 190340 224316 190352
rect 224368 190340 224374 190392
rect 218698 189116 218704 189168
rect 218756 189156 218762 189168
rect 226426 189156 226432 189168
rect 218756 189128 226432 189156
rect 218756 189116 218762 189128
rect 226426 189116 226432 189128
rect 226484 189116 226490 189168
rect 114462 189048 114468 189100
rect 114520 189088 114526 189100
rect 116394 189088 116400 189100
rect 114520 189060 116400 189088
rect 114520 189048 114526 189060
rect 116394 189048 116400 189060
rect 116452 189048 116458 189100
rect 214374 189048 214380 189100
rect 214432 189088 214438 189100
rect 226334 189088 226340 189100
rect 214432 189060 226340 189088
rect 214432 189048 214438 189060
rect 226334 189048 226340 189060
rect 226392 189048 226398 189100
rect 104802 188980 104808 189032
rect 104860 189020 104866 189032
rect 113266 189020 113272 189032
rect 104860 188992 113272 189020
rect 104860 188980 104866 188992
rect 113266 188980 113272 188992
rect 113324 188980 113330 189032
rect 213914 188980 213920 189032
rect 213972 189020 213978 189032
rect 224218 189020 224224 189032
rect 213972 188992 224224 189020
rect 213972 188980 213978 188992
rect 224218 188980 224224 188992
rect 224276 188980 224282 189032
rect 222930 187756 222936 187808
rect 222988 187796 222994 187808
rect 226426 187796 226432 187808
rect 222988 187768 226432 187796
rect 222988 187756 222994 187768
rect 226426 187756 226432 187768
rect 226484 187756 226490 187808
rect 114094 187688 114100 187740
rect 114152 187728 114158 187740
rect 116394 187728 116400 187740
rect 114152 187700 116400 187728
rect 114152 187688 114158 187700
rect 116394 187688 116400 187700
rect 116452 187688 116458 187740
rect 215938 187688 215944 187740
rect 215996 187728 216002 187740
rect 226334 187728 226340 187740
rect 215996 187700 226340 187728
rect 215996 187688 216002 187700
rect 226334 187688 226340 187700
rect 226392 187688 226398 187740
rect 104802 187620 104808 187672
rect 104860 187660 104866 187672
rect 114462 187660 114468 187672
rect 104860 187632 114468 187660
rect 104860 187620 104866 187632
rect 114462 187620 114468 187632
rect 114520 187620 114526 187672
rect 213914 186532 213920 186584
rect 213972 186572 213978 186584
rect 221458 186572 221464 186584
rect 213972 186544 221464 186572
rect 213972 186532 213978 186544
rect 221458 186532 221464 186544
rect 221516 186532 221522 186584
rect 224402 186396 224408 186448
rect 224460 186436 224466 186448
rect 226426 186436 226432 186448
rect 224460 186408 226432 186436
rect 224460 186396 224466 186408
rect 226426 186396 226432 186408
rect 226484 186396 226490 186448
rect 115934 186368 115940 186380
rect 114480 186340 115940 186368
rect 104710 186260 104716 186312
rect 104768 186300 104774 186312
rect 114480 186300 114508 186340
rect 115934 186328 115940 186340
rect 115992 186328 115998 186380
rect 214190 186328 214196 186380
rect 214248 186368 214254 186380
rect 226334 186368 226340 186380
rect 214248 186340 226340 186368
rect 214248 186328 214254 186340
rect 226334 186328 226340 186340
rect 226392 186328 226398 186380
rect 104768 186272 114508 186300
rect 104768 186260 104774 186272
rect 104802 186192 104808 186244
rect 104860 186232 104866 186244
rect 114094 186232 114100 186244
rect 104860 186204 114100 186232
rect 104860 186192 104866 186204
rect 114094 186192 114100 186204
rect 114152 186192 114158 186244
rect 213914 185036 213920 185088
rect 213972 185076 213978 185088
rect 220078 185076 220084 185088
rect 213972 185048 220084 185076
rect 213972 185036 213978 185048
rect 220078 185036 220084 185048
rect 220136 185036 220142 185088
rect 114462 184968 114468 185020
rect 114520 185008 114526 185020
rect 116394 185008 116400 185020
rect 114520 184980 116400 185008
rect 114520 184968 114526 184980
rect 116394 184968 116400 184980
rect 116452 184968 116458 185020
rect 220170 184968 220176 185020
rect 220228 185008 220234 185020
rect 226426 185008 226432 185020
rect 220228 184980 226432 185008
rect 220228 184968 220234 184980
rect 226426 184968 226432 184980
rect 226484 184968 226490 185020
rect 116026 184940 116032 184952
rect 114480 184912 116032 184940
rect 104802 184832 104808 184884
rect 104860 184872 104866 184884
rect 114480 184872 114508 184912
rect 116026 184900 116032 184912
rect 116084 184900 116090 184952
rect 214006 184900 214012 184952
rect 214064 184940 214070 184952
rect 226334 184940 226340 184952
rect 214064 184912 226340 184940
rect 214064 184900 214070 184912
rect 226334 184900 226340 184912
rect 226392 184900 226398 184952
rect 104860 184844 114508 184872
rect 104860 184832 104866 184844
rect 215294 184152 215300 184204
rect 215352 184192 215358 184204
rect 226518 184192 226524 184204
rect 215352 184164 226524 184192
rect 215352 184152 215358 184164
rect 226518 184152 226524 184164
rect 226576 184152 226582 184204
rect 114370 183540 114376 183592
rect 114428 183580 114434 183592
rect 116394 183580 116400 183592
rect 114428 183552 116400 183580
rect 114428 183540 114434 183552
rect 116394 183540 116400 183552
rect 116452 183540 116458 183592
rect 213914 183540 213920 183592
rect 213972 183580 213978 183592
rect 226334 183580 226340 183592
rect 213972 183552 226340 183580
rect 213972 183540 213978 183552
rect 226334 183540 226340 183552
rect 226392 183540 226398 183592
rect 104802 183472 104808 183524
rect 104860 183512 104866 183524
rect 114462 183512 114468 183524
rect 104860 183484 114468 183512
rect 104860 183472 104866 183484
rect 114462 183472 114468 183484
rect 114520 183472 114526 183524
rect 214466 182316 214472 182368
rect 214524 182356 214530 182368
rect 226426 182356 226432 182368
rect 214524 182328 226432 182356
rect 214524 182316 214530 182328
rect 226426 182316 226432 182328
rect 226484 182316 226490 182368
rect 215018 182248 215024 182300
rect 215076 182288 215082 182300
rect 226334 182288 226340 182300
rect 215076 182260 226340 182288
rect 215076 182248 215082 182260
rect 226334 182248 226340 182260
rect 226392 182248 226398 182300
rect 113174 182180 113180 182232
rect 113232 182220 113238 182232
rect 115934 182220 115940 182232
rect 113232 182192 115940 182220
rect 113232 182180 113238 182192
rect 115934 182180 115940 182192
rect 115992 182180 115998 182232
rect 104802 182112 104808 182164
rect 104860 182152 104866 182164
rect 114370 182152 114376 182164
rect 104860 182124 114376 182152
rect 104860 182112 104866 182124
rect 114370 182112 114376 182124
rect 114428 182112 114434 182164
rect 335998 182112 336004 182164
rect 336056 182152 336062 182164
rect 579982 182152 579988 182164
rect 336056 182124 579988 182152
rect 336056 182112 336062 182124
rect 579982 182112 579988 182124
rect 580040 182112 580046 182164
rect 221458 181228 221464 181280
rect 221516 181268 221522 181280
rect 226334 181268 226340 181280
rect 221516 181240 226340 181268
rect 221516 181228 221522 181240
rect 226334 181228 226340 181240
rect 226392 181228 226398 181280
rect 113266 181092 113272 181144
rect 113324 181132 113330 181144
rect 115934 181132 115940 181144
rect 113324 181104 115940 181132
rect 113324 181092 113330 181104
rect 115934 181092 115940 181104
rect 115992 181092 115998 181144
rect 215110 180820 215116 180872
rect 215168 180860 215174 180872
rect 226334 180860 226340 180872
rect 215168 180832 226340 180860
rect 215168 180820 215174 180832
rect 226334 180820 226340 180832
rect 226392 180820 226398 180872
rect 227714 180820 227720 180872
rect 227772 180860 227778 180872
rect 230842 180860 230848 180872
rect 227772 180832 230848 180860
rect 227772 180820 227778 180832
rect 230842 180820 230848 180832
rect 230900 180820 230906 180872
rect 104802 180752 104808 180804
rect 104860 180792 104866 180804
rect 113174 180792 113180 180804
rect 104860 180764 113180 180792
rect 104860 180752 104866 180764
rect 113174 180752 113180 180764
rect 113232 180752 113238 180804
rect 213914 180548 213920 180600
rect 213972 180588 213978 180600
rect 218698 180588 218704 180600
rect 213972 180560 218704 180588
rect 213972 180548 213978 180560
rect 218698 180548 218704 180560
rect 218756 180548 218762 180600
rect 214469 179571 214527 179577
rect 214469 179537 214481 179571
rect 214515 179568 214527 179571
rect 214834 179568 214840 179580
rect 214515 179540 214840 179568
rect 214515 179537 214527 179540
rect 214469 179531 214527 179537
rect 214834 179528 214840 179540
rect 214892 179528 214898 179580
rect 222838 179460 222844 179512
rect 222896 179500 222902 179512
rect 226426 179500 226432 179512
rect 222896 179472 226432 179500
rect 222896 179460 222902 179472
rect 226426 179460 226432 179472
rect 226484 179460 226490 179512
rect 113910 179392 113916 179444
rect 113968 179432 113974 179444
rect 116394 179432 116400 179444
rect 113968 179404 116400 179432
rect 113968 179392 113974 179404
rect 116394 179392 116400 179404
rect 116452 179392 116458 179444
rect 214834 179392 214840 179444
rect 214892 179432 214898 179444
rect 226334 179432 226340 179444
rect 214892 179404 226340 179432
rect 214892 179392 214898 179404
rect 226334 179392 226340 179404
rect 226392 179392 226398 179444
rect 104802 179324 104808 179376
rect 104860 179364 104866 179376
rect 113266 179364 113272 179376
rect 104860 179336 113272 179364
rect 104860 179324 104866 179336
rect 113266 179324 113272 179336
rect 113324 179324 113330 179376
rect 214006 179324 214012 179376
rect 214064 179364 214070 179376
rect 222930 179364 222936 179376
rect 214064 179336 222936 179364
rect 214064 179324 214070 179336
rect 222930 179324 222936 179336
rect 222988 179324 222994 179376
rect 213914 179052 213920 179104
rect 213972 179092 213978 179104
rect 215938 179092 215944 179104
rect 213972 179064 215944 179092
rect 213972 179052 213978 179064
rect 215938 179052 215944 179064
rect 215996 179052 216002 179104
rect 221550 178100 221556 178152
rect 221608 178140 221614 178152
rect 226426 178140 226432 178152
rect 221608 178112 226432 178140
rect 221608 178100 221614 178112
rect 226426 178100 226432 178112
rect 226484 178100 226490 178152
rect 114186 178032 114192 178084
rect 114244 178072 114250 178084
rect 115934 178072 115940 178084
rect 114244 178044 115940 178072
rect 114244 178032 114250 178044
rect 115934 178032 115940 178044
rect 115992 178032 115998 178084
rect 224310 178032 224316 178084
rect 224368 178072 224374 178084
rect 226334 178072 226340 178084
rect 224368 178044 226340 178072
rect 224368 178032 224374 178044
rect 226334 178032 226340 178044
rect 226392 178032 226398 178084
rect 104158 177964 104164 178016
rect 104216 178004 104222 178016
rect 113910 178004 113916 178016
rect 104216 177976 113916 178004
rect 104216 177964 104222 177976
rect 113910 177964 113916 177976
rect 113968 177964 113974 178016
rect 213914 177964 213920 178016
rect 213972 178004 213978 178016
rect 227070 178004 227076 178016
rect 213972 177976 227076 178004
rect 213972 177964 213978 177976
rect 227070 177964 227076 177976
rect 227128 177964 227134 178016
rect 114094 176740 114100 176792
rect 114152 176780 114158 176792
rect 115934 176780 115940 176792
rect 114152 176752 115940 176780
rect 114152 176740 114158 176752
rect 115934 176740 115940 176752
rect 115992 176740 115998 176792
rect 114462 176672 114468 176724
rect 114520 176712 114526 176724
rect 116394 176712 116400 176724
rect 114520 176684 116400 176712
rect 114520 176672 114526 176684
rect 116394 176672 116400 176684
rect 116452 176672 116458 176724
rect 218698 176672 218704 176724
rect 218756 176712 218762 176724
rect 226334 176712 226340 176724
rect 218756 176684 226340 176712
rect 218756 176672 218762 176684
rect 226334 176672 226340 176684
rect 226392 176672 226398 176724
rect 104158 176604 104164 176656
rect 104216 176644 104222 176656
rect 114186 176644 114192 176656
rect 104216 176616 114192 176644
rect 104216 176604 104222 176616
rect 114186 176604 114192 176616
rect 114244 176604 114250 176656
rect 214006 176604 214012 176656
rect 214064 176644 214070 176656
rect 224402 176644 224408 176656
rect 214064 176616 224408 176644
rect 214064 176604 214070 176616
rect 224402 176604 224408 176616
rect 224460 176604 224466 176656
rect 114278 175244 114284 175296
rect 114336 175284 114342 175296
rect 116394 175284 116400 175296
rect 114336 175256 116400 175284
rect 114336 175244 114342 175256
rect 116394 175244 116400 175256
rect 116452 175244 116458 175296
rect 224218 175244 224224 175296
rect 224276 175284 224282 175296
rect 226886 175284 226892 175296
rect 224276 175256 226892 175284
rect 224276 175244 224282 175256
rect 226886 175244 226892 175256
rect 226944 175244 226950 175296
rect 104802 175176 104808 175228
rect 104860 175216 104866 175228
rect 114094 175216 114100 175228
rect 104860 175188 114100 175216
rect 104860 175176 104866 175188
rect 114094 175176 114100 175188
rect 114152 175176 114158 175228
rect 104526 175108 104532 175160
rect 104584 175148 104590 175160
rect 114462 175148 114468 175160
rect 104584 175120 114468 175148
rect 104584 175108 104590 175120
rect 114462 175108 114468 175120
rect 114520 175108 114526 175160
rect 213914 174156 213920 174208
rect 213972 174196 213978 174208
rect 220170 174196 220176 174208
rect 213972 174168 220176 174196
rect 213972 174156 213978 174168
rect 220170 174156 220176 174168
rect 220228 174156 220234 174208
rect 223574 174088 223580 174140
rect 223632 174128 223638 174140
rect 227714 174128 227720 174140
rect 223632 174100 227720 174128
rect 223632 174088 223638 174100
rect 227714 174088 227720 174100
rect 227772 174088 227778 174140
rect 220078 174020 220084 174072
rect 220136 174060 220142 174072
rect 226426 174060 226432 174072
rect 220136 174032 226432 174060
rect 220136 174020 220142 174032
rect 226426 174020 226432 174032
rect 226484 174020 226490 174072
rect 114370 173884 114376 173936
rect 114428 173924 114434 173936
rect 115934 173924 115940 173936
rect 114428 173896 115940 173924
rect 114428 173884 114434 173896
rect 115934 173884 115940 173896
rect 115992 173884 115998 173936
rect 214466 173924 214472 173936
rect 214427 173896 214472 173924
rect 214466 173884 214472 173896
rect 214524 173884 214530 173936
rect 104802 173816 104808 173868
rect 104860 173856 104866 173868
rect 114278 173856 114284 173868
rect 104860 173828 114284 173856
rect 104860 173816 104866 173828
rect 114278 173816 114284 173828
rect 114336 173816 114342 173868
rect 213914 173816 213920 173868
rect 213972 173856 213978 173868
rect 226978 173856 226984 173868
rect 213972 173828 226984 173856
rect 213972 173816 213978 173828
rect 226978 173816 226984 173828
rect 227036 173816 227042 173868
rect 113174 172524 113180 172576
rect 113232 172564 113238 172576
rect 116394 172564 116400 172576
rect 113232 172536 116400 172564
rect 113232 172524 113238 172536
rect 116394 172524 116400 172536
rect 116452 172524 116458 172576
rect 104434 172456 104440 172508
rect 104492 172496 104498 172508
rect 114370 172496 114376 172508
rect 104492 172468 114376 172496
rect 104492 172456 104498 172468
rect 114370 172456 114376 172468
rect 114428 172456 114434 172508
rect 213914 172456 213920 172508
rect 213972 172496 213978 172508
rect 225690 172496 225696 172508
rect 213972 172468 225696 172496
rect 213972 172456 213978 172468
rect 225690 172456 225696 172468
rect 225748 172456 225754 172508
rect 218790 171776 218796 171828
rect 218848 171816 218854 171828
rect 223574 171816 223580 171828
rect 218848 171788 223580 171816
rect 218848 171776 218854 171788
rect 223574 171776 223580 171788
rect 223632 171776 223638 171828
rect 113266 171572 113272 171624
rect 113324 171612 113330 171624
rect 116118 171612 116124 171624
rect 113324 171584 116124 171612
rect 113324 171572 113330 171584
rect 116118 171572 116124 171584
rect 116176 171572 116182 171624
rect 104802 171028 104808 171080
rect 104860 171068 104866 171080
rect 113174 171068 113180 171080
rect 104860 171040 113180 171068
rect 104860 171028 104866 171040
rect 113174 171028 113180 171040
rect 113232 171028 113238 171080
rect 218054 170348 218060 170400
rect 218112 170388 218118 170400
rect 227438 170388 227444 170400
rect 218112 170360 227444 170388
rect 218112 170348 218118 170360
rect 227438 170348 227444 170360
rect 227496 170348 227502 170400
rect 113910 169804 113916 169856
rect 113968 169844 113974 169856
rect 116302 169844 116308 169856
rect 113968 169816 116308 169844
rect 113968 169804 113974 169816
rect 116302 169804 116308 169816
rect 116360 169804 116366 169856
rect 104250 169736 104256 169788
rect 104308 169776 104314 169788
rect 116394 169776 116400 169788
rect 104308 169748 116400 169776
rect 104308 169736 104314 169748
rect 116394 169736 116400 169748
rect 116452 169736 116458 169788
rect 104802 169668 104808 169720
rect 104860 169708 104866 169720
rect 113266 169708 113272 169720
rect 104860 169680 113272 169708
rect 104860 169668 104866 169680
rect 113266 169668 113272 169680
rect 113324 169668 113330 169720
rect 213914 169056 213920 169108
rect 213972 169096 213978 169108
rect 221458 169096 221464 169108
rect 213972 169068 221464 169096
rect 213972 169056 213978 169068
rect 221458 169056 221464 169068
rect 221516 169056 221522 169108
rect 104802 168376 104808 168428
rect 104860 168416 104866 168428
rect 116394 168416 116400 168428
rect 104860 168388 116400 168416
rect 104860 168376 104866 168388
rect 116394 168376 116400 168388
rect 116452 168376 116458 168428
rect 104158 168308 104164 168360
rect 104216 168348 104222 168360
rect 113910 168348 113916 168360
rect 104216 168320 113916 168348
rect 104216 168308 104222 168320
rect 113910 168308 113916 168320
rect 113968 168308 113974 168360
rect 213914 168308 213920 168360
rect 213972 168348 213978 168360
rect 222838 168348 222844 168360
rect 213972 168320 222844 168348
rect 213972 168308 213978 168320
rect 222838 168308 222844 168320
rect 222896 168308 222902 168360
rect 114462 167016 114468 167068
rect 114520 167056 114526 167068
rect 115934 167056 115940 167068
rect 114520 167028 115940 167056
rect 114520 167016 114526 167028
rect 115934 167016 115940 167028
rect 115992 167016 115998 167068
rect 213914 166948 213920 167000
rect 213972 166988 213978 167000
rect 224310 166988 224316 167000
rect 213972 166960 224316 166988
rect 213972 166948 213978 166960
rect 224310 166948 224316 166960
rect 224368 166948 224374 167000
rect 232222 166948 232228 167000
rect 232280 166988 232286 167000
rect 232590 166988 232596 167000
rect 232280 166960 232596 166988
rect 232280 166948 232286 166960
rect 232590 166948 232596 166960
rect 232648 166948 232654 167000
rect 214190 166880 214196 166932
rect 214248 166920 214254 166932
rect 214466 166920 214472 166932
rect 214248 166892 214472 166920
rect 214248 166880 214254 166892
rect 214466 166880 214472 166892
rect 214524 166880 214530 166932
rect 214006 166540 214012 166592
rect 214064 166580 214070 166592
rect 221550 166580 221556 166592
rect 214064 166552 221556 166580
rect 214064 166540 214070 166552
rect 221550 166540 221556 166552
rect 221608 166540 221614 166592
rect 113818 165588 113824 165640
rect 113876 165628 113882 165640
rect 115934 165628 115940 165640
rect 113876 165600 115940 165628
rect 113876 165588 113882 165600
rect 115934 165588 115940 165600
rect 115992 165588 115998 165640
rect 104618 165520 104624 165572
rect 104676 165560 104682 165572
rect 114462 165560 114468 165572
rect 104676 165532 114468 165560
rect 104676 165520 104682 165532
rect 114462 165520 114468 165532
rect 114520 165520 114526 165572
rect 213914 165520 213920 165572
rect 213972 165560 213978 165572
rect 225598 165560 225604 165572
rect 213972 165532 225604 165560
rect 213972 165520 213978 165532
rect 225598 165520 225604 165532
rect 225656 165520 225662 165572
rect 114462 164228 114468 164280
rect 114520 164268 114526 164280
rect 116118 164268 116124 164280
rect 114520 164240 116124 164268
rect 114520 164228 114526 164240
rect 116118 164228 116124 164240
rect 116176 164228 116182 164280
rect 104802 164160 104808 164212
rect 104860 164200 104866 164212
rect 113818 164200 113824 164212
rect 104860 164172 113824 164200
rect 104860 164160 104866 164172
rect 113818 164160 113824 164172
rect 113876 164160 113882 164212
rect 232314 164160 232320 164212
rect 232372 164200 232378 164212
rect 232590 164200 232596 164212
rect 232372 164172 232596 164200
rect 232372 164160 232378 164172
rect 232590 164160 232596 164172
rect 232648 164160 232654 164212
rect 213914 164092 213920 164144
rect 213972 164132 213978 164144
rect 218698 164132 218704 164144
rect 213972 164104 218704 164132
rect 213972 164092 213978 164104
rect 218698 164092 218704 164104
rect 218756 164092 218762 164144
rect 213914 163548 213920 163600
rect 213972 163588 213978 163600
rect 220078 163588 220084 163600
rect 213972 163560 220084 163588
rect 213972 163548 213978 163560
rect 220078 163548 220084 163560
rect 220136 163548 220142 163600
rect 113174 162868 113180 162920
rect 113232 162908 113238 162920
rect 116394 162908 116400 162920
rect 113232 162880 116400 162908
rect 113232 162868 113238 162880
rect 116394 162868 116400 162880
rect 116452 162868 116458 162920
rect 104802 162800 104808 162852
rect 104860 162840 104866 162852
rect 114462 162840 114468 162852
rect 104860 162812 114468 162840
rect 104860 162800 104866 162812
rect 114462 162800 114468 162812
rect 114520 162800 114526 162852
rect 213914 162800 213920 162852
rect 213972 162840 213978 162852
rect 224218 162840 224224 162852
rect 213972 162812 224224 162840
rect 213972 162800 213978 162812
rect 224218 162800 224224 162812
rect 224276 162800 224282 162852
rect 213914 162256 213920 162308
rect 213972 162296 213978 162308
rect 218054 162296 218060 162308
rect 213972 162268 218060 162296
rect 213972 162256 213978 162268
rect 218054 162256 218060 162268
rect 218112 162256 218118 162308
rect 113266 161984 113272 162036
rect 113324 162024 113330 162036
rect 116210 162024 116216 162036
rect 113324 161996 116216 162024
rect 113324 161984 113330 161996
rect 116210 161984 116216 161996
rect 116268 161984 116274 162036
rect 103698 161440 103704 161492
rect 103756 161480 103762 161492
rect 116394 161480 116400 161492
rect 103756 161452 116400 161480
rect 103756 161440 103762 161452
rect 116394 161440 116400 161452
rect 116452 161440 116458 161492
rect 104802 161372 104808 161424
rect 104860 161412 104866 161424
rect 113174 161412 113180 161424
rect 104860 161384 113180 161412
rect 104860 161372 104866 161384
rect 113174 161372 113180 161384
rect 113232 161372 113238 161424
rect 213914 161372 213920 161424
rect 213972 161412 213978 161424
rect 229738 161412 229744 161424
rect 213972 161384 229744 161412
rect 213972 161372 213978 161384
rect 229738 161372 229744 161384
rect 229796 161372 229802 161424
rect 213914 160828 213920 160880
rect 213972 160868 213978 160880
rect 218790 160868 218796 160880
rect 213972 160840 218796 160868
rect 213972 160828 213978 160840
rect 218790 160828 218796 160840
rect 218848 160828 218854 160880
rect 104250 160080 104256 160132
rect 104308 160120 104314 160132
rect 116394 160120 116400 160132
rect 104308 160092 116400 160120
rect 104308 160080 104314 160092
rect 116394 160080 116400 160092
rect 116452 160080 116458 160132
rect 104802 160012 104808 160064
rect 104860 160052 104866 160064
rect 113266 160052 113272 160064
rect 104860 160024 113272 160052
rect 104860 160012 104866 160024
rect 113266 160012 113272 160024
rect 113324 160012 113330 160064
rect 104802 158720 104808 158772
rect 104860 158760 104866 158772
rect 116394 158760 116400 158772
rect 104860 158732 116400 158760
rect 104860 158720 104866 158732
rect 116394 158720 116400 158732
rect 116452 158720 116458 158772
rect 104342 157360 104348 157412
rect 104400 157400 104406 157412
rect 116394 157400 116400 157412
rect 104400 157372 116400 157400
rect 104400 157360 104406 157372
rect 116394 157360 116400 157372
rect 116452 157360 116458 157412
rect 114278 155932 114284 155984
rect 114336 155972 114342 155984
rect 116026 155972 116032 155984
rect 114336 155944 116032 155972
rect 114336 155932 114342 155944
rect 116026 155932 116032 155944
rect 116084 155932 116090 155984
rect 213914 155932 213920 155984
rect 213972 155972 213978 155984
rect 224678 155972 224684 155984
rect 213972 155944 224684 155972
rect 213972 155932 213978 155944
rect 224678 155932 224684 155944
rect 224736 155932 224742 155984
rect 113450 154640 113456 154692
rect 113508 154680 113514 154692
rect 116026 154680 116032 154692
rect 113508 154652 116032 154680
rect 113508 154640 113514 154652
rect 116026 154640 116032 154652
rect 116084 154640 116090 154692
rect 104250 154572 104256 154624
rect 104308 154612 104314 154624
rect 116394 154612 116400 154624
rect 104308 154584 116400 154612
rect 104308 154572 104314 154584
rect 116394 154572 116400 154584
rect 116452 154572 116458 154624
rect 213914 154572 213920 154624
rect 213972 154612 213978 154624
rect 224770 154612 224776 154624
rect 213972 154584 224776 154612
rect 213972 154572 213978 154584
rect 224770 154572 224776 154584
rect 224828 154572 224834 154624
rect 104618 154504 104624 154556
rect 104676 154544 104682 154556
rect 114278 154544 114284 154556
rect 104676 154516 114284 154544
rect 104676 154504 104682 154516
rect 114278 154504 114284 154516
rect 114336 154504 114342 154556
rect 213914 153280 213920 153332
rect 213972 153320 213978 153332
rect 224586 153320 224592 153332
rect 213972 153292 224592 153320
rect 213972 153280 213978 153292
rect 224586 153280 224592 153292
rect 224644 153280 224650 153332
rect 103790 153212 103796 153264
rect 103848 153252 103854 153264
rect 115934 153252 115940 153264
rect 103848 153224 115940 153252
rect 103848 153212 103854 153224
rect 115934 153212 115940 153224
rect 115992 153212 115998 153264
rect 214006 153212 214012 153264
rect 214064 153252 214070 153264
rect 224862 153252 224868 153264
rect 214064 153224 224868 153252
rect 214064 153212 214070 153224
rect 224862 153212 224868 153224
rect 224920 153212 224926 153264
rect 104802 153144 104808 153196
rect 104860 153184 104866 153196
rect 113450 153184 113456 153196
rect 104860 153156 113456 153184
rect 104860 153144 104866 153156
rect 113450 153144 113456 153156
rect 113508 153144 113514 153196
rect 213914 151852 213920 151904
rect 213972 151892 213978 151904
rect 224494 151892 224500 151904
rect 213972 151864 224500 151892
rect 213972 151852 213978 151864
rect 224494 151852 224500 151864
rect 224552 151852 224558 151904
rect 103698 151784 103704 151836
rect 103756 151824 103762 151836
rect 116394 151824 116400 151836
rect 103756 151796 116400 151824
rect 103756 151784 103762 151796
rect 116394 151784 116400 151796
rect 116452 151784 116458 151836
rect 215938 151784 215944 151836
rect 215996 151824 216002 151836
rect 286134 151824 286140 151836
rect 215996 151796 286140 151824
rect 215996 151784 216002 151796
rect 286134 151784 286140 151796
rect 286192 151784 286198 151836
rect 213914 150832 213920 150884
rect 213972 150872 213978 150884
rect 216674 150872 216680 150884
rect 213972 150844 216680 150872
rect 213972 150832 213978 150844
rect 216674 150832 216680 150844
rect 216732 150832 216738 150884
rect 104342 150424 104348 150476
rect 104400 150464 104406 150476
rect 116394 150464 116400 150476
rect 104400 150436 116400 150464
rect 104400 150424 104406 150436
rect 116394 150424 116400 150436
rect 116452 150424 116458 150476
rect 213914 150424 213920 150476
rect 213972 150464 213978 150476
rect 224218 150464 224224 150476
rect 213972 150436 224224 150464
rect 213972 150424 213978 150436
rect 224218 150424 224224 150436
rect 224276 150424 224282 150476
rect 224678 150356 224684 150408
rect 224736 150396 224742 150408
rect 227438 150396 227444 150408
rect 224736 150368 227444 150396
rect 224736 150356 224742 150368
rect 227438 150356 227444 150368
rect 227496 150356 227502 150408
rect 232130 149676 232136 149728
rect 232188 149716 232194 149728
rect 232498 149716 232504 149728
rect 232188 149688 232504 149716
rect 232188 149676 232194 149688
rect 232498 149676 232504 149688
rect 232556 149676 232562 149728
rect 213914 149336 213920 149388
rect 213972 149376 213978 149388
rect 216766 149376 216772 149388
rect 213972 149348 216772 149376
rect 213972 149336 213978 149348
rect 216766 149336 216772 149348
rect 216824 149336 216830 149388
rect 104802 149064 104808 149116
rect 104860 149104 104866 149116
rect 116394 149104 116400 149116
rect 104860 149076 116400 149104
rect 104860 149064 104866 149076
rect 116394 149064 116400 149076
rect 116452 149064 116458 149116
rect 213914 149064 213920 149116
rect 213972 149104 213978 149116
rect 224126 149104 224132 149116
rect 213972 149076 224132 149104
rect 213972 149064 213978 149076
rect 224126 149064 224132 149076
rect 224184 149064 224190 149116
rect 214098 148996 214104 149048
rect 214156 149036 214162 149048
rect 227438 149036 227444 149048
rect 214156 149008 227444 149036
rect 214156 148996 214162 149008
rect 227438 148996 227444 149008
rect 227496 148996 227502 149048
rect 224770 148928 224776 148980
rect 224828 148968 224834 148980
rect 227530 148968 227536 148980
rect 224828 148940 227536 148968
rect 224828 148928 224834 148940
rect 227530 148928 227536 148940
rect 227588 148928 227594 148980
rect 214558 148316 214564 148368
rect 214616 148356 214622 148368
rect 214742 148356 214748 148368
rect 214616 148328 214748 148356
rect 214616 148316 214622 148328
rect 214742 148316 214748 148328
rect 214800 148316 214806 148368
rect 213914 147976 213920 148028
rect 213972 148016 213978 148028
rect 216858 148016 216864 148028
rect 213972 147988 216864 148016
rect 213972 147976 213978 147988
rect 216858 147976 216864 147988
rect 216916 147976 216922 148028
rect 104710 147636 104716 147688
rect 104768 147676 104774 147688
rect 116394 147676 116400 147688
rect 104768 147648 116400 147676
rect 104768 147636 104774 147648
rect 116394 147636 116400 147648
rect 116452 147636 116458 147688
rect 214926 147568 214932 147620
rect 214984 147608 214990 147620
rect 227438 147608 227444 147620
rect 214984 147580 227444 147608
rect 214984 147568 214990 147580
rect 227438 147568 227444 147580
rect 227496 147568 227502 147620
rect 224862 147500 224868 147552
rect 224920 147540 224926 147552
rect 226978 147540 226984 147552
rect 224920 147512 226984 147540
rect 224920 147500 224926 147512
rect 226978 147500 226984 147512
rect 227036 147500 227042 147552
rect 224586 147432 224592 147484
rect 224644 147472 224650 147484
rect 227530 147472 227536 147484
rect 224644 147444 227536 147472
rect 224644 147432 224650 147444
rect 227530 147432 227536 147444
rect 227588 147432 227594 147484
rect 113634 146344 113640 146396
rect 113692 146384 113698 146396
rect 115934 146384 115940 146396
rect 113692 146356 115940 146384
rect 113692 146344 113698 146356
rect 115934 146344 115940 146356
rect 115992 146344 115998 146396
rect 213914 146344 213920 146396
rect 213972 146384 213978 146396
rect 217594 146384 217600 146396
rect 213972 146356 217600 146384
rect 213972 146344 213978 146356
rect 217594 146344 217600 146356
rect 217652 146344 217658 146396
rect 104526 146276 104532 146328
rect 104584 146316 104590 146328
rect 116394 146316 116400 146328
rect 104584 146288 116400 146316
rect 104584 146276 104590 146288
rect 116394 146276 116400 146288
rect 116452 146276 116458 146328
rect 214006 146276 214012 146328
rect 214064 146316 214070 146328
rect 227622 146316 227628 146328
rect 214064 146288 227628 146316
rect 214064 146276 214070 146288
rect 227622 146276 227628 146288
rect 227680 146276 227686 146328
rect 216674 146208 216680 146260
rect 216732 146248 216738 146260
rect 226702 146248 226708 146260
rect 216732 146220 226708 146248
rect 216732 146208 216738 146220
rect 226702 146208 226708 146220
rect 226760 146208 226766 146260
rect 224494 146140 224500 146192
rect 224552 146180 224558 146192
rect 227438 146180 227444 146192
rect 224552 146152 227444 146180
rect 224552 146140 224558 146152
rect 227438 146140 227444 146152
rect 227496 146140 227502 146192
rect 213914 144984 213920 145036
rect 213972 145024 213978 145036
rect 217318 145024 217324 145036
rect 213972 144996 217324 145024
rect 213972 144984 213978 144996
rect 217318 144984 217324 144996
rect 217376 144984 217382 145036
rect 104158 144916 104164 144968
rect 104216 144956 104222 144968
rect 116026 144956 116032 144968
rect 104216 144928 116032 144956
rect 104216 144916 104222 144928
rect 116026 144916 116032 144928
rect 116084 144916 116090 144968
rect 214006 144916 214012 144968
rect 214064 144956 214070 144968
rect 227254 144956 227260 144968
rect 214064 144928 227260 144956
rect 214064 144916 214070 144928
rect 227254 144916 227260 144928
rect 227312 144916 227318 144968
rect 104618 144848 104624 144900
rect 104676 144888 104682 144900
rect 113634 144888 113640 144900
rect 104676 144860 113640 144888
rect 104676 144848 104682 144860
rect 113634 144848 113640 144860
rect 113692 144848 113698 144900
rect 216766 144848 216772 144900
rect 216824 144888 216830 144900
rect 226518 144888 226524 144900
rect 216824 144860 226524 144888
rect 216824 144848 216830 144860
rect 226518 144848 226524 144860
rect 226576 144848 226582 144900
rect 224218 144780 224224 144832
rect 224276 144820 224282 144832
rect 227438 144820 227444 144832
rect 224276 144792 227444 144820
rect 224276 144780 224282 144792
rect 227438 144780 227444 144792
rect 227496 144780 227502 144832
rect 213914 143624 213920 143676
rect 213972 143664 213978 143676
rect 216766 143664 216772 143676
rect 213972 143636 216772 143664
rect 213972 143624 213978 143636
rect 216766 143624 216772 143636
rect 216824 143624 216830 143676
rect 103514 143556 103520 143608
rect 103572 143596 103578 143608
rect 116394 143596 116400 143608
rect 103572 143568 116400 143596
rect 103572 143556 103578 143568
rect 116394 143556 116400 143568
rect 116452 143556 116458 143608
rect 214006 143556 214012 143608
rect 214064 143596 214070 143608
rect 227530 143596 227536 143608
rect 214064 143568 227536 143596
rect 214064 143556 214070 143568
rect 227530 143556 227536 143568
rect 227588 143556 227594 143608
rect 216858 143488 216864 143540
rect 216916 143528 216922 143540
rect 226886 143528 226892 143540
rect 216916 143500 226892 143528
rect 216916 143488 216922 143500
rect 226886 143488 226892 143500
rect 226944 143488 226950 143540
rect 214374 143420 214380 143472
rect 214432 143460 214438 143472
rect 214558 143460 214564 143472
rect 214432 143432 214564 143460
rect 214432 143420 214438 143432
rect 214558 143420 214564 143432
rect 214616 143420 214622 143472
rect 224126 143420 224132 143472
rect 224184 143460 224190 143472
rect 227438 143460 227444 143472
rect 224184 143432 227444 143460
rect 224184 143420 224190 143432
rect 227438 143420 227444 143432
rect 227496 143420 227502 143472
rect 213914 142196 213920 142248
rect 213972 142236 213978 142248
rect 216674 142236 216680 142248
rect 213972 142208 216680 142236
rect 213972 142196 213978 142208
rect 216674 142196 216680 142208
rect 216732 142196 216738 142248
rect 103698 142128 103704 142180
rect 103756 142168 103762 142180
rect 116394 142168 116400 142180
rect 103756 142140 116400 142168
rect 103756 142128 103762 142140
rect 116394 142128 116400 142140
rect 116452 142128 116458 142180
rect 214006 142128 214012 142180
rect 214064 142168 214070 142180
rect 227346 142168 227352 142180
rect 214064 142140 227352 142168
rect 214064 142128 214070 142140
rect 227346 142128 227352 142140
rect 227404 142128 227410 142180
rect 217594 142060 217600 142112
rect 217652 142100 217658 142112
rect 226702 142100 226708 142112
rect 217652 142072 226708 142100
rect 217652 142060 217658 142072
rect 226702 142060 226708 142072
rect 226760 142060 226766 142112
rect 104342 140768 104348 140820
rect 104400 140808 104406 140820
rect 116394 140808 116400 140820
rect 104400 140780 116400 140808
rect 104400 140768 104406 140780
rect 116394 140768 116400 140780
rect 116452 140768 116458 140820
rect 213914 140768 213920 140820
rect 213972 140808 213978 140820
rect 226702 140808 226708 140820
rect 213972 140780 226708 140808
rect 213972 140768 213978 140780
rect 226702 140768 226708 140780
rect 226760 140768 226766 140820
rect 217318 140700 217324 140752
rect 217376 140740 217382 140752
rect 227070 140740 227076 140752
rect 217376 140712 227076 140740
rect 217376 140700 217382 140712
rect 227070 140700 227076 140712
rect 227128 140700 227134 140752
rect 113542 139476 113548 139528
rect 113600 139516 113606 139528
rect 116302 139516 116308 139528
rect 113600 139488 116308 139516
rect 113600 139476 113606 139488
rect 116302 139476 116308 139488
rect 116360 139476 116366 139528
rect 213914 139476 213920 139528
rect 213972 139516 213978 139528
rect 226610 139516 226616 139528
rect 213972 139488 226616 139516
rect 213972 139476 213978 139488
rect 226610 139476 226616 139488
rect 226668 139476 226674 139528
rect 104802 139408 104808 139460
rect 104860 139448 104866 139460
rect 116394 139448 116400 139460
rect 104860 139420 116400 139448
rect 104860 139408 104866 139420
rect 116394 139408 116400 139420
rect 116452 139408 116458 139460
rect 214006 139408 214012 139460
rect 214064 139448 214070 139460
rect 226518 139448 226524 139460
rect 214064 139420 226524 139448
rect 214064 139408 214070 139420
rect 226518 139408 226524 139420
rect 226576 139408 226582 139460
rect 216766 139340 216772 139392
rect 216824 139380 216830 139392
rect 227438 139380 227444 139392
rect 216824 139352 227444 139380
rect 216824 139340 216830 139352
rect 227438 139340 227444 139352
rect 227496 139340 227502 139392
rect 214006 138048 214012 138100
rect 214064 138088 214070 138100
rect 226426 138088 226432 138100
rect 214064 138060 226432 138088
rect 214064 138048 214070 138060
rect 226426 138048 226432 138060
rect 226484 138048 226490 138100
rect 213914 137980 213920 138032
rect 213972 138020 213978 138032
rect 226794 138020 226800 138032
rect 213972 137992 226800 138020
rect 213972 137980 213978 137992
rect 226794 137980 226800 137992
rect 226852 137980 226858 138032
rect 216674 137912 216680 137964
rect 216732 137952 216738 137964
rect 227438 137952 227444 137964
rect 216732 137924 227444 137952
rect 216732 137912 216738 137924
rect 227438 137912 227444 137924
rect 227496 137912 227502 137964
rect 213914 136688 213920 136740
rect 213972 136728 213978 136740
rect 227070 136728 227076 136740
rect 213972 136700 227076 136728
rect 213972 136688 213978 136700
rect 227070 136688 227076 136700
rect 227128 136688 227134 136740
rect 104710 136620 104716 136672
rect 104768 136660 104774 136672
rect 116394 136660 116400 136672
rect 104768 136632 116400 136660
rect 104768 136620 104774 136632
rect 116394 136620 116400 136632
rect 116452 136620 116458 136672
rect 214006 136620 214012 136672
rect 214064 136660 214070 136672
rect 227438 136660 227444 136672
rect 214064 136632 227444 136660
rect 214064 136620 214070 136632
rect 227438 136620 227444 136632
rect 227496 136620 227502 136672
rect 104342 135260 104348 135312
rect 104400 135300 104406 135312
rect 115934 135300 115940 135312
rect 104400 135272 115940 135300
rect 104400 135260 104406 135272
rect 115934 135260 115940 135272
rect 115992 135260 115998 135312
rect 213914 135260 213920 135312
rect 213972 135300 213978 135312
rect 227622 135300 227628 135312
rect 213972 135272 227628 135300
rect 213972 135260 213978 135272
rect 227622 135260 227628 135272
rect 227680 135260 227686 135312
rect 104802 135192 104808 135244
rect 104860 135232 104866 135244
rect 113542 135232 113548 135244
rect 104860 135204 113548 135232
rect 104860 135192 104866 135204
rect 113542 135192 113548 135204
rect 113600 135192 113606 135244
rect 341518 135192 341524 135244
rect 341576 135232 341582 135244
rect 580166 135232 580172 135244
rect 341576 135204 580172 135232
rect 341576 135192 341582 135204
rect 580166 135192 580172 135204
rect 580224 135192 580230 135244
rect 214006 133968 214012 134020
rect 214064 134008 214070 134020
rect 227530 134008 227536 134020
rect 214064 133980 227536 134008
rect 214064 133968 214070 133980
rect 227530 133968 227536 133980
rect 227588 133968 227594 134020
rect 100478 133900 100484 133952
rect 100536 133940 100542 133952
rect 103606 133940 103612 133952
rect 100536 133912 103612 133940
rect 100536 133900 100542 133912
rect 103606 133900 103612 133912
rect 103664 133900 103670 133952
rect 109862 133900 109868 133952
rect 109920 133940 109926 133952
rect 116394 133940 116400 133952
rect 109920 133912 116400 133940
rect 109920 133900 109926 133912
rect 116394 133900 116400 133912
rect 116452 133900 116458 133952
rect 213914 133900 213920 133952
rect 213972 133940 213978 133952
rect 227346 133940 227352 133952
rect 213972 133912 227352 133940
rect 213972 133900 213978 133912
rect 227346 133900 227352 133912
rect 227404 133900 227410 133952
rect 104802 133832 104808 133884
rect 104860 133872 104866 133884
rect 115842 133872 115848 133884
rect 104860 133844 115848 133872
rect 104860 133832 104866 133844
rect 115842 133832 115848 133844
rect 115900 133832 115906 133884
rect 114554 132880 114560 132932
rect 114612 132920 114618 132932
rect 117130 132920 117136 132932
rect 114612 132892 117136 132920
rect 114612 132880 114618 132892
rect 117130 132880 117136 132892
rect 117188 132880 117194 132932
rect 213914 132540 213920 132592
rect 213972 132580 213978 132592
rect 226702 132580 226708 132592
rect 213972 132552 226708 132580
rect 213972 132540 213978 132552
rect 226702 132540 226708 132552
rect 226760 132540 226766 132592
rect 214006 132472 214012 132524
rect 214064 132512 214070 132524
rect 227438 132512 227444 132524
rect 214064 132484 227444 132512
rect 214064 132472 214070 132484
rect 227438 132472 227444 132484
rect 227496 132472 227502 132524
rect 113910 131180 113916 131232
rect 113968 131220 113974 131232
rect 116394 131220 116400 131232
rect 113968 131192 116400 131220
rect 113968 131180 113974 131192
rect 116394 131180 116400 131192
rect 116452 131180 116458 131232
rect 213914 131180 213920 131232
rect 213972 131220 213978 131232
rect 226518 131220 226524 131232
rect 213972 131192 226524 131220
rect 213972 131180 213978 131192
rect 226518 131180 226524 131192
rect 226576 131180 226582 131232
rect 100386 131112 100392 131164
rect 100444 131152 100450 131164
rect 115934 131152 115940 131164
rect 100444 131124 115940 131152
rect 100444 131112 100450 131124
rect 115934 131112 115940 131124
rect 115992 131112 115998 131164
rect 214006 131112 214012 131164
rect 214064 131152 214070 131164
rect 227070 131152 227076 131164
rect 214064 131124 227076 131152
rect 214064 131112 214070 131124
rect 227070 131112 227076 131124
rect 227128 131112 227134 131164
rect 103974 130704 103980 130756
rect 104032 130744 104038 130756
rect 109862 130744 109868 130756
rect 104032 130716 109868 130744
rect 104032 130704 104038 130716
rect 109862 130704 109868 130716
rect 109920 130704 109926 130756
rect 213914 129752 213920 129804
rect 213972 129792 213978 129804
rect 227530 129792 227536 129804
rect 213972 129764 227536 129792
rect 213972 129752 213978 129764
rect 227530 129752 227536 129764
rect 227588 129752 227594 129804
rect 104802 129684 104808 129736
rect 104860 129724 104866 129736
rect 114554 129724 114560 129736
rect 104860 129696 114560 129724
rect 104860 129684 104866 129696
rect 114554 129684 114560 129696
rect 114612 129684 114618 129736
rect 116394 129316 116400 129328
rect 10428 129288 116400 129316
rect 10428 129260 10456 129288
rect 116394 129276 116400 129288
rect 116452 129276 116458 129328
rect 10410 129208 10416 129260
rect 10468 129208 10474 129260
rect 213914 129004 213920 129056
rect 213972 129044 213978 129056
rect 227438 129044 227444 129056
rect 213972 129016 227444 129044
rect 213972 129004 213978 129016
rect 227438 129004 227444 129016
rect 227496 129004 227502 129056
rect 213914 128324 213920 128376
rect 213972 128364 213978 128376
rect 226334 128364 226340 128376
rect 213972 128336 226340 128364
rect 213972 128324 213978 128336
rect 226334 128324 226340 128336
rect 226392 128324 226398 128376
rect 9030 128256 9036 128308
rect 9088 128296 9094 128308
rect 116394 128296 116400 128308
rect 9088 128268 116400 128296
rect 9088 128256 9094 128268
rect 116394 128256 116400 128268
rect 116452 128256 116458 128308
rect 104802 128188 104808 128240
rect 104860 128228 104866 128240
rect 113910 128228 113916 128240
rect 104860 128200 113916 128228
rect 104860 128188 104866 128200
rect 113910 128188 113916 128200
rect 113968 128188 113974 128240
rect 103606 127576 103612 127628
rect 103664 127616 103670 127628
rect 116302 127616 116308 127628
rect 103664 127588 116308 127616
rect 103664 127576 103670 127588
rect 116302 127576 116308 127588
rect 116360 127576 116366 127628
rect 213914 127576 213920 127628
rect 213972 127616 213978 127628
rect 227438 127616 227444 127628
rect 213972 127588 227444 127616
rect 213972 127576 213978 127588
rect 227438 127576 227444 127588
rect 227496 127576 227502 127628
rect 213914 126964 213920 127016
rect 213972 127004 213978 127016
rect 227438 127004 227444 127016
rect 213972 126976 227444 127004
rect 213972 126964 213978 126976
rect 227438 126964 227444 126976
rect 227496 126964 227502 127016
rect 10318 126896 10324 126948
rect 10376 126936 10382 126948
rect 116394 126936 116400 126948
rect 10376 126908 116400 126936
rect 10376 126896 10382 126908
rect 116394 126896 116400 126908
rect 116452 126896 116458 126948
rect 213914 126216 213920 126268
rect 213972 126256 213978 126268
rect 227438 126256 227444 126268
rect 213972 126228 227444 126256
rect 213972 126216 213978 126228
rect 227438 126216 227444 126228
rect 227496 126216 227502 126268
rect 213914 125604 213920 125656
rect 213972 125644 213978 125656
rect 227438 125644 227444 125656
rect 213972 125616 227444 125644
rect 213972 125604 213978 125616
rect 227438 125604 227444 125616
rect 227496 125604 227502 125656
rect 8938 125536 8944 125588
rect 8996 125576 9002 125588
rect 116394 125576 116400 125588
rect 8996 125548 116400 125576
rect 8996 125536 9002 125548
rect 116394 125536 116400 125548
rect 116452 125536 116458 125588
rect 214374 125536 214380 125588
rect 214432 125576 214438 125588
rect 214466 125576 214472 125588
rect 214432 125548 214472 125576
rect 214432 125536 214438 125548
rect 214466 125536 214472 125548
rect 214524 125536 214530 125588
rect 78214 125468 78220 125520
rect 78272 125508 78278 125520
rect 100386 125508 100392 125520
rect 78272 125480 100392 125508
rect 78272 125468 78278 125480
rect 100386 125468 100392 125480
rect 100444 125468 100450 125520
rect 213914 124856 213920 124908
rect 213972 124896 213978 124908
rect 227254 124896 227260 124908
rect 213972 124868 227260 124896
rect 213972 124856 213978 124868
rect 227254 124856 227260 124868
rect 227312 124856 227318 124908
rect 213914 124108 213920 124160
rect 213972 124148 213978 124160
rect 227254 124148 227260 124160
rect 213972 124120 227260 124148
rect 213972 124108 213978 124120
rect 227254 124108 227260 124120
rect 227312 124108 227318 124160
rect 213914 123428 213920 123480
rect 213972 123468 213978 123480
rect 227254 123468 227260 123480
rect 213972 123440 227260 123468
rect 213972 123428 213978 123440
rect 227254 123428 227260 123440
rect 227312 123428 227318 123480
rect 213914 122748 213920 122800
rect 213972 122788 213978 122800
rect 227438 122788 227444 122800
rect 213972 122760 227444 122788
rect 213972 122748 213978 122760
rect 227438 122748 227444 122760
rect 227496 122748 227502 122800
rect 213914 122068 213920 122120
rect 213972 122108 213978 122120
rect 227438 122108 227444 122120
rect 213972 122080 227444 122108
rect 213972 122068 213978 122080
rect 227438 122068 227444 122080
rect 227496 122068 227502 122120
rect 50982 121456 50988 121508
rect 51040 121496 51046 121508
rect 116394 121496 116400 121508
rect 51040 121468 116400 121496
rect 51040 121456 51046 121468
rect 116394 121456 116400 121468
rect 116452 121456 116458 121508
rect 213914 121388 213920 121440
rect 213972 121428 213978 121440
rect 227438 121428 227444 121440
rect 213972 121400 227444 121428
rect 213972 121388 213978 121400
rect 227438 121388 227444 121400
rect 227496 121388 227502 121440
rect 213914 120708 213920 120760
rect 213972 120748 213978 120760
rect 227438 120748 227444 120760
rect 213972 120720 227444 120748
rect 213972 120708 213978 120720
rect 227438 120708 227444 120720
rect 227496 120708 227502 120760
rect 94498 120096 94504 120148
rect 94556 120136 94562 120148
rect 116394 120136 116400 120148
rect 94556 120108 116400 120136
rect 94556 120096 94562 120108
rect 116394 120096 116400 120108
rect 116452 120096 116458 120148
rect 213914 120028 213920 120080
rect 213972 120068 213978 120080
rect 227438 120068 227444 120080
rect 213972 120040 227444 120068
rect 213972 120028 213978 120040
rect 227438 120028 227444 120040
rect 227496 120028 227502 120080
rect 94682 118668 94688 118720
rect 94740 118708 94746 118720
rect 116394 118708 116400 118720
rect 94740 118680 116400 118708
rect 94740 118668 94746 118680
rect 116394 118668 116400 118680
rect 116452 118668 116458 118720
rect 213914 118600 213920 118652
rect 213972 118640 213978 118652
rect 226426 118640 226432 118652
rect 213972 118612 226432 118640
rect 213972 118600 213978 118612
rect 226426 118600 226432 118612
rect 226484 118600 226490 118652
rect 214006 118532 214012 118584
rect 214064 118572 214070 118584
rect 226334 118572 226340 118584
rect 214064 118544 226340 118572
rect 214064 118532 214070 118544
rect 226334 118532 226340 118544
rect 226392 118532 226398 118584
rect 94590 117308 94596 117360
rect 94648 117348 94654 117360
rect 116394 117348 116400 117360
rect 94648 117320 116400 117348
rect 94648 117308 94654 117320
rect 116394 117308 116400 117320
rect 116452 117308 116458 117360
rect 214006 117240 214012 117292
rect 214064 117280 214070 117292
rect 227438 117280 227444 117292
rect 214064 117252 227444 117280
rect 214064 117240 214070 117252
rect 227438 117240 227444 117252
rect 227496 117240 227502 117292
rect 213914 117172 213920 117224
rect 213972 117212 213978 117224
rect 226242 117212 226248 117224
rect 213972 117184 226248 117212
rect 213972 117172 213978 117184
rect 226242 117172 226248 117184
rect 226300 117172 226306 117224
rect 94958 116016 94964 116068
rect 95016 116056 95022 116068
rect 116118 116056 116124 116068
rect 95016 116028 116124 116056
rect 95016 116016 95022 116028
rect 116118 116016 116124 116028
rect 116176 116016 116182 116068
rect 94774 115948 94780 116000
rect 94832 115988 94838 116000
rect 116394 115988 116400 116000
rect 94832 115960 116400 115988
rect 94832 115948 94838 115960
rect 116394 115948 116400 115960
rect 116452 115948 116458 116000
rect 214006 115880 214012 115932
rect 214064 115920 214070 115932
rect 227438 115920 227444 115932
rect 214064 115892 227444 115920
rect 214064 115880 214070 115892
rect 227438 115880 227444 115892
rect 227496 115880 227502 115932
rect 213914 115812 213920 115864
rect 213972 115852 213978 115864
rect 226150 115852 226156 115864
rect 213972 115824 226156 115852
rect 213972 115812 213978 115824
rect 226150 115812 226156 115824
rect 226208 115812 226214 115864
rect 94866 114520 94872 114572
rect 94924 114560 94930 114572
rect 116394 114560 116400 114572
rect 94924 114532 116400 114560
rect 94924 114520 94930 114532
rect 116394 114520 116400 114532
rect 116452 114520 116458 114572
rect 214006 114452 214012 114504
rect 214064 114492 214070 114504
rect 227070 114492 227076 114504
rect 214064 114464 227076 114492
rect 214064 114452 214070 114464
rect 227070 114452 227076 114464
rect 227128 114452 227134 114504
rect 213914 114384 213920 114436
rect 213972 114424 213978 114436
rect 226242 114424 226248 114436
rect 213972 114396 226248 114424
rect 213972 114384 213978 114396
rect 226242 114384 226248 114396
rect 226300 114384 226306 114436
rect 97258 113160 97264 113212
rect 97316 113200 97322 113212
rect 116394 113200 116400 113212
rect 97316 113172 116400 113200
rect 97316 113160 97322 113172
rect 116394 113160 116400 113172
rect 116452 113160 116458 113212
rect 213914 113092 213920 113144
rect 213972 113132 213978 113144
rect 226150 113132 226156 113144
rect 213972 113104 226156 113132
rect 213972 113092 213978 113104
rect 226150 113092 226156 113104
rect 226208 113092 226214 113144
rect 94406 111800 94412 111852
rect 94464 111840 94470 111852
rect 116394 111840 116400 111852
rect 94464 111812 116400 111840
rect 94464 111800 94470 111812
rect 116394 111800 116400 111812
rect 116452 111800 116458 111852
rect 214006 111732 214012 111784
rect 214064 111772 214070 111784
rect 226242 111772 226248 111784
rect 214064 111744 226248 111772
rect 214064 111732 214070 111744
rect 226242 111732 226248 111744
rect 226300 111732 226306 111784
rect 213914 111664 213920 111716
rect 213972 111704 213978 111716
rect 226058 111704 226064 111716
rect 213972 111676 226064 111704
rect 213972 111664 213978 111676
rect 226058 111664 226064 111676
rect 226116 111664 226122 111716
rect 95878 110440 95884 110492
rect 95936 110480 95942 110492
rect 116394 110480 116400 110492
rect 95936 110452 116400 110480
rect 95936 110440 95942 110452
rect 116394 110440 116400 110452
rect 116452 110440 116458 110492
rect 214006 110372 214012 110424
rect 214064 110412 214070 110424
rect 226150 110412 226156 110424
rect 214064 110384 226156 110412
rect 214064 110372 214070 110384
rect 226150 110372 226156 110384
rect 226208 110372 226214 110424
rect 213914 110304 213920 110356
rect 213972 110344 213978 110356
rect 225966 110344 225972 110356
rect 213972 110316 225972 110344
rect 213972 110304 213978 110316
rect 225966 110304 225972 110316
rect 226024 110304 226030 110356
rect 95142 109012 95148 109064
rect 95200 109052 95206 109064
rect 116394 109052 116400 109064
rect 95200 109024 116400 109052
rect 95200 109012 95206 109024
rect 116394 109012 116400 109024
rect 116452 109012 116458 109064
rect 214006 108944 214012 108996
rect 214064 108984 214070 108996
rect 226242 108984 226248 108996
rect 214064 108956 226248 108984
rect 214064 108944 214070 108956
rect 226242 108944 226248 108956
rect 226300 108944 226306 108996
rect 213914 108876 213920 108928
rect 213972 108916 213978 108928
rect 225874 108916 225880 108928
rect 213972 108888 225880 108916
rect 213972 108876 213978 108888
rect 225874 108876 225880 108888
rect 225932 108876 225938 108928
rect 102778 107720 102784 107772
rect 102836 107760 102842 107772
rect 116302 107760 116308 107772
rect 102836 107732 116308 107760
rect 102836 107720 102842 107732
rect 116302 107720 116308 107732
rect 116360 107720 116366 107772
rect 95050 107652 95056 107704
rect 95108 107692 95114 107704
rect 116394 107692 116400 107704
rect 95108 107664 116400 107692
rect 95108 107652 95114 107664
rect 116394 107652 116400 107664
rect 116452 107652 116458 107704
rect 213914 107584 213920 107636
rect 213972 107624 213978 107636
rect 226058 107624 226064 107636
rect 213972 107596 226064 107624
rect 213972 107584 213978 107596
rect 226058 107584 226064 107596
rect 226116 107584 226122 107636
rect 98638 106292 98644 106344
rect 98696 106332 98702 106344
rect 116394 106332 116400 106344
rect 98696 106304 116400 106332
rect 98696 106292 98702 106304
rect 116394 106292 116400 106304
rect 116452 106292 116458 106344
rect 213914 106224 213920 106276
rect 213972 106264 213978 106276
rect 225782 106264 225788 106276
rect 213972 106236 225788 106264
rect 213972 106224 213978 106236
rect 225782 106224 225788 106236
rect 225840 106224 225846 106276
rect 214006 106156 214012 106208
rect 214064 106196 214070 106208
rect 226242 106196 226248 106208
rect 214064 106168 226248 106196
rect 214064 106156 214070 106168
rect 226242 106156 226248 106168
rect 226300 106156 226306 106208
rect 94314 104864 94320 104916
rect 94372 104904 94378 104916
rect 116394 104904 116400 104916
rect 94372 104876 116400 104904
rect 94372 104864 94378 104876
rect 116394 104864 116400 104876
rect 116452 104864 116458 104916
rect 224770 104864 224776 104916
rect 224828 104904 224834 104916
rect 227438 104904 227444 104916
rect 224828 104876 227444 104904
rect 224828 104864 224834 104876
rect 227438 104864 227444 104876
rect 227496 104864 227502 104916
rect 214006 104796 214012 104848
rect 214064 104836 214070 104848
rect 226150 104836 226156 104848
rect 214064 104808 226156 104836
rect 214064 104796 214070 104808
rect 226150 104796 226156 104808
rect 226208 104796 226214 104848
rect 213914 104728 213920 104780
rect 213972 104768 213978 104780
rect 225598 104768 225604 104780
rect 213972 104740 225604 104768
rect 213972 104728 213978 104740
rect 225598 104728 225604 104740
rect 225656 104728 225662 104780
rect 224862 103640 224868 103692
rect 224920 103680 224926 103692
rect 227438 103680 227444 103692
rect 224920 103652 227444 103680
rect 224920 103640 224926 103652
rect 227438 103640 227444 103652
rect 227496 103640 227502 103692
rect 101398 103504 101404 103556
rect 101456 103544 101462 103556
rect 116394 103544 116400 103556
rect 101456 103516 116400 103544
rect 101456 103504 101462 103516
rect 116394 103504 116400 103516
rect 116452 103504 116458 103556
rect 214006 103436 214012 103488
rect 214064 103476 214070 103488
rect 225966 103476 225972 103488
rect 214064 103448 225972 103476
rect 214064 103436 214070 103448
rect 225966 103436 225972 103448
rect 226024 103436 226030 103488
rect 213914 103368 213920 103420
rect 213972 103408 213978 103420
rect 225690 103408 225696 103420
rect 213972 103380 225696 103408
rect 213972 103368 213978 103380
rect 225690 103368 225696 103380
rect 225748 103368 225754 103420
rect 94222 102144 94228 102196
rect 94280 102184 94286 102196
rect 116302 102184 116308 102196
rect 94280 102156 116308 102184
rect 94280 102144 94286 102156
rect 116302 102144 116308 102156
rect 116360 102144 116366 102196
rect 213914 102076 213920 102128
rect 213972 102116 213978 102128
rect 225874 102116 225880 102128
rect 213972 102088 225880 102116
rect 213972 102076 213978 102088
rect 225874 102076 225880 102088
rect 225932 102076 225938 102128
rect 314194 102076 314200 102128
rect 314252 102116 314258 102128
rect 338390 102116 338396 102128
rect 314252 102088 338396 102116
rect 314252 102076 314258 102088
rect 338390 102076 338396 102088
rect 338448 102076 338454 102128
rect 105538 100784 105544 100836
rect 105596 100824 105602 100836
rect 116394 100824 116400 100836
rect 105596 100796 116400 100824
rect 105596 100784 105602 100796
rect 116394 100784 116400 100796
rect 116452 100784 116458 100836
rect 104158 100716 104164 100768
rect 104216 100756 104222 100768
rect 116302 100756 116308 100768
rect 104216 100728 116308 100756
rect 104216 100716 104222 100728
rect 116302 100716 116308 100728
rect 116360 100716 116366 100768
rect 213914 100648 213920 100700
rect 213972 100688 213978 100700
rect 226150 100688 226156 100700
rect 213972 100660 226156 100688
rect 213972 100648 213978 100660
rect 226150 100648 226156 100660
rect 226208 100648 226214 100700
rect 232130 100648 232136 100700
rect 232188 100688 232194 100700
rect 258074 100688 258080 100700
rect 232188 100660 258080 100688
rect 232188 100648 232194 100660
rect 258074 100648 258080 100660
rect 258132 100648 258138 100700
rect 214006 100580 214012 100632
rect 214064 100620 214070 100632
rect 226058 100620 226064 100632
rect 214064 100592 226064 100620
rect 214064 100580 214070 100592
rect 226058 100580 226064 100592
rect 226116 100580 226122 100632
rect 97350 99356 97356 99408
rect 97408 99396 97414 99408
rect 116394 99396 116400 99408
rect 97408 99368 116400 99396
rect 97408 99356 97414 99368
rect 116394 99356 116400 99368
rect 116452 99356 116458 99408
rect 214650 99288 214656 99340
rect 214708 99328 214714 99340
rect 226242 99328 226248 99340
rect 214708 99300 226248 99328
rect 214708 99288 214714 99300
rect 226242 99288 226248 99300
rect 226300 99288 226306 99340
rect 232130 99288 232136 99340
rect 232188 99328 232194 99340
rect 232498 99328 232504 99340
rect 232188 99300 232504 99328
rect 232188 99288 232194 99300
rect 232498 99288 232504 99300
rect 232556 99288 232562 99340
rect 215110 99220 215116 99272
rect 215168 99260 215174 99272
rect 224770 99260 224776 99272
rect 215168 99232 224776 99260
rect 215168 99220 215174 99232
rect 224770 99220 224776 99232
rect 224828 99220 224834 99272
rect 94130 97996 94136 98048
rect 94188 98036 94194 98048
rect 116394 98036 116400 98048
rect 94188 98008 116400 98036
rect 94188 97996 94194 98008
rect 116394 97996 116400 98008
rect 116452 97996 116458 98048
rect 214098 97928 214104 97980
rect 214156 97968 214162 97980
rect 224862 97968 224868 97980
rect 214156 97940 224868 97968
rect 214156 97928 214162 97940
rect 224862 97928 224868 97940
rect 224920 97928 224926 97980
rect 213914 97588 213920 97640
rect 213972 97628 213978 97640
rect 215938 97628 215944 97640
rect 213972 97600 215944 97628
rect 213972 97588 213978 97600
rect 215938 97588 215944 97600
rect 215996 97588 216002 97640
rect 100018 96636 100024 96688
rect 100076 96676 100082 96688
rect 116394 96676 116400 96688
rect 100076 96648 116400 96676
rect 100076 96636 100082 96648
rect 116394 96636 116400 96648
rect 116452 96636 116458 96688
rect 94682 95208 94688 95260
rect 94740 95248 94746 95260
rect 116302 95248 116308 95260
rect 94740 95220 116308 95248
rect 94740 95208 94746 95220
rect 116302 95208 116308 95220
rect 116360 95208 116366 95260
rect 215110 95140 215116 95192
rect 215168 95180 215174 95192
rect 576118 95180 576124 95192
rect 215168 95152 576124 95180
rect 215168 95140 215174 95152
rect 576118 95140 576124 95152
rect 576176 95140 576182 95192
rect 94498 93848 94504 93900
rect 94556 93888 94562 93900
rect 116394 93888 116400 93900
rect 94556 93860 116400 93888
rect 94556 93848 94562 93860
rect 116394 93848 116400 93860
rect 116452 93848 116458 93900
rect 215202 93780 215208 93832
rect 215260 93820 215266 93832
rect 578878 93820 578884 93832
rect 215260 93792 578884 93820
rect 215260 93780 215266 93792
rect 578878 93780 578884 93792
rect 578936 93780 578942 93832
rect 215110 93712 215116 93764
rect 215168 93752 215174 93764
rect 577498 93752 577504 93764
rect 215168 93724 577504 93752
rect 215168 93712 215174 93724
rect 577498 93712 577504 93724
rect 577556 93712 577562 93764
rect 95142 93508 95148 93560
rect 95200 93548 95206 93560
rect 97258 93548 97264 93560
rect 95200 93520 97264 93548
rect 95200 93508 95206 93520
rect 97258 93508 97264 93520
rect 97316 93508 97322 93560
rect 95970 92488 95976 92540
rect 96028 92528 96034 92540
rect 116394 92528 116400 92540
rect 96028 92500 116400 92528
rect 96028 92488 96034 92500
rect 116394 92488 116400 92500
rect 116452 92488 116458 92540
rect 94590 91808 94596 91860
rect 94648 91848 94654 91860
rect 95878 91848 95884 91860
rect 94648 91820 95884 91848
rect 94648 91808 94654 91820
rect 95878 91808 95884 91820
rect 95936 91808 95942 91860
rect 94590 91060 94596 91112
rect 94648 91100 94654 91112
rect 116394 91100 116400 91112
rect 94648 91072 116400 91100
rect 94648 91060 94654 91072
rect 116394 91060 116400 91072
rect 116452 91060 116458 91112
rect 94774 90992 94780 91044
rect 94832 91032 94838 91044
rect 102778 91032 102784 91044
rect 94832 91004 102784 91032
rect 94832 90992 94838 91004
rect 102778 90992 102784 91004
rect 102836 90992 102842 91044
rect 98730 90312 98736 90364
rect 98788 90352 98794 90364
rect 116486 90352 116492 90364
rect 98788 90324 116492 90352
rect 98788 90312 98794 90324
rect 116486 90312 116492 90324
rect 116544 90312 116550 90364
rect 102870 89700 102876 89752
rect 102928 89740 102934 89752
rect 116394 89740 116400 89752
rect 102928 89712 116400 89740
rect 102928 89700 102934 89712
rect 116394 89700 116400 89712
rect 116452 89700 116458 89752
rect 94958 88340 94964 88392
rect 95016 88380 95022 88392
rect 115934 88380 115940 88392
rect 95016 88352 115940 88380
rect 95016 88340 95022 88352
rect 115934 88340 115940 88352
rect 115992 88340 115998 88392
rect 340138 88272 340144 88324
rect 340196 88312 340202 88324
rect 580166 88312 580172 88324
rect 340196 88284 580172 88312
rect 340196 88272 340202 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 95142 88204 95148 88256
rect 95200 88244 95206 88256
rect 98638 88244 98644 88256
rect 95200 88216 98644 88244
rect 95200 88204 95206 88216
rect 98638 88204 98644 88216
rect 98696 88204 98702 88256
rect 97258 86980 97264 87032
rect 97316 87020 97322 87032
rect 116394 87020 116400 87032
rect 97316 86992 116400 87020
rect 97316 86980 97322 86992
rect 116394 86980 116400 86992
rect 116452 86980 116458 87032
rect 94406 86572 94412 86624
rect 94464 86612 94470 86624
rect 101398 86612 101404 86624
rect 94464 86584 101404 86612
rect 94464 86572 94470 86584
rect 101398 86572 101404 86584
rect 101456 86572 101462 86624
rect 101490 85620 101496 85672
rect 101548 85660 101554 85672
rect 116394 85660 116400 85672
rect 101548 85632 116400 85660
rect 101548 85620 101554 85632
rect 116394 85620 116400 85632
rect 116452 85620 116458 85672
rect 94774 85552 94780 85604
rect 94832 85592 94838 85604
rect 116302 85592 116308 85604
rect 94832 85564 116308 85592
rect 94832 85552 94838 85564
rect 116302 85552 116308 85564
rect 116360 85552 116366 85604
rect 215110 85552 215116 85604
rect 215168 85592 215174 85604
rect 224218 85592 224224 85604
rect 215168 85564 224224 85592
rect 215168 85552 215174 85564
rect 224218 85552 224224 85564
rect 224276 85552 224282 85604
rect 95142 85484 95148 85536
rect 95200 85524 95206 85536
rect 104158 85524 104164 85536
rect 95200 85496 104164 85524
rect 95200 85484 95206 85496
rect 104158 85484 104164 85496
rect 104216 85484 104222 85536
rect 94866 84192 94872 84244
rect 94924 84232 94930 84244
rect 116394 84232 116400 84244
rect 94924 84204 116400 84232
rect 94924 84192 94930 84204
rect 116394 84192 116400 84204
rect 116452 84192 116458 84244
rect 215110 84192 215116 84244
rect 215168 84232 215174 84244
rect 225598 84232 225604 84244
rect 215168 84204 225604 84232
rect 215168 84192 215174 84204
rect 225598 84192 225604 84204
rect 225656 84192 225662 84244
rect 95142 84124 95148 84176
rect 95200 84164 95206 84176
rect 105538 84164 105544 84176
rect 95200 84136 105544 84164
rect 95200 84124 95206 84136
rect 105538 84124 105544 84136
rect 105596 84124 105602 84176
rect 214006 83512 214012 83564
rect 214064 83552 214070 83564
rect 214374 83552 214380 83564
rect 214064 83524 214380 83552
rect 214064 83512 214070 83524
rect 214374 83512 214380 83524
rect 214432 83512 214438 83564
rect 284478 83512 284484 83564
rect 284536 83552 284542 83564
rect 413278 83552 413284 83564
rect 284536 83524 413284 83552
rect 284536 83512 284542 83524
rect 413278 83512 413284 83524
rect 413336 83512 413342 83564
rect 320818 83444 320824 83496
rect 320876 83484 320882 83496
rect 580258 83484 580264 83496
rect 320876 83456 580264 83484
rect 320876 83444 320882 83456
rect 580258 83444 580264 83456
rect 580316 83444 580322 83496
rect 94222 83376 94228 83428
rect 94280 83416 94286 83428
rect 97350 83416 97356 83428
rect 94280 83388 97356 83416
rect 94280 83376 94286 83388
rect 97350 83376 97356 83388
rect 97408 83376 97414 83428
rect 95878 82832 95884 82884
rect 95936 82872 95942 82884
rect 116394 82872 116400 82884
rect 95936 82844 116400 82872
rect 95936 82832 95942 82844
rect 116394 82832 116400 82844
rect 116452 82832 116458 82884
rect 215938 82832 215944 82884
rect 215996 82872 216002 82884
rect 248138 82872 248144 82884
rect 215996 82844 248144 82872
rect 215996 82832 216002 82844
rect 248138 82832 248144 82844
rect 248196 82832 248202 82884
rect 95050 81404 95056 81456
rect 95108 81444 95114 81456
rect 115934 81444 115940 81456
rect 95108 81416 115940 81444
rect 95108 81404 95114 81416
rect 115934 81404 115940 81416
rect 115992 81404 115998 81456
rect 214190 81404 214196 81456
rect 214248 81444 214254 81456
rect 226978 81444 226984 81456
rect 214248 81416 226984 81444
rect 214248 81404 214254 81416
rect 226978 81404 226984 81416
rect 227036 81404 227042 81456
rect 215018 81336 215024 81388
rect 215076 81376 215082 81388
rect 227346 81376 227352 81388
rect 215076 81348 227352 81376
rect 215076 81336 215082 81348
rect 227346 81336 227352 81348
rect 227404 81336 227410 81388
rect 94406 81268 94412 81320
rect 94464 81308 94470 81320
rect 100018 81308 100024 81320
rect 94464 81280 100024 81308
rect 94464 81268 94470 81280
rect 100018 81268 100024 81280
rect 100076 81268 100082 81320
rect 214834 81268 214840 81320
rect 214892 81308 214898 81320
rect 227438 81308 227444 81320
rect 214892 81280 227444 81308
rect 214892 81268 214898 81280
rect 227438 81268 227444 81280
rect 227496 81268 227502 81320
rect 215110 80112 215116 80164
rect 215168 80152 215174 80164
rect 220170 80152 220176 80164
rect 215168 80124 220176 80152
rect 215168 80112 215174 80124
rect 220170 80112 220176 80124
rect 220228 80112 220234 80164
rect 232406 80152 232412 80164
rect 232332 80124 232412 80152
rect 98638 80044 98644 80096
rect 98696 80084 98702 80096
rect 116394 80084 116400 80096
rect 98696 80056 116400 80084
rect 98696 80044 98702 80056
rect 116394 80044 116400 80056
rect 116452 80044 116458 80096
rect 232332 80028 232360 80124
rect 232406 80112 232412 80124
rect 232464 80112 232470 80164
rect 94406 79976 94412 80028
rect 94464 80016 94470 80028
rect 98730 80016 98736 80028
rect 94464 79988 98736 80016
rect 94464 79976 94470 79988
rect 98730 79976 98736 79988
rect 98788 79976 98794 80028
rect 214282 79976 214288 80028
rect 214340 80016 214346 80028
rect 227530 80016 227536 80028
rect 214340 79988 227536 80016
rect 214340 79976 214346 79988
rect 227530 79976 227536 79988
rect 227588 79976 227594 80028
rect 232314 79976 232320 80028
rect 232372 79976 232378 80028
rect 214558 79908 214564 79960
rect 214616 79948 214622 79960
rect 227438 79948 227444 79960
rect 214616 79920 227444 79948
rect 214616 79908 214622 79920
rect 227438 79908 227444 79920
rect 227496 79908 227502 79960
rect 100018 78752 100024 78804
rect 100076 78792 100082 78804
rect 116394 78792 116400 78804
rect 100076 78764 116400 78792
rect 100076 78752 100082 78764
rect 116394 78752 116400 78764
rect 116452 78752 116458 78804
rect 213914 78752 213920 78804
rect 213972 78792 213978 78804
rect 220814 78792 220820 78804
rect 213972 78764 220820 78792
rect 213972 78752 213978 78764
rect 220814 78752 220820 78764
rect 220872 78752 220878 78804
rect 95142 78684 95148 78736
rect 95200 78724 95206 78736
rect 116210 78724 116216 78736
rect 95200 78696 116216 78724
rect 95200 78684 95206 78696
rect 116210 78684 116216 78696
rect 116268 78684 116274 78736
rect 214006 78616 214012 78668
rect 214064 78656 214070 78668
rect 227530 78656 227536 78668
rect 214064 78628 227536 78656
rect 214064 78616 214070 78628
rect 227530 78616 227536 78628
rect 227588 78616 227594 78668
rect 214742 78548 214748 78600
rect 214800 78588 214806 78600
rect 227438 78588 227444 78600
rect 214800 78560 227444 78588
rect 214800 78548 214806 78560
rect 227438 78548 227444 78560
rect 227496 78548 227502 78600
rect 94222 78208 94228 78260
rect 94280 78248 94286 78260
rect 95970 78248 95976 78260
rect 94280 78220 95976 78248
rect 94280 78208 94286 78220
rect 95970 78208 95976 78220
rect 96028 78208 96034 78260
rect 94682 77256 94688 77308
rect 94740 77296 94746 77308
rect 116394 77296 116400 77308
rect 94740 77268 116400 77296
rect 94740 77256 94746 77268
rect 116394 77256 116400 77268
rect 116452 77256 116458 77308
rect 213914 77256 213920 77308
rect 213972 77296 213978 77308
rect 218790 77296 218796 77308
rect 213972 77268 218796 77296
rect 213972 77256 213978 77268
rect 218790 77256 218796 77268
rect 218848 77256 218854 77308
rect 214650 77188 214656 77240
rect 214708 77228 214714 77240
rect 227438 77228 227444 77240
rect 214708 77200 227444 77228
rect 214708 77188 214714 77200
rect 227438 77188 227444 77200
rect 227496 77188 227502 77240
rect 214466 77120 214472 77172
rect 214524 77160 214530 77172
rect 227530 77160 227536 77172
rect 214524 77132 227536 77160
rect 214524 77120 214530 77132
rect 227530 77120 227536 77132
rect 227588 77120 227594 77172
rect 213914 76032 213920 76084
rect 213972 76072 213978 76084
rect 219434 76072 219440 76084
rect 213972 76044 219440 76072
rect 213972 76032 213978 76044
rect 219434 76032 219440 76044
rect 219492 76032 219498 76084
rect 97350 75896 97356 75948
rect 97408 75936 97414 75948
rect 116394 75936 116400 75948
rect 97408 75908 116400 75936
rect 97408 75896 97414 75908
rect 116394 75896 116400 75908
rect 116452 75896 116458 75948
rect 224218 75828 224224 75880
rect 224276 75868 224282 75880
rect 227438 75868 227444 75880
rect 224276 75840 227444 75868
rect 224276 75828 224282 75840
rect 227438 75828 227444 75840
rect 227496 75828 227502 75880
rect 94590 75692 94596 75744
rect 94648 75732 94654 75744
rect 102870 75732 102876 75744
rect 94648 75704 102876 75732
rect 94648 75692 94654 75704
rect 102870 75692 102876 75704
rect 102928 75692 102934 75744
rect 214190 75692 214196 75744
rect 214248 75732 214254 75744
rect 227438 75732 227444 75744
rect 214248 75704 227444 75732
rect 214248 75692 214254 75704
rect 227438 75692 227444 75704
rect 227496 75692 227502 75744
rect 213914 74604 213920 74656
rect 213972 74644 213978 74656
rect 216030 74644 216036 74656
rect 213972 74616 216036 74644
rect 213972 74604 213978 74616
rect 216030 74604 216036 74616
rect 216088 74604 216094 74656
rect 94498 74536 94504 74588
rect 94556 74576 94562 74588
rect 116394 74576 116400 74588
rect 94556 74548 116400 74576
rect 94556 74536 94562 74548
rect 116394 74536 116400 74548
rect 116452 74536 116458 74588
rect 215220 74548 215432 74576
rect 214374 74400 214380 74452
rect 214432 74440 214438 74452
rect 215220 74440 215248 74548
rect 215404 74508 215432 74548
rect 227438 74508 227444 74520
rect 215404 74480 227444 74508
rect 227438 74468 227444 74480
rect 227496 74468 227502 74520
rect 214432 74412 215248 74440
rect 214432 74400 214438 74412
rect 94590 74264 94596 74316
rect 94648 74304 94654 74316
rect 97258 74304 97264 74316
rect 94648 74276 97264 74304
rect 94648 74264 94654 74276
rect 97258 74264 97264 74276
rect 97316 74264 97322 74316
rect 95970 73176 95976 73228
rect 96028 73216 96034 73228
rect 116394 73216 116400 73228
rect 96028 73188 116400 73216
rect 96028 73176 96034 73188
rect 116394 73176 116400 73188
rect 116452 73176 116458 73228
rect 213914 73176 213920 73228
rect 213972 73216 213978 73228
rect 218054 73216 218060 73228
rect 213972 73188 218060 73216
rect 213972 73176 213978 73188
rect 218054 73176 218060 73188
rect 218112 73176 218118 73228
rect 215202 73108 215208 73160
rect 215260 73148 215266 73160
rect 227438 73148 227444 73160
rect 215260 73120 227444 73148
rect 215260 73108 215266 73120
rect 227438 73108 227444 73120
rect 227496 73108 227502 73160
rect 220170 73040 220176 73092
rect 220228 73080 220234 73092
rect 227530 73080 227536 73092
rect 220228 73052 227536 73080
rect 220228 73040 220234 73052
rect 227530 73040 227536 73052
rect 227588 73040 227594 73092
rect 94406 72904 94412 72956
rect 94464 72944 94470 72956
rect 101490 72944 101496 72956
rect 94464 72916 101496 72944
rect 94464 72904 94470 72916
rect 101490 72904 101496 72916
rect 101548 72904 101554 72956
rect 94958 71748 94964 71800
rect 95016 71788 95022 71800
rect 116394 71788 116400 71800
rect 95016 71760 116400 71788
rect 95016 71748 95022 71760
rect 116394 71748 116400 71760
rect 116452 71748 116458 71800
rect 214926 71680 214932 71732
rect 214984 71720 214990 71732
rect 227438 71720 227444 71732
rect 214984 71692 227444 71720
rect 214984 71680 214990 71692
rect 227438 71680 227444 71692
rect 227496 71680 227502 71732
rect 220814 71612 220820 71664
rect 220872 71652 220878 71664
rect 227530 71652 227536 71664
rect 220872 71624 227536 71652
rect 220872 71612 220878 71624
rect 227530 71612 227536 71624
rect 227588 71612 227594 71664
rect 214006 70456 214012 70508
rect 214064 70496 214070 70508
rect 224494 70496 224500 70508
rect 214064 70468 224500 70496
rect 214064 70456 214070 70468
rect 224494 70456 224500 70468
rect 224552 70456 224558 70508
rect 94590 70388 94596 70440
rect 94648 70428 94654 70440
rect 116394 70428 116400 70440
rect 94648 70400 116400 70428
rect 94648 70388 94654 70400
rect 116394 70388 116400 70400
rect 116452 70388 116458 70440
rect 213914 70388 213920 70440
rect 213972 70428 213978 70440
rect 224402 70428 224408 70440
rect 213972 70400 224408 70428
rect 213972 70388 213978 70400
rect 224402 70388 224408 70400
rect 224460 70388 224466 70440
rect 214834 70320 214840 70372
rect 214892 70360 214898 70372
rect 227438 70360 227444 70372
rect 214892 70332 227444 70360
rect 214892 70320 214898 70332
rect 227438 70320 227444 70332
rect 227496 70320 227502 70372
rect 94866 70252 94872 70304
rect 94924 70292 94930 70304
rect 95878 70292 95884 70304
rect 94924 70264 95884 70292
rect 94924 70252 94930 70264
rect 95878 70252 95884 70264
rect 95936 70252 95942 70304
rect 218790 70252 218796 70304
rect 218848 70292 218854 70304
rect 226518 70292 226524 70304
rect 218848 70264 226524 70292
rect 218848 70252 218854 70264
rect 226518 70252 226524 70264
rect 226576 70252 226582 70304
rect 215110 69096 215116 69148
rect 215168 69136 215174 69148
rect 224218 69136 224224 69148
rect 215168 69108 224224 69136
rect 215168 69096 215174 69108
rect 224218 69096 224224 69108
rect 224276 69096 224282 69148
rect 94406 69028 94412 69080
rect 94464 69068 94470 69080
rect 116394 69068 116400 69080
rect 94464 69040 116400 69068
rect 94464 69028 94470 69040
rect 116394 69028 116400 69040
rect 116452 69028 116458 69080
rect 214650 69028 214656 69080
rect 214708 69068 214714 69080
rect 224126 69068 224132 69080
rect 214708 69040 224132 69068
rect 214708 69028 214714 69040
rect 224126 69028 224132 69040
rect 224184 69028 224190 69080
rect 215018 68960 215024 69012
rect 215076 69000 215082 69012
rect 227438 69000 227444 69012
rect 215076 68972 227444 69000
rect 215076 68960 215082 68972
rect 227438 68960 227444 68972
rect 227496 68960 227502 69012
rect 219434 68892 219440 68944
rect 219492 68932 219498 68944
rect 227530 68932 227536 68944
rect 219492 68904 227536 68932
rect 219492 68892 219498 68904
rect 227530 68892 227536 68904
rect 227588 68892 227594 68944
rect 93854 68484 93860 68536
rect 93912 68524 93918 68536
rect 98638 68524 98644 68536
rect 93912 68496 98644 68524
rect 93912 68484 93918 68496
rect 98638 68484 98644 68496
rect 98696 68484 98702 68536
rect 214466 67668 214472 67720
rect 214524 67708 214530 67720
rect 224678 67708 224684 67720
rect 214524 67680 224684 67708
rect 214524 67668 214530 67680
rect 224678 67668 224684 67680
rect 224736 67668 224742 67720
rect 94866 67600 94872 67652
rect 94924 67640 94930 67652
rect 116394 67640 116400 67652
rect 94924 67612 116400 67640
rect 94924 67600 94930 67612
rect 116394 67600 116400 67612
rect 116452 67600 116458 67652
rect 215110 67600 215116 67652
rect 215168 67640 215174 67652
rect 224862 67640 224868 67652
rect 215168 67612 224868 67640
rect 215168 67600 215174 67612
rect 224862 67600 224868 67612
rect 224920 67600 224926 67652
rect 214742 67532 214748 67584
rect 214800 67572 214806 67584
rect 227438 67572 227444 67584
rect 214800 67544 227444 67572
rect 214800 67532 214806 67544
rect 227438 67532 227444 67544
rect 227496 67532 227502 67584
rect 216030 67464 216036 67516
rect 216088 67504 216094 67516
rect 227530 67504 227536 67516
rect 216088 67476 227536 67504
rect 216088 67464 216094 67476
rect 227530 67464 227536 67476
rect 227588 67464 227594 67516
rect 95142 66852 95148 66904
rect 95200 66892 95206 66904
rect 100018 66892 100024 66904
rect 95200 66864 100024 66892
rect 95200 66852 95206 66864
rect 100018 66852 100024 66864
rect 100076 66852 100082 66904
rect 94774 66240 94780 66292
rect 94832 66280 94838 66292
rect 116394 66280 116400 66292
rect 94832 66252 116400 66280
rect 94832 66240 94838 66252
rect 116394 66240 116400 66252
rect 116452 66240 116458 66292
rect 215110 66240 215116 66292
rect 215168 66280 215174 66292
rect 224310 66280 224316 66292
rect 215168 66252 224316 66280
rect 215168 66240 215174 66252
rect 224310 66240 224316 66252
rect 224368 66240 224374 66292
rect 214098 66172 214104 66224
rect 214156 66212 214162 66224
rect 227438 66212 227444 66224
rect 214156 66184 227444 66212
rect 214156 66172 214162 66184
rect 227438 66172 227444 66184
rect 227496 66172 227502 66224
rect 218054 66104 218060 66156
rect 218112 66144 218118 66156
rect 227530 66144 227536 66156
rect 218112 66116 227536 66144
rect 218112 66104 218118 66116
rect 227530 66104 227536 66116
rect 227588 66104 227594 66156
rect 214374 65492 214380 65544
rect 214432 65532 214438 65544
rect 216766 65532 216772 65544
rect 214432 65504 216772 65532
rect 214432 65492 214438 65504
rect 216766 65492 216772 65504
rect 216824 65492 216830 65544
rect 94682 65288 94688 65340
rect 94740 65328 94746 65340
rect 97350 65328 97356 65340
rect 94740 65300 97356 65328
rect 94740 65288 94746 65300
rect 97350 65288 97356 65300
rect 97408 65288 97414 65340
rect 94314 64880 94320 64932
rect 94372 64920 94378 64932
rect 116394 64920 116400 64932
rect 94372 64892 116400 64920
rect 94372 64880 94378 64892
rect 116394 64880 116400 64892
rect 116452 64880 116458 64932
rect 214006 64880 214012 64932
rect 214064 64920 214070 64932
rect 224586 64920 224592 64932
rect 214064 64892 224592 64920
rect 214064 64880 214070 64892
rect 224586 64880 224592 64892
rect 224644 64880 224650 64932
rect 214558 64812 214564 64864
rect 214616 64852 214622 64864
rect 227438 64852 227444 64864
rect 214616 64824 227444 64852
rect 214616 64812 214622 64824
rect 227438 64812 227444 64824
rect 227496 64812 227502 64864
rect 224494 64472 224500 64524
rect 224552 64512 224558 64524
rect 227438 64512 227444 64524
rect 224552 64484 227444 64512
rect 224552 64472 224558 64484
rect 227438 64472 227444 64484
rect 227496 64472 227502 64524
rect 224402 64268 224408 64320
rect 224460 64308 224466 64320
rect 227530 64308 227536 64320
rect 224460 64280 227536 64308
rect 224460 64268 224466 64280
rect 227530 64268 227536 64280
rect 227588 64268 227594 64320
rect 94222 63656 94228 63708
rect 94280 63696 94286 63708
rect 94774 63696 94780 63708
rect 94280 63668 94780 63696
rect 94280 63656 94286 63668
rect 94774 63656 94780 63668
rect 94832 63656 94838 63708
rect 214558 63588 214564 63640
rect 214616 63628 214622 63640
rect 216950 63628 216956 63640
rect 214616 63600 216956 63628
rect 214616 63588 214622 63600
rect 216950 63588 216956 63600
rect 217008 63588 217014 63640
rect 95142 63520 95148 63572
rect 95200 63560 95206 63572
rect 115934 63560 115940 63572
rect 95200 63532 115940 63560
rect 95200 63520 95206 63532
rect 115934 63520 115940 63532
rect 115992 63520 115998 63572
rect 215110 63520 215116 63572
rect 215168 63560 215174 63572
rect 224034 63560 224040 63572
rect 215168 63532 224040 63560
rect 215168 63520 215174 63532
rect 224034 63520 224040 63532
rect 224092 63520 224098 63572
rect 94866 63452 94872 63504
rect 94924 63492 94930 63504
rect 95970 63492 95976 63504
rect 94924 63464 95976 63492
rect 94924 63452 94930 63464
rect 95970 63452 95976 63464
rect 96028 63452 96034 63504
rect 224126 63452 224132 63504
rect 224184 63492 224190 63504
rect 227438 63492 227444 63504
rect 224184 63464 227444 63492
rect 224184 63452 224190 63464
rect 227438 63452 227444 63464
rect 227496 63452 227502 63504
rect 224218 63384 224224 63436
rect 224276 63424 224282 63436
rect 227530 63424 227536 63436
rect 224276 63396 227536 63424
rect 224276 63384 224282 63396
rect 227530 63384 227536 63396
rect 227588 63384 227594 63436
rect 487614 62772 487620 62824
rect 487672 62812 487678 62824
rect 576210 62812 576216 62824
rect 487672 62784 576216 62812
rect 487672 62772 487678 62784
rect 576210 62772 576216 62784
rect 576268 62772 576274 62824
rect 94682 62160 94688 62212
rect 94740 62200 94746 62212
rect 116210 62200 116216 62212
rect 94740 62172 116216 62200
rect 94740 62160 94746 62172
rect 116210 62160 116216 62172
rect 116268 62160 116274 62212
rect 214650 62160 214656 62212
rect 214708 62200 214714 62212
rect 216674 62200 216680 62212
rect 214708 62172 216680 62200
rect 214708 62160 214714 62172
rect 216674 62160 216680 62172
rect 216732 62160 216738 62212
rect 94498 62092 94504 62144
rect 94556 62132 94562 62144
rect 116394 62132 116400 62144
rect 94556 62104 116400 62132
rect 94556 62092 94562 62104
rect 116394 62092 116400 62104
rect 116452 62092 116458 62144
rect 215110 62092 215116 62144
rect 215168 62132 215174 62144
rect 224126 62132 224132 62144
rect 215168 62104 224132 62132
rect 215168 62092 215174 62104
rect 224126 62092 224132 62104
rect 224184 62092 224190 62144
rect 93946 62024 93952 62076
rect 94004 62064 94010 62076
rect 116578 62064 116584 62076
rect 94004 62036 116584 62064
rect 94004 62024 94010 62036
rect 116578 62024 116584 62036
rect 116636 62024 116642 62076
rect 224678 62024 224684 62076
rect 224736 62064 224742 62076
rect 227530 62064 227536 62076
rect 224736 62036 227536 62064
rect 224736 62024 224742 62036
rect 227530 62024 227536 62036
rect 227588 62024 227594 62076
rect 224862 61956 224868 62008
rect 224920 61996 224926 62008
rect 226702 61996 226708 62008
rect 224920 61968 226708 61996
rect 224920 61956 224926 61968
rect 226702 61956 226708 61968
rect 226760 61956 226766 62008
rect 214558 61208 214564 61260
rect 214616 61248 214622 61260
rect 216858 61248 216864 61260
rect 214616 61220 216864 61248
rect 214616 61208 214622 61220
rect 216858 61208 216864 61220
rect 216916 61208 216922 61260
rect 94958 60732 94964 60784
rect 95016 60772 95022 60784
rect 116394 60772 116400 60784
rect 95016 60744 116400 60772
rect 95016 60732 95022 60744
rect 116394 60732 116400 60744
rect 116452 60732 116458 60784
rect 215110 60732 215116 60784
rect 215168 60772 215174 60784
rect 224218 60772 224224 60784
rect 215168 60744 224224 60772
rect 215168 60732 215174 60744
rect 224218 60732 224224 60744
rect 224276 60732 224282 60784
rect 216766 60664 216772 60716
rect 216824 60704 216830 60716
rect 227438 60704 227444 60716
rect 216824 60676 227444 60704
rect 216824 60664 216830 60676
rect 227438 60664 227444 60676
rect 227496 60664 227502 60716
rect 224310 60596 224316 60648
rect 224368 60636 224374 60648
rect 227070 60636 227076 60648
rect 224368 60608 227076 60636
rect 224368 60596 224374 60608
rect 227070 60596 227076 60608
rect 227128 60596 227134 60648
rect 95050 59372 95056 59424
rect 95108 59412 95114 59424
rect 116394 59412 116400 59424
rect 95108 59384 116400 59412
rect 95108 59372 95114 59384
rect 116394 59372 116400 59384
rect 116452 59372 116458 59424
rect 214558 59372 214564 59424
rect 214616 59412 214622 59424
rect 217594 59412 217600 59424
rect 214616 59384 217600 59412
rect 214616 59372 214622 59384
rect 217594 59372 217600 59384
rect 217652 59372 217658 59424
rect 216950 59304 216956 59356
rect 217008 59344 217014 59356
rect 227530 59344 227536 59356
rect 217008 59316 227536 59344
rect 217008 59304 217014 59316
rect 227530 59304 227536 59316
rect 227588 59304 227594 59356
rect 224586 59236 224592 59288
rect 224644 59276 224650 59288
rect 227438 59276 227444 59288
rect 224644 59248 227444 59276
rect 224644 59236 224650 59248
rect 227438 59236 227444 59248
rect 227496 59236 227502 59288
rect 214098 58012 214104 58064
rect 214156 58052 214162 58064
rect 217502 58052 217508 58064
rect 214156 58024 217508 58052
rect 214156 58012 214162 58024
rect 217502 58012 217508 58024
rect 217560 58012 217566 58064
rect 94406 57944 94412 57996
rect 94464 57984 94470 57996
rect 116394 57984 116400 57996
rect 94464 57956 116400 57984
rect 94464 57944 94470 57956
rect 116394 57944 116400 57956
rect 116452 57944 116458 57996
rect 214190 57944 214196 57996
rect 214248 57984 214254 57996
rect 217410 57984 217416 57996
rect 214248 57956 217416 57984
rect 214248 57944 214254 57956
rect 217410 57944 217416 57956
rect 217468 57944 217474 57996
rect 216674 57876 216680 57928
rect 216732 57916 216738 57928
rect 227438 57916 227444 57928
rect 216732 57888 227444 57916
rect 216732 57876 216738 57888
rect 227438 57876 227444 57888
rect 227496 57876 227502 57928
rect 224034 57808 224040 57860
rect 224092 57848 224098 57860
rect 227254 57848 227260 57860
rect 224092 57820 227260 57848
rect 224092 57808 224098 57820
rect 227254 57808 227260 57820
rect 227312 57808 227318 57860
rect 213914 56652 213920 56704
rect 213972 56692 213978 56704
rect 216766 56692 216772 56704
rect 213972 56664 216772 56692
rect 213972 56652 213978 56664
rect 216766 56652 216772 56664
rect 216824 56652 216830 56704
rect 93854 56584 93860 56636
rect 93912 56624 93918 56636
rect 116302 56624 116308 56636
rect 93912 56596 116308 56624
rect 93912 56584 93918 56596
rect 116302 56584 116308 56596
rect 116360 56584 116366 56636
rect 214006 56584 214012 56636
rect 214064 56624 214070 56636
rect 216674 56624 216680 56636
rect 214064 56596 216680 56624
rect 214064 56584 214070 56596
rect 216674 56584 216680 56596
rect 216732 56584 216738 56636
rect 216858 56516 216864 56568
rect 216916 56556 216922 56568
rect 227438 56556 227444 56568
rect 216916 56528 227444 56556
rect 216916 56516 216922 56528
rect 227438 56516 227444 56528
rect 227496 56516 227502 56568
rect 224126 56448 224132 56500
rect 224184 56488 224190 56500
rect 227254 56488 227260 56500
rect 224184 56460 227260 56488
rect 224184 56448 224190 56460
rect 227254 56448 227260 56460
rect 227312 56448 227318 56500
rect 94038 55292 94044 55344
rect 94096 55332 94102 55344
rect 116394 55332 116400 55344
rect 94096 55304 116400 55332
rect 94096 55292 94102 55304
rect 116394 55292 116400 55304
rect 116452 55292 116458 55344
rect 93946 55224 93952 55276
rect 94004 55264 94010 55276
rect 116302 55264 116308 55276
rect 94004 55236 116308 55264
rect 94004 55224 94010 55236
rect 116302 55224 116308 55236
rect 116360 55224 116366 55276
rect 215110 55224 215116 55276
rect 215168 55264 215174 55276
rect 227530 55264 227536 55276
rect 215168 55236 227536 55264
rect 215168 55224 215174 55236
rect 227530 55224 227536 55236
rect 227588 55224 227594 55276
rect 217594 55156 217600 55208
rect 217652 55196 217658 55208
rect 217652 55168 224172 55196
rect 217652 55156 217658 55168
rect 224144 55060 224172 55168
rect 224218 55156 224224 55208
rect 224276 55196 224282 55208
rect 227438 55196 227444 55208
rect 224276 55168 227444 55196
rect 224276 55156 224282 55168
rect 227438 55156 227444 55168
rect 227496 55156 227502 55208
rect 226518 55060 226524 55072
rect 224144 55032 226524 55060
rect 226518 55020 226524 55032
rect 226576 55020 226582 55072
rect 215110 53864 215116 53916
rect 215168 53904 215174 53916
rect 226978 53904 226984 53916
rect 215168 53876 226984 53904
rect 215168 53864 215174 53876
rect 226978 53864 226984 53876
rect 227036 53864 227042 53916
rect 94774 53796 94780 53848
rect 94832 53836 94838 53848
rect 116394 53836 116400 53848
rect 94832 53808 116400 53836
rect 94832 53796 94838 53808
rect 116394 53796 116400 53808
rect 116452 53796 116458 53848
rect 214742 53796 214748 53848
rect 214800 53836 214806 53848
rect 226610 53836 226616 53848
rect 214800 53808 226616 53836
rect 214800 53796 214806 53808
rect 226610 53796 226616 53808
rect 226668 53796 226674 53848
rect 217502 53728 217508 53780
rect 217560 53768 217566 53780
rect 227438 53768 227444 53780
rect 217560 53740 227444 53768
rect 217560 53728 217566 53740
rect 227438 53728 227444 53740
rect 227496 53728 227502 53780
rect 217410 53660 217416 53712
rect 217468 53700 217474 53712
rect 226518 53700 226524 53712
rect 217468 53672 226524 53700
rect 217468 53660 217474 53672
rect 226518 53660 226524 53672
rect 226576 53660 226582 53712
rect 215110 52504 215116 52556
rect 215168 52544 215174 52556
rect 226794 52544 226800 52556
rect 215168 52516 226800 52544
rect 215168 52504 215174 52516
rect 226794 52504 226800 52516
rect 226852 52504 226858 52556
rect 95142 52436 95148 52488
rect 95200 52476 95206 52488
rect 116394 52476 116400 52488
rect 95200 52448 116400 52476
rect 95200 52436 95206 52448
rect 116394 52436 116400 52448
rect 116452 52436 116458 52488
rect 214742 52436 214748 52488
rect 214800 52476 214806 52488
rect 226702 52476 226708 52488
rect 214800 52448 226708 52476
rect 214800 52436 214806 52448
rect 226702 52436 226708 52448
rect 226760 52436 226766 52488
rect 216674 52368 216680 52420
rect 216732 52408 216738 52420
rect 227438 52408 227444 52420
rect 216732 52380 227444 52408
rect 216732 52368 216738 52380
rect 227438 52368 227444 52380
rect 227496 52368 227502 52420
rect 216766 52300 216772 52352
rect 216824 52340 216830 52352
rect 227254 52340 227260 52352
rect 216824 52312 227260 52340
rect 216824 52300 216830 52312
rect 227254 52300 227260 52312
rect 227312 52300 227318 52352
rect 215110 51144 215116 51196
rect 215168 51184 215174 51196
rect 226334 51184 226340 51196
rect 215168 51156 226340 51184
rect 215168 51144 215174 51156
rect 226334 51144 226340 51156
rect 226392 51144 226398 51196
rect 94222 51076 94228 51128
rect 94280 51116 94286 51128
rect 115934 51116 115940 51128
rect 94280 51088 115940 51116
rect 94280 51076 94286 51088
rect 115934 51076 115940 51088
rect 115992 51076 115998 51128
rect 214098 51076 214104 51128
rect 214156 51116 214162 51128
rect 226518 51116 226524 51128
rect 214156 51088 226524 51116
rect 214156 51076 214162 51088
rect 226518 51076 226524 51088
rect 226576 51076 226582 51128
rect 215110 49784 215116 49836
rect 215168 49824 215174 49836
rect 227622 49824 227628 49836
rect 215168 49796 227628 49824
rect 215168 49784 215174 49796
rect 227622 49784 227628 49796
rect 227680 49784 227686 49836
rect 95050 49716 95056 49768
rect 95108 49756 95114 49768
rect 116394 49756 116400 49768
rect 95108 49728 116400 49756
rect 95108 49716 95114 49728
rect 116394 49716 116400 49728
rect 116452 49716 116458 49768
rect 215202 49716 215208 49768
rect 215260 49756 215266 49768
rect 227530 49756 227536 49768
rect 215260 49728 227536 49756
rect 215260 49716 215266 49728
rect 227530 49716 227536 49728
rect 227588 49716 227594 49768
rect 94498 48356 94504 48408
rect 94556 48396 94562 48408
rect 116118 48396 116124 48408
rect 94556 48368 116124 48396
rect 94556 48356 94562 48368
rect 116118 48356 116124 48368
rect 116176 48356 116182 48408
rect 94406 48288 94412 48340
rect 94464 48328 94470 48340
rect 116394 48328 116400 48340
rect 94464 48300 116400 48328
rect 94464 48288 94470 48300
rect 116394 48288 116400 48300
rect 116452 48288 116458 48340
rect 215110 48288 215116 48340
rect 215168 48328 215174 48340
rect 227346 48328 227352 48340
rect 215168 48300 227352 48328
rect 215168 48288 215174 48300
rect 227346 48288 227352 48300
rect 227404 48288 227410 48340
rect 214742 46996 214748 47048
rect 214800 47036 214806 47048
rect 227438 47036 227444 47048
rect 214800 47008 227444 47036
rect 214800 46996 214806 47008
rect 227438 46996 227444 47008
rect 227496 46996 227502 47048
rect 94130 46928 94136 46980
rect 94188 46968 94194 46980
rect 116394 46968 116400 46980
rect 94188 46940 116400 46968
rect 94188 46928 94194 46940
rect 116394 46928 116400 46940
rect 116452 46928 116458 46980
rect 214006 46928 214012 46980
rect 214064 46968 214070 46980
rect 226702 46968 226708 46980
rect 214064 46940 226708 46968
rect 214064 46928 214070 46940
rect 226702 46928 226708 46940
rect 226760 46928 226766 46980
rect 215110 45636 215116 45688
rect 215168 45676 215174 45688
rect 227254 45676 227260 45688
rect 215168 45648 227260 45676
rect 215168 45636 215174 45648
rect 227254 45636 227260 45648
rect 227312 45636 227318 45688
rect 93946 45568 93952 45620
rect 94004 45608 94010 45620
rect 116394 45608 116400 45620
rect 94004 45580 116400 45608
rect 94004 45568 94010 45580
rect 116394 45568 116400 45580
rect 116452 45568 116458 45620
rect 215202 45568 215208 45620
rect 215260 45608 215266 45620
rect 227070 45608 227076 45620
rect 215260 45580 227076 45608
rect 215260 45568 215266 45580
rect 227070 45568 227076 45580
rect 227128 45568 227134 45620
rect 215202 44208 215208 44260
rect 215260 44248 215266 44260
rect 227438 44248 227444 44260
rect 215260 44220 227444 44248
rect 215260 44208 215266 44220
rect 227438 44208 227444 44220
rect 227496 44208 227502 44260
rect 94774 44140 94780 44192
rect 94832 44180 94838 44192
rect 116394 44180 116400 44192
rect 94832 44152 116400 44180
rect 94832 44140 94838 44152
rect 116394 44140 116400 44152
rect 116452 44140 116458 44192
rect 215110 44140 215116 44192
rect 215168 44180 215174 44192
rect 227530 44180 227536 44192
rect 215168 44152 227536 44180
rect 215168 44140 215174 44152
rect 227530 44140 227536 44152
rect 227588 44140 227594 44192
rect 94590 42780 94596 42832
rect 94648 42820 94654 42832
rect 115934 42820 115940 42832
rect 94648 42792 115940 42820
rect 94648 42780 94654 42792
rect 115934 42780 115940 42792
rect 115992 42780 115998 42832
rect 214374 42780 214380 42832
rect 214432 42820 214438 42832
rect 226426 42820 226432 42832
rect 214432 42792 226432 42820
rect 214432 42780 214438 42792
rect 226426 42780 226432 42792
rect 226484 42780 226490 42832
rect 215110 41488 215116 41540
rect 215168 41528 215174 41540
rect 226610 41528 226616 41540
rect 215168 41500 226616 41528
rect 215168 41488 215174 41500
rect 226610 41488 226616 41500
rect 226668 41488 226674 41540
rect 95142 41420 95148 41472
rect 95200 41460 95206 41472
rect 116394 41460 116400 41472
rect 95200 41432 116400 41460
rect 95200 41420 95206 41432
rect 116394 41420 116400 41432
rect 116452 41420 116458 41472
rect 214098 41420 214104 41472
rect 214156 41460 214162 41472
rect 226334 41460 226340 41472
rect 214156 41432 226340 41460
rect 214156 41420 214162 41432
rect 226334 41420 226340 41432
rect 226392 41420 226398 41472
rect 560938 41352 560944 41404
rect 560996 41392 561002 41404
rect 580166 41392 580172 41404
rect 560996 41364 580172 41392
rect 560996 41352 561002 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 94498 40128 94504 40180
rect 94556 40168 94562 40180
rect 116302 40168 116308 40180
rect 94556 40140 116308 40168
rect 94556 40128 94562 40140
rect 116302 40128 116308 40140
rect 116360 40128 116366 40180
rect 215110 40128 215116 40180
rect 215168 40168 215174 40180
rect 227438 40168 227444 40180
rect 215168 40140 227444 40168
rect 215168 40128 215174 40140
rect 227438 40128 227444 40140
rect 227496 40128 227502 40180
rect 95050 40060 95056 40112
rect 95108 40100 95114 40112
rect 116394 40100 116400 40112
rect 95108 40072 116400 40100
rect 95108 40060 95114 40072
rect 116394 40060 116400 40072
rect 116452 40060 116458 40112
rect 214650 40060 214656 40112
rect 214708 40100 214714 40112
rect 227070 40100 227076 40112
rect 214708 40072 227076 40100
rect 214708 40060 214714 40072
rect 227070 40060 227076 40072
rect 227128 40060 227134 40112
rect 215110 38700 215116 38752
rect 215168 38740 215174 38752
rect 227530 38740 227536 38752
rect 215168 38712 227536 38740
rect 215168 38700 215174 38712
rect 227530 38700 227536 38712
rect 227588 38700 227594 38752
rect 94590 38632 94596 38684
rect 94648 38672 94654 38684
rect 116394 38672 116400 38684
rect 94648 38644 116400 38672
rect 94648 38632 94654 38644
rect 116394 38632 116400 38644
rect 116452 38632 116458 38684
rect 214558 38632 214564 38684
rect 214616 38672 214622 38684
rect 226702 38672 226708 38684
rect 214616 38644 226708 38672
rect 214616 38632 214622 38644
rect 226702 38632 226708 38644
rect 226760 38632 226766 38684
rect 93854 37272 93860 37324
rect 93912 37312 93918 37324
rect 116394 37312 116400 37324
rect 93912 37284 116400 37312
rect 93912 37272 93918 37284
rect 116394 37272 116400 37284
rect 116452 37272 116458 37324
rect 215110 37272 215116 37324
rect 215168 37312 215174 37324
rect 227438 37312 227444 37324
rect 215168 37284 227444 37312
rect 215168 37272 215174 37284
rect 227438 37272 227444 37284
rect 227496 37272 227502 37324
rect 214098 35980 214104 36032
rect 214156 36020 214162 36032
rect 226702 36020 226708 36032
rect 214156 35992 226708 36020
rect 214156 35980 214162 35992
rect 226702 35980 226708 35992
rect 226760 35980 226766 36032
rect 93946 35912 93952 35964
rect 94004 35952 94010 35964
rect 116394 35952 116400 35964
rect 94004 35924 116400 35952
rect 94004 35912 94010 35924
rect 116394 35912 116400 35924
rect 116452 35912 116458 35964
rect 215110 35912 215116 35964
rect 215168 35952 215174 35964
rect 227438 35952 227444 35964
rect 215168 35924 227444 35952
rect 215168 35912 215174 35924
rect 227438 35912 227444 35924
rect 227496 35912 227502 35964
rect 215110 34552 215116 34604
rect 215168 34592 215174 34604
rect 227346 34592 227352 34604
rect 215168 34564 227352 34592
rect 215168 34552 215174 34564
rect 227346 34552 227352 34564
rect 227404 34552 227410 34604
rect 95142 34484 95148 34536
rect 95200 34524 95206 34536
rect 116394 34524 116400 34536
rect 95200 34496 116400 34524
rect 95200 34484 95206 34496
rect 116394 34484 116400 34496
rect 116452 34484 116458 34536
rect 214650 34484 214656 34536
rect 214708 34524 214714 34536
rect 227438 34524 227444 34536
rect 214708 34496 227444 34524
rect 214708 34484 214714 34496
rect 227438 34484 227444 34496
rect 227496 34484 227502 34536
rect 214558 33192 214564 33244
rect 214616 33232 214622 33244
rect 227438 33232 227444 33244
rect 214616 33204 227444 33232
rect 214616 33192 214622 33204
rect 227438 33192 227444 33204
rect 227496 33192 227502 33244
rect 95142 33124 95148 33176
rect 95200 33164 95206 33176
rect 116302 33164 116308 33176
rect 95200 33136 116308 33164
rect 95200 33124 95206 33136
rect 116302 33124 116308 33136
rect 116360 33124 116366 33176
rect 215110 33124 215116 33176
rect 215168 33164 215174 33176
rect 227530 33164 227536 33176
rect 215168 33136 227536 33164
rect 215168 33124 215174 33136
rect 227530 33124 227536 33136
rect 227588 33124 227594 33176
rect 213914 32512 213920 32564
rect 213972 32552 213978 32564
rect 215938 32552 215944 32564
rect 213972 32524 215944 32552
rect 213972 32512 213978 32524
rect 215938 32512 215944 32524
rect 215996 32512 216002 32564
rect 95142 32376 95148 32428
rect 95200 32416 95206 32428
rect 116394 32416 116400 32428
rect 95200 32388 116400 32416
rect 95200 32376 95206 32388
rect 116394 32376 116400 32388
rect 116452 32376 116458 32428
rect 215110 32376 215116 32428
rect 215168 32416 215174 32428
rect 227438 32416 227444 32428
rect 215168 32388 227444 32416
rect 215168 32376 215174 32388
rect 227438 32376 227444 32388
rect 227496 32376 227502 32428
rect 71682 31764 71688 31816
rect 71740 31804 71746 31816
rect 116394 31804 116400 31816
rect 71740 31776 116400 31804
rect 71740 31764 71746 31776
rect 116394 31764 116400 31776
rect 116452 31764 116458 31816
rect 29914 31288 29920 31340
rect 29972 31328 29978 31340
rect 32306 31328 32312 31340
rect 29972 31300 32312 31328
rect 29972 31288 29978 31300
rect 32306 31288 32312 31300
rect 32364 31328 32370 31340
rect 38565 31331 38623 31337
rect 38565 31328 38577 31331
rect 32364 31300 38577 31328
rect 32364 31288 32370 31300
rect 38565 31297 38577 31300
rect 38611 31297 38623 31331
rect 38565 31291 38623 31297
rect 105538 30268 105544 30320
rect 105596 30308 105602 30320
rect 195422 30308 195428 30320
rect 105596 30280 195428 30308
rect 105596 30268 105602 30280
rect 195422 30268 195428 30280
rect 195480 30268 195486 30320
rect 95878 30200 95884 30252
rect 95936 30240 95942 30252
rect 185026 30240 185032 30252
rect 95936 30212 185032 30240
rect 95936 30200 95942 30212
rect 185026 30200 185032 30212
rect 185084 30200 185090 30252
rect 50338 30132 50344 30184
rect 50396 30172 50402 30184
rect 133141 30175 133199 30181
rect 133141 30172 133153 30175
rect 50396 30144 133153 30172
rect 50396 30132 50402 30144
rect 133141 30141 133153 30144
rect 133187 30141 133199 30175
rect 133141 30135 133199 30141
rect 163498 30132 163504 30184
rect 163556 30172 163562 30184
rect 174630 30172 174636 30184
rect 163556 30144 174636 30172
rect 163556 30132 163562 30144
rect 174630 30132 174636 30144
rect 174688 30132 174694 30184
rect 82078 30064 82084 30116
rect 82136 30104 82142 30116
rect 177206 30104 177212 30116
rect 82136 30076 177212 30104
rect 82136 30064 82142 30076
rect 177206 30064 177212 30076
rect 177264 30064 177270 30116
rect 53098 29996 53104 30048
rect 53156 30036 53162 30048
rect 148594 30036 148600 30048
rect 53156 30008 148600 30036
rect 53156 29996 53162 30008
rect 148594 29996 148600 30008
rect 148652 29996 148658 30048
rect 164878 29996 164884 30048
rect 164936 30036 164942 30048
rect 179782 30036 179788 30048
rect 164936 30008 179788 30036
rect 164936 29996 164942 30008
rect 179782 29996 179788 30008
rect 179840 29996 179846 30048
rect 75178 29928 75184 29980
rect 75236 29968 75242 29980
rect 172054 29968 172060 29980
rect 75236 29940 172060 29968
rect 75236 29928 75242 29940
rect 172054 29928 172060 29940
rect 172112 29928 172118 29980
rect 31018 29860 31024 29912
rect 31076 29900 31082 29912
rect 127710 29900 127716 29912
rect 31076 29872 127716 29900
rect 31076 29860 31082 29872
rect 127710 29860 127716 29872
rect 127768 29860 127774 29912
rect 133141 29903 133199 29909
rect 133141 29869 133153 29903
rect 133187 29900 133199 29903
rect 143350 29900 143356 29912
rect 133187 29872 143356 29900
rect 133187 29869 133199 29872
rect 133141 29863 133199 29869
rect 143350 29860 143356 29872
rect 143408 29860 143414 29912
rect 166258 29860 166264 29912
rect 166316 29900 166322 29912
rect 182450 29900 182456 29912
rect 166316 29872 182456 29900
rect 166316 29860 166322 29872
rect 182450 29860 182456 29872
rect 182508 29860 182514 29912
rect 66898 29792 66904 29844
rect 66956 29832 66962 29844
rect 166810 29832 166816 29844
rect 66956 29804 166816 29832
rect 66956 29792 66962 29804
rect 166810 29792 166816 29804
rect 166868 29792 166874 29844
rect 169110 29792 169116 29844
rect 169168 29832 169174 29844
rect 187602 29832 187608 29844
rect 169168 29804 187608 29832
rect 169168 29792 169174 29804
rect 187602 29792 187608 29804
rect 187660 29792 187666 29844
rect 25498 29724 25504 29776
rect 25556 29764 25562 29776
rect 126882 29764 126888 29776
rect 25556 29736 126888 29764
rect 25556 29724 25562 29736
rect 126882 29724 126888 29736
rect 126940 29724 126946 29776
rect 169018 29724 169024 29776
rect 169076 29764 169082 29776
rect 192846 29764 192852 29776
rect 169076 29736 192852 29764
rect 169076 29724 169082 29736
rect 192846 29724 192852 29736
rect 192904 29724 192910 29776
rect 59998 29656 60004 29708
rect 60056 29696 60062 29708
rect 161566 29696 161572 29708
rect 60056 29668 161572 29696
rect 60056 29656 60062 29668
rect 161566 29656 161572 29668
rect 161624 29656 161630 29708
rect 171778 29656 171784 29708
rect 171836 29696 171842 29708
rect 198090 29696 198096 29708
rect 171836 29668 198096 29696
rect 171836 29656 171842 29668
rect 198090 29656 198096 29668
rect 198148 29656 198154 29708
rect 28258 29588 28264 29640
rect 28316 29628 28322 29640
rect 130378 29628 130384 29640
rect 28316 29600 130384 29628
rect 28316 29588 28322 29600
rect 130378 29588 130384 29600
rect 130436 29588 130442 29640
rect 173158 29588 173164 29640
rect 173216 29628 173222 29640
rect 205818 29628 205824 29640
rect 173216 29600 205824 29628
rect 173216 29588 173222 29600
rect 205818 29588 205824 29600
rect 205876 29588 205882 29640
rect 89717 29563 89775 29569
rect 89717 29560 89729 29563
rect 89640 29532 89729 29560
rect 80057 29495 80115 29501
rect 80057 29461 80069 29495
rect 80103 29492 80115 29495
rect 89640 29492 89668 29532
rect 89717 29529 89729 29532
rect 89763 29529 89775 29563
rect 89717 29523 89775 29529
rect 111702 29520 111708 29572
rect 111760 29560 111766 29572
rect 200666 29560 200672 29572
rect 111760 29532 200672 29560
rect 111760 29520 111766 29532
rect 200666 29520 200672 29532
rect 200724 29520 200730 29572
rect 80103 29464 89668 29492
rect 102612 29464 102824 29492
rect 80103 29461 80115 29464
rect 80057 29455 80115 29461
rect 46198 29384 46204 29436
rect 46256 29424 46262 29436
rect 102612 29424 102640 29464
rect 46256 29396 102640 29424
rect 102796 29424 102824 29464
rect 115842 29452 115848 29504
rect 115900 29492 115906 29504
rect 203242 29492 203248 29504
rect 115900 29464 203248 29492
rect 115900 29452 115906 29464
rect 203242 29452 203248 29464
rect 203300 29452 203306 29504
rect 133782 29424 133788 29436
rect 102796 29396 133788 29424
rect 46256 29384 46262 29396
rect 133782 29384 133788 29396
rect 133840 29384 133846 29436
rect 57977 29359 58035 29365
rect 57977 29356 57989 29359
rect 51000 29328 57989 29356
rect 51000 29152 51028 29328
rect 57977 29325 57989 29328
rect 58023 29325 58035 29359
rect 80057 29359 80115 29365
rect 80057 29356 80069 29359
rect 57977 29319 58035 29325
rect 74552 29328 80069 29356
rect 74445 29291 74503 29297
rect 74445 29257 74457 29291
rect 74491 29288 74503 29291
rect 74552 29288 74580 29328
rect 80057 29325 80069 29328
rect 80103 29325 80115 29359
rect 80057 29319 80115 29325
rect 89717 29359 89775 29365
rect 89717 29325 89729 29359
rect 89763 29356 89775 29359
rect 89763 29328 102732 29356
rect 89763 29325 89775 29328
rect 89717 29319 89775 29325
rect 74491 29260 74580 29288
rect 102704 29288 102732 29328
rect 102778 29316 102784 29368
rect 102836 29356 102842 29368
rect 190270 29356 190276 29368
rect 102836 29328 190276 29356
rect 102836 29316 102842 29328
rect 190270 29316 190276 29328
rect 190328 29316 190334 29368
rect 109957 29291 110015 29297
rect 109957 29288 109969 29291
rect 102704 29260 109969 29288
rect 74491 29257 74503 29260
rect 74445 29251 74503 29257
rect 109957 29257 109969 29260
rect 110003 29257 110015 29291
rect 109957 29251 110015 29257
rect 117958 29248 117964 29300
rect 118016 29288 118022 29300
rect 121457 29291 121515 29297
rect 121457 29288 121469 29291
rect 118016 29260 121469 29288
rect 118016 29248 118022 29260
rect 121457 29257 121469 29260
rect 121503 29257 121515 29291
rect 121457 29251 121515 29257
rect 122742 29248 122748 29300
rect 122800 29288 122806 29300
rect 208486 29288 208492 29300
rect 122800 29260 208492 29288
rect 122800 29248 122806 29260
rect 208486 29248 208492 29260
rect 208544 29248 208550 29300
rect 68002 29180 68008 29232
rect 68060 29220 68066 29232
rect 74537 29223 74595 29229
rect 74537 29220 74549 29223
rect 68060 29192 74549 29220
rect 68060 29180 68066 29192
rect 74537 29189 74549 29192
rect 74583 29189 74595 29223
rect 74537 29183 74595 29189
rect 83001 29223 83059 29229
rect 83001 29189 83013 29223
rect 83047 29220 83059 29223
rect 94225 29223 94283 29229
rect 94225 29220 94237 29223
rect 83047 29192 94237 29220
rect 83047 29189 83059 29192
rect 83001 29183 83059 29189
rect 94225 29189 94237 29192
rect 94271 29189 94283 29223
rect 94225 29183 94283 29189
rect 104161 29223 104219 29229
rect 104161 29189 104173 29223
rect 104207 29220 104219 29223
rect 123386 29220 123392 29232
rect 104207 29192 123392 29220
rect 104207 29189 104219 29192
rect 104161 29183 104219 29189
rect 123386 29180 123392 29192
rect 123444 29180 123450 29232
rect 125502 29180 125508 29232
rect 125560 29220 125566 29232
rect 211062 29220 211068 29232
rect 125560 29192 211068 29220
rect 125560 29180 125566 29192
rect 211062 29180 211068 29192
rect 211120 29180 211126 29232
rect 42628 29124 51028 29152
rect 38565 29087 38623 29093
rect 38565 29053 38577 29087
rect 38611 29084 38623 29087
rect 41325 29087 41383 29093
rect 41325 29084 41337 29087
rect 38611 29056 41337 29084
rect 38611 29053 38623 29056
rect 38565 29047 38623 29053
rect 41325 29053 41337 29056
rect 41371 29053 41383 29087
rect 41325 29047 41383 29053
rect 41417 29087 41475 29093
rect 41417 29053 41429 29087
rect 41463 29084 41475 29087
rect 42628 29084 42656 29124
rect 57238 29112 57244 29164
rect 57296 29152 57302 29164
rect 131206 29152 131212 29164
rect 57296 29124 131212 29152
rect 57296 29112 57302 29124
rect 131206 29112 131212 29124
rect 131264 29112 131270 29164
rect 41463 29056 42656 29084
rect 41463 29053 41475 29056
rect 41417 29047 41475 29053
rect 61378 29044 61384 29096
rect 61436 29084 61442 29096
rect 134702 29084 134708 29096
rect 61436 29056 134708 29084
rect 61436 29044 61442 29056
rect 134702 29044 134708 29056
rect 134760 29044 134766 29096
rect 162118 29044 162124 29096
rect 162176 29084 162182 29096
rect 162176 29056 164464 29084
rect 162176 29044 162182 29056
rect 57977 29019 58035 29025
rect 57977 28985 57989 29019
rect 58023 29016 58035 29019
rect 74445 29019 74503 29025
rect 74445 29016 74457 29019
rect 58023 28988 74457 29016
rect 58023 28985 58035 28988
rect 57977 28979 58035 28985
rect 74445 28985 74457 28988
rect 74491 28985 74503 29019
rect 74445 28979 74503 28985
rect 74537 29019 74595 29025
rect 74537 28985 74549 29019
rect 74583 29016 74595 29019
rect 83001 29019 83059 29025
rect 83001 29016 83013 29019
rect 74583 28988 83013 29016
rect 74583 28985 74595 28988
rect 74537 28979 74595 28985
rect 83001 28985 83013 28988
rect 83047 28985 83059 29019
rect 83001 28979 83059 28985
rect 94225 29019 94283 29025
rect 94225 28985 94237 29019
rect 94271 29016 94283 29019
rect 104161 29019 104219 29025
rect 104161 29016 104173 29019
rect 94271 28988 104173 29016
rect 94271 28985 94283 28988
rect 94225 28979 94283 28985
rect 104161 28985 104173 28988
rect 104207 28985 104219 29019
rect 104161 28979 104219 28985
rect 109957 29019 110015 29025
rect 109957 28985 109969 29019
rect 110003 29016 110015 29019
rect 119982 29016 119988 29028
rect 110003 28988 119988 29016
rect 110003 28985 110015 28988
rect 109957 28979 110015 28985
rect 119982 28976 119988 28988
rect 120040 28976 120046 29028
rect 121457 29019 121515 29025
rect 121457 28985 121469 29019
rect 121503 29016 121515 29019
rect 124306 29016 124312 29028
rect 121503 28988 124312 29016
rect 121503 28985 121515 28988
rect 121457 28979 121515 28985
rect 124306 28976 124312 28988
rect 124364 28976 124370 29028
rect 152458 28976 152464 29028
rect 152516 29016 152522 29028
rect 156414 29016 156420 29028
rect 152516 28988 156420 29016
rect 152516 28976 152522 28988
rect 156414 28976 156420 28988
rect 156472 28976 156478 29028
rect 156598 28976 156604 29028
rect 156656 29016 156662 29028
rect 158990 29016 158996 29028
rect 156656 28988 158996 29016
rect 156656 28976 156662 28988
rect 158990 28976 158996 28988
rect 159048 28976 159054 29028
rect 159358 28976 159364 29028
rect 159416 29016 159422 29028
rect 164234 29016 164240 29028
rect 159416 28988 164240 29016
rect 159416 28976 159422 28988
rect 164234 28976 164240 28988
rect 164292 28976 164298 29028
rect 164436 29016 164464 29056
rect 169386 29016 169392 29028
rect 164436 28988 169392 29016
rect 169386 28976 169392 28988
rect 169444 28976 169450 29028
rect 68002 28948 68008 28960
rect 67963 28920 68008 28948
rect 68002 28908 68008 28920
rect 68060 28908 68066 28960
rect 103422 28364 103428 28416
rect 103480 28404 103486 28416
rect 194594 28404 194600 28416
rect 103480 28376 194600 28404
rect 103480 28364 103486 28376
rect 194594 28364 194600 28376
rect 194652 28364 194658 28416
rect 60642 28296 60648 28348
rect 60700 28336 60706 28348
rect 163314 28336 163320 28348
rect 60700 28308 163320 28336
rect 60700 28296 60706 28308
rect 163314 28296 163320 28308
rect 163372 28296 163378 28348
rect 10318 28228 10324 28280
rect 10376 28268 10382 28280
rect 121638 28268 121644 28280
rect 10376 28240 121644 28268
rect 10376 28228 10382 28240
rect 121638 28228 121644 28240
rect 121696 28228 121702 28280
rect 3418 27548 3424 27600
rect 3476 27588 3482 27600
rect 411254 27588 411260 27600
rect 3476 27560 411260 27588
rect 3476 27548 3482 27560
rect 411254 27548 411260 27560
rect 411312 27548 411318 27600
rect 110322 26868 110328 26920
rect 110380 26908 110386 26920
rect 199746 26908 199752 26920
rect 110380 26880 199752 26908
rect 110380 26868 110386 26880
rect 199746 26868 199752 26880
rect 199804 26868 199810 26920
rect 138106 26732 138112 26784
rect 138164 26772 138170 26784
rect 138750 26772 138756 26784
rect 138164 26744 138756 26772
rect 138164 26732 138170 26744
rect 138750 26732 138756 26744
rect 138808 26732 138814 26784
rect 144914 26732 144920 26784
rect 144972 26772 144978 26784
rect 145742 26772 145748 26784
rect 144972 26744 145748 26772
rect 144972 26732 144978 26744
rect 145742 26732 145748 26744
rect 145800 26732 145806 26784
rect 149054 26732 149060 26784
rect 149112 26772 149118 26784
rect 149974 26772 149980 26784
rect 149112 26744 149980 26772
rect 149112 26732 149118 26744
rect 149974 26732 149980 26744
rect 150032 26732 150038 26784
rect 154574 26732 154580 26784
rect 154632 26772 154638 26784
rect 155126 26772 155132 26784
rect 154632 26744 155132 26772
rect 154632 26732 154638 26744
rect 155126 26732 155132 26744
rect 155184 26732 155190 26784
rect 183557 26231 183615 26237
rect 183557 26197 183569 26231
rect 183603 26228 183615 26231
rect 197170 26228 197176 26240
rect 183603 26200 197176 26228
rect 183603 26197 183615 26200
rect 183557 26191 183615 26197
rect 197170 26188 197176 26200
rect 197228 26188 197234 26240
rect 172517 25891 172575 25897
rect 172517 25857 172529 25891
rect 172563 25888 172575 25891
rect 182085 25891 182143 25897
rect 182085 25888 182097 25891
rect 172563 25860 182097 25888
rect 172563 25857 172575 25860
rect 172517 25851 172575 25857
rect 182085 25857 182097 25860
rect 182131 25857 182143 25891
rect 182085 25851 182143 25857
rect 144733 25823 144791 25829
rect 144733 25820 144745 25823
rect 135272 25792 144745 25820
rect 115845 25755 115903 25761
rect 115845 25721 115857 25755
rect 115891 25721 115903 25755
rect 115845 25715 115903 25721
rect 128357 25755 128415 25761
rect 128357 25721 128369 25755
rect 128403 25752 128415 25755
rect 135272 25752 135300 25792
rect 144733 25789 144745 25792
rect 144779 25789 144791 25823
rect 144733 25783 144791 25789
rect 183557 25823 183615 25829
rect 183557 25789 183569 25823
rect 183603 25789 183615 25823
rect 183557 25783 183615 25789
rect 128403 25724 135300 25752
rect 144825 25755 144883 25761
rect 128403 25721 128415 25724
rect 128357 25715 128415 25721
rect 144825 25721 144837 25755
rect 144871 25721 144883 25755
rect 144825 25715 144883 25721
rect 169021 25755 169079 25761
rect 169021 25721 169033 25755
rect 169067 25752 169079 25755
rect 172517 25755 172575 25761
rect 172517 25752 172529 25755
rect 169067 25724 172529 25752
rect 169067 25721 169079 25724
rect 169021 25715 169079 25721
rect 172517 25721 172529 25724
rect 172563 25721 172575 25755
rect 172517 25715 172575 25721
rect 182085 25755 182143 25761
rect 182085 25721 182097 25755
rect 182131 25752 182143 25755
rect 183572 25752 183600 25783
rect 182131 25724 183600 25752
rect 182131 25721 182143 25724
rect 182085 25715 182143 25721
rect 115860 25684 115888 25715
rect 128265 25687 128323 25693
rect 128265 25684 128277 25687
rect 115860 25656 128277 25684
rect 128265 25653 128277 25656
rect 128311 25653 128323 25687
rect 144840 25684 144868 25715
rect 164237 25687 164295 25693
rect 164237 25684 164249 25687
rect 144840 25656 164249 25684
rect 128265 25647 128323 25653
rect 164237 25653 164249 25656
rect 164283 25653 164295 25687
rect 164237 25647 164295 25653
rect 67542 25576 67548 25628
rect 67600 25616 67606 25628
rect 168558 25616 168564 25628
rect 67600 25588 168564 25616
rect 67600 25576 67606 25588
rect 168558 25576 168564 25588
rect 168616 25576 168622 25628
rect 11698 25508 11704 25560
rect 11756 25548 11762 25560
rect 125134 25548 125140 25560
rect 11756 25520 125140 25548
rect 11756 25508 11762 25520
rect 125134 25508 125140 25520
rect 125192 25508 125198 25560
rect 164237 25483 164295 25489
rect 164237 25449 164249 25483
rect 164283 25480 164295 25483
rect 169021 25483 169079 25489
rect 169021 25480 169033 25483
rect 164283 25452 169033 25480
rect 164283 25449 164295 25452
rect 164237 25443 164295 25449
rect 169021 25449 169033 25452
rect 169067 25449 169079 25483
rect 169021 25443 169079 25449
rect 114462 24216 114468 24268
rect 114520 24256 114526 24268
rect 202414 24256 202420 24268
rect 114520 24228 202420 24256
rect 114520 24216 114526 24228
rect 202414 24216 202420 24228
rect 202472 24216 202478 24268
rect 74442 24148 74448 24200
rect 74500 24188 74506 24200
rect 173710 24188 173716 24200
rect 74500 24160 173716 24188
rect 74500 24148 74506 24160
rect 173710 24148 173716 24160
rect 173768 24148 173774 24200
rect 52362 24080 52368 24132
rect 52420 24120 52426 24132
rect 157242 24120 157248 24132
rect 52420 24092 157248 24120
rect 52420 24080 52426 24092
rect 157242 24080 157248 24092
rect 157300 24080 157306 24132
rect 125410 22856 125416 22908
rect 125468 22896 125474 22908
rect 210234 22896 210240 22908
rect 125468 22868 210240 22896
rect 125468 22856 125474 22868
rect 210234 22856 210240 22868
rect 210292 22856 210298 22908
rect 85482 22788 85488 22840
rect 85540 22828 85546 22840
rect 181530 22828 181536 22840
rect 85540 22800 181536 22828
rect 85540 22788 85546 22800
rect 181530 22788 181536 22800
rect 181588 22788 181594 22840
rect 63402 22720 63408 22772
rect 63460 22760 63466 22772
rect 165062 22760 165068 22772
rect 63460 22732 165068 22760
rect 63460 22720 63466 22732
rect 165062 22720 165068 22732
rect 165120 22720 165126 22772
rect 121454 22448 121460 22500
rect 121512 22488 121518 22500
rect 122190 22488 122196 22500
rect 121512 22460 122196 22488
rect 121512 22448 121518 22460
rect 122190 22448 122196 22460
rect 122248 22448 122254 22500
rect 203058 22108 203064 22160
rect 203116 22148 203122 22160
rect 203886 22148 203892 22160
rect 203116 22120 203892 22148
rect 203116 22108 203122 22120
rect 203886 22108 203892 22120
rect 203944 22108 203950 22160
rect 121454 22040 121460 22092
rect 121512 22080 121518 22092
rect 121638 22080 121644 22092
rect 121512 22052 121644 22080
rect 121512 22040 121518 22052
rect 121638 22040 121644 22052
rect 121696 22040 121702 22092
rect 96522 21428 96528 21480
rect 96580 21468 96586 21480
rect 189166 21468 189172 21480
rect 96580 21440 189172 21468
rect 96580 21428 96586 21440
rect 189166 21428 189172 21440
rect 189224 21428 189230 21480
rect 59262 21360 59268 21412
rect 59320 21400 59326 21412
rect 161566 21400 161572 21412
rect 59320 21372 161572 21400
rect 59320 21360 59326 21372
rect 161566 21360 161572 21372
rect 161624 21360 161630 21412
rect 107562 20680 107568 20732
rect 107620 20720 107626 20732
rect 115845 20723 115903 20729
rect 115845 20720 115857 20723
rect 107620 20692 115857 20720
rect 107620 20680 107626 20692
rect 115845 20689 115857 20692
rect 115891 20689 115903 20723
rect 115845 20683 115903 20689
rect 99190 20000 99196 20052
rect 99248 20040 99254 20052
rect 191926 20040 191932 20052
rect 99248 20012 191932 20040
rect 99248 20000 99254 20012
rect 191926 20000 191932 20012
rect 191984 20000 191990 20052
rect 66162 19932 66168 19984
rect 66220 19972 66226 19984
rect 166994 19972 167000 19984
rect 66220 19944 167000 19972
rect 66220 19932 66226 19944
rect 166994 19932 167000 19944
rect 167052 19932 167058 19984
rect 68005 19363 68063 19369
rect 68005 19329 68017 19363
rect 68051 19360 68063 19363
rect 68094 19360 68100 19372
rect 68051 19332 68100 19360
rect 68051 19329 68063 19332
rect 68005 19323 68063 19329
rect 68094 19320 68100 19332
rect 68152 19320 68158 19372
rect 65981 19295 66039 19301
rect 65981 19261 65993 19295
rect 66027 19292 66039 19295
rect 66162 19292 66168 19304
rect 66027 19264 66168 19292
rect 66027 19261 66039 19264
rect 65981 19255 66039 19261
rect 66162 19252 66168 19264
rect 66220 19252 66226 19304
rect 121638 19292 121644 19304
rect 121599 19264 121644 19292
rect 121638 19252 121644 19264
rect 121696 19252 121702 19304
rect 182177 19295 182235 19301
rect 182177 19261 182189 19295
rect 182223 19292 182235 19295
rect 182266 19292 182272 19304
rect 182223 19264 182272 19292
rect 182223 19261 182235 19264
rect 182177 19255 182235 19261
rect 182266 19252 182272 19264
rect 182324 19252 182330 19304
rect 184566 19252 184572 19304
rect 184624 19292 184630 19304
rect 185026 19292 185032 19304
rect 184624 19264 185032 19292
rect 184624 19252 184630 19264
rect 185026 19252 185032 19264
rect 185084 19252 185090 19304
rect 117130 18708 117136 18760
rect 117188 18748 117194 18760
rect 204254 18748 204260 18760
rect 117188 18720 204260 18748
rect 117188 18708 117194 18720
rect 204254 18708 204260 18720
rect 204312 18708 204318 18760
rect 89622 18640 89628 18692
rect 89680 18680 89686 18692
rect 183554 18680 183560 18692
rect 89680 18652 183560 18680
rect 89680 18640 89686 18652
rect 183554 18640 183560 18652
rect 183612 18640 183618 18692
rect 53742 18572 53748 18624
rect 53800 18612 53806 18624
rect 157334 18612 157340 18624
rect 53800 18584 157340 18612
rect 53800 18572 53806 18584
rect 157334 18572 157340 18584
rect 157392 18572 157398 18624
rect 121362 17348 121368 17400
rect 121420 17388 121426 17400
rect 207014 17388 207020 17400
rect 121420 17360 207020 17388
rect 121420 17348 121426 17360
rect 207014 17348 207020 17360
rect 207072 17348 207078 17400
rect 92382 17280 92388 17332
rect 92440 17320 92446 17332
rect 186406 17320 186412 17332
rect 92440 17292 186412 17320
rect 92440 17280 92446 17292
rect 186406 17280 186412 17292
rect 186464 17280 186470 17332
rect 56502 17212 56508 17264
rect 56560 17252 56566 17264
rect 158806 17252 158812 17264
rect 56560 17224 158812 17252
rect 56560 17212 56566 17224
rect 158806 17212 158812 17224
rect 158864 17212 158870 17264
rect 492858 16396 492864 16448
rect 492916 16436 492922 16448
rect 493594 16436 493600 16448
rect 492916 16408 493600 16436
rect 492916 16396 492922 16408
rect 493594 16396 493600 16408
rect 493652 16396 493658 16448
rect 378042 16328 378048 16380
rect 378100 16368 378106 16380
rect 494790 16368 494796 16380
rect 378100 16340 494796 16368
rect 378100 16328 378106 16340
rect 494790 16328 494796 16340
rect 494848 16328 494854 16380
rect 318058 16260 318064 16312
rect 318116 16300 318122 16312
rect 458358 16300 458364 16312
rect 318116 16272 458364 16300
rect 318116 16260 318122 16272
rect 458358 16260 458364 16272
rect 458416 16260 458422 16312
rect 300118 16192 300124 16244
rect 300176 16232 300182 16244
rect 456334 16232 456340 16244
rect 300176 16204 456340 16232
rect 300176 16192 300182 16204
rect 456334 16192 456340 16204
rect 456392 16192 456398 16244
rect 286318 16124 286324 16176
rect 286376 16164 286382 16176
rect 452838 16164 452844 16176
rect 286376 16136 452844 16164
rect 286376 16124 286382 16136
rect 452838 16124 452844 16136
rect 452896 16124 452902 16176
rect 296622 16056 296628 16108
rect 296680 16096 296686 16108
rect 468570 16096 468576 16108
rect 296680 16068 468576 16096
rect 296680 16056 296686 16068
rect 468570 16056 468576 16068
rect 468628 16056 468634 16108
rect 285582 15988 285588 16040
rect 285640 16028 285646 16040
rect 465166 16028 465172 16040
rect 285640 16000 465172 16028
rect 285640 15988 285646 16000
rect 465166 15988 465172 16000
rect 465224 15988 465230 16040
rect 82722 15920 82728 15972
rect 82780 15960 82786 15972
rect 178126 15960 178132 15972
rect 82780 15932 178132 15960
rect 82780 15920 82786 15932
rect 178126 15920 178132 15932
rect 178184 15920 178190 15972
rect 280062 15920 280068 15972
rect 280120 15960 280126 15972
rect 463602 15960 463608 15972
rect 280120 15932 463608 15960
rect 280120 15920 280126 15932
rect 463602 15920 463608 15932
rect 463660 15920 463666 15972
rect 48222 15852 48228 15904
rect 48280 15892 48286 15904
rect 154666 15892 154672 15904
rect 48280 15864 154672 15892
rect 48280 15852 48286 15864
rect 154666 15852 154672 15864
rect 154724 15852 154730 15904
rect 278682 15852 278688 15904
rect 278740 15892 278746 15904
rect 462866 15892 462872 15904
rect 278740 15864 462872 15892
rect 278740 15852 278746 15864
rect 462866 15852 462872 15864
rect 462924 15852 462930 15904
rect 273162 15784 273168 15836
rect 273220 15824 273226 15836
rect 461302 15824 461308 15836
rect 273220 15796 461308 15824
rect 273220 15784 273226 15796
rect 461302 15784 461308 15796
rect 461360 15784 461366 15836
rect 266262 15716 266268 15768
rect 266320 15756 266326 15768
rect 459002 15756 459008 15768
rect 266320 15728 459008 15756
rect 266320 15716 266326 15728
rect 459002 15716 459008 15728
rect 459060 15716 459066 15768
rect 259362 15648 259368 15700
rect 259420 15688 259426 15700
rect 456702 15688 456708 15700
rect 259420 15660 456708 15688
rect 259420 15648 259426 15660
rect 456702 15648 456708 15660
rect 456760 15648 456766 15700
rect 240042 15580 240048 15632
rect 240100 15620 240106 15632
rect 450538 15620 450544 15632
rect 240100 15592 450544 15620
rect 240100 15580 240106 15592
rect 450538 15580 450544 15592
rect 450596 15580 450602 15632
rect 233142 15512 233148 15564
rect 233200 15552 233206 15564
rect 448238 15552 448244 15564
rect 233200 15524 448244 15552
rect 233200 15512 233206 15524
rect 448238 15512 448244 15524
rect 448296 15512 448302 15564
rect 222102 15444 222108 15496
rect 222160 15484 222166 15496
rect 444834 15484 444840 15496
rect 222160 15456 444840 15484
rect 222160 15444 222166 15456
rect 444834 15444 444840 15456
rect 444892 15444 444898 15496
rect 202782 15376 202788 15428
rect 202840 15416 202846 15428
rect 438670 15416 438676 15428
rect 202840 15388 438676 15416
rect 202840 15376 202846 15388
rect 438670 15376 438676 15388
rect 438728 15376 438734 15428
rect 204162 15308 204168 15360
rect 204220 15348 204226 15360
rect 439038 15348 439044 15360
rect 204220 15320 439044 15348
rect 204220 15308 204226 15320
rect 439038 15308 439044 15320
rect 439096 15308 439102 15360
rect 195882 15240 195888 15292
rect 195940 15280 195946 15292
rect 436370 15280 436376 15292
rect 195940 15252 436376 15280
rect 195940 15240 195946 15252
rect 436370 15240 436376 15252
rect 436428 15240 436434 15292
rect 188982 15172 188988 15224
rect 189040 15212 189046 15224
rect 434070 15212 434076 15224
rect 189040 15184 434076 15212
rect 189040 15172 189046 15184
rect 434070 15172 434076 15184
rect 434128 15172 434134 15224
rect 456978 15172 456984 15224
rect 457036 15212 457042 15224
rect 457438 15212 457444 15224
rect 457036 15184 457444 15212
rect 457036 15172 457042 15184
rect 457438 15172 457444 15184
rect 457496 15172 457502 15224
rect 354582 15104 354588 15156
rect 354640 15144 354646 15156
rect 487338 15144 487344 15156
rect 354640 15116 487344 15144
rect 354640 15104 354646 15116
rect 487338 15104 487344 15116
rect 487396 15104 487402 15156
rect 503622 15104 503628 15156
rect 503680 15144 503686 15156
rect 535638 15144 535644 15156
rect 503680 15116 535644 15144
rect 503680 15104 503686 15116
rect 535638 15104 535644 15116
rect 535696 15104 535702 15156
rect 538122 15104 538128 15156
rect 538180 15144 538186 15156
rect 546770 15144 546776 15156
rect 538180 15116 546776 15144
rect 538180 15104 538186 15116
rect 546770 15104 546776 15116
rect 546828 15104 546834 15156
rect 340782 15036 340788 15088
rect 340840 15076 340846 15088
rect 482738 15076 482744 15088
rect 340840 15048 482744 15076
rect 340840 15036 340846 15048
rect 482738 15036 482744 15048
rect 482796 15036 482802 15088
rect 489822 15036 489828 15088
rect 489880 15076 489886 15088
rect 531038 15076 531044 15088
rect 489880 15048 531044 15076
rect 489880 15036 489886 15048
rect 531038 15036 531044 15048
rect 531096 15036 531102 15088
rect 535362 15036 535368 15088
rect 535420 15076 535426 15088
rect 545666 15076 545672 15088
rect 535420 15048 545672 15076
rect 535420 15036 535426 15048
rect 545666 15036 545672 15048
rect 545724 15036 545730 15088
rect 332502 14968 332508 15020
rect 332560 15008 332566 15020
rect 480438 15008 480444 15020
rect 332560 14980 480444 15008
rect 332560 14968 332566 14980
rect 480438 14968 480444 14980
rect 480496 14968 480502 15020
rect 496722 14968 496728 15020
rect 496780 15008 496786 15020
rect 533338 15008 533344 15020
rect 496780 14980 533344 15008
rect 496780 14968 496786 14980
rect 533338 14968 533344 14980
rect 533396 14968 533402 15020
rect 533982 14968 533988 15020
rect 534040 15008 534046 15020
rect 545298 15008 545304 15020
rect 534040 14980 545304 15008
rect 534040 14968 534046 14980
rect 545298 14968 545304 14980
rect 545356 14968 545362 15020
rect 325602 14900 325608 14952
rect 325660 14940 325666 14952
rect 478138 14940 478144 14952
rect 325660 14912 478144 14940
rect 325660 14900 325666 14912
rect 478138 14900 478144 14912
rect 478196 14900 478202 14952
rect 487062 14900 487068 14952
rect 487120 14940 487126 14952
rect 529934 14940 529940 14952
rect 487120 14912 529940 14940
rect 487120 14900 487126 14912
rect 529934 14900 529940 14912
rect 529992 14900 529998 14952
rect 531222 14900 531228 14952
rect 531280 14940 531286 14952
rect 544470 14940 544476 14952
rect 531280 14912 544476 14940
rect 531280 14900 531286 14912
rect 544470 14900 544476 14912
rect 544528 14900 544534 14952
rect 555234 14900 555240 14952
rect 555292 14940 555298 14952
rect 563054 14940 563060 14952
rect 555292 14912 563060 14940
rect 555292 14900 555298 14912
rect 563054 14900 563060 14912
rect 563112 14900 563118 14952
rect 318702 14832 318708 14884
rect 318760 14872 318766 14884
rect 475838 14872 475844 14884
rect 318760 14844 475844 14872
rect 318760 14832 318766 14844
rect 475838 14832 475844 14844
rect 475896 14832 475902 14884
rect 482922 14832 482928 14884
rect 482980 14872 482986 14884
rect 528738 14872 528744 14884
rect 482980 14844 528744 14872
rect 482980 14832 482986 14844
rect 528738 14832 528744 14844
rect 528796 14832 528802 14884
rect 532602 14832 532608 14884
rect 532660 14872 532666 14884
rect 544838 14872 544844 14884
rect 532660 14844 544844 14872
rect 532660 14832 532666 14844
rect 544838 14832 544844 14844
rect 544896 14832 544902 14884
rect 311802 14764 311808 14816
rect 311860 14804 311866 14816
rect 473538 14804 473544 14816
rect 311860 14776 473544 14804
rect 311860 14764 311866 14776
rect 473538 14764 473544 14776
rect 473596 14764 473602 14816
rect 478782 14764 478788 14816
rect 478840 14804 478846 14816
rect 527266 14804 527272 14816
rect 478840 14776 527272 14804
rect 478840 14764 478846 14776
rect 527266 14764 527272 14776
rect 527324 14764 527330 14816
rect 529842 14764 529848 14816
rect 529900 14804 529906 14816
rect 543734 14804 543740 14816
rect 529900 14776 543740 14804
rect 529900 14764 529906 14776
rect 543734 14764 543740 14776
rect 543792 14764 543798 14816
rect 304994 14696 305000 14748
rect 305052 14736 305058 14748
rect 468938 14736 468944 14748
rect 305052 14708 468944 14736
rect 305052 14696 305058 14708
rect 468938 14696 468944 14708
rect 468996 14696 469002 14748
rect 476022 14696 476028 14748
rect 476080 14736 476086 14748
rect 526438 14736 526444 14748
rect 476080 14708 526444 14736
rect 476080 14696 476086 14708
rect 526438 14696 526444 14708
rect 526496 14696 526502 14748
rect 526622 14696 526628 14748
rect 526680 14736 526686 14748
rect 542538 14736 542544 14748
rect 526680 14708 542544 14736
rect 526680 14696 526686 14708
rect 542538 14696 542544 14708
rect 542596 14696 542602 14748
rect 302234 14628 302240 14680
rect 302292 14668 302298 14680
rect 466638 14668 466644 14680
rect 302292 14640 466644 14668
rect 302292 14628 302298 14640
rect 466638 14628 466644 14640
rect 466696 14628 466702 14680
rect 469030 14628 469036 14680
rect 469088 14668 469094 14680
rect 469088 14640 519492 14668
rect 469088 14628 469094 14640
rect 214558 14560 214564 14612
rect 214616 14600 214622 14612
rect 424134 14600 424140 14612
rect 214616 14572 424140 14600
rect 214616 14560 214622 14572
rect 424134 14560 424140 14572
rect 424192 14560 424198 14612
rect 447778 14560 447784 14612
rect 447836 14600 447842 14612
rect 517238 14600 517244 14612
rect 447836 14572 517244 14600
rect 447836 14560 447842 14572
rect 517238 14560 517244 14572
rect 517296 14560 517302 14612
rect 519464 14600 519492 14640
rect 523678 14628 523684 14680
rect 523736 14668 523742 14680
rect 540238 14668 540244 14680
rect 523736 14640 540244 14668
rect 523736 14628 523742 14640
rect 540238 14628 540244 14640
rect 540296 14628 540302 14680
rect 524138 14600 524144 14612
rect 519464 14572 524144 14600
rect 524138 14560 524144 14572
rect 524196 14560 524202 14612
rect 524322 14560 524328 14612
rect 524380 14600 524386 14612
rect 542170 14600 542176 14612
rect 524380 14572 542176 14600
rect 524380 14560 524386 14572
rect 542170 14560 542176 14572
rect 542228 14560 542234 14612
rect 204898 14492 204904 14544
rect 204956 14532 204962 14544
rect 422938 14532 422944 14544
rect 204956 14504 422944 14532
rect 204956 14492 204962 14504
rect 422938 14492 422944 14504
rect 422996 14492 423002 14544
rect 443822 14492 443828 14544
rect 443880 14532 443886 14544
rect 514938 14532 514944 14544
rect 443880 14504 514944 14532
rect 443880 14492 443886 14504
rect 514938 14492 514944 14504
rect 514996 14492 515002 14544
rect 521562 14492 521568 14544
rect 521620 14532 521626 14544
rect 541066 14532 541072 14544
rect 521620 14504 541072 14532
rect 521620 14492 521626 14504
rect 541066 14492 541072 14504
rect 541124 14492 541130 14544
rect 546310 14492 546316 14544
rect 546368 14532 546374 14544
rect 549070 14532 549076 14544
rect 546368 14504 549076 14532
rect 546368 14492 546374 14504
rect 549070 14492 549076 14504
rect 549128 14492 549134 14544
rect 554866 14492 554872 14544
rect 554924 14532 554930 14544
rect 563146 14532 563152 14544
rect 554924 14504 563152 14532
rect 554924 14492 554930 14504
rect 563146 14492 563152 14504
rect 563204 14492 563210 14544
rect 13722 14424 13728 14476
rect 13780 14464 13786 14476
rect 128538 14464 128544 14476
rect 13780 14436 128544 14464
rect 13780 14424 13786 14436
rect 128538 14424 128544 14436
rect 128596 14424 128602 14476
rect 174170 14424 174176 14476
rect 174228 14464 174234 14476
rect 421834 14464 421840 14476
rect 174228 14436 421840 14464
rect 174228 14424 174234 14436
rect 421834 14424 421840 14436
rect 421892 14424 421898 14476
rect 428921 14467 428979 14473
rect 428921 14433 428933 14467
rect 428967 14464 428979 14467
rect 511534 14464 511540 14476
rect 428967 14436 511540 14464
rect 428967 14433 428979 14436
rect 428921 14427 428979 14433
rect 511534 14424 511540 14436
rect 511592 14424 511598 14476
rect 513558 14424 513564 14476
rect 513616 14464 513622 14476
rect 514018 14464 514024 14476
rect 513616 14436 514024 14464
rect 513616 14424 513622 14436
rect 514018 14424 514024 14436
rect 514076 14424 514082 14476
rect 517422 14424 517428 14476
rect 517480 14464 517486 14476
rect 539870 14464 539876 14476
rect 517480 14436 539876 14464
rect 517480 14424 517486 14436
rect 539870 14424 539876 14436
rect 539928 14424 539934 14476
rect 547782 14424 547788 14476
rect 547840 14464 547846 14476
rect 549898 14464 549904 14476
rect 547840 14436 549904 14464
rect 547840 14424 547846 14436
rect 549898 14424 549904 14436
rect 549956 14424 549962 14476
rect 361482 14356 361488 14408
rect 361540 14396 361546 14408
rect 489638 14396 489644 14408
rect 361540 14368 489644 14396
rect 361540 14356 361546 14368
rect 489638 14356 489644 14368
rect 489696 14356 489702 14408
rect 502518 14356 502524 14408
rect 502576 14396 502582 14408
rect 503162 14396 503168 14408
rect 502576 14368 503168 14396
rect 502576 14356 502582 14368
rect 503162 14356 503168 14368
rect 503220 14356 503226 14408
rect 507762 14356 507768 14408
rect 507820 14396 507826 14408
rect 536834 14396 536840 14408
rect 507820 14368 536840 14396
rect 507820 14356 507826 14368
rect 536834 14356 536840 14368
rect 536892 14356 536898 14408
rect 544378 14356 544384 14408
rect 544436 14396 544442 14408
rect 546402 14396 546408 14408
rect 544436 14368 546408 14396
rect 544436 14356 544442 14368
rect 546402 14356 546408 14368
rect 546460 14356 546466 14408
rect 547690 14356 547696 14408
rect 547748 14396 547754 14408
rect 549438 14396 549444 14408
rect 547748 14368 549444 14396
rect 547748 14356 547754 14368
rect 549438 14356 549444 14368
rect 549496 14356 549502 14408
rect 551370 14356 551376 14408
rect 551428 14396 551434 14408
rect 551922 14396 551928 14408
rect 551428 14368 551928 14396
rect 551428 14356 551434 14368
rect 551922 14356 551928 14368
rect 551980 14356 551986 14408
rect 368382 14288 368388 14340
rect 368440 14328 368446 14340
rect 491938 14328 491944 14340
rect 368440 14300 491944 14328
rect 368440 14288 368446 14300
rect 491938 14288 491944 14300
rect 491996 14288 492002 14340
rect 514018 14288 514024 14340
rect 514076 14328 514082 14340
rect 521838 14328 521844 14340
rect 514076 14300 521844 14328
rect 514076 14288 514082 14300
rect 521838 14288 521844 14300
rect 521896 14288 521902 14340
rect 522298 14288 522304 14340
rect 522356 14328 522362 14340
rect 539134 14328 539140 14340
rect 522356 14300 539140 14328
rect 522356 14288 522362 14300
rect 539134 14288 539140 14300
rect 539192 14288 539198 14340
rect 545669 14331 545727 14337
rect 545669 14297 545681 14331
rect 545715 14328 545727 14331
rect 548334 14328 548340 14340
rect 545715 14300 548340 14328
rect 545715 14297 545727 14300
rect 545669 14291 545727 14297
rect 548334 14288 548340 14300
rect 548392 14288 548398 14340
rect 375190 14220 375196 14272
rect 375248 14260 375254 14272
rect 494238 14260 494244 14272
rect 375248 14232 494244 14260
rect 375248 14220 375254 14232
rect 494238 14220 494244 14232
rect 494296 14220 494302 14272
rect 520918 14220 520924 14272
rect 520976 14260 520982 14272
rect 537938 14260 537944 14272
rect 520976 14232 537944 14260
rect 520976 14220 520982 14232
rect 537938 14220 537944 14232
rect 537996 14220 538002 14272
rect 546034 14260 546040 14272
rect 542188 14232 546040 14260
rect 383562 14152 383568 14204
rect 383620 14192 383626 14204
rect 496538 14192 496544 14204
rect 383620 14164 496544 14192
rect 383620 14152 383626 14164
rect 496538 14152 496544 14164
rect 496596 14152 496602 14204
rect 525150 14152 525156 14204
rect 525208 14192 525214 14204
rect 541434 14192 541440 14204
rect 525208 14164 541440 14192
rect 525208 14152 525214 14164
rect 541434 14152 541440 14164
rect 541492 14152 541498 14204
rect 390462 14084 390468 14136
rect 390520 14124 390526 14136
rect 498838 14124 498844 14136
rect 390520 14096 498844 14124
rect 390520 14084 390526 14096
rect 498838 14084 498844 14096
rect 498896 14084 498902 14136
rect 519722 14084 519728 14136
rect 519780 14124 519786 14136
rect 534534 14124 534540 14136
rect 519780 14096 534540 14124
rect 519780 14084 519786 14096
rect 534534 14084 534540 14096
rect 534592 14084 534598 14136
rect 536742 14084 536748 14136
rect 536800 14124 536806 14136
rect 542188 14124 542216 14232
rect 546034 14220 546040 14232
rect 546092 14220 546098 14272
rect 553670 14220 553676 14272
rect 553728 14260 553734 14272
rect 556982 14260 556988 14272
rect 553728 14232 556988 14260
rect 553728 14220 553734 14232
rect 556982 14220 556988 14232
rect 557040 14220 557046 14272
rect 543642 14152 543648 14204
rect 543700 14192 543706 14204
rect 545669 14195 545727 14201
rect 545669 14192 545681 14195
rect 543700 14164 545681 14192
rect 543700 14152 543706 14164
rect 545669 14161 545681 14164
rect 545715 14161 545727 14195
rect 545669 14155 545727 14161
rect 545758 14152 545764 14204
rect 545816 14192 545822 14204
rect 547138 14192 547144 14204
rect 545816 14164 547144 14192
rect 545816 14152 545822 14164
rect 547138 14152 547144 14164
rect 547196 14152 547202 14204
rect 554038 14152 554044 14204
rect 554096 14192 554102 14204
rect 556890 14192 556896 14204
rect 554096 14164 556896 14192
rect 554096 14152 554102 14164
rect 556890 14152 556896 14164
rect 556948 14152 556954 14204
rect 536800 14096 542216 14124
rect 536800 14084 536806 14096
rect 552566 14084 552572 14136
rect 552624 14124 552630 14136
rect 555234 14124 555240 14136
rect 552624 14096 555240 14124
rect 552624 14084 552630 14096
rect 555234 14084 555240 14096
rect 555292 14084 555298 14136
rect 313274 14016 313280 14068
rect 313332 14056 313338 14068
rect 420638 14056 420644 14068
rect 313332 14028 420644 14056
rect 313332 14016 313338 14028
rect 420638 14016 420644 14028
rect 420696 14016 420702 14068
rect 420822 14016 420828 14068
rect 420880 14056 420886 14068
rect 508038 14056 508044 14068
rect 420880 14028 508044 14056
rect 420880 14016 420886 14028
rect 508038 14016 508044 14028
rect 508096 14016 508102 14068
rect 528462 14016 528468 14068
rect 528520 14056 528526 14068
rect 543366 14056 543372 14068
rect 528520 14028 543372 14056
rect 528520 14016 528526 14028
rect 543366 14016 543372 14028
rect 543424 14016 543430 14068
rect 545022 14016 545028 14068
rect 545080 14056 545086 14068
rect 548702 14056 548708 14068
rect 545080 14028 548708 14056
rect 545080 14016 545086 14028
rect 548702 14016 548708 14028
rect 548760 14016 548766 14068
rect 552934 14016 552940 14068
rect 552992 14056 552998 14068
rect 555418 14056 555424 14068
rect 552992 14028 555424 14056
rect 552992 14016 552998 14028
rect 555418 14016 555424 14028
rect 555476 14016 555482 14068
rect 397362 13948 397368 14000
rect 397420 13988 397426 14000
rect 501138 13988 501144 14000
rect 397420 13960 501144 13988
rect 397420 13948 397426 13960
rect 501138 13948 501144 13960
rect 501196 13948 501202 14000
rect 509878 13948 509884 14000
rect 509936 13988 509942 14000
rect 512638 13988 512644 14000
rect 509936 13960 512644 13988
rect 509936 13948 509942 13960
rect 512638 13948 512644 13960
rect 512696 13948 512702 14000
rect 518342 13948 518348 14000
rect 518400 13988 518406 14000
rect 532234 13988 532240 14000
rect 518400 13960 532240 13988
rect 518400 13948 518406 13960
rect 532234 13948 532240 13960
rect 532292 13948 532298 14000
rect 553302 13948 553308 14000
rect 553360 13988 553366 14000
rect 555510 13988 555516 14000
rect 553360 13960 555516 13988
rect 553360 13948 553366 13960
rect 555510 13948 555516 13960
rect 555568 13948 555574 14000
rect 408402 13880 408408 13932
rect 408460 13920 408466 13932
rect 504634 13920 504640 13932
rect 408460 13892 504640 13920
rect 408460 13880 408466 13892
rect 504634 13880 504640 13892
rect 504692 13880 504698 13932
rect 511258 13880 511264 13932
rect 511316 13920 511322 13932
rect 513834 13920 513840 13932
rect 511316 13892 513840 13920
rect 511316 13880 511322 13892
rect 513834 13880 513840 13892
rect 513892 13880 513898 13932
rect 555602 13880 555608 13932
rect 555660 13920 555666 13932
rect 555970 13920 555976 13932
rect 555660 13892 555976 13920
rect 555660 13880 555666 13892
rect 555970 13880 555976 13892
rect 556028 13880 556034 13932
rect 556338 13880 556344 13932
rect 556396 13920 556402 13932
rect 557350 13920 557356 13932
rect 556396 13892 557356 13920
rect 556396 13880 556402 13892
rect 557350 13880 557356 13892
rect 557408 13880 557414 13932
rect 557534 13880 557540 13932
rect 557592 13920 557598 13932
rect 558822 13920 558828 13932
rect 557592 13892 558828 13920
rect 557592 13880 557598 13892
rect 558822 13880 558828 13892
rect 558880 13880 558886 13932
rect 559098 13880 559104 13932
rect 559156 13920 559162 13932
rect 560110 13920 560116 13932
rect 559156 13892 560116 13920
rect 559156 13880 559162 13892
rect 560110 13880 560116 13892
rect 560168 13880 560174 13932
rect 330294 13812 330300 13864
rect 330352 13852 330358 13864
rect 425238 13852 425244 13864
rect 330352 13824 425244 13852
rect 330352 13812 330358 13824
rect 425238 13812 425244 13824
rect 425296 13812 425302 13864
rect 425422 13812 425428 13864
rect 425480 13852 425486 13864
rect 425480 13824 432000 13852
rect 425480 13812 425486 13824
rect 268378 13744 268384 13796
rect 268436 13784 268442 13796
rect 287057 13787 287115 13793
rect 287057 13784 287069 13787
rect 268436 13756 287069 13784
rect 268436 13744 268442 13756
rect 287057 13753 287069 13756
rect 287103 13753 287115 13787
rect 287057 13747 287115 13753
rect 296625 13787 296683 13793
rect 296625 13753 296637 13787
rect 296671 13784 296683 13787
rect 306377 13787 306435 13793
rect 306377 13784 306389 13787
rect 296671 13756 306389 13784
rect 296671 13753 296683 13756
rect 296625 13747 296683 13753
rect 306377 13753 306389 13756
rect 306423 13753 306435 13787
rect 306377 13747 306435 13753
rect 315945 13787 316003 13793
rect 315945 13753 315957 13787
rect 315991 13784 316003 13787
rect 325697 13787 325755 13793
rect 325697 13784 325709 13787
rect 315991 13756 325709 13784
rect 315991 13753 316003 13756
rect 315945 13747 316003 13753
rect 325697 13753 325709 13756
rect 325743 13753 325755 13787
rect 325697 13747 325755 13753
rect 335265 13787 335323 13793
rect 335265 13753 335277 13787
rect 335311 13784 335323 13787
rect 384209 13787 384267 13793
rect 384209 13784 384221 13787
rect 335311 13756 384221 13784
rect 335311 13753 335323 13756
rect 335265 13747 335323 13753
rect 384209 13753 384221 13756
rect 384255 13753 384267 13787
rect 384209 13747 384267 13753
rect 393225 13787 393283 13793
rect 393225 13753 393237 13787
rect 393271 13784 393283 13787
rect 402977 13787 403035 13793
rect 402977 13784 402989 13787
rect 393271 13756 402989 13784
rect 393271 13753 393283 13756
rect 393225 13747 393283 13753
rect 402977 13753 402989 13756
rect 403023 13753 403035 13787
rect 402977 13747 403035 13753
rect 403069 13787 403127 13793
rect 403069 13753 403081 13787
rect 403115 13784 403127 13787
rect 412453 13787 412511 13793
rect 412453 13784 412465 13787
rect 403115 13756 412465 13784
rect 403115 13753 403127 13756
rect 403069 13747 403127 13753
rect 412453 13753 412465 13756
rect 412499 13753 412511 13787
rect 412453 13747 412511 13753
rect 412545 13787 412603 13793
rect 412545 13753 412557 13787
rect 412591 13784 412603 13787
rect 422294 13784 422300 13796
rect 412591 13756 422300 13784
rect 412591 13753 412603 13756
rect 412545 13747 412603 13753
rect 422294 13744 422300 13756
rect 422352 13744 422358 13796
rect 431972 13793 432000 13824
rect 457438 13812 457444 13864
rect 457496 13852 457502 13864
rect 519538 13852 519544 13864
rect 457496 13824 519544 13852
rect 457496 13812 457502 13824
rect 519538 13812 519544 13824
rect 519596 13812 519602 13864
rect 551738 13812 551744 13864
rect 551796 13852 551802 13864
rect 553394 13852 553400 13864
rect 551796 13824 553400 13852
rect 551796 13812 551802 13824
rect 553394 13812 553400 13824
rect 553452 13812 553458 13864
rect 554498 13812 554504 13864
rect 554556 13852 554562 13864
rect 556706 13852 556712 13864
rect 554556 13824 556712 13852
rect 554556 13812 554562 13824
rect 556706 13812 556712 13824
rect 556764 13812 556770 13864
rect 556798 13812 556804 13864
rect 556856 13852 556862 13864
rect 557442 13852 557448 13864
rect 556856 13824 557448 13852
rect 556856 13812 556862 13824
rect 557442 13812 557448 13824
rect 557500 13812 557506 13864
rect 557902 13812 557908 13864
rect 557960 13852 557966 13864
rect 558638 13852 558644 13864
rect 557960 13824 558644 13852
rect 557960 13812 557966 13824
rect 558638 13812 558644 13824
rect 558696 13812 558702 13864
rect 559834 13812 559840 13864
rect 559892 13852 559898 13864
rect 560202 13852 560208 13864
rect 559892 13824 560208 13852
rect 559892 13812 559898 13824
rect 560202 13812 560208 13824
rect 560260 13812 560266 13864
rect 560570 13812 560576 13864
rect 560628 13852 560634 13864
rect 561490 13852 561496 13864
rect 560628 13824 561496 13852
rect 560628 13812 560634 13824
rect 561490 13812 561496 13824
rect 561548 13812 561554 13864
rect 422389 13787 422447 13793
rect 422389 13753 422401 13787
rect 422435 13784 422447 13787
rect 431773 13787 431831 13793
rect 431773 13784 431785 13787
rect 422435 13756 431785 13784
rect 422435 13753 422447 13756
rect 422389 13747 422447 13753
rect 431773 13753 431785 13756
rect 431819 13753 431831 13787
rect 431773 13747 431831 13753
rect 431957 13787 432015 13793
rect 431957 13753 431969 13787
rect 432003 13753 432015 13787
rect 431957 13747 432015 13753
rect 436189 13787 436247 13793
rect 436189 13753 436201 13787
rect 436235 13784 436247 13787
rect 463234 13784 463240 13796
rect 436235 13756 463240 13784
rect 436235 13753 436247 13756
rect 436189 13747 436247 13753
rect 463234 13744 463240 13756
rect 463292 13744 463298 13796
rect 261478 13676 261484 13728
rect 261536 13716 261542 13728
rect 366821 13719 366879 13725
rect 366821 13716 366833 13719
rect 261536 13688 366833 13716
rect 261536 13676 261542 13688
rect 366821 13685 366833 13688
rect 366867 13685 366879 13719
rect 366821 13679 366879 13685
rect 367005 13719 367063 13725
rect 367005 13685 367017 13719
rect 367051 13716 367063 13719
rect 433702 13716 433708 13728
rect 367051 13688 433708 13716
rect 367051 13685 367063 13688
rect 367005 13679 367063 13685
rect 433702 13676 433708 13688
rect 433760 13676 433766 13728
rect 433978 13676 433984 13728
rect 434036 13716 434042 13728
rect 470134 13716 470140 13728
rect 434036 13688 470140 13716
rect 434036 13676 434042 13688
rect 470134 13676 470140 13688
rect 470192 13676 470198 13728
rect 257338 13608 257344 13660
rect 257396 13648 257402 13660
rect 431402 13648 431408 13660
rect 257396 13620 431408 13648
rect 257396 13608 257402 13620
rect 431402 13608 431408 13620
rect 431460 13608 431466 13660
rect 431957 13651 432015 13657
rect 431957 13617 431969 13651
rect 432003 13648 432015 13651
rect 436002 13648 436008 13660
rect 432003 13620 436008 13648
rect 432003 13617 432015 13620
rect 431957 13611 432015 13617
rect 436002 13608 436008 13620
rect 436060 13608 436066 13660
rect 438854 13608 438860 13660
rect 438912 13648 438918 13660
rect 439314 13648 439320 13660
rect 438912 13620 439320 13648
rect 438912 13608 438918 13620
rect 439314 13608 439320 13620
rect 439372 13608 439378 13660
rect 474734 13648 474740 13660
rect 445496 13620 474740 13648
rect 211062 13540 211068 13592
rect 211120 13580 211126 13592
rect 441338 13580 441344 13592
rect 211120 13552 441344 13580
rect 211120 13540 211126 13552
rect 441338 13540 441344 13552
rect 441396 13540 441402 13592
rect 219250 13472 219256 13524
rect 219308 13512 219314 13524
rect 366545 13515 366603 13521
rect 366545 13512 366557 13515
rect 219308 13484 366557 13512
rect 219308 13472 219314 13484
rect 366545 13481 366557 13484
rect 366591 13481 366603 13515
rect 366545 13475 366603 13481
rect 366729 13515 366787 13521
rect 366729 13481 366741 13515
rect 366775 13512 366787 13515
rect 443638 13512 443644 13524
rect 366775 13484 443644 13512
rect 366775 13481 366787 13484
rect 366729 13475 366787 13481
rect 443638 13472 443644 13484
rect 443696 13472 443702 13524
rect 208302 13404 208308 13456
rect 208360 13444 208366 13456
rect 366637 13447 366695 13453
rect 366637 13444 366649 13447
rect 208360 13416 366649 13444
rect 208360 13404 208366 13416
rect 366637 13413 366649 13416
rect 366683 13413 366695 13447
rect 366637 13407 366695 13413
rect 366913 13447 366971 13453
rect 366913 13413 366925 13447
rect 366959 13444 366971 13447
rect 440234 13444 440240 13456
rect 366959 13416 440240 13444
rect 366959 13413 366971 13416
rect 366913 13407 366971 13413
rect 440234 13404 440240 13416
rect 440292 13404 440298 13456
rect 191742 13336 191748 13388
rect 191800 13376 191806 13388
rect 434898 13376 434904 13388
rect 191800 13348 434904 13376
rect 191800 13336 191806 13348
rect 434898 13336 434904 13348
rect 434956 13336 434962 13388
rect 435358 13336 435364 13388
rect 435416 13376 435422 13388
rect 445496 13376 445524 13620
rect 474734 13608 474740 13620
rect 474792 13608 474798 13660
rect 464246 13472 464252 13524
rect 464304 13512 464310 13524
rect 500034 13512 500040 13524
rect 464304 13484 500040 13512
rect 464304 13472 464310 13484
rect 500034 13472 500040 13484
rect 500092 13472 500098 13524
rect 445662 13404 445668 13456
rect 445720 13444 445726 13456
rect 451921 13447 451979 13453
rect 451921 13444 451933 13447
rect 445720 13416 451933 13444
rect 445720 13404 445726 13416
rect 451921 13413 451933 13416
rect 451967 13413 451979 13447
rect 451921 13407 451979 13413
rect 461578 13404 461584 13456
rect 461636 13444 461642 13456
rect 490834 13444 490840 13456
rect 461636 13416 490840 13444
rect 461636 13404 461642 13416
rect 490834 13404 490840 13416
rect 490892 13404 490898 13456
rect 491202 13404 491208 13456
rect 491260 13444 491266 13456
rect 531498 13444 531504 13456
rect 491260 13416 531504 13444
rect 491260 13404 491266 13416
rect 531498 13404 531504 13416
rect 531556 13404 531562 13456
rect 435416 13348 445524 13376
rect 435416 13336 435422 13348
rect 461026 13336 461032 13388
rect 461084 13376 461090 13388
rect 461670 13376 461676 13388
rect 461084 13348 461676 13376
rect 461084 13336 461090 13348
rect 461670 13336 461676 13348
rect 461728 13336 461734 13388
rect 467742 13336 467748 13388
rect 467800 13376 467806 13388
rect 523770 13376 523776 13388
rect 467800 13348 523776 13376
rect 467800 13336 467806 13348
rect 523770 13336 523776 13348
rect 523828 13336 523834 13388
rect 184845 13311 184903 13317
rect 184845 13277 184857 13311
rect 184891 13308 184903 13311
rect 366821 13311 366879 13317
rect 366821 13308 366833 13311
rect 184891 13280 366833 13308
rect 184891 13277 184903 13280
rect 184845 13271 184903 13277
rect 366821 13277 366833 13280
rect 366867 13277 366879 13311
rect 366821 13271 366879 13277
rect 366913 13311 366971 13317
rect 366913 13277 366925 13311
rect 366959 13308 366971 13311
rect 432598 13308 432604 13320
rect 366959 13280 432604 13308
rect 366959 13277 366971 13280
rect 366913 13271 366971 13277
rect 432598 13268 432604 13280
rect 432656 13268 432662 13320
rect 439314 13268 439320 13320
rect 439372 13308 439378 13320
rect 506934 13308 506940 13320
rect 439372 13280 506940 13308
rect 439372 13268 439378 13280
rect 506934 13268 506940 13280
rect 506992 13268 506998 13320
rect 131022 13200 131028 13252
rect 131080 13240 131086 13252
rect 415302 13240 415308 13252
rect 131080 13212 415308 13240
rect 131080 13200 131086 13212
rect 415302 13200 415308 13212
rect 415360 13200 415366 13252
rect 419442 13200 419448 13252
rect 419500 13240 419506 13252
rect 508498 13240 508504 13252
rect 419500 13212 508504 13240
rect 419500 13200 419506 13212
rect 508498 13200 508504 13212
rect 508556 13200 508562 13252
rect 516042 13200 516048 13252
rect 516100 13240 516106 13252
rect 539502 13240 539508 13252
rect 516100 13212 539508 13240
rect 516100 13200 516106 13212
rect 539502 13200 539508 13212
rect 539560 13200 539566 13252
rect 46842 13132 46848 13184
rect 46900 13172 46906 13184
rect 152090 13172 152096 13184
rect 46900 13144 152096 13172
rect 46900 13132 46906 13144
rect 152090 13132 152096 13144
rect 152148 13132 152154 13184
rect 173802 13132 173808 13184
rect 173860 13172 173866 13184
rect 366545 13175 366603 13181
rect 366545 13172 366557 13175
rect 173860 13144 366557 13172
rect 173860 13132 173866 13144
rect 366545 13141 366557 13144
rect 366591 13141 366603 13175
rect 366545 13135 366603 13141
rect 366821 13175 366879 13181
rect 366821 13141 366833 13175
rect 366867 13172 366879 13175
rect 429102 13172 429108 13184
rect 366867 13144 429108 13172
rect 366867 13141 366879 13144
rect 366821 13135 366879 13141
rect 429102 13132 429108 13144
rect 429160 13132 429166 13184
rect 429194 13132 429200 13184
rect 429252 13172 429258 13184
rect 436189 13175 436247 13181
rect 436189 13172 436201 13175
rect 429252 13144 436201 13172
rect 429252 13132 429258 13144
rect 436189 13141 436201 13144
rect 436235 13141 436247 13175
rect 436189 13135 436247 13141
rect 437566 13132 437572 13184
rect 437624 13172 437630 13184
rect 437934 13172 437940 13184
rect 437624 13144 437940 13172
rect 437624 13132 437630 13144
rect 437934 13132 437940 13144
rect 437992 13132 437998 13184
rect 451921 13175 451979 13181
rect 451921 13141 451933 13175
rect 451967 13172 451979 13175
rect 516870 13172 516876 13184
rect 451967 13144 516876 13172
rect 451967 13141 451979 13144
rect 451921 13135 451979 13141
rect 516870 13132 516876 13144
rect 516928 13132 516934 13184
rect 126882 13064 126888 13116
rect 126940 13104 126946 13116
rect 366637 13107 366695 13113
rect 366637 13104 366649 13107
rect 126940 13076 366649 13104
rect 126940 13064 126946 13076
rect 366637 13073 366649 13076
rect 366683 13073 366695 13107
rect 366637 13067 366695 13073
rect 366913 13107 366971 13113
rect 366913 13073 366925 13107
rect 366959 13104 366971 13107
rect 414198 13104 414204 13116
rect 366959 13076 414204 13104
rect 366959 13073 366971 13076
rect 366913 13067 366971 13073
rect 414198 13064 414204 13076
rect 414256 13064 414262 13116
rect 416682 13064 416688 13116
rect 416740 13104 416746 13116
rect 507302 13104 507308 13116
rect 416740 13076 507308 13104
rect 416740 13064 416746 13076
rect 507302 13064 507308 13076
rect 507360 13064 507366 13116
rect 510522 13064 510528 13116
rect 510580 13104 510586 13116
rect 537570 13104 537576 13116
rect 510580 13076 537576 13104
rect 510580 13064 510586 13076
rect 537570 13064 537576 13076
rect 537628 13064 537634 13116
rect 287057 13039 287115 13045
rect 287057 13005 287069 13039
rect 287103 13036 287115 13039
rect 296625 13039 296683 13045
rect 296625 13036 296637 13039
rect 287103 13008 296637 13036
rect 287103 13005 287115 13008
rect 287057 12999 287115 13005
rect 296625 13005 296637 13008
rect 296671 13005 296683 13039
rect 296625 12999 296683 13005
rect 304258 12996 304264 13048
rect 304316 13036 304322 13048
rect 454034 13036 454040 13048
rect 304316 13008 454040 13036
rect 304316 12996 304322 13008
rect 454034 12996 454040 13008
rect 454092 12996 454098 13048
rect 456797 13039 456855 13045
rect 456797 13005 456809 13039
rect 456843 13036 456855 13039
rect 461489 13039 461547 13045
rect 461489 13036 461501 13039
rect 456843 13008 461501 13036
rect 456843 13005 456855 13008
rect 456797 12999 456855 13005
rect 461489 13005 461501 13008
rect 461535 13005 461547 13039
rect 461489 12999 461547 13005
rect 461765 13039 461823 13045
rect 461765 13005 461777 13039
rect 461811 13036 461823 13039
rect 475381 13039 475439 13045
rect 475381 13036 475393 13039
rect 461811 13008 475393 13036
rect 461811 13005 461823 13008
rect 461765 12999 461823 13005
rect 475381 13005 475393 13008
rect 475427 13005 475439 13039
rect 475381 12999 475439 13005
rect 306377 12971 306435 12977
rect 306377 12937 306389 12971
rect 306423 12968 306435 12971
rect 315945 12971 316003 12977
rect 315945 12968 315957 12971
rect 306423 12940 315957 12968
rect 306423 12937 306435 12940
rect 306377 12931 306435 12937
rect 315945 12937 315957 12940
rect 315991 12937 316003 12971
rect 315945 12931 316003 12937
rect 325697 12971 325755 12977
rect 325697 12937 325709 12971
rect 325743 12968 325755 12971
rect 335265 12971 335323 12977
rect 335265 12968 335277 12971
rect 325743 12940 335277 12968
rect 325743 12937 325755 12940
rect 325697 12931 325755 12937
rect 335265 12937 335277 12940
rect 335311 12937 335323 12971
rect 335265 12931 335323 12937
rect 349062 12928 349068 12980
rect 349120 12968 349126 12980
rect 485498 12968 485504 12980
rect 349120 12940 485504 12968
rect 349120 12928 349126 12940
rect 485498 12928 485504 12940
rect 485556 12928 485562 12980
rect 351822 12860 351828 12912
rect 351880 12900 351886 12912
rect 366913 12903 366971 12909
rect 366913 12900 366925 12903
rect 351880 12872 366925 12900
rect 351880 12860 351886 12872
rect 366913 12869 366925 12872
rect 366959 12869 366971 12903
rect 366913 12863 366971 12869
rect 367005 12903 367063 12909
rect 367005 12869 367017 12903
rect 367051 12900 367063 12903
rect 382369 12903 382427 12909
rect 382369 12900 382381 12903
rect 367051 12872 382381 12900
rect 367051 12869 367063 12872
rect 367005 12863 367063 12869
rect 382369 12869 382381 12872
rect 382415 12869 382427 12903
rect 382369 12863 382427 12869
rect 393222 12860 393228 12912
rect 393280 12900 393286 12912
rect 402974 12900 402980 12912
rect 393280 12872 402980 12900
rect 393280 12860 393286 12872
rect 402974 12860 402980 12872
rect 403032 12860 403038 12912
rect 412542 12860 412548 12912
rect 412600 12900 412606 12912
rect 422294 12900 422300 12912
rect 412600 12872 422300 12900
rect 412600 12860 412606 12872
rect 422294 12860 422300 12872
rect 422352 12860 422358 12912
rect 431862 12860 431868 12912
rect 431920 12900 431926 12912
rect 461673 12903 461731 12909
rect 431920 12872 461624 12900
rect 431920 12860 431926 12872
rect 393133 12835 393191 12841
rect 393133 12801 393145 12835
rect 393179 12832 393191 12835
rect 403069 12835 403127 12841
rect 403069 12832 403081 12835
rect 393179 12804 403081 12832
rect 393179 12801 393191 12804
rect 393133 12795 393191 12801
rect 403069 12801 403081 12804
rect 403115 12801 403127 12835
rect 403069 12795 403127 12801
rect 412453 12835 412511 12841
rect 412453 12801 412465 12835
rect 412499 12832 412511 12835
rect 422389 12835 422447 12841
rect 422389 12832 422401 12835
rect 412499 12804 422401 12832
rect 412499 12801 412511 12804
rect 412453 12795 412511 12801
rect 422389 12801 422401 12804
rect 422435 12801 422447 12835
rect 422389 12795 422447 12801
rect 431773 12835 431831 12841
rect 431773 12801 431785 12835
rect 431819 12832 431831 12835
rect 456797 12835 456855 12841
rect 456797 12832 456809 12835
rect 431819 12804 456809 12832
rect 431819 12801 431831 12804
rect 431773 12795 431831 12801
rect 456797 12801 456809 12804
rect 456843 12801 456855 12835
rect 461596 12832 461624 12872
rect 461673 12869 461685 12903
rect 461719 12900 461731 12903
rect 475381 12903 475439 12909
rect 461719 12872 470548 12900
rect 461719 12869 461731 12872
rect 461673 12863 461731 12869
rect 461765 12835 461823 12841
rect 461765 12832 461777 12835
rect 461596 12804 461777 12832
rect 456797 12795 456855 12801
rect 461765 12801 461777 12804
rect 461811 12801 461823 12835
rect 470520 12832 470548 12872
rect 475381 12869 475393 12903
rect 475427 12900 475439 12903
rect 486602 12900 486608 12912
rect 475427 12872 486608 12900
rect 475427 12869 475439 12872
rect 475381 12863 475439 12869
rect 486602 12860 486608 12872
rect 486660 12860 486666 12912
rect 488902 12832 488908 12844
rect 470520 12804 488908 12832
rect 461765 12795 461823 12801
rect 488902 12792 488908 12804
rect 488960 12792 488966 12844
rect 367005 12767 367063 12773
rect 367005 12764 367017 12767
rect 360396 12736 367017 12764
rect 358722 12656 358728 12708
rect 358780 12696 358786 12708
rect 360396 12696 360424 12736
rect 367005 12733 367017 12736
rect 367051 12733 367063 12767
rect 367005 12727 367063 12733
rect 375285 12767 375343 12773
rect 375285 12733 375297 12767
rect 375331 12764 375343 12767
rect 379517 12767 379575 12773
rect 379517 12764 379529 12767
rect 375331 12736 379529 12764
rect 375331 12733 375343 12736
rect 375285 12727 375343 12733
rect 379517 12733 379529 12736
rect 379563 12733 379575 12767
rect 379517 12727 379575 12733
rect 387702 12724 387708 12776
rect 387760 12764 387766 12776
rect 498102 12764 498108 12776
rect 387760 12736 498108 12764
rect 387760 12724 387766 12736
rect 498102 12724 498108 12736
rect 498160 12724 498166 12776
rect 358780 12668 360424 12696
rect 358780 12656 358786 12668
rect 364978 12656 364984 12708
rect 365036 12696 365042 12708
rect 464338 12696 464344 12708
rect 365036 12668 464344 12696
rect 365036 12656 365042 12668
rect 464338 12656 464344 12668
rect 464396 12656 464402 12708
rect 384209 12631 384267 12637
rect 384209 12597 384221 12631
rect 384255 12628 384267 12631
rect 393225 12631 393283 12637
rect 393225 12628 393237 12631
rect 384255 12600 393237 12628
rect 384255 12597 384267 12600
rect 384209 12591 384267 12597
rect 393225 12597 393237 12600
rect 393271 12597 393283 12631
rect 393225 12591 393283 12597
rect 409782 12588 409788 12640
rect 409840 12628 409846 12640
rect 505002 12628 505008 12640
rect 409840 12600 505008 12628
rect 409840 12588 409846 12600
rect 505002 12588 505008 12600
rect 505060 12588 505066 12640
rect 367005 12563 367063 12569
rect 367005 12529 367017 12563
rect 367051 12560 367063 12563
rect 375285 12563 375343 12569
rect 375285 12560 375297 12563
rect 367051 12532 375297 12560
rect 367051 12529 367063 12532
rect 367005 12523 367063 12529
rect 375285 12529 375297 12532
rect 375331 12529 375343 12563
rect 375285 12523 375343 12529
rect 379517 12563 379575 12569
rect 379517 12529 379529 12563
rect 379563 12560 379575 12563
rect 393133 12563 393191 12569
rect 393133 12560 393145 12563
rect 379563 12532 393145 12560
rect 379563 12529 379575 12532
rect 379517 12523 379575 12529
rect 393133 12529 393145 12532
rect 393179 12529 393191 12563
rect 393133 12523 393191 12529
rect 402977 12563 403035 12569
rect 402977 12529 402989 12563
rect 403023 12560 403035 12563
rect 412545 12563 412603 12569
rect 412545 12560 412557 12563
rect 403023 12532 412557 12560
rect 403023 12529 403035 12532
rect 402977 12523 403035 12529
rect 412545 12529 412557 12532
rect 412591 12529 412603 12563
rect 412545 12523 412603 12529
rect 423582 12520 423588 12572
rect 423640 12560 423646 12572
rect 509602 12560 509608 12572
rect 423640 12532 509608 12560
rect 423640 12520 423646 12532
rect 509602 12520 509608 12532
rect 509660 12520 509666 12572
rect 528830 12520 528836 12572
rect 528888 12560 528894 12572
rect 529290 12560 529296 12572
rect 528888 12532 529296 12560
rect 528888 12520 528894 12532
rect 529290 12520 529296 12532
rect 529348 12520 529354 12572
rect 67177 12495 67235 12501
rect 67177 12461 67189 12495
rect 67223 12492 67235 12495
rect 67542 12492 67548 12504
rect 67223 12464 67548 12492
rect 67223 12461 67235 12464
rect 67177 12455 67235 12461
rect 67542 12452 67548 12464
rect 67600 12452 67606 12504
rect 179417 12495 179475 12501
rect 179417 12461 179429 12495
rect 179463 12492 179475 12495
rect 179506 12492 179512 12504
rect 179463 12464 179512 12492
rect 179463 12461 179475 12464
rect 179417 12455 179475 12461
rect 179506 12452 179512 12464
rect 179564 12452 179570 12504
rect 382369 12495 382427 12501
rect 382369 12461 382381 12495
rect 382415 12492 382427 12495
rect 393222 12492 393228 12504
rect 382415 12464 393228 12492
rect 382415 12461 382427 12464
rect 382369 12455 382427 12461
rect 393222 12452 393228 12464
rect 393280 12452 393286 12504
rect 403066 12452 403072 12504
rect 403124 12492 403130 12504
rect 410426 12492 410432 12504
rect 403124 12464 410432 12492
rect 403124 12452 403130 12464
rect 410426 12452 410432 12464
rect 410484 12452 410490 12504
rect 410518 12452 410524 12504
rect 410576 12492 410582 12504
rect 460934 12492 460940 12504
rect 410576 12464 460940 12492
rect 410576 12452 410582 12464
rect 460934 12452 460940 12464
rect 460992 12452 460998 12504
rect 121638 12424 121644 12436
rect 121599 12396 121644 12424
rect 121638 12384 121644 12396
rect 121696 12384 121702 12436
rect 208673 12427 208731 12433
rect 208673 12393 208685 12427
rect 208719 12424 208731 12427
rect 219345 12427 219403 12433
rect 219345 12424 219357 12427
rect 208719 12396 219357 12424
rect 208719 12393 208731 12396
rect 208673 12387 208731 12393
rect 219345 12393 219357 12396
rect 219391 12393 219403 12427
rect 219345 12387 219403 12393
rect 229189 12427 229247 12433
rect 229189 12393 229201 12427
rect 229235 12424 229247 12427
rect 238573 12427 238631 12433
rect 238573 12424 238585 12427
rect 229235 12396 238585 12424
rect 229235 12393 229247 12396
rect 229189 12387 229247 12393
rect 238573 12393 238585 12396
rect 238619 12393 238631 12427
rect 238573 12387 238631 12393
rect 248509 12427 248567 12433
rect 248509 12393 248521 12427
rect 248555 12424 248567 12427
rect 257893 12427 257951 12433
rect 257893 12424 257905 12427
rect 248555 12396 257905 12424
rect 248555 12393 248567 12396
rect 248509 12387 248567 12393
rect 257893 12393 257905 12396
rect 257939 12393 257951 12427
rect 257893 12387 257951 12393
rect 275278 12384 275284 12436
rect 275336 12424 275342 12436
rect 445938 12424 445944 12436
rect 275336 12396 445944 12424
rect 275336 12384 275342 12396
rect 445938 12384 445944 12396
rect 445996 12384 446002 12436
rect 497090 12384 497096 12436
rect 497148 12424 497154 12436
rect 497734 12424 497740 12436
rect 497148 12396 497740 12424
rect 497148 12384 497154 12396
rect 497734 12384 497740 12396
rect 497792 12384 497798 12436
rect 555234 12384 555240 12436
rect 555292 12424 555298 12436
rect 555878 12424 555884 12436
rect 555292 12396 555884 12424
rect 555292 12384 555298 12396
rect 555878 12384 555884 12396
rect 555936 12384 555942 12436
rect 210421 12359 210479 12365
rect 210421 12325 210433 12359
rect 210467 12356 210479 12359
rect 219253 12359 219311 12365
rect 219253 12356 219265 12359
rect 210467 12328 219265 12356
rect 210467 12325 210479 12328
rect 210421 12319 210479 12325
rect 219253 12325 219265 12328
rect 219299 12325 219311 12359
rect 219253 12319 219311 12325
rect 225598 12316 225604 12368
rect 225656 12356 225662 12368
rect 427538 12356 427544 12368
rect 225656 12328 427544 12356
rect 225656 12316 225662 12328
rect 427538 12316 427544 12328
rect 427596 12316 427602 12368
rect 428918 12356 428924 12368
rect 428879 12328 428924 12356
rect 428918 12316 428924 12328
rect 428976 12316 428982 12368
rect 431678 12316 431684 12368
rect 431736 12356 431742 12368
rect 467834 12356 467840 12368
rect 431736 12328 467840 12356
rect 431736 12316 431742 12328
rect 467834 12316 467840 12328
rect 467892 12316 467898 12368
rect 196802 12248 196808 12300
rect 196860 12288 196866 12300
rect 436738 12288 436744 12300
rect 196860 12260 436744 12288
rect 196860 12248 196866 12260
rect 436738 12248 436744 12260
rect 436796 12248 436802 12300
rect 194502 12180 194508 12232
rect 194560 12220 194566 12232
rect 435634 12220 435640 12232
rect 194560 12192 435640 12220
rect 194560 12180 194566 12192
rect 435634 12180 435640 12192
rect 435692 12180 435698 12232
rect 190362 12112 190368 12164
rect 190420 12152 190426 12164
rect 208673 12155 208731 12161
rect 208673 12152 208685 12155
rect 190420 12124 208685 12152
rect 190420 12112 190426 12124
rect 208673 12121 208685 12124
rect 208719 12121 208731 12155
rect 208673 12115 208731 12121
rect 219345 12155 219403 12161
rect 219345 12121 219357 12155
rect 219391 12152 219403 12155
rect 229094 12152 229100 12164
rect 219391 12124 229100 12152
rect 219391 12121 219403 12124
rect 219345 12115 219403 12121
rect 229094 12112 229100 12124
rect 229152 12112 229158 12164
rect 238662 12112 238668 12164
rect 238720 12152 238726 12164
rect 248414 12152 248420 12164
rect 238720 12124 248420 12152
rect 238720 12112 238726 12124
rect 248414 12112 248420 12124
rect 248472 12112 248478 12164
rect 257982 12112 257988 12164
rect 258040 12152 258046 12164
rect 267734 12152 267740 12164
rect 258040 12124 267740 12152
rect 258040 12112 258046 12124
rect 267734 12112 267740 12124
rect 267792 12112 267798 12164
rect 277302 12112 277308 12164
rect 277360 12152 277366 12164
rect 287054 12152 287060 12164
rect 277360 12124 287060 12152
rect 277360 12112 277366 12124
rect 287054 12112 287060 12124
rect 287112 12112 287118 12164
rect 296625 12155 296683 12161
rect 296625 12121 296637 12155
rect 296671 12152 296683 12155
rect 306374 12152 306380 12164
rect 296671 12124 306380 12152
rect 296671 12121 296683 12124
rect 296625 12115 296683 12121
rect 306374 12112 306380 12124
rect 306432 12112 306438 12164
rect 315942 12112 315948 12164
rect 316000 12152 316006 12164
rect 325694 12152 325700 12164
rect 316000 12124 325700 12152
rect 316000 12112 316006 12124
rect 325694 12112 325700 12124
rect 325752 12112 325758 12164
rect 335262 12112 335268 12164
rect 335320 12152 335326 12164
rect 383657 12155 383715 12161
rect 383657 12152 383669 12155
rect 335320 12124 383669 12152
rect 335320 12112 335326 12124
rect 383657 12121 383669 12124
rect 383703 12121 383715 12155
rect 383657 12115 383715 12121
rect 393225 12155 393283 12161
rect 393225 12121 393237 12155
rect 393271 12152 393283 12155
rect 402977 12155 403035 12161
rect 402977 12152 402989 12155
rect 393271 12124 402989 12152
rect 393271 12121 393283 12124
rect 393225 12115 393283 12121
rect 402977 12121 402989 12124
rect 403023 12121 403035 12155
rect 402977 12115 403035 12121
rect 412545 12155 412603 12161
rect 412545 12121 412557 12155
rect 412591 12152 412603 12155
rect 419445 12155 419503 12161
rect 419445 12152 419457 12155
rect 412591 12124 419457 12152
rect 412591 12121 412603 12124
rect 412545 12115 412603 12121
rect 419445 12121 419457 12124
rect 419491 12121 419503 12155
rect 433334 12152 433340 12164
rect 419445 12115 419503 12121
rect 419552 12124 433340 12152
rect 186222 12044 186228 12096
rect 186280 12084 186286 12096
rect 210421 12087 210479 12093
rect 210421 12084 210433 12087
rect 186280 12056 210433 12084
rect 186280 12044 186286 12056
rect 210421 12053 210433 12056
rect 210467 12053 210479 12087
rect 210421 12047 210479 12053
rect 219253 12087 219311 12093
rect 219253 12053 219265 12087
rect 219299 12084 219311 12087
rect 229189 12087 229247 12093
rect 229189 12084 229201 12087
rect 219299 12056 229201 12084
rect 219299 12053 219311 12056
rect 219253 12047 219311 12053
rect 229189 12053 229201 12056
rect 229235 12053 229247 12087
rect 229189 12047 229247 12053
rect 238573 12087 238631 12093
rect 238573 12053 238585 12087
rect 238619 12084 238631 12087
rect 248509 12087 248567 12093
rect 248509 12084 248521 12087
rect 238619 12056 248521 12084
rect 238619 12053 238631 12056
rect 238573 12047 238631 12053
rect 248509 12053 248521 12056
rect 248555 12053 248567 12087
rect 248509 12047 248567 12053
rect 257893 12087 257951 12093
rect 257893 12053 257905 12087
rect 257939 12084 257951 12087
rect 267829 12087 267887 12093
rect 267829 12084 267841 12087
rect 257939 12056 267841 12084
rect 257939 12053 257951 12056
rect 257893 12047 257951 12053
rect 267829 12053 267841 12056
rect 267875 12053 267887 12087
rect 267829 12047 267887 12053
rect 277213 12087 277271 12093
rect 277213 12053 277225 12087
rect 277259 12084 277271 12087
rect 287149 12087 287207 12093
rect 287149 12084 287161 12087
rect 277259 12056 287161 12084
rect 277259 12053 277271 12056
rect 277213 12047 277271 12053
rect 287149 12053 287161 12056
rect 287195 12053 287207 12087
rect 287149 12047 287207 12053
rect 296533 12087 296591 12093
rect 296533 12053 296545 12087
rect 296579 12084 296591 12087
rect 306469 12087 306527 12093
rect 306469 12084 306481 12087
rect 296579 12056 306481 12084
rect 296579 12053 296591 12056
rect 296533 12047 296591 12053
rect 306469 12053 306481 12056
rect 306515 12053 306527 12087
rect 306469 12047 306527 12053
rect 315853 12087 315911 12093
rect 315853 12053 315865 12087
rect 315899 12084 315911 12087
rect 325789 12087 325847 12093
rect 325789 12084 325801 12087
rect 315899 12056 325801 12084
rect 315899 12053 315911 12056
rect 315853 12047 315911 12053
rect 325789 12053 325801 12056
rect 325835 12053 325847 12087
rect 325789 12047 325847 12053
rect 335173 12087 335231 12093
rect 335173 12053 335185 12087
rect 335219 12084 335231 12087
rect 383749 12087 383807 12093
rect 383749 12084 383761 12087
rect 335219 12056 383761 12084
rect 335219 12053 335231 12056
rect 335173 12047 335231 12053
rect 383749 12053 383761 12056
rect 383795 12053 383807 12087
rect 383749 12047 383807 12053
rect 393133 12087 393191 12093
rect 393133 12053 393145 12087
rect 393179 12084 393191 12087
rect 403069 12087 403127 12093
rect 403069 12084 403081 12087
rect 393179 12056 403081 12084
rect 393179 12053 393191 12056
rect 393133 12047 393191 12053
rect 403069 12053 403081 12056
rect 403115 12053 403127 12087
rect 403069 12047 403127 12053
rect 412453 12087 412511 12093
rect 412453 12053 412465 12087
rect 412499 12084 412511 12087
rect 419552 12084 419580 12124
rect 433334 12112 433340 12124
rect 433392 12112 433398 12164
rect 465534 12152 465540 12164
rect 460952 12124 465540 12152
rect 432138 12084 432144 12096
rect 412499 12056 419580 12084
rect 419644 12056 432144 12084
rect 412499 12053 412511 12056
rect 412453 12047 412511 12053
rect 182542 11976 182548 12028
rect 182600 12016 182606 12028
rect 210329 12019 210387 12025
rect 210329 12016 210341 12019
rect 182600 11988 210341 12016
rect 182600 11976 182606 11988
rect 210329 11985 210341 11988
rect 210375 11985 210387 12019
rect 210329 11979 210387 11985
rect 219345 12019 219403 12025
rect 219345 11985 219357 12019
rect 219391 12016 219403 12019
rect 229097 12019 229155 12025
rect 229097 12016 229109 12019
rect 219391 11988 229109 12016
rect 219391 11985 219403 11988
rect 219345 11979 219403 11985
rect 229097 11985 229109 11988
rect 229143 11985 229155 12019
rect 229097 11979 229155 11985
rect 238665 12019 238723 12025
rect 238665 11985 238677 12019
rect 238711 12016 238723 12019
rect 248417 12019 248475 12025
rect 248417 12016 248429 12019
rect 238711 11988 248429 12016
rect 238711 11985 238723 11988
rect 238665 11979 238723 11985
rect 248417 11985 248429 11988
rect 248463 11985 248475 12019
rect 248417 11979 248475 11985
rect 257985 12019 258043 12025
rect 257985 11985 257997 12019
rect 258031 12016 258043 12019
rect 267737 12019 267795 12025
rect 267737 12016 267749 12019
rect 258031 11988 267749 12016
rect 258031 11985 258043 11988
rect 257985 11979 258043 11985
rect 267737 11985 267749 11988
rect 267783 11985 267795 12019
rect 267737 11979 267795 11985
rect 277305 12019 277363 12025
rect 277305 11985 277317 12019
rect 277351 12016 277363 12019
rect 287057 12019 287115 12025
rect 287057 12016 287069 12019
rect 277351 11988 287069 12016
rect 277351 11985 277363 11988
rect 277305 11979 277363 11985
rect 287057 11985 287069 11988
rect 287103 11985 287115 12019
rect 287057 11979 287115 11985
rect 296625 12019 296683 12025
rect 296625 11985 296637 12019
rect 296671 12016 296683 12019
rect 306377 12019 306435 12025
rect 306377 12016 306389 12019
rect 296671 11988 306389 12016
rect 296671 11985 296683 11988
rect 296625 11979 296683 11985
rect 306377 11985 306389 11988
rect 306423 11985 306435 12019
rect 306377 11979 306435 11985
rect 315945 12019 316003 12025
rect 315945 11985 315957 12019
rect 315991 12016 316003 12019
rect 325697 12019 325755 12025
rect 325697 12016 325709 12019
rect 315991 11988 325709 12016
rect 315991 11985 316003 11988
rect 315945 11979 316003 11985
rect 325697 11985 325709 11988
rect 325743 11985 325755 12019
rect 325697 11979 325755 11985
rect 335265 12019 335323 12025
rect 335265 11985 335277 12019
rect 335311 12016 335323 12019
rect 383657 12019 383715 12025
rect 383657 12016 383669 12019
rect 335311 11988 383669 12016
rect 335311 11985 335323 11988
rect 335265 11979 335323 11985
rect 383657 11985 383669 11988
rect 383703 11985 383715 12019
rect 383657 11979 383715 11985
rect 383841 12019 383899 12025
rect 383841 11985 383853 12019
rect 383887 12016 383899 12019
rect 393041 12019 393099 12025
rect 393041 12016 393053 12019
rect 383887 11988 393053 12016
rect 383887 11985 383899 11988
rect 383841 11979 383899 11985
rect 393041 11985 393053 11988
rect 393087 11985 393099 12019
rect 393041 11979 393099 11985
rect 393225 12019 393283 12025
rect 393225 11985 393237 12019
rect 393271 12016 393283 12019
rect 402977 12019 403035 12025
rect 402977 12016 402989 12019
rect 393271 11988 402989 12016
rect 393271 11985 393283 11988
rect 393225 11979 393283 11985
rect 402977 11985 402989 11988
rect 403023 11985 403035 12019
rect 402977 11979 403035 11985
rect 403161 12019 403219 12025
rect 403161 11985 403173 12019
rect 403207 12016 403219 12019
rect 412361 12019 412419 12025
rect 412361 12016 412373 12019
rect 403207 11988 412373 12016
rect 403207 11985 403219 11988
rect 403161 11979 403219 11985
rect 412361 11985 412373 11988
rect 412407 11985 412419 12019
rect 412361 11979 412419 11985
rect 412545 12019 412603 12025
rect 412545 11985 412557 12019
rect 412591 12016 412603 12019
rect 419644 12016 419672 12056
rect 432138 12044 432144 12056
rect 432196 12044 432202 12096
rect 433426 12044 433432 12096
rect 433484 12084 433490 12096
rect 438213 12087 438271 12093
rect 438213 12084 438225 12087
rect 433484 12056 438225 12084
rect 433484 12044 433490 12056
rect 438213 12053 438225 12056
rect 438259 12053 438271 12087
rect 438213 12047 438271 12053
rect 441706 12044 441712 12096
rect 441764 12084 441770 12096
rect 442626 12084 442632 12096
rect 441764 12056 442632 12084
rect 441764 12044 441770 12056
rect 442626 12044 442632 12056
rect 442684 12044 442690 12096
rect 456886 12044 456892 12096
rect 456944 12084 456950 12096
rect 457622 12084 457628 12096
rect 456944 12056 457628 12084
rect 456944 12044 456950 12056
rect 457622 12044 457628 12056
rect 457680 12044 457686 12096
rect 431034 12016 431040 12028
rect 412591 11988 419672 12016
rect 422864 11988 431040 12016
rect 412591 11985 412603 11988
rect 412545 11979 412603 11985
rect 179322 11908 179328 11960
rect 179380 11948 179386 11960
rect 422864 11948 422892 11988
rect 431034 11976 431040 11988
rect 431092 11976 431098 12028
rect 460952 12016 460980 12124
rect 465534 12112 465540 12124
rect 465592 12112 465598 12164
rect 431144 11988 460980 12016
rect 429562 11948 429568 11960
rect 179380 11920 422892 11948
rect 422956 11920 429568 11948
rect 179380 11908 179386 11920
rect 175458 11840 175464 11892
rect 175516 11880 175522 11892
rect 422956 11880 422984 11920
rect 429562 11908 429568 11920
rect 429620 11908 429626 11960
rect 430482 11908 430488 11960
rect 430540 11948 430546 11960
rect 431144 11948 431172 11988
rect 463786 11976 463792 12028
rect 463844 12016 463850 12028
rect 464430 12016 464436 12028
rect 463844 11988 464436 12016
rect 463844 11976 463850 11988
rect 464430 11976 464436 11988
rect 464488 11976 464494 12028
rect 469398 11976 469404 12028
rect 469456 12016 469462 12028
rect 470226 12016 470232 12028
rect 469456 11988 470232 12016
rect 469456 11976 469462 11988
rect 470226 11976 470232 11988
rect 470284 11976 470290 12028
rect 470597 12019 470655 12025
rect 470597 11985 470609 12019
rect 470643 12016 470655 12019
rect 479334 12016 479340 12028
rect 470643 11988 479340 12016
rect 470643 11985 470655 11988
rect 470597 11979 470655 11985
rect 479334 11976 479340 11988
rect 479392 11976 479398 12028
rect 430540 11920 431172 11948
rect 430540 11908 430546 11920
rect 436094 11908 436100 11960
rect 436152 11948 436158 11960
rect 438213 11951 438271 11957
rect 436152 11920 438164 11948
rect 436152 11908 436158 11920
rect 434438 11880 434444 11892
rect 175516 11852 422984 11880
rect 423048 11852 434444 11880
rect 175516 11840 175522 11852
rect 38562 11772 38568 11824
rect 38620 11812 38626 11824
rect 147766 11812 147772 11824
rect 38620 11784 147772 11812
rect 38620 11772 38626 11784
rect 147766 11772 147772 11784
rect 147824 11772 147830 11824
rect 160002 11772 160008 11824
rect 160060 11812 160066 11824
rect 419353 11815 419411 11821
rect 419353 11812 419365 11815
rect 160060 11784 419365 11812
rect 160060 11772 160066 11784
rect 419353 11781 419365 11784
rect 419399 11781 419411 11815
rect 419353 11775 419411 11781
rect 419445 11815 419503 11821
rect 419445 11781 419457 11815
rect 419491 11812 419503 11815
rect 423048 11812 423076 11852
rect 434438 11840 434444 11852
rect 434496 11840 434502 11892
rect 437474 11840 437480 11892
rect 437532 11880 437538 11892
rect 438026 11880 438032 11892
rect 437532 11852 438032 11880
rect 437532 11840 437538 11852
rect 438026 11840 438032 11852
rect 438084 11840 438090 11892
rect 438136 11880 438164 11920
rect 438213 11917 438225 11951
rect 438259 11948 438271 11951
rect 472434 11948 472440 11960
rect 438259 11920 472440 11948
rect 438259 11917 438271 11920
rect 438213 11911 438271 11917
rect 472434 11908 472440 11920
rect 472492 11908 472498 11960
rect 485038 11948 485044 11960
rect 482664 11920 485044 11948
rect 470597 11883 470655 11889
rect 470597 11880 470609 11883
rect 438136 11852 470609 11880
rect 470597 11849 470609 11852
rect 470643 11849 470655 11883
rect 470597 11843 470655 11849
rect 470686 11840 470692 11892
rect 470744 11880 470750 11892
rect 471422 11880 471428 11892
rect 470744 11852 471428 11880
rect 470744 11840 470750 11852
rect 471422 11840 471428 11852
rect 471480 11840 471486 11892
rect 419491 11784 423076 11812
rect 419491 11781 419503 11784
rect 419445 11775 419503 11781
rect 426434 11772 426440 11824
rect 426492 11812 426498 11824
rect 482664 11812 482692 11920
rect 485038 11908 485044 11920
rect 485096 11908 485102 11960
rect 503530 11840 503536 11892
rect 503588 11880 503594 11892
rect 535270 11880 535276 11892
rect 503588 11852 535276 11880
rect 503588 11840 503594 11852
rect 535270 11840 535276 11852
rect 535328 11840 535334 11892
rect 426492 11784 482692 11812
rect 426492 11772 426498 11784
rect 483106 11772 483112 11824
rect 483164 11812 483170 11824
rect 484026 11812 484032 11824
rect 483164 11784 484032 11812
rect 483164 11772 483170 11784
rect 484026 11772 484032 11784
rect 484084 11772 484090 11824
rect 502242 11772 502248 11824
rect 502300 11812 502306 11824
rect 534902 11812 534908 11824
rect 502300 11784 534908 11812
rect 502300 11772 502306 11784
rect 534902 11772 534908 11784
rect 534960 11772 534966 11824
rect 132494 11704 132500 11756
rect 132552 11744 132558 11756
rect 416038 11744 416044 11756
rect 132552 11716 416044 11744
rect 132552 11704 132558 11716
rect 416038 11704 416044 11716
rect 416096 11704 416102 11756
rect 417970 11704 417976 11756
rect 418028 11744 418034 11756
rect 507670 11744 507676 11756
rect 418028 11716 507676 11744
rect 418028 11704 418034 11716
rect 507670 11704 507676 11716
rect 507728 11704 507734 11756
rect 524414 11704 524420 11756
rect 524472 11744 524478 11756
rect 524690 11744 524696 11756
rect 524472 11716 524696 11744
rect 524472 11704 524478 11716
rect 524690 11704 524696 11716
rect 524748 11704 524754 11756
rect 534718 11704 534724 11756
rect 534776 11744 534782 11756
rect 541802 11744 541808 11756
rect 534776 11716 541808 11744
rect 534776 11704 534782 11716
rect 541802 11704 541808 11716
rect 541860 11704 541866 11756
rect 210329 11679 210387 11685
rect 210329 11645 210341 11679
rect 210375 11676 210387 11679
rect 219345 11679 219403 11685
rect 219345 11676 219357 11679
rect 210375 11648 219357 11676
rect 210375 11645 210387 11648
rect 210329 11639 210387 11645
rect 219345 11645 219357 11648
rect 219391 11645 219403 11679
rect 219345 11639 219403 11645
rect 229097 11679 229155 11685
rect 229097 11645 229109 11679
rect 229143 11676 229155 11679
rect 238665 11679 238723 11685
rect 238665 11676 238677 11679
rect 229143 11648 238677 11676
rect 229143 11645 229155 11648
rect 229097 11639 229155 11645
rect 238665 11645 238677 11648
rect 238711 11645 238723 11679
rect 238665 11639 238723 11645
rect 248417 11679 248475 11685
rect 248417 11645 248429 11679
rect 248463 11676 248475 11679
rect 257985 11679 258043 11685
rect 257985 11676 257997 11679
rect 248463 11648 257997 11676
rect 248463 11645 248475 11648
rect 248417 11639 248475 11645
rect 257985 11645 257997 11648
rect 258031 11645 258043 11679
rect 257985 11639 258043 11645
rect 267737 11679 267795 11685
rect 267737 11645 267749 11679
rect 267783 11676 267795 11679
rect 277305 11679 277363 11685
rect 277305 11676 277317 11679
rect 267783 11648 277317 11676
rect 267783 11645 267795 11648
rect 267737 11639 267795 11645
rect 277305 11645 277317 11648
rect 277351 11645 277363 11679
rect 277305 11639 277363 11645
rect 287057 11679 287115 11685
rect 287057 11645 287069 11679
rect 287103 11676 287115 11679
rect 296625 11679 296683 11685
rect 296625 11676 296637 11679
rect 287103 11648 296637 11676
rect 287103 11645 287115 11648
rect 287057 11639 287115 11645
rect 296625 11645 296637 11648
rect 296671 11645 296683 11679
rect 296625 11639 296683 11645
rect 306377 11679 306435 11685
rect 306377 11645 306389 11679
rect 306423 11676 306435 11679
rect 315945 11679 316003 11685
rect 315945 11676 315957 11679
rect 306423 11648 315957 11676
rect 306423 11645 306435 11648
rect 306377 11639 306435 11645
rect 315945 11645 315957 11648
rect 315991 11645 316003 11679
rect 315945 11639 316003 11645
rect 325697 11679 325755 11685
rect 325697 11645 325709 11679
rect 325743 11676 325755 11679
rect 335265 11679 335323 11685
rect 335265 11676 335277 11679
rect 325743 11648 335277 11676
rect 325743 11645 325755 11648
rect 325697 11639 325755 11645
rect 335265 11645 335277 11648
rect 335311 11645 335323 11679
rect 335265 11639 335323 11645
rect 382182 11636 382188 11688
rect 382240 11676 382246 11688
rect 496170 11676 496176 11688
rect 382240 11648 496176 11676
rect 382240 11636 382246 11648
rect 496170 11636 496176 11648
rect 496228 11636 496234 11688
rect 507854 11636 507860 11688
rect 507912 11676 507918 11688
rect 508682 11676 508688 11688
rect 507912 11648 508688 11676
rect 507912 11636 507918 11648
rect 508682 11636 508688 11648
rect 508740 11636 508746 11688
rect 510706 11636 510712 11688
rect 510764 11676 510770 11688
rect 511626 11676 511632 11688
rect 510764 11648 511632 11676
rect 510764 11636 510770 11648
rect 511626 11636 511632 11648
rect 511684 11636 511690 11688
rect 524598 11636 524604 11688
rect 524656 11676 524662 11688
rect 525426 11676 525432 11688
rect 524656 11648 525432 11676
rect 524656 11636 524662 11648
rect 525426 11636 525432 11648
rect 525484 11636 525490 11688
rect 527266 11636 527272 11688
rect 527324 11676 527330 11688
rect 527726 11676 527732 11688
rect 527324 11648 527732 11676
rect 527324 11636 527330 11648
rect 527726 11636 527732 11648
rect 527784 11636 527790 11688
rect 267829 11611 267887 11617
rect 267829 11577 267841 11611
rect 267875 11608 267887 11611
rect 277213 11611 277271 11617
rect 277213 11608 277225 11611
rect 267875 11580 277225 11608
rect 267875 11577 267887 11580
rect 267829 11571 267887 11577
rect 277213 11577 277225 11580
rect 277259 11577 277271 11611
rect 277213 11571 277271 11577
rect 287149 11611 287207 11617
rect 287149 11577 287161 11611
rect 287195 11608 287207 11611
rect 296533 11611 296591 11617
rect 296533 11608 296545 11611
rect 287195 11580 296545 11608
rect 287195 11577 287207 11580
rect 287149 11571 287207 11577
rect 296533 11577 296545 11580
rect 296579 11577 296591 11611
rect 296533 11571 296591 11577
rect 306469 11611 306527 11617
rect 306469 11577 306481 11611
rect 306515 11608 306527 11611
rect 315853 11611 315911 11617
rect 315853 11608 315865 11611
rect 306515 11580 315865 11608
rect 306515 11577 306527 11580
rect 306469 11571 306527 11577
rect 315853 11577 315865 11580
rect 315899 11577 315911 11611
rect 315853 11571 315911 11577
rect 325789 11611 325847 11617
rect 325789 11577 325801 11611
rect 325835 11608 325847 11611
rect 335173 11611 335231 11617
rect 335173 11608 335185 11611
rect 325835 11580 335185 11608
rect 325835 11577 325847 11580
rect 325789 11571 325847 11577
rect 335173 11577 335185 11580
rect 335219 11577 335231 11611
rect 335173 11571 335231 11577
rect 384942 11568 384948 11620
rect 385000 11608 385006 11620
rect 497366 11608 497372 11620
rect 385000 11580 497372 11608
rect 385000 11568 385006 11580
rect 497366 11568 497372 11580
rect 497424 11568 497430 11620
rect 229094 11500 229100 11552
rect 229152 11540 229158 11552
rect 238662 11540 238668 11552
rect 229152 11512 238668 11540
rect 229152 11500 229158 11512
rect 238662 11500 238668 11512
rect 238720 11500 238726 11552
rect 248414 11500 248420 11552
rect 248472 11540 248478 11552
rect 257982 11540 257988 11552
rect 248472 11512 257988 11540
rect 248472 11500 248478 11512
rect 257982 11500 257988 11512
rect 258040 11500 258046 11552
rect 267734 11500 267740 11552
rect 267792 11540 267798 11552
rect 277302 11540 277308 11552
rect 267792 11512 277308 11540
rect 267792 11500 267798 11512
rect 277302 11500 277308 11512
rect 277360 11500 277366 11552
rect 287054 11500 287060 11552
rect 287112 11540 287118 11552
rect 296441 11543 296499 11549
rect 296441 11540 296453 11543
rect 287112 11512 296453 11540
rect 287112 11500 287118 11512
rect 296441 11509 296453 11512
rect 296487 11509 296499 11543
rect 296441 11503 296499 11509
rect 306374 11500 306380 11552
rect 306432 11540 306438 11552
rect 315942 11540 315948 11552
rect 306432 11512 315948 11540
rect 306432 11500 306438 11512
rect 315942 11500 315948 11512
rect 316000 11500 316006 11552
rect 325694 11500 325700 11552
rect 325752 11540 325758 11552
rect 335262 11540 335268 11552
rect 325752 11512 335268 11540
rect 325752 11500 325758 11512
rect 335262 11500 335268 11512
rect 335320 11500 335326 11552
rect 389082 11500 389088 11552
rect 389140 11540 389146 11552
rect 498470 11540 498476 11552
rect 389140 11512 498476 11540
rect 389140 11500 389146 11512
rect 498470 11500 498476 11512
rect 498528 11500 498534 11552
rect 391842 11432 391848 11484
rect 391900 11472 391906 11484
rect 499666 11472 499672 11484
rect 391900 11444 499672 11472
rect 391900 11432 391906 11444
rect 499666 11432 499672 11444
rect 499724 11432 499730 11484
rect 383657 11407 383715 11413
rect 383657 11373 383669 11407
rect 383703 11404 383715 11407
rect 393225 11407 393283 11413
rect 393225 11404 393237 11407
rect 383703 11376 393237 11404
rect 383703 11373 383715 11376
rect 383657 11367 383715 11373
rect 393225 11373 393237 11376
rect 393271 11373 393283 11407
rect 393225 11367 393283 11373
rect 395982 11364 395988 11416
rect 396040 11404 396046 11416
rect 500770 11404 500776 11416
rect 396040 11376 500776 11404
rect 396040 11364 396046 11376
rect 500770 11364 500776 11376
rect 500828 11364 500834 11416
rect 383749 11339 383807 11345
rect 383749 11305 383761 11339
rect 383795 11336 383807 11339
rect 393133 11339 393191 11345
rect 393133 11336 393145 11339
rect 383795 11308 393145 11336
rect 383795 11305 383807 11308
rect 383749 11299 383807 11305
rect 393133 11305 393145 11308
rect 393179 11305 393191 11339
rect 393133 11299 393191 11305
rect 400122 11296 400128 11348
rect 400180 11336 400186 11348
rect 501966 11336 501972 11348
rect 400180 11308 501972 11336
rect 400180 11296 400186 11308
rect 501966 11296 501972 11308
rect 502024 11296 502030 11348
rect 552198 11296 552204 11348
rect 552256 11336 552262 11348
rect 554958 11336 554964 11348
rect 552256 11308 554964 11336
rect 552256 11296 552262 11308
rect 554958 11296 554964 11308
rect 555016 11296 555022 11348
rect 407022 11228 407028 11280
rect 407080 11268 407086 11280
rect 504266 11268 504272 11280
rect 407080 11240 504272 11268
rect 407080 11228 407086 11240
rect 504266 11228 504272 11240
rect 504324 11228 504330 11280
rect 409690 11160 409696 11212
rect 409748 11200 409754 11212
rect 505370 11200 505376 11212
rect 409748 11172 505376 11200
rect 409748 11160 409754 11172
rect 505370 11160 505376 11172
rect 505428 11160 505434 11212
rect 402977 11135 403035 11141
rect 402977 11101 402989 11135
rect 403023 11132 403035 11135
rect 412545 11135 412603 11141
rect 412545 11132 412557 11135
rect 403023 11104 412557 11132
rect 403023 11101 403035 11104
rect 402977 11095 403035 11101
rect 412545 11101 412557 11104
rect 412591 11101 412603 11135
rect 412545 11095 412603 11101
rect 413922 11092 413928 11144
rect 413980 11132 413986 11144
rect 506566 11132 506572 11144
rect 413980 11104 506572 11132
rect 413980 11092 413986 11104
rect 506566 11092 506572 11104
rect 506624 11092 506630 11144
rect 403069 11067 403127 11073
rect 403069 11033 403081 11067
rect 403115 11064 403127 11067
rect 412453 11067 412511 11073
rect 412453 11064 412465 11067
rect 403115 11036 412465 11064
rect 403115 11033 403127 11036
rect 403069 11027 403127 11033
rect 412453 11033 412465 11036
rect 412499 11033 412511 11067
rect 412453 11027 412511 11033
rect 415486 11024 415492 11076
rect 415544 11064 415550 11076
rect 416314 11064 416320 11076
rect 415544 11036 416320 11064
rect 415544 11024 415550 11036
rect 416314 11024 416320 11036
rect 416372 11024 416378 11076
rect 419353 11067 419411 11073
rect 419353 11033 419365 11067
rect 419399 11064 419411 11067
rect 424870 11064 424876 11076
rect 419399 11036 424876 11064
rect 419399 11033 419411 11036
rect 419353 11027 419411 11033
rect 424870 11024 424876 11036
rect 424928 11024 424934 11076
rect 425054 11024 425060 11076
rect 425112 11064 425118 11076
rect 462038 11064 462044 11076
rect 425112 11036 462044 11064
rect 425112 11024 425118 11036
rect 462038 11024 462044 11036
rect 462096 11024 462102 11076
rect 465350 11024 465356 11076
rect 465408 11064 465414 11076
rect 466178 11064 466184 11076
rect 465408 11036 466184 11064
rect 465408 11024 465414 11036
rect 466178 11024 466184 11036
rect 466236 11024 466242 11076
rect 339402 10956 339408 11008
rect 339460 10996 339466 11008
rect 482370 10996 482376 11008
rect 339460 10968 482376 10996
rect 339460 10956 339466 10968
rect 482370 10956 482376 10968
rect 482428 10956 482434 11008
rect 335262 10888 335268 10940
rect 335320 10928 335326 10940
rect 481266 10928 481272 10940
rect 335320 10900 481272 10928
rect 335320 10888 335326 10900
rect 481266 10888 481272 10900
rect 481324 10888 481330 10940
rect 328362 10820 328368 10872
rect 328420 10860 328426 10872
rect 478966 10860 478972 10872
rect 328420 10832 478972 10860
rect 328420 10820 328426 10832
rect 478966 10820 478972 10832
rect 479024 10820 479030 10872
rect 324222 10752 324228 10804
rect 324280 10792 324286 10804
rect 477770 10792 477776 10804
rect 324280 10764 477776 10792
rect 324280 10752 324286 10764
rect 477770 10752 477776 10764
rect 477828 10752 477834 10804
rect 321462 10684 321468 10736
rect 321520 10724 321526 10736
rect 476666 10724 476672 10736
rect 321520 10696 476672 10724
rect 321520 10684 321526 10696
rect 476666 10684 476672 10696
rect 476724 10684 476730 10736
rect 298002 10616 298008 10668
rect 298060 10656 298066 10668
rect 304994 10656 305000 10668
rect 298060 10628 305000 10656
rect 298060 10616 298066 10628
rect 304994 10616 305000 10628
rect 305052 10616 305058 10668
rect 317322 10616 317328 10668
rect 317380 10656 317386 10668
rect 475470 10656 475476 10668
rect 317380 10628 475476 10656
rect 317380 10616 317386 10628
rect 475470 10616 475476 10628
rect 475528 10616 475534 10668
rect 485038 10616 485044 10668
rect 485096 10656 485102 10668
rect 510338 10656 510344 10668
rect 485096 10628 510344 10656
rect 485096 10616 485102 10628
rect 510338 10616 510344 10628
rect 510396 10616 510402 10668
rect 310422 10548 310428 10600
rect 310480 10588 310486 10600
rect 473170 10588 473176 10600
rect 310480 10560 473176 10588
rect 310480 10548 310486 10560
rect 473170 10548 473176 10560
rect 473228 10548 473234 10600
rect 479518 10548 479524 10600
rect 479576 10588 479582 10600
rect 505738 10588 505744 10600
rect 479576 10560 505744 10588
rect 479576 10548 479582 10560
rect 505738 10548 505744 10560
rect 505796 10548 505802 10600
rect 306282 10480 306288 10532
rect 306340 10520 306346 10532
rect 472066 10520 472072 10532
rect 306340 10492 472072 10520
rect 306340 10480 306346 10492
rect 472066 10480 472072 10492
rect 472124 10480 472130 10532
rect 499482 10480 499488 10532
rect 499540 10520 499546 10532
rect 534166 10520 534172 10532
rect 499540 10492 534172 10520
rect 499540 10480 499546 10492
rect 534166 10480 534172 10492
rect 534224 10480 534230 10532
rect 146846 10412 146852 10464
rect 146904 10452 146910 10464
rect 313274 10452 313280 10464
rect 146904 10424 313280 10452
rect 146904 10412 146910 10424
rect 313274 10412 313280 10424
rect 313332 10412 313338 10464
rect 314562 10412 314568 10464
rect 314620 10452 314626 10464
rect 474366 10452 474372 10464
rect 314620 10424 474372 10452
rect 314620 10412 314626 10424
rect 474366 10412 474372 10424
rect 474424 10412 474430 10464
rect 498102 10412 498108 10464
rect 498160 10452 498166 10464
rect 533798 10452 533804 10464
rect 498160 10424 533804 10452
rect 498160 10412 498166 10424
rect 533798 10412 533804 10424
rect 533856 10412 533862 10464
rect 289722 10344 289728 10396
rect 289780 10384 289786 10396
rect 302234 10384 302240 10396
rect 289780 10356 302240 10384
rect 289780 10344 289786 10356
rect 302234 10344 302240 10356
rect 302292 10344 302298 10396
rect 303522 10344 303528 10396
rect 303580 10384 303586 10396
rect 470870 10384 470876 10396
rect 303580 10356 470876 10384
rect 303580 10344 303586 10356
rect 470870 10344 470876 10356
rect 470928 10344 470934 10396
rect 486970 10344 486976 10396
rect 487028 10384 487034 10396
rect 530302 10384 530308 10396
rect 487028 10356 530308 10384
rect 487028 10344 487034 10356
rect 530302 10344 530308 10356
rect 530360 10344 530366 10396
rect 10410 10276 10416 10328
rect 10468 10316 10474 10328
rect 120074 10316 120080 10328
rect 10468 10288 120080 10316
rect 10468 10276 10474 10288
rect 120074 10276 120080 10288
rect 120132 10276 120138 10328
rect 161382 10276 161388 10328
rect 161440 10316 161446 10328
rect 330294 10316 330300 10328
rect 161440 10288 330300 10316
rect 161440 10276 161446 10288
rect 330294 10276 330300 10288
rect 330352 10276 330358 10328
rect 332410 10276 332416 10328
rect 332468 10316 332474 10328
rect 480070 10316 480076 10328
rect 332468 10288 480076 10316
rect 332468 10276 332474 10288
rect 480070 10276 480076 10288
rect 480128 10276 480134 10328
rect 481542 10276 481548 10328
rect 481600 10316 481606 10328
rect 528370 10316 528376 10328
rect 481600 10288 528376 10316
rect 481600 10276 481606 10288
rect 528370 10276 528376 10288
rect 528428 10276 528434 10328
rect 342162 10208 342168 10260
rect 342220 10248 342226 10260
rect 483566 10248 483572 10260
rect 342220 10220 483572 10248
rect 342220 10208 342226 10220
rect 483566 10208 483572 10220
rect 483624 10208 483630 10260
rect 346302 10140 346308 10192
rect 346360 10180 346366 10192
rect 484670 10180 484676 10192
rect 346360 10152 484676 10180
rect 346360 10140 346366 10152
rect 484670 10140 484676 10152
rect 484728 10140 484734 10192
rect 348970 10072 348976 10124
rect 349028 10112 349034 10124
rect 485866 10112 485872 10124
rect 349028 10084 485872 10112
rect 349028 10072 349034 10084
rect 485866 10072 485872 10084
rect 485924 10072 485930 10124
rect 353202 10004 353208 10056
rect 353260 10044 353266 10056
rect 486694 10044 486700 10056
rect 353260 10016 486700 10044
rect 353260 10004 353266 10016
rect 486694 10004 486700 10016
rect 486752 10004 486758 10056
rect 357342 9936 357348 9988
rect 357400 9976 357406 9988
rect 488166 9976 488172 9988
rect 357400 9948 488172 9976
rect 357400 9936 357406 9948
rect 488166 9936 488172 9948
rect 488224 9936 488230 9988
rect 360102 9868 360108 9920
rect 360160 9908 360166 9920
rect 489270 9908 489276 9920
rect 360160 9880 489276 9908
rect 360160 9868 360166 9880
rect 489270 9868 489276 9880
rect 489328 9868 489334 9920
rect 363322 9800 363328 9852
rect 363380 9840 363386 9852
rect 490466 9840 490472 9852
rect 363380 9812 490472 9840
rect 363380 9800 363386 9812
rect 490466 9800 490472 9812
rect 490524 9800 490530 9852
rect 367002 9732 367008 9784
rect 367060 9772 367066 9784
rect 491570 9772 491576 9784
rect 367060 9744 491576 9772
rect 367060 9732 367066 9744
rect 491570 9732 491576 9744
rect 491628 9732 491634 9784
rect 65978 9704 65984 9716
rect 65939 9676 65984 9704
rect 65978 9664 65984 9676
rect 66036 9664 66042 9716
rect 67174 9704 67180 9716
rect 67135 9676 67180 9704
rect 67174 9664 67180 9676
rect 67232 9664 67238 9716
rect 179414 9704 179420 9716
rect 179375 9676 179420 9704
rect 179414 9664 179420 9676
rect 179472 9664 179478 9716
rect 182174 9704 182180 9716
rect 182135 9676 182180 9704
rect 182174 9664 182180 9676
rect 182232 9664 182238 9716
rect 184842 9704 184848 9716
rect 184803 9676 184848 9704
rect 184842 9664 184848 9676
rect 184900 9664 184906 9716
rect 205726 9664 205732 9716
rect 205784 9704 205790 9716
rect 206002 9704 206008 9716
rect 205784 9676 206008 9704
rect 205784 9664 205790 9676
rect 206002 9664 206008 9676
rect 206060 9664 206066 9716
rect 208486 9664 208492 9716
rect 208544 9704 208550 9716
rect 208854 9704 208860 9716
rect 208544 9676 208860 9704
rect 208544 9664 208550 9676
rect 208854 9664 208860 9676
rect 208912 9664 208918 9716
rect 403618 9664 403624 9716
rect 403676 9704 403682 9716
rect 502334 9704 502340 9716
rect 403676 9676 502340 9704
rect 403676 9664 403682 9676
rect 502334 9664 502340 9676
rect 502392 9664 502398 9716
rect 530118 9664 530124 9716
rect 530176 9704 530182 9716
rect 530670 9704 530676 9716
rect 530176 9676 530676 9704
rect 530176 9664 530182 9676
rect 530670 9664 530676 9676
rect 530728 9664 530734 9716
rect 548886 9664 548892 9716
rect 548944 9704 548950 9716
rect 550266 9704 550272 9716
rect 548944 9676 550272 9704
rect 548944 9664 548950 9676
rect 550266 9664 550272 9676
rect 550324 9664 550330 9716
rect 126609 9639 126667 9645
rect 126609 9605 126621 9639
rect 126655 9636 126667 9639
rect 126882 9636 126888 9648
rect 126655 9608 126888 9636
rect 126655 9605 126667 9608
rect 126609 9599 126667 9605
rect 126882 9596 126888 9608
rect 126940 9596 126946 9648
rect 202782 9636 202788 9648
rect 202743 9608 202788 9636
rect 202782 9596 202788 9608
rect 202840 9596 202846 9648
rect 245562 9596 245568 9648
rect 245620 9636 245626 9648
rect 451921 9639 451979 9645
rect 245620 9608 451412 9636
rect 245620 9596 245626 9608
rect 241974 9528 241980 9580
rect 242032 9568 242038 9580
rect 451274 9568 451280 9580
rect 242032 9540 451280 9568
rect 242032 9528 242038 9540
rect 451274 9528 451280 9540
rect 451332 9528 451338 9580
rect 451384 9568 451412 9608
rect 451921 9605 451933 9639
rect 451967 9636 451979 9639
rect 477034 9636 477040 9648
rect 451967 9608 477040 9636
rect 451967 9605 451979 9608
rect 451921 9599 451979 9605
rect 477034 9596 477040 9608
rect 477092 9596 477098 9648
rect 452470 9568 452476 9580
rect 451384 9540 452476 9568
rect 452470 9528 452476 9540
rect 452528 9528 452534 9580
rect 452654 9528 452660 9580
rect 452712 9568 452718 9580
rect 486234 9568 486240 9580
rect 452712 9540 486240 9568
rect 452712 9528 452718 9540
rect 486234 9528 486240 9540
rect 486292 9528 486298 9580
rect 238386 9460 238392 9512
rect 238444 9500 238450 9512
rect 443181 9503 443239 9509
rect 443181 9500 443193 9503
rect 238444 9472 443193 9500
rect 238444 9460 238450 9472
rect 443181 9469 443193 9472
rect 443227 9469 443239 9503
rect 448790 9500 448796 9512
rect 443181 9463 443239 9469
rect 443288 9472 448796 9500
rect 234798 9392 234804 9444
rect 234856 9432 234862 9444
rect 443288 9432 443316 9472
rect 448790 9460 448796 9472
rect 448848 9460 448854 9512
rect 451182 9460 451188 9512
rect 451240 9500 451246 9512
rect 483934 9500 483940 9512
rect 451240 9472 483940 9500
rect 451240 9460 451246 9472
rect 483934 9460 483940 9472
rect 483992 9460 483998 9512
rect 447870 9432 447876 9444
rect 234856 9404 443316 9432
rect 443380 9404 447876 9432
rect 234856 9392 234862 9404
rect 231302 9324 231308 9376
rect 231360 9364 231366 9376
rect 443380 9364 443408 9404
rect 447870 9392 447876 9404
rect 447928 9392 447934 9444
rect 458542 9392 458548 9444
rect 458600 9432 458606 9444
rect 493134 9432 493140 9444
rect 458600 9404 493140 9432
rect 458600 9392 458606 9404
rect 493134 9392 493140 9404
rect 493192 9392 493198 9444
rect 494238 9392 494244 9444
rect 494296 9432 494302 9444
rect 532326 9432 532332 9444
rect 494296 9404 532332 9432
rect 494296 9392 494302 9404
rect 532326 9392 532332 9404
rect 532384 9392 532390 9444
rect 446766 9364 446772 9376
rect 231360 9336 443408 9364
rect 443472 9336 446772 9364
rect 231360 9324 231366 9336
rect 227714 9256 227720 9308
rect 227772 9296 227778 9308
rect 443472 9296 443500 9336
rect 446766 9324 446772 9336
rect 446824 9324 446830 9376
rect 452746 9324 452752 9376
rect 452804 9364 452810 9376
rect 488534 9364 488540 9376
rect 452804 9336 488540 9364
rect 452804 9324 452810 9336
rect 488534 9324 488540 9336
rect 488592 9324 488598 9376
rect 495342 9324 495348 9376
rect 495400 9364 495406 9376
rect 532970 9364 532976 9376
rect 495400 9336 532976 9364
rect 495400 9324 495406 9336
rect 532970 9324 532976 9336
rect 533028 9324 533034 9376
rect 445570 9296 445576 9308
rect 227772 9268 443500 9296
rect 443564 9268 445576 9296
rect 227772 9256 227778 9268
rect 224126 9188 224132 9240
rect 224184 9228 224190 9240
rect 443564 9228 443592 9268
rect 445570 9256 445576 9268
rect 445628 9256 445634 9308
rect 446214 9256 446220 9308
rect 446272 9296 446278 9308
rect 481634 9296 481640 9308
rect 446272 9268 481640 9296
rect 446272 9256 446278 9268
rect 481634 9256 481640 9268
rect 481692 9256 481698 9308
rect 483474 9256 483480 9308
rect 483532 9296 483538 9308
rect 529198 9296 529204 9308
rect 483532 9268 529204 9296
rect 483532 9256 483538 9268
rect 529198 9256 529204 9268
rect 529256 9256 529262 9308
rect 224184 9200 443592 9228
rect 224184 9188 224190 9200
rect 445294 9188 445300 9240
rect 445352 9228 445358 9240
rect 451921 9231 451979 9237
rect 451921 9228 451933 9231
rect 445352 9200 451933 9228
rect 445352 9188 445358 9200
rect 451921 9197 451933 9200
rect 451967 9197 451979 9231
rect 451921 9191 451979 9197
rect 463234 9188 463240 9240
rect 463292 9228 463298 9240
rect 522666 9228 522672 9240
rect 463292 9200 522672 9228
rect 463292 9188 463298 9200
rect 522666 9188 522672 9200
rect 522724 9188 522730 9240
rect 220538 9120 220544 9172
rect 220596 9160 220602 9172
rect 444466 9160 444472 9172
rect 220596 9132 444472 9160
rect 220596 9120 220602 9132
rect 444466 9120 444472 9132
rect 444524 9120 444530 9172
rect 459738 9120 459744 9172
rect 459796 9160 459802 9172
rect 521470 9160 521476 9172
rect 459796 9132 521476 9160
rect 459796 9120 459802 9132
rect 521470 9120 521476 9132
rect 521528 9120 521534 9172
rect 217042 9052 217048 9104
rect 217100 9092 217106 9104
rect 442994 9092 443000 9104
rect 217100 9064 443000 9092
rect 217100 9052 217106 9064
rect 442994 9052 443000 9064
rect 443052 9052 443058 9104
rect 443181 9095 443239 9101
rect 443181 9061 443193 9095
rect 443227 9092 443239 9095
rect 450170 9092 450176 9104
rect 443227 9064 450176 9092
rect 443227 9061 443239 9064
rect 443181 9055 443239 9061
rect 450170 9052 450176 9064
rect 450228 9052 450234 9104
rect 456058 9052 456064 9104
rect 456116 9092 456122 9104
rect 520274 9092 520280 9104
rect 456116 9064 520280 9092
rect 456116 9052 456122 9064
rect 520274 9052 520280 9064
rect 520332 9052 520338 9104
rect 150618 8984 150624 9036
rect 150676 9024 150682 9036
rect 174170 9024 174176 9036
rect 150676 8996 174176 9024
rect 150676 8984 150682 8996
rect 174170 8984 174176 8996
rect 174228 8984 174234 9036
rect 213454 8984 213460 9036
rect 213512 9024 213518 9036
rect 442166 9024 442172 9036
rect 213512 8996 442172 9024
rect 213512 8984 213518 8996
rect 442166 8984 442172 8996
rect 442224 8984 442230 9036
rect 452470 8984 452476 9036
rect 452528 9024 452534 9036
rect 518986 9024 518992 9036
rect 452528 8996 518992 9024
rect 452528 8984 452534 8996
rect 518986 8984 518992 8996
rect 519044 8984 519050 9036
rect 18322 8916 18328 8968
rect 18380 8956 18386 8968
rect 132586 8956 132592 8968
rect 18380 8928 132592 8956
rect 18380 8916 18386 8928
rect 132586 8916 132592 8928
rect 132644 8916 132650 8968
rect 153930 8916 153936 8968
rect 153988 8956 153994 8968
rect 204898 8956 204904 8968
rect 153988 8928 204904 8956
rect 153988 8916 153994 8928
rect 204898 8916 204904 8928
rect 204956 8916 204962 8968
rect 209866 8916 209872 8968
rect 209924 8956 209930 8968
rect 440970 8956 440976 8968
rect 209924 8928 440976 8956
rect 209924 8916 209930 8928
rect 440970 8916 440976 8928
rect 441028 8916 441034 8968
rect 448977 8959 449035 8965
rect 448977 8925 448989 8959
rect 449023 8956 449035 8959
rect 518066 8956 518072 8968
rect 449023 8928 518072 8956
rect 449023 8925 449035 8928
rect 448977 8919 449035 8925
rect 518066 8916 518072 8928
rect 518124 8916 518130 8968
rect 533246 8916 533252 8968
rect 533304 8956 533310 8968
rect 542998 8956 543004 8968
rect 533304 8928 543004 8956
rect 533304 8916 533310 8928
rect 542998 8916 543004 8928
rect 543056 8916 543062 8968
rect 249150 8848 249156 8900
rect 249208 8888 249214 8900
rect 453666 8888 453672 8900
rect 249208 8860 453672 8888
rect 249208 8848 249214 8860
rect 453666 8848 453672 8860
rect 453724 8848 453730 8900
rect 252646 8780 252652 8832
rect 252704 8820 252710 8832
rect 454770 8820 454776 8832
rect 252704 8792 454776 8820
rect 252704 8780 252710 8792
rect 454770 8780 454776 8792
rect 454828 8780 454834 8832
rect 256234 8712 256240 8764
rect 256292 8752 256298 8764
rect 455966 8752 455972 8764
rect 256292 8724 455972 8752
rect 256292 8712 256298 8724
rect 455966 8712 455972 8724
rect 456024 8712 456030 8764
rect 259822 8644 259828 8696
rect 259880 8684 259886 8696
rect 457070 8684 457076 8696
rect 259880 8656 457076 8684
rect 259880 8644 259886 8656
rect 457070 8644 457076 8656
rect 457128 8644 457134 8696
rect 263410 8576 263416 8628
rect 263468 8616 263474 8628
rect 458266 8616 458272 8628
rect 263468 8588 458272 8616
rect 263468 8576 263474 8588
rect 458266 8576 458272 8588
rect 458324 8576 458330 8628
rect 266998 8508 267004 8560
rect 267056 8548 267062 8560
rect 459370 8548 459376 8560
rect 267056 8520 459376 8548
rect 267056 8508 267062 8520
rect 459370 8508 459376 8520
rect 459428 8508 459434 8560
rect 270494 8440 270500 8492
rect 270552 8480 270558 8492
rect 460566 8480 460572 8492
rect 270552 8452 460572 8480
rect 270552 8440 270558 8452
rect 460566 8440 460572 8452
rect 460624 8440 460630 8492
rect 370406 8372 370412 8424
rect 370464 8412 370470 8424
rect 492766 8412 492772 8424
rect 370464 8384 492772 8412
rect 370464 8372 370470 8384
rect 492766 8372 492772 8384
rect 492824 8372 492830 8424
rect 402514 8304 402520 8356
rect 402572 8344 402578 8356
rect 503070 8344 503076 8356
rect 402572 8316 503076 8344
rect 402572 8304 402578 8316
rect 503070 8304 503076 8316
rect 503128 8304 503134 8356
rect 372798 8236 372804 8288
rect 372856 8276 372862 8288
rect 493502 8276 493508 8288
rect 372856 8248 493508 8276
rect 372856 8236 372862 8248
rect 493502 8236 493508 8248
rect 493560 8236 493566 8288
rect 369210 8168 369216 8220
rect 369268 8208 369274 8220
rect 492398 8208 492404 8220
rect 369268 8180 492404 8208
rect 369268 8168 369274 8180
rect 492398 8168 492404 8180
rect 492456 8168 492462 8220
rect 365714 8100 365720 8152
rect 365772 8140 365778 8152
rect 490926 8140 490932 8152
rect 365772 8112 490932 8140
rect 365772 8100 365778 8112
rect 490926 8100 490932 8112
rect 490984 8100 490990 8152
rect 292298 8032 292304 8084
rect 292356 8072 292362 8084
rect 459554 8072 459560 8084
rect 292356 8044 459560 8072
rect 292356 8032 292362 8044
rect 459554 8032 459560 8044
rect 459612 8032 459618 8084
rect 220814 7964 220820 8016
rect 220872 8004 220878 8016
rect 432966 8004 432972 8016
rect 220872 7976 432972 8004
rect 220872 7964 220878 7976
rect 432966 7964 432972 7976
rect 433024 7964 433030 8016
rect 195514 7896 195520 7948
rect 195572 7936 195578 7948
rect 431770 7936 431776 7948
rect 195572 7908 431776 7936
rect 195572 7896 195578 7908
rect 431770 7896 431776 7908
rect 431828 7896 431834 7948
rect 186225 7871 186283 7877
rect 186225 7837 186237 7871
rect 186271 7868 186283 7871
rect 428366 7868 428372 7880
rect 186271 7840 428372 7868
rect 186271 7837 186283 7840
rect 186225 7831 186283 7837
rect 428366 7828 428372 7840
rect 428424 7828 428430 7880
rect 441890 7828 441896 7880
rect 441948 7868 441954 7880
rect 515766 7868 515772 7880
rect 441948 7840 515772 7868
rect 441948 7828 441954 7840
rect 515766 7828 515772 7840
rect 515824 7828 515830 7880
rect 177758 7760 177764 7812
rect 177816 7800 177822 7812
rect 430666 7800 430672 7812
rect 177816 7772 430672 7800
rect 177816 7760 177822 7772
rect 430666 7760 430672 7772
rect 430724 7760 430730 7812
rect 438210 7760 438216 7812
rect 438268 7800 438274 7812
rect 514570 7800 514576 7812
rect 438268 7772 514576 7800
rect 438268 7760 438274 7772
rect 514570 7760 514576 7772
rect 514628 7760 514634 7812
rect 174170 7692 174176 7744
rect 174228 7732 174234 7744
rect 429470 7732 429476 7744
rect 174228 7704 429476 7732
rect 174228 7692 174234 7704
rect 429470 7692 429476 7704
rect 429528 7692 429534 7744
rect 434622 7692 434628 7744
rect 434680 7732 434686 7744
rect 513466 7732 513472 7744
rect 434680 7704 513472 7732
rect 434680 7692 434686 7704
rect 513466 7692 513472 7704
rect 513524 7692 513530 7744
rect 167086 7624 167092 7676
rect 167144 7664 167150 7676
rect 427170 7664 427176 7676
rect 167144 7636 427176 7664
rect 167144 7624 167150 7636
rect 427170 7624 427176 7636
rect 427228 7624 427234 7676
rect 431126 7624 431132 7676
rect 431184 7664 431190 7676
rect 512270 7664 512276 7676
rect 431184 7636 512276 7664
rect 431184 7624 431190 7636
rect 512270 7624 512276 7636
rect 512328 7624 512334 7676
rect 513190 7624 513196 7676
rect 513248 7664 513254 7676
rect 538766 7664 538772 7676
rect 513248 7636 538772 7664
rect 513248 7624 513254 7636
rect 538766 7624 538772 7636
rect 538824 7624 538830 7676
rect 31478 7556 31484 7608
rect 31536 7596 31542 7608
rect 142246 7596 142252 7608
rect 31536 7568 142252 7596
rect 31536 7556 31542 7568
rect 142246 7556 142252 7568
rect 142304 7556 142310 7608
rect 143258 7556 143264 7608
rect 143316 7596 143322 7608
rect 144178 7596 144184 7608
rect 143316 7568 144184 7596
rect 143316 7556 143322 7568
rect 144178 7556 144184 7568
rect 144236 7556 144242 7608
rect 163498 7556 163504 7608
rect 163556 7596 163562 7608
rect 426066 7596 426072 7608
rect 163556 7568 426072 7596
rect 163556 7556 163562 7568
rect 426066 7556 426072 7568
rect 426124 7556 426130 7608
rect 427538 7556 427544 7608
rect 427596 7596 427602 7608
rect 511166 7596 511172 7608
rect 427596 7568 511172 7596
rect 427596 7556 427602 7568
rect 511166 7556 511172 7568
rect 511224 7556 511230 7608
rect 511994 7556 512000 7608
rect 512052 7596 512058 7608
rect 538398 7596 538404 7608
rect 512052 7568 538404 7596
rect 512052 7556 512058 7568
rect 538398 7556 538404 7568
rect 538456 7556 538462 7608
rect 376386 7488 376392 7540
rect 376444 7528 376450 7540
rect 494698 7528 494704 7540
rect 376444 7500 494704 7528
rect 376444 7488 376450 7500
rect 494698 7488 494704 7500
rect 494756 7488 494762 7540
rect 379974 7420 379980 7472
rect 380032 7460 380038 7472
rect 495802 7460 495808 7472
rect 380032 7432 495808 7460
rect 380032 7420 380038 7432
rect 495802 7420 495808 7432
rect 495860 7420 495866 7472
rect 383470 7352 383476 7404
rect 383528 7392 383534 7404
rect 496998 7392 497004 7404
rect 383528 7364 497004 7392
rect 383528 7352 383534 7364
rect 496998 7352 497004 7364
rect 497056 7352 497062 7404
rect 390646 7284 390652 7336
rect 390704 7324 390710 7336
rect 499298 7324 499304 7336
rect 390704 7296 499304 7324
rect 390704 7284 390710 7296
rect 499298 7284 499304 7296
rect 499356 7284 499362 7336
rect 394234 7216 394240 7268
rect 394292 7256 394298 7268
rect 500402 7256 500408 7268
rect 394292 7228 500408 7256
rect 394292 7216 394298 7228
rect 500402 7216 500408 7228
rect 500460 7216 500466 7268
rect 397822 7148 397828 7200
rect 397880 7188 397886 7200
rect 501598 7188 501604 7200
rect 397880 7160 501604 7188
rect 397880 7148 397886 7160
rect 501598 7148 501604 7160
rect 501656 7148 501662 7200
rect 401318 7080 401324 7132
rect 401376 7120 401382 7132
rect 502702 7120 502708 7132
rect 401376 7092 502708 7120
rect 401376 7080 401382 7092
rect 502702 7080 502708 7092
rect 502760 7080 502766 7132
rect 404906 7012 404912 7064
rect 404964 7052 404970 7064
rect 503898 7052 503904 7064
rect 404964 7024 503904 7052
rect 404964 7012 404970 7024
rect 503898 7012 503904 7024
rect 503956 7012 503962 7064
rect 412082 6944 412088 6996
rect 412140 6984 412146 6996
rect 506198 6984 506204 6996
rect 412140 6956 506204 6984
rect 412140 6944 412146 6956
rect 506198 6944 506204 6956
rect 506256 6944 506262 6996
rect 539594 6876 539600 6928
rect 539652 6916 539658 6928
rect 540514 6916 540520 6928
rect 539652 6888 540520 6916
rect 539652 6876 539658 6888
rect 540514 6876 540520 6888
rect 540572 6876 540578 6928
rect 77846 6808 77852 6860
rect 77904 6848 77910 6860
rect 175366 6848 175372 6860
rect 77904 6820 175372 6848
rect 77904 6808 77910 6820
rect 175366 6808 175372 6820
rect 175424 6808 175430 6860
rect 315758 6808 315764 6860
rect 315816 6848 315822 6860
rect 474918 6848 474924 6860
rect 315816 6820 474924 6848
rect 315816 6808 315822 6820
rect 474918 6808 474924 6820
rect 474976 6808 474982 6860
rect 70670 6740 70676 6792
rect 70728 6780 70734 6792
rect 171226 6780 171232 6792
rect 70728 6752 171232 6780
rect 70728 6740 70734 6752
rect 171226 6740 171232 6752
rect 171284 6740 171290 6792
rect 312170 6740 312176 6792
rect 312228 6780 312234 6792
rect 473446 6780 473452 6792
rect 312228 6752 473452 6780
rect 312228 6740 312234 6752
rect 473446 6740 473452 6752
rect 473504 6740 473510 6792
rect 63586 6672 63592 6724
rect 63644 6712 63650 6724
rect 165706 6712 165712 6724
rect 63644 6684 165712 6712
rect 63644 6672 63650 6684
rect 165706 6672 165712 6684
rect 165764 6672 165770 6724
rect 308582 6672 308588 6724
rect 308640 6712 308646 6724
rect 472158 6712 472164 6724
rect 308640 6684 472164 6712
rect 308640 6672 308646 6684
rect 472158 6672 472164 6684
rect 472216 6672 472222 6724
rect 56410 6604 56416 6656
rect 56468 6644 56474 6656
rect 160094 6644 160100 6656
rect 56468 6616 160100 6644
rect 56468 6604 56474 6616
rect 160094 6604 160100 6616
rect 160152 6604 160158 6656
rect 304994 6604 305000 6656
rect 305052 6644 305058 6656
rect 470686 6644 470692 6656
rect 305052 6616 470692 6644
rect 305052 6604 305058 6616
rect 470686 6604 470692 6616
rect 470744 6604 470750 6656
rect 476114 6604 476120 6656
rect 476172 6644 476178 6656
rect 496906 6644 496912 6656
rect 476172 6616 496912 6644
rect 476172 6604 476178 6616
rect 496906 6604 496912 6616
rect 496964 6604 496970 6656
rect 49326 6536 49332 6588
rect 49384 6576 49390 6588
rect 154574 6576 154580 6588
rect 49384 6548 154580 6576
rect 49384 6536 49390 6548
rect 154574 6536 154580 6548
rect 154632 6536 154638 6588
rect 301406 6536 301412 6588
rect 301464 6576 301470 6588
rect 469398 6576 469404 6588
rect 301464 6548 469404 6576
rect 301464 6536 301470 6548
rect 469398 6536 469404 6548
rect 469456 6536 469462 6588
rect 480714 6536 480720 6588
rect 480772 6576 480778 6588
rect 509326 6576 509332 6588
rect 480772 6548 509332 6576
rect 480772 6536 480778 6548
rect 509326 6536 509332 6548
rect 509384 6536 509390 6588
rect 44542 6468 44548 6520
rect 44600 6508 44606 6520
rect 151814 6508 151820 6520
rect 44600 6480 151820 6508
rect 44600 6468 44606 6480
rect 151814 6468 151820 6480
rect 151872 6468 151878 6520
rect 297910 6468 297916 6520
rect 297968 6508 297974 6520
rect 469306 6508 469312 6520
rect 297968 6480 469312 6508
rect 297968 6468 297974 6480
rect 469306 6468 469312 6480
rect 469364 6468 469370 6520
rect 471882 6468 471888 6520
rect 471940 6508 471946 6520
rect 495618 6508 495624 6520
rect 471940 6480 495624 6508
rect 471940 6468 471946 6480
rect 495618 6468 495624 6480
rect 495676 6468 495682 6520
rect 506014 6468 506020 6520
rect 506072 6508 506078 6520
rect 535638 6508 535644 6520
rect 506072 6480 535644 6508
rect 506072 6468 506078 6480
rect 535638 6468 535644 6480
rect 535696 6468 535702 6520
rect 40954 6400 40960 6452
rect 41012 6440 41018 6452
rect 149146 6440 149152 6452
rect 41012 6412 149152 6440
rect 41012 6400 41018 6412
rect 149146 6400 149152 6412
rect 149204 6400 149210 6452
rect 294322 6400 294328 6452
rect 294380 6440 294386 6452
rect 468018 6440 468024 6452
rect 294380 6412 468024 6440
rect 294380 6400 294386 6412
rect 468018 6400 468024 6412
rect 468076 6400 468082 6452
rect 477586 6400 477592 6452
rect 477644 6440 477650 6452
rect 502518 6440 502524 6452
rect 477644 6412 502524 6440
rect 477644 6400 477650 6412
rect 502518 6400 502524 6412
rect 502576 6400 502582 6452
rect 504818 6400 504824 6452
rect 504876 6440 504882 6452
rect 535546 6440 535552 6452
rect 504876 6412 535552 6440
rect 504876 6400 504882 6412
rect 535546 6400 535552 6412
rect 535604 6400 535610 6452
rect 37366 6332 37372 6384
rect 37424 6372 37430 6384
rect 146294 6372 146300 6384
rect 37424 6344 146300 6372
rect 37424 6332 37430 6344
rect 146294 6332 146300 6344
rect 146352 6332 146358 6384
rect 290734 6332 290740 6384
rect 290792 6372 290798 6384
rect 466546 6372 466552 6384
rect 290792 6344 466552 6372
rect 290792 6332 290798 6344
rect 466546 6332 466552 6344
rect 466604 6332 466610 6384
rect 473906 6332 473912 6384
rect 473964 6372 473970 6384
rect 525886 6372 525892 6384
rect 473964 6344 525892 6372
rect 473964 6332 473970 6344
rect 525886 6332 525892 6344
rect 525944 6332 525950 6384
rect 33870 6264 33876 6316
rect 33928 6304 33934 6316
rect 143534 6304 143540 6316
rect 33928 6276 143540 6304
rect 33928 6264 33934 6276
rect 143534 6264 143540 6276
rect 143592 6264 143598 6316
rect 287146 6264 287152 6316
rect 287204 6304 287210 6316
rect 465166 6304 465172 6316
rect 287204 6276 465172 6304
rect 287204 6264 287210 6276
rect 465166 6264 465172 6276
rect 465224 6264 465230 6316
rect 470318 6264 470324 6316
rect 470376 6304 470382 6316
rect 524414 6304 524420 6316
rect 470376 6276 524420 6304
rect 470376 6264 470382 6276
rect 524414 6264 524420 6276
rect 524472 6264 524478 6316
rect 8846 6196 8852 6248
rect 8904 6236 8910 6248
rect 125686 6236 125692 6248
rect 8904 6208 125692 6236
rect 8904 6196 8910 6208
rect 125686 6196 125692 6208
rect 125744 6196 125750 6248
rect 149238 6196 149244 6248
rect 149296 6236 149302 6248
rect 421190 6236 421196 6248
rect 149296 6208 421196 6236
rect 149296 6196 149302 6208
rect 421190 6196 421196 6208
rect 421248 6196 421254 6248
rect 423950 6196 423956 6248
rect 424008 6236 424014 6248
rect 509510 6236 509516 6248
rect 424008 6208 509516 6236
rect 424008 6196 424014 6208
rect 509510 6196 509516 6208
rect 509568 6196 509574 6248
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 121638 6168 121644 6180
rect 4120 6140 121644 6168
rect 4120 6128 4126 6140
rect 121638 6128 121644 6140
rect 121696 6128 121702 6180
rect 144454 6128 144460 6180
rect 144512 6168 144518 6180
rect 419718 6168 419724 6180
rect 144512 6140 419724 6168
rect 144512 6128 144518 6140
rect 419718 6128 419724 6140
rect 419776 6128 419782 6180
rect 420362 6128 420368 6180
rect 420420 6168 420426 6180
rect 507854 6168 507860 6180
rect 420420 6140 507860 6168
rect 420420 6128 420426 6140
rect 507854 6128 507860 6140
rect 507912 6128 507918 6180
rect 519078 6128 519084 6180
rect 519136 6168 519142 6180
rect 539594 6168 539600 6180
rect 519136 6140 539600 6168
rect 519136 6128 519142 6140
rect 539594 6128 539600 6140
rect 539652 6128 539658 6180
rect 319254 6060 319260 6112
rect 319312 6100 319318 6112
rect 476206 6100 476212 6112
rect 319312 6072 476212 6100
rect 319312 6060 319318 6072
rect 476206 6060 476212 6072
rect 476264 6060 476270 6112
rect 322842 5992 322848 6044
rect 322900 6032 322906 6044
rect 476298 6032 476304 6044
rect 322900 6004 476304 6032
rect 322900 5992 322906 6004
rect 476298 5992 476304 6004
rect 476356 5992 476362 6044
rect 326430 5924 326436 5976
rect 326488 5964 326494 5976
rect 477494 5964 477500 5976
rect 326488 5936 477500 5964
rect 326488 5924 326494 5936
rect 477494 5924 477500 5936
rect 477552 5924 477558 5976
rect 330018 5856 330024 5908
rect 330076 5896 330082 5908
rect 479058 5896 479064 5908
rect 330076 5868 479064 5896
rect 330076 5856 330082 5868
rect 479058 5856 479064 5868
rect 479116 5856 479122 5908
rect 333606 5788 333612 5840
rect 333664 5828 333670 5840
rect 480346 5828 480352 5840
rect 333664 5800 480352 5828
rect 333664 5788 333670 5800
rect 480346 5788 480352 5800
rect 480404 5788 480410 5840
rect 337102 5720 337108 5772
rect 337160 5760 337166 5772
rect 481818 5760 481824 5772
rect 337160 5732 481824 5760
rect 337160 5720 337166 5732
rect 481818 5720 481824 5732
rect 481876 5720 481882 5772
rect 340690 5652 340696 5704
rect 340748 5692 340754 5704
rect 483290 5692 483296 5704
rect 340748 5664 483296 5692
rect 340748 5652 340754 5664
rect 483290 5652 483296 5664
rect 483348 5652 483354 5704
rect 344278 5584 344284 5636
rect 344336 5624 344342 5636
rect 483106 5624 483112 5636
rect 344336 5596 483112 5624
rect 344336 5584 344342 5596
rect 483106 5584 483112 5596
rect 483164 5584 483170 5636
rect 385770 5516 385776 5568
rect 385828 5556 385834 5568
rect 470870 5556 470876 5568
rect 385828 5528 470876 5556
rect 385828 5516 385834 5528
rect 470870 5516 470876 5528
rect 470928 5516 470934 5568
rect 90910 5448 90916 5500
rect 90968 5488 90974 5500
rect 184750 5488 184756 5500
rect 90968 5460 184756 5488
rect 90968 5448 90974 5460
rect 184750 5448 184756 5460
rect 184808 5448 184814 5500
rect 240778 5448 240784 5500
rect 240836 5488 240842 5500
rect 450630 5488 450636 5500
rect 240836 5460 450636 5488
rect 240836 5448 240842 5460
rect 450630 5448 450636 5460
rect 450688 5448 450694 5500
rect 469122 5448 469128 5500
rect 469180 5488 469186 5500
rect 524506 5488 524512 5500
rect 469180 5460 524512 5488
rect 469180 5448 469186 5460
rect 524506 5448 524512 5460
rect 524564 5448 524570 5500
rect 87322 5380 87328 5432
rect 87380 5420 87386 5432
rect 182174 5420 182180 5432
rect 87380 5392 182180 5420
rect 87380 5380 87386 5392
rect 182174 5380 182180 5392
rect 182232 5380 182238 5432
rect 237190 5380 237196 5432
rect 237248 5420 237254 5432
rect 449526 5420 449532 5432
rect 237248 5392 449532 5420
rect 237248 5380 237254 5392
rect 449526 5380 449532 5392
rect 449584 5380 449590 5432
rect 465626 5380 465632 5432
rect 465684 5420 465690 5432
rect 523310 5420 523316 5432
rect 465684 5392 523316 5420
rect 465684 5380 465690 5392
rect 523310 5380 523316 5392
rect 523368 5380 523374 5432
rect 83826 5312 83832 5364
rect 83884 5352 83890 5364
rect 179414 5352 179420 5364
rect 83884 5324 179420 5352
rect 83884 5312 83890 5324
rect 179414 5312 179420 5324
rect 179472 5312 179478 5364
rect 233694 5312 233700 5364
rect 233752 5352 233758 5364
rect 448698 5352 448704 5364
rect 233752 5324 448704 5352
rect 233752 5312 233758 5324
rect 448698 5312 448704 5324
rect 448756 5312 448762 5364
rect 462038 5312 462044 5364
rect 462096 5352 462102 5364
rect 521930 5352 521936 5364
rect 462096 5324 521936 5352
rect 462096 5312 462102 5324
rect 521930 5312 521936 5324
rect 521988 5312 521994 5364
rect 80238 5244 80244 5296
rect 80296 5284 80302 5296
rect 178034 5284 178040 5296
rect 80296 5256 178040 5284
rect 80296 5244 80302 5256
rect 178034 5244 178040 5256
rect 178092 5244 178098 5296
rect 230106 5244 230112 5296
rect 230164 5284 230170 5296
rect 447318 5284 447324 5296
rect 230164 5256 447324 5284
rect 230164 5244 230170 5256
rect 447318 5244 447324 5256
rect 447376 5244 447382 5296
rect 458450 5244 458456 5296
rect 458508 5284 458514 5296
rect 520826 5284 520832 5296
rect 458508 5256 520832 5284
rect 458508 5244 458514 5256
rect 520826 5244 520832 5256
rect 520884 5244 520890 5296
rect 76650 5176 76656 5228
rect 76708 5216 76714 5228
rect 175274 5216 175280 5228
rect 76708 5188 175280 5216
rect 76708 5176 76714 5188
rect 175274 5176 175280 5188
rect 175332 5176 175338 5228
rect 226518 5176 226524 5228
rect 226576 5216 226582 5228
rect 445846 5216 445852 5228
rect 226576 5188 445852 5216
rect 226576 5176 226582 5188
rect 445846 5176 445852 5188
rect 445904 5176 445910 5228
rect 454862 5176 454868 5228
rect 454920 5216 454926 5228
rect 519630 5216 519636 5228
rect 454920 5188 519636 5216
rect 454920 5176 454926 5188
rect 519630 5176 519636 5188
rect 519688 5176 519694 5228
rect 69474 5108 69480 5160
rect 69532 5148 69538 5160
rect 169754 5148 169760 5160
rect 69532 5120 169760 5148
rect 69532 5108 69538 5120
rect 169754 5108 169760 5120
rect 169812 5108 169818 5160
rect 222930 5108 222936 5160
rect 222988 5148 222994 5160
rect 444466 5148 444472 5160
rect 222988 5120 444472 5148
rect 222988 5108 222994 5120
rect 444466 5108 444472 5120
rect 444524 5108 444530 5160
rect 451274 5108 451280 5160
rect 451332 5148 451338 5160
rect 518526 5148 518532 5160
rect 451332 5120 518532 5148
rect 451332 5108 451338 5120
rect 518526 5108 518532 5120
rect 518584 5108 518590 5160
rect 73062 5040 73068 5092
rect 73120 5080 73126 5092
rect 172514 5080 172520 5092
rect 73120 5052 172520 5080
rect 73120 5040 73126 5052
rect 172514 5040 172520 5052
rect 172572 5040 172578 5092
rect 219342 5040 219348 5092
rect 219400 5080 219406 5092
rect 443178 5080 443184 5092
rect 219400 5052 443184 5080
rect 219400 5040 219406 5052
rect 443178 5040 443184 5052
rect 443236 5040 443242 5092
rect 447870 5040 447876 5092
rect 447928 5080 447934 5092
rect 517698 5080 517704 5092
rect 447928 5052 517704 5080
rect 447928 5040 447934 5052
rect 517698 5040 517704 5052
rect 517756 5040 517762 5092
rect 30282 4972 30288 5024
rect 30340 5012 30346 5024
rect 140866 5012 140872 5024
rect 30340 4984 140872 5012
rect 30340 4972 30346 4984
rect 140866 4972 140872 4984
rect 140924 4972 140930 5024
rect 215846 4972 215852 5024
rect 215904 5012 215910 5024
rect 441706 5012 441712 5024
rect 215904 4984 441712 5012
rect 215904 4972 215910 4984
rect 441706 4972 441712 4984
rect 441764 4972 441770 5024
rect 444190 4972 444196 5024
rect 444248 5012 444254 5024
rect 516318 5012 516324 5024
rect 444248 4984 516324 5012
rect 444248 4972 444254 4984
rect 516318 4972 516324 4984
rect 516376 4972 516382 5024
rect 26694 4904 26700 4956
rect 26752 4944 26758 4956
rect 138106 4944 138112 4956
rect 26752 4916 138112 4944
rect 26752 4904 26758 4916
rect 138106 4904 138112 4916
rect 138164 4904 138170 4956
rect 183833 4947 183891 4953
rect 183833 4913 183845 4947
rect 183879 4944 183891 4947
rect 416774 4944 416780 4956
rect 183879 4916 416780 4944
rect 183879 4913 183891 4916
rect 183833 4907 183891 4913
rect 416774 4904 416780 4916
rect 416832 4904 416838 4956
rect 426342 4904 426348 4956
rect 426400 4944 426406 4956
rect 510890 4944 510896 4956
rect 426400 4916 510896 4944
rect 426400 4904 426406 4916
rect 510890 4904 510896 4916
rect 510948 4904 510954 4956
rect 17218 4836 17224 4888
rect 17276 4876 17282 4888
rect 131206 4876 131212 4888
rect 17276 4848 131212 4876
rect 17276 4836 17282 4848
rect 131206 4836 131212 4848
rect 131264 4836 131270 4888
rect 208670 4836 208676 4888
rect 208728 4876 208734 4888
rect 440418 4876 440424 4888
rect 208728 4848 440424 4876
rect 208728 4836 208734 4848
rect 440418 4836 440424 4848
rect 440476 4836 440482 4888
rect 440602 4836 440608 4888
rect 440660 4876 440666 4888
rect 515122 4876 515128 4888
rect 440660 4848 515128 4876
rect 440660 4836 440666 4848
rect 515122 4836 515128 4848
rect 515180 4836 515186 4888
rect 21910 4768 21916 4820
rect 21968 4808 21974 4820
rect 135346 4808 135352 4820
rect 21968 4780 135352 4808
rect 21968 4768 21974 4780
rect 135346 4768 135352 4780
rect 135404 4768 135410 4820
rect 197998 4768 198004 4820
rect 198056 4808 198062 4820
rect 436830 4808 436836 4820
rect 198056 4780 436836 4808
rect 198056 4768 198062 4780
rect 436830 4768 436836 4780
rect 436888 4768 436894 4820
rect 437014 4768 437020 4820
rect 437072 4808 437078 4820
rect 513558 4808 513564 4820
rect 437072 4780 513564 4808
rect 437072 4768 437078 4780
rect 513558 4768 513564 4780
rect 513616 4768 513622 4820
rect 94498 4700 94504 4752
rect 94556 4740 94562 4752
rect 187694 4740 187700 4752
rect 94556 4712 187700 4740
rect 94556 4700 94562 4712
rect 187694 4700 187700 4712
rect 187752 4700 187758 4752
rect 244366 4700 244372 4752
rect 244424 4740 244430 4752
rect 451826 4740 451832 4752
rect 244424 4712 451832 4740
rect 244424 4700 244430 4712
rect 451826 4700 451832 4712
rect 451884 4700 451890 4752
rect 472710 4700 472716 4752
rect 472768 4740 472774 4752
rect 524598 4740 524604 4752
rect 472768 4712 524604 4740
rect 472768 4700 472774 4712
rect 524598 4700 524604 4712
rect 524656 4700 524662 4752
rect 98086 4632 98092 4684
rect 98144 4672 98150 4684
rect 190454 4672 190460 4684
rect 98144 4644 190460 4672
rect 98144 4632 98150 4644
rect 190454 4632 190460 4644
rect 190512 4632 190518 4684
rect 247954 4632 247960 4684
rect 248012 4672 248018 4684
rect 452930 4672 452936 4684
rect 248012 4644 452936 4672
rect 248012 4632 248018 4644
rect 452930 4632 452936 4644
rect 452988 4632 452994 4684
rect 476298 4632 476304 4684
rect 476356 4672 476362 4684
rect 525978 4672 525984 4684
rect 476356 4644 525984 4672
rect 476356 4632 476362 4644
rect 525978 4632 525984 4644
rect 526036 4632 526042 4684
rect 101582 4564 101588 4616
rect 101640 4604 101646 4616
rect 193214 4604 193220 4616
rect 101640 4576 193220 4604
rect 101640 4564 101646 4576
rect 193214 4564 193220 4576
rect 193272 4564 193278 4616
rect 251450 4564 251456 4616
rect 251508 4604 251514 4616
rect 454126 4604 454132 4616
rect 251508 4576 454132 4604
rect 251508 4564 251514 4576
rect 454126 4564 454132 4576
rect 454184 4564 454190 4616
rect 479886 4564 479892 4616
rect 479944 4604 479950 4616
rect 527266 4604 527272 4616
rect 479944 4576 527272 4604
rect 479944 4564 479950 4576
rect 527266 4564 527272 4576
rect 527324 4564 527330 4616
rect 108758 4496 108764 4548
rect 108816 4536 108822 4548
rect 198734 4536 198740 4548
rect 108816 4508 198740 4536
rect 108816 4496 108822 4508
rect 198734 4496 198740 4508
rect 198792 4496 198798 4548
rect 255038 4496 255044 4548
rect 255096 4536 255102 4548
rect 455414 4536 455420 4548
rect 255096 4508 455420 4536
rect 255096 4496 255102 4508
rect 455414 4496 455420 4508
rect 455472 4496 455478 4548
rect 484578 4496 484584 4548
rect 484636 4536 484642 4548
rect 528738 4536 528744 4548
rect 484636 4508 528744 4536
rect 484636 4496 484642 4508
rect 528738 4496 528744 4508
rect 528796 4496 528802 4548
rect 105170 4428 105176 4480
rect 105228 4468 105234 4480
rect 195974 4468 195980 4480
rect 105228 4440 195980 4468
rect 105228 4428 105234 4440
rect 195974 4428 195980 4440
rect 196032 4428 196038 4480
rect 291930 4428 291936 4480
rect 291988 4468 291994 4480
rect 466730 4468 466736 4480
rect 291988 4440 466736 4468
rect 291988 4428 291994 4440
rect 466730 4428 466736 4440
rect 466788 4428 466794 4480
rect 488166 4428 488172 4480
rect 488224 4468 488230 4480
rect 530118 4468 530124 4480
rect 488224 4440 530124 4468
rect 488224 4428 488230 4440
rect 530118 4428 530124 4440
rect 530176 4428 530182 4480
rect 112346 4360 112352 4412
rect 112404 4400 112410 4412
rect 201402 4400 201408 4412
rect 112404 4372 201408 4400
rect 112404 4360 112410 4372
rect 201402 4360 201408 4372
rect 201460 4360 201466 4412
rect 354950 4360 354956 4412
rect 355008 4400 355014 4412
rect 487246 4400 487252 4412
rect 355008 4372 487252 4400
rect 355008 4360 355014 4372
rect 487246 4360 487252 4372
rect 487304 4360 487310 4412
rect 491754 4360 491760 4412
rect 491812 4400 491818 4412
rect 531498 4400 531504 4412
rect 491812 4372 531504 4400
rect 491812 4360 491818 4372
rect 531498 4360 531504 4372
rect 531556 4360 531562 4412
rect 119430 4292 119436 4344
rect 119488 4332 119494 4344
rect 122926 4332 122932 4344
rect 119488 4304 122932 4332
rect 119488 4292 119494 4304
rect 122926 4292 122932 4304
rect 122984 4292 122990 4344
rect 123018 4292 123024 4344
rect 123076 4332 123082 4344
rect 125597 4335 125655 4341
rect 125597 4332 125609 4335
rect 123076 4304 125609 4332
rect 123076 4292 123082 4304
rect 125597 4301 125609 4304
rect 125643 4301 125655 4335
rect 125597 4295 125655 4301
rect 125686 4292 125692 4344
rect 125744 4332 125750 4344
rect 206002 4332 206008 4344
rect 125744 4304 206008 4332
rect 125744 4292 125750 4304
rect 206002 4292 206008 4304
rect 206060 4292 206066 4344
rect 373994 4292 374000 4344
rect 374052 4332 374058 4344
rect 492858 4332 492864 4344
rect 374052 4304 492864 4332
rect 374052 4292 374058 4304
rect 492858 4292 492864 4304
rect 492916 4292 492922 4344
rect 508406 4292 508412 4344
rect 508464 4332 508470 4344
rect 537018 4332 537024 4344
rect 508464 4304 537024 4332
rect 508464 4292 508470 4304
rect 537018 4292 537024 4304
rect 537076 4292 537082 4344
rect 115934 4224 115940 4276
rect 115992 4264 115998 4276
rect 203058 4264 203064 4276
rect 115992 4236 203064 4264
rect 115992 4224 115998 4236
rect 203058 4224 203064 4236
rect 203116 4224 203122 4276
rect 429930 4224 429936 4276
rect 429988 4264 429994 4276
rect 510706 4264 510712 4276
rect 429988 4236 510712 4264
rect 429988 4224 429994 4236
rect 510706 4224 510712 4236
rect 510764 4224 510770 4276
rect 93857 4199 93915 4205
rect 93857 4165 93869 4199
rect 93903 4196 93915 4199
rect 103425 4199 103483 4205
rect 103425 4196 103437 4199
rect 93903 4168 103437 4196
rect 93903 4165 93915 4168
rect 93857 4159 93915 4165
rect 103425 4165 103437 4168
rect 103471 4165 103483 4199
rect 103425 4159 103483 4165
rect 113177 4199 113235 4205
rect 113177 4165 113189 4199
rect 113223 4196 113235 4199
rect 125505 4199 125563 4205
rect 125505 4196 125517 4199
rect 113223 4168 125517 4196
rect 113223 4165 113235 4168
rect 113177 4159 113235 4165
rect 125505 4165 125517 4168
rect 125551 4165 125563 4199
rect 125505 4159 125563 4165
rect 125597 4199 125655 4205
rect 125597 4165 125609 4199
rect 125643 4196 125655 4199
rect 208854 4196 208860 4208
rect 125643 4168 208860 4196
rect 125643 4165 125655 4168
rect 125597 4159 125655 4165
rect 208854 4156 208860 4168
rect 208912 4156 208918 4208
rect 383286 4156 383292 4208
rect 383344 4196 383350 4208
rect 383562 4196 383568 4208
rect 383344 4168 383568 4196
rect 383344 4156 383350 4168
rect 383562 4156 383568 4168
rect 383620 4156 383626 4208
rect 418062 4156 418068 4208
rect 418120 4196 418126 4208
rect 420822 4196 420828 4208
rect 418120 4168 420828 4196
rect 418120 4156 418126 4168
rect 420822 4156 420828 4168
rect 420880 4156 420886 4208
rect 433518 4156 433524 4208
rect 433576 4196 433582 4208
rect 512086 4196 512092 4208
rect 433576 4168 512092 4196
rect 433576 4156 433582 4168
rect 512086 4156 512092 4168
rect 512144 4156 512150 4208
rect 35897 4131 35955 4137
rect 35897 4097 35909 4131
rect 35943 4128 35955 4131
rect 45462 4128 45468 4140
rect 35943 4100 45468 4128
rect 35943 4097 35955 4100
rect 35897 4091 35955 4097
rect 45462 4088 45468 4100
rect 45520 4088 45526 4140
rect 45649 4131 45707 4137
rect 45649 4097 45661 4131
rect 45695 4128 45707 4131
rect 50338 4128 50344 4140
rect 45695 4100 50344 4128
rect 45695 4097 45707 4100
rect 45649 4091 45707 4097
rect 50338 4088 50344 4100
rect 50396 4088 50402 4140
rect 57606 4088 57612 4140
rect 57664 4128 57670 4140
rect 59998 4128 60004 4140
rect 57664 4100 60004 4128
rect 57664 4088 57670 4100
rect 59998 4088 60004 4100
rect 60056 4088 60062 4140
rect 60093 4131 60151 4137
rect 60093 4097 60105 4131
rect 60139 4128 60151 4131
rect 60139 4100 139624 4128
rect 60139 4097 60151 4100
rect 60093 4091 60151 4097
rect 19518 4020 19524 4072
rect 19576 4060 19582 4072
rect 46198 4060 46204 4072
rect 19576 4032 46204 4060
rect 19576 4020 19582 4032
rect 46198 4020 46204 4032
rect 46256 4020 46262 4072
rect 46934 4020 46940 4072
rect 46992 4060 46998 4072
rect 139489 4063 139547 4069
rect 139489 4060 139501 4063
rect 46992 4032 139501 4060
rect 46992 4020 46998 4032
rect 139489 4029 139501 4032
rect 139535 4029 139547 4063
rect 139596 4060 139624 4100
rect 139670 4088 139676 4140
rect 139728 4128 139734 4140
rect 140682 4128 140688 4140
rect 139728 4100 140688 4128
rect 139728 4088 139734 4100
rect 140682 4088 140688 4100
rect 140740 4088 140746 4140
rect 147677 4131 147735 4137
rect 147677 4097 147689 4131
rect 147723 4128 147735 4131
rect 147723 4100 157380 4128
rect 147723 4097 147735 4100
rect 147677 4091 147735 4097
rect 152458 4060 152464 4072
rect 139596 4032 152464 4060
rect 139489 4023 139547 4029
rect 152458 4020 152464 4032
rect 152516 4020 152522 4072
rect 43346 3952 43352 4004
rect 43404 3992 43410 4004
rect 150434 3992 150440 4004
rect 43404 3964 150440 3992
rect 43404 3952 43410 3964
rect 150434 3952 150440 3964
rect 150492 3952 150498 4004
rect 157352 3992 157380 4100
rect 172974 4088 172980 4140
rect 173032 4128 173038 4140
rect 173802 4128 173808 4140
rect 173032 4100 173808 4128
rect 173032 4088 173038 4100
rect 173802 4088 173808 4100
rect 173860 4088 173866 4140
rect 195241 4131 195299 4137
rect 195241 4097 195253 4131
rect 195287 4128 195299 4131
rect 220814 4128 220820 4140
rect 195287 4100 220820 4128
rect 195287 4097 195299 4100
rect 195241 4091 195299 4097
rect 220814 4088 220820 4100
rect 220872 4088 220878 4140
rect 360930 4088 360936 4140
rect 360988 4128 360994 4140
rect 361482 4128 361488 4140
rect 360988 4100 361488 4128
rect 360988 4088 360994 4100
rect 361482 4088 361488 4100
rect 361540 4088 361546 4140
rect 364518 4088 364524 4140
rect 364576 4128 364582 4140
rect 461578 4128 461584 4140
rect 364576 4100 461584 4128
rect 364576 4088 364582 4100
rect 461578 4088 461584 4100
rect 461636 4088 461642 4140
rect 500126 4088 500132 4140
rect 500184 4128 500190 4140
rect 502334 4128 502340 4140
rect 500184 4100 502340 4128
rect 500184 4088 500190 4100
rect 502334 4088 502340 4100
rect 502392 4088 502398 4140
rect 502518 4088 502524 4140
rect 502576 4128 502582 4140
rect 515493 4131 515551 4137
rect 515493 4128 515505 4131
rect 502576 4100 515505 4128
rect 502576 4088 502582 4100
rect 515493 4097 515505 4100
rect 515539 4097 515551 4131
rect 515493 4091 515551 4097
rect 515582 4088 515588 4140
rect 515640 4128 515646 4140
rect 516042 4128 516048 4140
rect 515640 4100 516048 4128
rect 515640 4088 515646 4100
rect 516042 4088 516048 4100
rect 516100 4088 516106 4140
rect 516778 4088 516784 4140
rect 516836 4128 516842 4140
rect 517422 4128 517428 4140
rect 516836 4100 517428 4128
rect 516836 4088 516842 4100
rect 517422 4088 517428 4100
rect 517480 4088 517486 4140
rect 518342 4128 518348 4140
rect 517532 4100 518348 4128
rect 157518 4020 157524 4072
rect 157576 4060 157582 4072
rect 204073 4063 204131 4069
rect 204073 4060 204085 4063
rect 157576 4032 204085 4060
rect 157576 4020 157582 4032
rect 204073 4029 204085 4032
rect 204119 4029 204131 4063
rect 204073 4023 204131 4029
rect 207474 4020 207480 4072
rect 207532 4060 207538 4072
rect 208302 4060 208308 4072
rect 207532 4032 208308 4060
rect 207532 4020 207538 4032
rect 208302 4020 208308 4032
rect 208360 4020 208366 4072
rect 225322 4020 225328 4072
rect 225380 4060 225386 4072
rect 275278 4060 275284 4072
rect 225380 4032 275284 4060
rect 225380 4020 225386 4032
rect 275278 4020 275284 4032
rect 275336 4020 275342 4072
rect 350258 4020 350264 4072
rect 350316 4060 350322 4072
rect 441617 4063 441675 4069
rect 441617 4060 441629 4063
rect 350316 4032 441629 4060
rect 350316 4020 350322 4032
rect 441617 4029 441629 4032
rect 441663 4029 441675 4063
rect 441617 4023 441675 4029
rect 492950 4020 492956 4072
rect 493008 4060 493014 4072
rect 502429 4063 502487 4069
rect 502429 4060 502441 4063
rect 493008 4032 502441 4060
rect 493008 4020 493014 4032
rect 502429 4029 502441 4032
rect 502475 4029 502487 4063
rect 502429 4023 502487 4029
rect 502613 4063 502671 4069
rect 502613 4029 502625 4063
rect 502659 4060 502671 4063
rect 517532 4060 517560 4100
rect 518342 4088 518348 4100
rect 518400 4088 518406 4140
rect 520274 4088 520280 4140
rect 520332 4128 520338 4140
rect 521562 4128 521568 4140
rect 520332 4100 521568 4128
rect 520332 4088 520338 4100
rect 521562 4088 521568 4100
rect 521620 4088 521626 4140
rect 523862 4088 523868 4140
rect 523920 4128 523926 4140
rect 524322 4128 524328 4140
rect 523920 4100 524328 4128
rect 523920 4088 523926 4100
rect 524322 4088 524328 4100
rect 524380 4088 524386 4140
rect 550082 4088 550088 4140
rect 550140 4128 550146 4140
rect 550542 4128 550548 4140
rect 550140 4100 550548 4128
rect 550140 4088 550146 4100
rect 550542 4088 550548 4100
rect 550600 4088 550606 4140
rect 551922 4088 551928 4140
rect 551980 4128 551986 4140
rect 552382 4128 552388 4140
rect 551980 4100 552388 4128
rect 551980 4088 551986 4100
rect 552382 4088 552388 4100
rect 552440 4088 552446 4140
rect 555418 4088 555424 4140
rect 555476 4128 555482 4140
rect 557166 4128 557172 4140
rect 555476 4100 557172 4128
rect 555476 4088 555482 4100
rect 557166 4088 557172 4100
rect 557224 4088 557230 4140
rect 558638 4088 558644 4140
rect 558696 4128 558702 4140
rect 572622 4128 572628 4140
rect 558696 4100 572628 4128
rect 558696 4088 558702 4100
rect 572622 4088 572628 4100
rect 572680 4088 572686 4140
rect 502659 4032 517560 4060
rect 502659 4029 502671 4032
rect 502613 4023 502671 4029
rect 517882 4020 517888 4072
rect 517940 4060 517946 4072
rect 523678 4060 523684 4072
rect 517940 4032 523684 4060
rect 517940 4020 517946 4032
rect 523678 4020 523684 4032
rect 523736 4020 523742 4072
rect 556982 4020 556988 4072
rect 557040 4060 557046 4072
rect 559558 4060 559564 4072
rect 557040 4032 559564 4060
rect 557040 4020 557046 4032
rect 559558 4020 559564 4032
rect 559616 4020 559622 4072
rect 570230 4060 570236 4072
rect 559760 4032 570236 4060
rect 162857 3995 162915 4001
rect 162857 3992 162869 3995
rect 157352 3964 162869 3992
rect 162857 3961 162869 3964
rect 162903 3961 162915 3995
rect 162857 3955 162915 3961
rect 168190 3952 168196 4004
rect 168248 3992 168254 4004
rect 225598 3992 225604 4004
rect 168248 3964 225604 3992
rect 168248 3952 168254 3964
rect 225598 3952 225604 3964
rect 225656 3952 225662 4004
rect 246758 3952 246764 4004
rect 246816 3992 246822 4004
rect 286318 3992 286324 4004
rect 246816 3964 286324 3992
rect 246816 3952 246822 3964
rect 286318 3952 286324 3964
rect 286376 3952 286382 4004
rect 343082 3952 343088 4004
rect 343140 3992 343146 4004
rect 451182 3992 451188 4004
rect 343140 3964 451188 3992
rect 343140 3952 343146 3964
rect 451182 3952 451188 3964
rect 451240 3952 451246 4004
rect 463513 3995 463571 4001
rect 463513 3992 463525 3995
rect 454052 3964 463525 3992
rect 42150 3884 42156 3936
rect 42208 3924 42214 3936
rect 149054 3924 149060 3936
rect 42208 3896 149060 3924
rect 42208 3884 42214 3896
rect 149054 3884 149060 3896
rect 149112 3884 149118 3936
rect 168009 3927 168067 3933
rect 168009 3893 168021 3927
rect 168055 3924 168067 3927
rect 232498 3924 232504 3936
rect 168055 3896 232504 3924
rect 168055 3893 168067 3896
rect 168009 3887 168067 3893
rect 232498 3884 232504 3896
rect 232556 3884 232562 3936
rect 257430 3884 257436 3936
rect 257488 3924 257494 3936
rect 300118 3924 300124 3936
rect 257488 3896 300124 3924
rect 257488 3884 257494 3896
rect 300118 3884 300124 3896
rect 300176 3884 300182 3936
rect 328822 3884 328828 3936
rect 328880 3924 328886 3936
rect 436094 3924 436100 3936
rect 328880 3896 436100 3924
rect 328880 3884 328886 3896
rect 436094 3884 436100 3896
rect 436152 3884 436158 3936
rect 439406 3884 439412 3936
rect 439464 3924 439470 3936
rect 443546 3924 443552 3936
rect 439464 3896 443552 3924
rect 439464 3884 439470 3896
rect 443546 3884 443552 3896
rect 443604 3884 443610 3936
rect 36170 3816 36176 3868
rect 36228 3856 36234 3868
rect 55217 3859 55275 3865
rect 55217 3856 55229 3859
rect 36228 3828 55229 3856
rect 36228 3816 36234 3828
rect 55217 3825 55229 3828
rect 55263 3825 55275 3859
rect 55217 3819 55275 3825
rect 64782 3816 64788 3868
rect 64840 3856 64846 3868
rect 66898 3856 66904 3868
rect 64840 3828 66904 3856
rect 64840 3816 64846 3828
rect 66898 3816 66904 3828
rect 66956 3816 66962 3868
rect 66993 3859 67051 3865
rect 66993 3825 67005 3859
rect 67039 3856 67051 3859
rect 74537 3859 74595 3865
rect 74537 3856 74549 3859
rect 67039 3828 74549 3856
rect 67039 3825 67051 3828
rect 66993 3819 67051 3825
rect 74537 3825 74549 3828
rect 74583 3825 74595 3859
rect 74537 3819 74595 3825
rect 84105 3859 84163 3865
rect 84105 3825 84117 3859
rect 84151 3856 84163 3859
rect 93857 3859 93915 3865
rect 93857 3856 93869 3859
rect 84151 3828 93869 3856
rect 84151 3825 84163 3828
rect 84105 3819 84163 3825
rect 93857 3825 93869 3828
rect 93903 3825 93915 3859
rect 93857 3819 93915 3825
rect 103425 3859 103483 3865
rect 103425 3825 103437 3859
rect 103471 3856 103483 3859
rect 113174 3856 113180 3868
rect 103471 3828 113180 3856
rect 103471 3825 103483 3828
rect 103425 3819 103483 3825
rect 113174 3816 113180 3828
rect 113232 3816 113238 3868
rect 118694 3816 118700 3868
rect 118752 3856 118758 3868
rect 130105 3859 130163 3865
rect 130105 3856 130117 3859
rect 118752 3828 130117 3856
rect 118752 3816 118758 3828
rect 130105 3825 130117 3828
rect 130151 3825 130163 3859
rect 130105 3819 130163 3825
rect 130194 3816 130200 3868
rect 130252 3856 130258 3868
rect 131022 3856 131028 3868
rect 130252 3828 131028 3856
rect 130252 3816 130258 3828
rect 131022 3816 131028 3828
rect 131080 3816 131086 3868
rect 133141 3859 133199 3865
rect 133141 3825 133153 3859
rect 133187 3856 133199 3859
rect 142801 3859 142859 3865
rect 133187 3828 138704 3856
rect 133187 3825 133199 3828
rect 133141 3819 133199 3825
rect 11238 3748 11244 3800
rect 11296 3788 11302 3800
rect 31018 3788 31024 3800
rect 11296 3760 31024 3788
rect 11296 3748 11302 3760
rect 31018 3748 31024 3760
rect 31076 3748 31082 3800
rect 34974 3748 34980 3800
rect 35032 3788 35038 3800
rect 138569 3791 138627 3797
rect 138569 3788 138581 3791
rect 35032 3760 138581 3788
rect 35032 3748 35038 3760
rect 138569 3757 138581 3760
rect 138615 3757 138627 3791
rect 138676 3788 138704 3828
rect 142801 3825 142813 3859
rect 142847 3856 142859 3859
rect 147677 3859 147735 3865
rect 147677 3856 147689 3859
rect 142847 3828 147689 3856
rect 142847 3825 142859 3828
rect 142801 3819 142859 3825
rect 147677 3825 147689 3828
rect 147723 3825 147735 3859
rect 147677 3819 147735 3825
rect 162857 3859 162915 3865
rect 162857 3825 162869 3859
rect 162903 3856 162915 3859
rect 166905 3859 166963 3865
rect 166905 3856 166917 3859
rect 162903 3828 166917 3856
rect 162903 3825 162915 3828
rect 162857 3819 162915 3825
rect 166905 3825 166917 3828
rect 166951 3825 166963 3859
rect 166905 3819 166963 3825
rect 166997 3859 167055 3865
rect 166997 3825 167009 3859
rect 167043 3856 167055 3859
rect 167043 3828 180656 3856
rect 167043 3825 167055 3828
rect 166997 3819 167055 3825
rect 139394 3788 139400 3800
rect 138676 3760 139400 3788
rect 138569 3751 138627 3757
rect 139394 3748 139400 3760
rect 139452 3748 139458 3800
rect 139489 3791 139547 3797
rect 139489 3757 139501 3791
rect 139535 3788 139547 3791
rect 153194 3788 153200 3800
rect 139535 3760 153200 3788
rect 139535 3757 139547 3760
rect 139489 3751 139547 3757
rect 153194 3748 153200 3760
rect 153252 3748 153258 3800
rect 180628 3788 180656 3828
rect 184750 3816 184756 3868
rect 184808 3856 184814 3868
rect 195241 3859 195299 3865
rect 195241 3856 195253 3859
rect 184808 3828 195253 3856
rect 184808 3816 184814 3828
rect 195241 3825 195253 3828
rect 195287 3825 195299 3859
rect 195241 3819 195299 3825
rect 195333 3859 195391 3865
rect 195333 3825 195345 3859
rect 195379 3856 195391 3859
rect 268378 3856 268384 3868
rect 195379 3828 268384 3856
rect 195379 3825 195391 3828
rect 195333 3819 195391 3825
rect 268378 3816 268384 3828
rect 268436 3816 268442 3868
rect 331214 3816 331220 3868
rect 331272 3856 331278 3868
rect 332410 3856 332416 3868
rect 331272 3828 332416 3856
rect 331272 3816 331278 3828
rect 332410 3816 332416 3828
rect 332468 3816 332474 3868
rect 335906 3816 335912 3868
rect 335964 3856 335970 3868
rect 446214 3856 446220 3868
rect 335964 3828 446220 3856
rect 335964 3816 335970 3828
rect 446214 3816 446220 3828
rect 446272 3816 446278 3868
rect 453945 3859 454003 3865
rect 453945 3825 453957 3859
rect 453991 3856 454003 3859
rect 454052 3856 454080 3964
rect 463513 3961 463525 3964
rect 463559 3961 463571 3995
rect 463513 3955 463571 3961
rect 463697 3995 463755 4001
rect 463697 3961 463709 3995
rect 463743 3992 463755 3995
rect 473265 3995 473323 4001
rect 473265 3992 473277 3995
rect 463743 3964 473277 3992
rect 463743 3961 463755 3964
rect 463697 3955 463755 3961
rect 473265 3961 473277 3964
rect 473311 3961 473323 3995
rect 473265 3955 473323 3961
rect 478690 3952 478696 4004
rect 478748 3992 478754 4004
rect 502521 3995 502579 4001
rect 502521 3992 502533 3995
rect 478748 3964 502533 3992
rect 478748 3952 478754 3964
rect 502521 3961 502533 3964
rect 502567 3961 502579 3995
rect 502521 3955 502579 3961
rect 502705 3995 502763 4001
rect 502705 3961 502717 3995
rect 502751 3992 502763 3995
rect 527358 3992 527364 4004
rect 502751 3964 527364 3992
rect 502751 3961 502763 3964
rect 502705 3955 502763 3961
rect 527358 3952 527364 3964
rect 527416 3952 527422 4004
rect 555510 3952 555516 4004
rect 555568 3992 555574 4004
rect 558362 3992 558368 4004
rect 555568 3964 558368 3992
rect 555568 3952 555574 3964
rect 558362 3952 558368 3964
rect 558420 3952 558426 4004
rect 471514 3884 471520 3936
rect 471572 3924 471578 3936
rect 502337 3927 502395 3933
rect 502337 3924 502349 3927
rect 471572 3896 502349 3924
rect 471572 3884 471578 3896
rect 502337 3893 502349 3896
rect 502383 3893 502395 3927
rect 502337 3887 502395 3893
rect 502613 3927 502671 3933
rect 502613 3893 502625 3927
rect 502659 3924 502671 3927
rect 524690 3924 524696 3936
rect 502659 3896 524696 3924
rect 502659 3893 502671 3896
rect 502613 3887 502671 3893
rect 524690 3884 524696 3896
rect 524748 3884 524754 3936
rect 557258 3884 557264 3936
rect 557316 3924 557322 3936
rect 559760 3924 559788 4032
rect 570230 4020 570236 4032
rect 570288 4020 570294 4072
rect 559837 3995 559895 4001
rect 559837 3961 559849 3995
rect 559883 3992 559895 3995
rect 573818 3992 573824 4004
rect 559883 3964 573824 3992
rect 559883 3961 559895 3964
rect 559837 3955 559895 3961
rect 573818 3952 573824 3964
rect 573876 3952 573882 4004
rect 557316 3896 559788 3924
rect 557316 3884 557322 3896
rect 560110 3884 560116 3936
rect 560168 3924 560174 3936
rect 576210 3924 576216 3936
rect 560168 3896 576216 3924
rect 560168 3884 560174 3896
rect 576210 3884 576216 3896
rect 576268 3884 576274 3936
rect 453991 3828 454080 3856
rect 453991 3825 454003 3828
rect 453945 3819 454003 3825
rect 460842 3816 460848 3868
rect 460900 3856 460906 3868
rect 483017 3859 483075 3865
rect 483017 3856 483029 3859
rect 460900 3828 483029 3856
rect 460900 3816 460906 3828
rect 483017 3825 483029 3828
rect 483063 3825 483075 3859
rect 483017 3819 483075 3825
rect 483201 3859 483259 3865
rect 483201 3825 483213 3859
rect 483247 3856 483259 3859
rect 514018 3856 514024 3868
rect 483247 3828 514024 3856
rect 483247 3825 483259 3828
rect 483201 3819 483259 3825
rect 514018 3816 514024 3828
rect 514076 3816 514082 3868
rect 515493 3859 515551 3865
rect 515493 3825 515505 3859
rect 515539 3856 515551 3859
rect 519722 3856 519728 3868
rect 515539 3828 519728 3856
rect 515539 3825 515551 3828
rect 515493 3819 515551 3825
rect 519722 3816 519728 3828
rect 519780 3816 519786 3868
rect 545298 3816 545304 3868
rect 545356 3856 545362 3868
rect 546310 3856 546316 3868
rect 545356 3828 546316 3856
rect 545356 3816 545362 3828
rect 546310 3816 546316 3828
rect 546368 3816 546374 3868
rect 558730 3816 558736 3868
rect 558788 3856 558794 3868
rect 575014 3856 575020 3868
rect 558788 3828 575020 3856
rect 558788 3816 558794 3828
rect 575014 3816 575020 3828
rect 575072 3816 575078 3868
rect 183833 3791 183891 3797
rect 183833 3788 183845 3791
rect 180628 3760 183845 3788
rect 183833 3757 183845 3760
rect 183879 3757 183891 3791
rect 183833 3751 183891 3757
rect 187234 3748 187240 3800
rect 187292 3788 187298 3800
rect 261478 3788 261484 3800
rect 187292 3760 261484 3788
rect 187292 3748 187298 3760
rect 261478 3748 261484 3760
rect 261536 3748 261542 3800
rect 314470 3748 314476 3800
rect 314528 3788 314534 3800
rect 435358 3788 435364 3800
rect 314528 3760 435364 3788
rect 314528 3748 314534 3760
rect 435358 3748 435364 3760
rect 435416 3748 435422 3800
rect 441617 3791 441675 3797
rect 441617 3757 441629 3791
rect 441663 3788 441675 3791
rect 452654 3788 452660 3800
rect 441663 3760 452660 3788
rect 441663 3757 441675 3760
rect 441617 3751 441675 3757
rect 452654 3748 452660 3760
rect 452712 3748 452718 3800
rect 464430 3748 464436 3800
rect 464488 3788 464494 3800
rect 483109 3791 483167 3797
rect 483109 3788 483121 3791
rect 464488 3760 483121 3788
rect 464488 3748 464494 3760
rect 483109 3757 483121 3760
rect 483155 3757 483167 3791
rect 483109 3751 483167 3757
rect 483293 3791 483351 3797
rect 483293 3757 483305 3791
rect 483339 3788 483351 3791
rect 502429 3791 502487 3797
rect 502429 3788 502441 3791
rect 483339 3760 502441 3788
rect 483339 3757 483351 3760
rect 483293 3751 483351 3757
rect 502429 3757 502441 3760
rect 502475 3757 502487 3791
rect 502429 3751 502487 3757
rect 502613 3791 502671 3797
rect 502613 3757 502625 3791
rect 502659 3788 502671 3791
rect 523218 3788 523224 3800
rect 502659 3760 523224 3788
rect 502659 3757 502671 3760
rect 502613 3751 502671 3757
rect 523218 3748 523224 3760
rect 523276 3748 523282 3800
rect 559742 3748 559748 3800
rect 559800 3788 559806 3800
rect 577406 3788 577412 3800
rect 559800 3760 577412 3788
rect 559800 3748 559806 3760
rect 577406 3748 577412 3760
rect 577464 3748 577470 3800
rect 2866 3680 2872 3732
rect 2924 3720 2930 3732
rect 10318 3720 10324 3732
rect 2924 3692 10324 3720
rect 2924 3680 2930 3692
rect 10318 3680 10324 3692
rect 10376 3680 10382 3732
rect 14826 3680 14832 3732
rect 14884 3720 14890 3732
rect 28258 3720 28264 3732
rect 14884 3692 28264 3720
rect 14884 3680 14890 3692
rect 28258 3680 28264 3692
rect 28316 3680 28322 3732
rect 29086 3680 29092 3732
rect 29144 3720 29150 3732
rect 35897 3723 35955 3729
rect 35897 3720 35909 3723
rect 29144 3692 35909 3720
rect 29144 3680 29150 3692
rect 35897 3689 35909 3692
rect 35943 3689 35955 3723
rect 35897 3683 35955 3689
rect 45462 3680 45468 3732
rect 45520 3720 45526 3732
rect 55217 3723 55275 3729
rect 55217 3720 55229 3723
rect 45520 3692 55229 3720
rect 45520 3680 45526 3692
rect 55217 3689 55229 3692
rect 55263 3689 55275 3723
rect 55217 3683 55275 3689
rect 62301 3723 62359 3729
rect 62301 3689 62313 3723
rect 62347 3720 62359 3723
rect 74537 3723 74595 3729
rect 74537 3720 74549 3723
rect 62347 3692 74549 3720
rect 62347 3689 62359 3692
rect 62301 3683 62359 3689
rect 74537 3689 74549 3692
rect 74583 3689 74595 3723
rect 74537 3683 74595 3689
rect 84105 3723 84163 3729
rect 84105 3689 84117 3723
rect 84151 3720 84163 3723
rect 93857 3723 93915 3729
rect 93857 3720 93869 3723
rect 84151 3692 93869 3720
rect 84151 3689 84163 3692
rect 84105 3683 84163 3689
rect 93857 3689 93869 3692
rect 93903 3689 93915 3723
rect 93857 3683 93915 3689
rect 103425 3723 103483 3729
rect 103425 3689 103437 3723
rect 103471 3720 103483 3723
rect 113177 3723 113235 3729
rect 113177 3720 113189 3723
rect 103471 3692 113189 3720
rect 103471 3689 103483 3692
rect 103425 3683 103483 3689
rect 113177 3689 113189 3692
rect 113223 3689 113235 3723
rect 113177 3683 113235 3689
rect 120626 3680 120632 3732
rect 120684 3720 120690 3732
rect 121362 3720 121368 3732
rect 120684 3692 121368 3720
rect 120684 3680 120690 3692
rect 121362 3680 121368 3692
rect 121420 3680 121426 3732
rect 121822 3680 121828 3732
rect 121880 3720 121886 3732
rect 122742 3720 122748 3732
rect 121880 3692 122748 3720
rect 121880 3680 121886 3692
rect 122742 3680 122748 3692
rect 122800 3680 122806 3732
rect 124214 3680 124220 3732
rect 124272 3720 124278 3732
rect 125410 3720 125416 3732
rect 124272 3692 125416 3720
rect 124272 3680 124278 3692
rect 125410 3680 125416 3692
rect 125468 3680 125474 3732
rect 125505 3723 125563 3729
rect 125505 3689 125517 3723
rect 125551 3720 125563 3723
rect 130013 3723 130071 3729
rect 130013 3720 130025 3723
rect 125551 3692 130025 3720
rect 125551 3689 125563 3692
rect 125505 3683 125563 3689
rect 130013 3689 130025 3692
rect 130059 3689 130071 3723
rect 130013 3683 130071 3689
rect 130105 3723 130163 3729
rect 130105 3689 130117 3723
rect 130151 3720 130163 3723
rect 144914 3720 144920 3732
rect 130151 3692 144920 3720
rect 130151 3689 130163 3692
rect 130105 3683 130163 3689
rect 144914 3680 144920 3692
rect 144972 3680 144978 3732
rect 176470 3680 176476 3732
rect 176528 3720 176534 3732
rect 250438 3720 250444 3732
rect 176528 3692 250444 3720
rect 176528 3680 176534 3692
rect 250438 3680 250444 3692
rect 250496 3680 250502 3732
rect 264606 3680 264612 3732
rect 264664 3720 264670 3732
rect 318058 3720 318064 3732
rect 264664 3692 318064 3720
rect 264664 3680 264670 3692
rect 318058 3680 318064 3692
rect 318116 3680 318122 3732
rect 321646 3680 321652 3732
rect 321704 3720 321710 3732
rect 445294 3720 445300 3732
rect 321704 3692 445300 3720
rect 321704 3680 321710 3692
rect 445294 3680 445300 3692
rect 445352 3680 445358 3732
rect 457254 3680 457260 3732
rect 457312 3720 457318 3732
rect 483017 3723 483075 3729
rect 483017 3720 483029 3723
rect 457312 3692 483029 3720
rect 457312 3680 457318 3692
rect 483017 3689 483029 3692
rect 483063 3689 483075 3723
rect 483017 3683 483075 3689
rect 483201 3723 483259 3729
rect 483201 3689 483213 3723
rect 483247 3720 483259 3723
rect 520550 3720 520556 3732
rect 483247 3692 502472 3720
rect 483247 3689 483259 3692
rect 483201 3683 483259 3689
rect 10042 3612 10048 3664
rect 10100 3652 10106 3664
rect 25498 3652 25504 3664
rect 10100 3624 25504 3652
rect 10100 3612 10106 3624
rect 25498 3612 25504 3624
rect 25556 3612 25562 3664
rect 27890 3612 27896 3664
rect 27948 3652 27954 3664
rect 133141 3655 133199 3661
rect 133141 3652 133153 3655
rect 27948 3624 133153 3652
rect 27948 3612 27954 3624
rect 133141 3621 133153 3624
rect 133187 3621 133199 3655
rect 133141 3615 133199 3621
rect 133230 3612 133236 3664
rect 133288 3652 133294 3664
rect 136634 3652 136640 3664
rect 133288 3624 136640 3652
rect 133288 3612 133294 3624
rect 136634 3612 136640 3624
rect 136692 3612 136698 3664
rect 137278 3612 137284 3664
rect 137336 3652 137342 3664
rect 142801 3655 142859 3661
rect 142801 3652 142813 3655
rect 137336 3624 142813 3652
rect 137336 3612 137342 3624
rect 142801 3621 142813 3624
rect 142847 3621 142859 3655
rect 142801 3615 142859 3621
rect 169386 3612 169392 3664
rect 169444 3652 169450 3664
rect 182269 3655 182327 3661
rect 182269 3652 182281 3655
rect 169444 3624 182281 3652
rect 169444 3612 169450 3624
rect 182269 3621 182281 3624
rect 182315 3621 182327 3655
rect 182269 3615 182327 3621
rect 182545 3655 182603 3661
rect 182545 3621 182557 3655
rect 182591 3652 182603 3655
rect 243538 3652 243544 3664
rect 182591 3624 243544 3652
rect 182591 3621 182603 3624
rect 182545 3615 182603 3621
rect 243538 3612 243544 3624
rect 243596 3612 243602 3664
rect 250346 3612 250352 3664
rect 250404 3652 250410 3664
rect 304258 3652 304264 3664
rect 250404 3624 304264 3652
rect 250404 3612 250410 3624
rect 304258 3612 304264 3624
rect 304316 3612 304322 3664
rect 307386 3612 307392 3664
rect 307444 3652 307450 3664
rect 430761 3655 430819 3661
rect 430761 3652 430773 3655
rect 307444 3624 430773 3652
rect 307444 3612 307450 3624
rect 430761 3621 430773 3624
rect 430807 3621 430819 3655
rect 433978 3652 433984 3664
rect 430761 3615 430819 3621
rect 430868 3624 433984 3652
rect 6454 3544 6460 3596
rect 6512 3584 6518 3596
rect 113450 3584 113456 3596
rect 6512 3556 113456 3584
rect 6512 3544 6518 3556
rect 113450 3544 113456 3556
rect 113508 3544 113514 3596
rect 113542 3544 113548 3596
rect 113600 3584 113606 3596
rect 114462 3584 114468 3596
rect 113600 3556 114468 3584
rect 113600 3544 113606 3556
rect 114462 3544 114468 3556
rect 114520 3544 114526 3596
rect 114738 3544 114744 3596
rect 114796 3584 114802 3596
rect 115842 3584 115848 3596
rect 114796 3556 115848 3584
rect 114796 3544 114802 3556
rect 115842 3544 115848 3556
rect 115900 3544 115906 3596
rect 116026 3544 116032 3596
rect 116084 3584 116090 3596
rect 117958 3584 117964 3596
rect 116084 3556 117964 3584
rect 116084 3544 116090 3556
rect 117958 3544 117964 3556
rect 118016 3544 118022 3596
rect 118234 3544 118240 3596
rect 118292 3584 118298 3596
rect 173158 3584 173164 3596
rect 118292 3556 173164 3584
rect 118292 3544 118298 3556
rect 173158 3544 173164 3556
rect 173216 3544 173222 3596
rect 180150 3544 180156 3596
rect 180208 3584 180214 3596
rect 182174 3584 182180 3596
rect 180208 3556 182180 3584
rect 180208 3544 180214 3556
rect 182174 3544 182180 3556
rect 182232 3544 182238 3596
rect 182634 3544 182640 3596
rect 182692 3584 182698 3596
rect 257338 3584 257344 3596
rect 182692 3556 257344 3584
rect 182692 3544 182698 3556
rect 257338 3544 257344 3556
rect 257396 3544 257402 3596
rect 268102 3544 268108 3596
rect 268160 3584 268166 3596
rect 292298 3584 292304 3596
rect 268160 3556 292304 3584
rect 268160 3544 268166 3556
rect 292298 3544 292304 3556
rect 292356 3544 292362 3596
rect 295518 3544 295524 3596
rect 295576 3584 295582 3596
rect 296622 3584 296628 3596
rect 295576 3556 296628 3584
rect 295576 3544 295582 3556
rect 296622 3544 296628 3556
rect 296680 3544 296686 3596
rect 296714 3544 296720 3596
rect 296772 3584 296778 3596
rect 298002 3584 298008 3596
rect 296772 3556 298008 3584
rect 296772 3544 296778 3556
rect 298002 3544 298008 3556
rect 298060 3544 298066 3596
rect 302602 3544 302608 3596
rect 302660 3584 302666 3596
rect 303522 3584 303528 3596
rect 302660 3556 303528 3584
rect 302660 3544 302666 3556
rect 303522 3544 303528 3556
rect 303580 3544 303586 3596
rect 303617 3587 303675 3593
rect 303617 3553 303629 3587
rect 303663 3584 303675 3587
rect 430868 3584 430896 3624
rect 433978 3612 433984 3624
rect 434036 3612 434042 3664
rect 442994 3612 443000 3664
rect 443052 3652 443058 3664
rect 463513 3655 463571 3661
rect 443052 3624 451964 3652
rect 443052 3612 443058 3624
rect 303663 3556 430896 3584
rect 430945 3587 431003 3593
rect 303663 3553 303675 3556
rect 303617 3547 303675 3553
rect 430945 3553 430957 3587
rect 430991 3584 431003 3587
rect 432601 3587 432659 3593
rect 432601 3584 432613 3587
rect 430991 3556 432613 3584
rect 430991 3553 431003 3556
rect 430945 3547 431003 3553
rect 432601 3553 432613 3556
rect 432647 3553 432659 3587
rect 439314 3584 439320 3596
rect 432601 3547 432659 3553
rect 432800 3556 439320 3584
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 10410 3516 10416 3528
rect 1728 3488 10416 3516
rect 1728 3476 1734 3488
rect 10410 3476 10416 3488
rect 10468 3476 10474 3528
rect 24302 3476 24308 3528
rect 24360 3516 24366 3528
rect 129826 3516 129832 3528
rect 24360 3488 129832 3516
rect 24360 3476 24366 3488
rect 129826 3476 129832 3488
rect 129884 3476 129890 3528
rect 135438 3516 135444 3528
rect 129936 3488 135444 3516
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 9122 3448 9128 3460
rect 624 3420 9128 3448
rect 624 3408 630 3420
rect 9122 3408 9128 3420
rect 9180 3408 9186 3460
rect 23106 3408 23112 3460
rect 23164 3448 23170 3460
rect 129936 3448 129964 3488
rect 135438 3476 135444 3488
rect 135496 3476 135502 3528
rect 138569 3519 138627 3525
rect 138569 3485 138581 3519
rect 138615 3516 138627 3519
rect 145006 3516 145012 3528
rect 138615 3488 145012 3516
rect 138615 3485 138627 3488
rect 138569 3479 138627 3485
rect 145006 3476 145012 3488
rect 145064 3476 145070 3528
rect 152734 3476 152740 3528
rect 152792 3516 152798 3528
rect 152792 3488 157380 3516
rect 152792 3476 152798 3488
rect 23164 3420 129964 3448
rect 130013 3451 130071 3457
rect 23164 3408 23170 3420
rect 130013 3417 130025 3451
rect 130059 3448 130071 3451
rect 140774 3448 140780 3460
rect 130059 3420 140780 3448
rect 130059 3417 130071 3420
rect 130013 3411 130071 3417
rect 140774 3408 140780 3420
rect 140832 3408 140838 3460
rect 7650 3340 7656 3392
rect 7708 3380 7714 3392
rect 11698 3380 11704 3392
rect 7708 3352 11704 3380
rect 7708 3340 7714 3352
rect 11698 3340 11704 3352
rect 11756 3340 11762 3392
rect 32674 3340 32680 3392
rect 32732 3380 32738 3392
rect 45649 3383 45707 3389
rect 45649 3380 45661 3383
rect 32732 3352 45661 3380
rect 32732 3340 32738 3352
rect 45649 3349 45661 3352
rect 45695 3349 45707 3383
rect 45649 3343 45707 3349
rect 45738 3340 45744 3392
rect 45796 3380 45802 3392
rect 46842 3380 46848 3392
rect 45796 3352 46848 3380
rect 45796 3340 45802 3352
rect 46842 3340 46848 3352
rect 46900 3340 46906 3392
rect 51626 3340 51632 3392
rect 51684 3380 51690 3392
rect 52362 3380 52368 3392
rect 51684 3352 52368 3380
rect 51684 3340 51690 3352
rect 52362 3340 52368 3352
rect 52420 3340 52426 3392
rect 52822 3340 52828 3392
rect 52880 3380 52886 3392
rect 53742 3380 53748 3392
rect 52880 3352 53748 3380
rect 52880 3340 52886 3352
rect 53742 3340 53748 3352
rect 53800 3340 53806 3392
rect 54018 3340 54024 3392
rect 54076 3380 54082 3392
rect 156598 3380 156604 3392
rect 54076 3352 156604 3380
rect 54076 3340 54082 3352
rect 156598 3340 156604 3352
rect 156656 3340 156662 3392
rect 157352 3380 157380 3488
rect 162302 3476 162308 3528
rect 162360 3516 162366 3528
rect 182269 3519 182327 3525
rect 182269 3516 182281 3519
rect 162360 3488 182281 3516
rect 162360 3476 162366 3488
rect 182269 3485 182281 3488
rect 182315 3485 182327 3519
rect 182269 3479 182327 3485
rect 182361 3519 182419 3525
rect 182361 3485 182373 3519
rect 182407 3516 182419 3519
rect 239398 3516 239404 3528
rect 182407 3488 239404 3516
rect 182407 3485 182419 3488
rect 182361 3479 182419 3485
rect 239398 3476 239404 3488
rect 239456 3476 239462 3528
rect 239582 3476 239588 3528
rect 239640 3516 239646 3528
rect 240042 3516 240048 3528
rect 239640 3488 240048 3516
rect 239640 3476 239646 3488
rect 240042 3476 240048 3488
rect 240100 3476 240106 3528
rect 258626 3476 258632 3528
rect 258684 3516 258690 3528
rect 259362 3516 259368 3528
rect 258684 3488 259368 3516
rect 258684 3476 258690 3488
rect 259362 3476 259368 3488
rect 259420 3476 259426 3528
rect 265802 3476 265808 3528
rect 265860 3516 265866 3528
rect 266262 3516 266268 3528
rect 265860 3488 266268 3516
rect 265860 3476 265866 3488
rect 266262 3476 266268 3488
rect 266320 3476 266326 3528
rect 271690 3476 271696 3528
rect 271748 3516 271754 3528
rect 406013 3519 406071 3525
rect 406013 3516 406025 3519
rect 271748 3488 406025 3516
rect 271748 3476 271754 3488
rect 406013 3485 406025 3488
rect 406059 3485 406071 3519
rect 406013 3479 406071 3485
rect 406102 3476 406108 3528
rect 406160 3516 406166 3528
rect 407022 3516 407028 3528
rect 406160 3488 407028 3516
rect 406160 3476 406166 3488
rect 407022 3476 407028 3488
rect 407080 3476 407086 3528
rect 407298 3476 407304 3528
rect 407356 3516 407362 3528
rect 408402 3516 408408 3528
rect 407356 3488 408408 3516
rect 407356 3476 407362 3488
rect 408402 3476 408408 3488
rect 408460 3476 408466 3528
rect 408494 3476 408500 3528
rect 408552 3516 408558 3528
rect 409782 3516 409788 3528
rect 408552 3488 409788 3516
rect 408552 3476 408558 3488
rect 409782 3476 409788 3488
rect 409840 3476 409846 3528
rect 413278 3476 413284 3528
rect 413336 3516 413342 3528
rect 413922 3516 413928 3528
rect 413336 3488 413928 3516
rect 413336 3476 413342 3488
rect 413922 3476 413928 3488
rect 413980 3476 413986 3528
rect 415670 3476 415676 3528
rect 415728 3516 415734 3528
rect 416682 3516 416688 3528
rect 415728 3488 416688 3516
rect 415728 3476 415734 3488
rect 416682 3476 416688 3488
rect 416740 3476 416746 3528
rect 416866 3476 416872 3528
rect 416924 3516 416930 3528
rect 417970 3516 417976 3528
rect 416924 3488 417976 3516
rect 416924 3476 416930 3488
rect 417970 3476 417976 3488
rect 418028 3476 418034 3528
rect 418065 3519 418123 3525
rect 418065 3485 418077 3519
rect 418111 3516 418123 3519
rect 421374 3516 421380 3528
rect 418111 3488 421380 3516
rect 418111 3485 418123 3488
rect 418065 3479 418123 3485
rect 421374 3476 421380 3488
rect 421432 3476 421438 3528
rect 421469 3519 421527 3525
rect 421469 3485 421481 3519
rect 421515 3516 421527 3519
rect 422665 3519 422723 3525
rect 422665 3516 422677 3519
rect 421515 3488 422677 3516
rect 421515 3485 421527 3488
rect 421469 3479 421527 3485
rect 422665 3485 422677 3488
rect 422711 3485 422723 3519
rect 422665 3479 422723 3485
rect 422754 3476 422760 3528
rect 422812 3516 422818 3528
rect 423582 3516 423588 3528
rect 422812 3488 423588 3516
rect 422812 3476 422818 3488
rect 423582 3476 423588 3488
rect 423640 3476 423646 3528
rect 423677 3519 423735 3525
rect 423677 3485 423689 3519
rect 423723 3516 423735 3519
rect 426434 3516 426440 3528
rect 423723 3488 426440 3516
rect 423723 3485 423735 3488
rect 423677 3479 423735 3485
rect 426434 3476 426440 3488
rect 426492 3476 426498 3528
rect 426526 3476 426532 3528
rect 426584 3516 426590 3528
rect 432800 3516 432828 3556
rect 439314 3544 439320 3556
rect 439372 3544 439378 3596
rect 446582 3544 446588 3596
rect 446640 3584 446646 3596
rect 447778 3584 447784 3596
rect 446640 3556 447784 3584
rect 446640 3544 446646 3556
rect 447778 3544 447784 3556
rect 447836 3544 447842 3596
rect 451936 3584 451964 3624
rect 463513 3621 463525 3655
rect 463559 3652 463571 3655
rect 463697 3655 463755 3661
rect 463697 3652 463709 3655
rect 463559 3624 463709 3652
rect 463559 3621 463571 3624
rect 463513 3615 463571 3621
rect 463697 3621 463709 3624
rect 463743 3621 463755 3655
rect 463697 3615 463755 3621
rect 473265 3655 473323 3661
rect 473265 3621 473277 3655
rect 473311 3652 473323 3655
rect 483109 3655 483167 3661
rect 483109 3652 483121 3655
rect 473311 3624 483121 3652
rect 473311 3621 473323 3624
rect 473265 3615 473323 3621
rect 483109 3621 483121 3624
rect 483155 3621 483167 3655
rect 483109 3615 483167 3621
rect 483293 3655 483351 3661
rect 483293 3621 483305 3655
rect 483339 3652 483351 3655
rect 492677 3655 492735 3661
rect 492677 3652 492689 3655
rect 483339 3624 492689 3652
rect 483339 3621 483351 3624
rect 483293 3615 483351 3621
rect 492677 3621 492689 3624
rect 492723 3621 492735 3655
rect 492677 3615 492735 3621
rect 502245 3655 502303 3661
rect 502245 3621 502257 3655
rect 502291 3652 502303 3655
rect 502337 3655 502395 3661
rect 502337 3652 502349 3655
rect 502291 3624 502349 3652
rect 502291 3621 502303 3624
rect 502245 3615 502303 3621
rect 502337 3621 502349 3624
rect 502383 3621 502395 3655
rect 502444 3652 502472 3692
rect 502536 3692 520556 3720
rect 502536 3652 502564 3692
rect 520550 3680 520556 3692
rect 520608 3680 520614 3732
rect 544102 3680 544108 3732
rect 544160 3720 544166 3732
rect 545022 3720 545028 3732
rect 544160 3692 545028 3720
rect 544160 3680 544166 3692
rect 545022 3680 545028 3692
rect 545080 3680 545086 3732
rect 558546 3680 558552 3732
rect 558604 3720 558610 3732
rect 559837 3723 559895 3729
rect 559837 3720 559849 3723
rect 558604 3692 559849 3720
rect 558604 3680 558610 3692
rect 559837 3689 559849 3692
rect 559883 3689 559895 3723
rect 559837 3683 559895 3689
rect 560202 3680 560208 3732
rect 560260 3720 560266 3732
rect 578602 3720 578608 3732
rect 560260 3692 578608 3720
rect 560260 3680 560266 3692
rect 578602 3680 578608 3692
rect 578660 3680 578666 3732
rect 502444 3624 502564 3652
rect 502613 3655 502671 3661
rect 502337 3615 502395 3621
rect 502613 3621 502625 3655
rect 502659 3652 502671 3655
rect 518158 3652 518164 3664
rect 502659 3624 518164 3652
rect 502659 3621 502671 3624
rect 502613 3615 502671 3621
rect 518158 3612 518164 3624
rect 518216 3612 518222 3664
rect 556890 3612 556896 3664
rect 556948 3652 556954 3664
rect 560754 3652 560760 3664
rect 556948 3624 560760 3652
rect 556948 3612 556954 3624
rect 560754 3612 560760 3624
rect 560812 3612 560818 3664
rect 561582 3612 561588 3664
rect 561640 3652 561646 3664
rect 582190 3652 582196 3664
rect 561640 3624 582196 3652
rect 561640 3612 561646 3624
rect 582190 3612 582196 3624
rect 582248 3612 582254 3664
rect 463789 3587 463847 3593
rect 463789 3584 463801 3587
rect 451936 3556 463801 3584
rect 463789 3553 463801 3556
rect 463835 3553 463847 3587
rect 463789 3547 463847 3553
rect 463881 3587 463939 3593
rect 463881 3553 463893 3587
rect 463927 3584 463939 3587
rect 473354 3584 473360 3596
rect 463927 3556 473360 3584
rect 463927 3553 463939 3556
rect 463881 3547 463939 3553
rect 473354 3544 473360 3556
rect 473412 3544 473418 3596
rect 473446 3544 473452 3596
rect 473504 3584 473510 3596
rect 483201 3587 483259 3593
rect 483201 3584 483213 3587
rect 473504 3556 483213 3584
rect 473504 3544 473510 3556
rect 483201 3553 483213 3556
rect 483247 3553 483259 3587
rect 483201 3547 483259 3553
rect 483385 3587 483443 3593
rect 483385 3553 483397 3587
rect 483431 3584 483443 3587
rect 516226 3584 516232 3596
rect 483431 3556 516232 3584
rect 483431 3553 483443 3556
rect 483385 3547 483443 3553
rect 516226 3544 516232 3556
rect 516284 3544 516290 3596
rect 526254 3544 526260 3596
rect 526312 3584 526318 3596
rect 533246 3584 533252 3596
rect 526312 3556 533252 3584
rect 526312 3544 526318 3556
rect 533246 3544 533252 3556
rect 533304 3544 533310 3596
rect 536926 3544 536932 3596
rect 536984 3584 536990 3596
rect 544378 3584 544384 3596
rect 536984 3556 544384 3584
rect 536984 3544 536990 3556
rect 544378 3544 544384 3556
rect 544436 3544 544442 3596
rect 556706 3544 556712 3596
rect 556764 3584 556770 3596
rect 561950 3584 561956 3596
rect 556764 3556 561956 3584
rect 556764 3544 556770 3556
rect 561950 3544 561956 3556
rect 562008 3544 562014 3596
rect 563698 3544 563704 3596
rect 563756 3584 563762 3596
rect 583386 3584 583392 3596
rect 563756 3556 583392 3584
rect 563756 3544 563762 3556
rect 583386 3544 583392 3556
rect 583444 3544 583450 3596
rect 426584 3488 432828 3516
rect 432877 3519 432935 3525
rect 426584 3476 426590 3488
rect 432877 3485 432889 3519
rect 432923 3516 432935 3519
rect 433426 3516 433432 3528
rect 432923 3488 433432 3516
rect 432923 3485 432935 3488
rect 432877 3479 432935 3485
rect 433426 3476 433432 3488
rect 433484 3476 433490 3528
rect 435818 3476 435824 3528
rect 435876 3516 435882 3528
rect 483017 3519 483075 3525
rect 483017 3516 483029 3519
rect 435876 3488 483029 3516
rect 435876 3476 435882 3488
rect 483017 3485 483029 3488
rect 483063 3485 483075 3519
rect 483017 3479 483075 3485
rect 483293 3519 483351 3525
rect 483293 3485 483305 3519
rect 483339 3516 483351 3519
rect 501141 3519 501199 3525
rect 501141 3516 501153 3519
rect 483339 3488 501153 3516
rect 483339 3485 483351 3488
rect 483293 3479 483351 3485
rect 501141 3485 501153 3488
rect 501187 3485 501199 3519
rect 501141 3479 501199 3485
rect 501230 3476 501236 3528
rect 501288 3516 501294 3528
rect 502242 3516 502248 3528
rect 501288 3488 502248 3516
rect 501288 3476 501294 3488
rect 502242 3476 502248 3488
rect 502300 3476 502306 3528
rect 502426 3476 502432 3528
rect 502484 3516 502490 3528
rect 503530 3516 503536 3528
rect 502484 3488 503536 3516
rect 502484 3476 502490 3488
rect 503530 3476 503536 3488
rect 503588 3476 503594 3528
rect 507210 3476 507216 3528
rect 507268 3516 507274 3528
rect 507762 3516 507768 3528
rect 507268 3488 507768 3516
rect 507268 3476 507274 3488
rect 507762 3476 507768 3488
rect 507820 3476 507826 3528
rect 509602 3476 509608 3528
rect 509660 3516 509666 3528
rect 510522 3516 510528 3528
rect 509660 3488 510528 3516
rect 509660 3476 509666 3488
rect 510522 3476 510528 3488
rect 510580 3476 510586 3528
rect 525058 3476 525064 3528
rect 525116 3516 525122 3528
rect 526346 3516 526352 3528
rect 525116 3488 526352 3516
rect 525116 3476 525122 3488
rect 526346 3476 526352 3488
rect 526404 3476 526410 3528
rect 526548 3488 528600 3516
rect 180705 3451 180763 3457
rect 180705 3417 180717 3451
rect 180751 3448 180763 3451
rect 182177 3451 182235 3457
rect 182177 3448 182189 3451
rect 180751 3420 182189 3448
rect 180751 3417 180763 3420
rect 180705 3411 180763 3417
rect 182177 3417 182189 3420
rect 182223 3417 182235 3451
rect 182177 3411 182235 3417
rect 193125 3451 193183 3457
rect 193125 3417 193137 3451
rect 193171 3448 193183 3451
rect 201497 3451 201555 3457
rect 201497 3448 201509 3451
rect 193171 3420 201509 3448
rect 193171 3417 193183 3420
rect 193125 3411 193183 3417
rect 201497 3417 201509 3420
rect 201543 3417 201555 3451
rect 246298 3448 246304 3460
rect 201497 3411 201555 3417
rect 203076 3420 246304 3448
rect 162857 3383 162915 3389
rect 162857 3380 162869 3383
rect 157352 3352 162869 3380
rect 162857 3349 162869 3352
rect 162903 3349 162915 3383
rect 162857 3343 162915 3349
rect 170582 3340 170588 3392
rect 170640 3380 170646 3392
rect 186225 3383 186283 3389
rect 186225 3380 186237 3383
rect 170640 3352 186237 3380
rect 170640 3340 170646 3352
rect 186225 3349 186237 3352
rect 186271 3349 186283 3383
rect 186225 3343 186283 3349
rect 186317 3383 186375 3389
rect 186317 3349 186329 3383
rect 186363 3380 186375 3383
rect 186363 3352 189120 3380
rect 186363 3349 186375 3352
rect 186317 3343 186375 3349
rect 16022 3272 16028 3324
rect 16080 3312 16086 3324
rect 50341 3315 50399 3321
rect 50341 3312 50353 3315
rect 16080 3284 50353 3312
rect 16080 3272 16086 3284
rect 50341 3281 50353 3284
rect 50387 3281 50399 3315
rect 50341 3275 50399 3281
rect 50522 3272 50528 3324
rect 50580 3312 50586 3324
rect 50580 3284 58756 3312
rect 50580 3272 50586 3284
rect 20714 3204 20720 3256
rect 20772 3244 20778 3256
rect 57977 3247 58035 3253
rect 57977 3244 57989 3247
rect 20772 3216 57989 3244
rect 20772 3204 20778 3216
rect 57977 3213 57989 3216
rect 58023 3213 58035 3247
rect 58728 3244 58756 3284
rect 58802 3272 58808 3324
rect 58860 3312 58866 3324
rect 59262 3312 59268 3324
rect 58860 3284 59268 3312
rect 58860 3272 58866 3284
rect 59262 3272 59268 3284
rect 59320 3272 59326 3324
rect 59998 3272 60004 3324
rect 60056 3312 60062 3324
rect 60642 3312 60648 3324
rect 60056 3284 60648 3312
rect 60056 3272 60062 3284
rect 60642 3272 60648 3284
rect 60700 3272 60706 3324
rect 61194 3272 61200 3324
rect 61252 3312 61258 3324
rect 159358 3312 159364 3324
rect 61252 3284 159364 3312
rect 61252 3272 61258 3284
rect 159358 3272 159364 3284
rect 159416 3272 159422 3324
rect 188430 3272 188436 3324
rect 188488 3312 188494 3324
rect 188982 3312 188988 3324
rect 188488 3284 188988 3312
rect 188488 3272 188494 3284
rect 188982 3272 188988 3284
rect 189040 3272 189046 3324
rect 189092 3312 189120 3352
rect 189626 3340 189632 3392
rect 189684 3380 189690 3392
rect 190362 3380 190368 3392
rect 189684 3352 190368 3380
rect 189684 3340 189690 3352
rect 190362 3340 190368 3352
rect 190420 3340 190426 3392
rect 190822 3340 190828 3392
rect 190880 3380 190886 3392
rect 191742 3380 191748 3392
rect 190880 3352 191748 3380
rect 190880 3340 190886 3352
rect 191742 3340 191748 3352
rect 191800 3340 191806 3392
rect 194410 3340 194416 3392
rect 194468 3380 194474 3392
rect 195333 3383 195391 3389
rect 195333 3380 195345 3383
rect 194468 3352 195345 3380
rect 194468 3340 194474 3352
rect 195333 3349 195345 3352
rect 195379 3349 195391 3383
rect 195333 3343 195391 3349
rect 195514 3312 195520 3324
rect 189092 3284 195520 3312
rect 195514 3272 195520 3284
rect 195572 3272 195578 3324
rect 201497 3315 201555 3321
rect 201497 3281 201509 3315
rect 201543 3312 201555 3315
rect 203076 3312 203104 3420
rect 246298 3408 246304 3420
rect 246356 3408 246362 3460
rect 419721 3451 419779 3457
rect 419721 3448 419733 3451
rect 277596 3420 419733 3448
rect 204073 3383 204131 3389
rect 204073 3349 204085 3383
rect 204119 3380 204131 3383
rect 214558 3380 214564 3392
rect 204119 3352 214564 3380
rect 204119 3349 204131 3352
rect 204073 3343 204131 3349
rect 214558 3340 214564 3352
rect 214616 3340 214622 3392
rect 218146 3340 218152 3392
rect 218204 3380 218210 3392
rect 219250 3380 219256 3392
rect 218204 3352 219256 3380
rect 218204 3340 218210 3352
rect 219250 3340 219256 3352
rect 219308 3340 219314 3392
rect 232498 3340 232504 3392
rect 232556 3380 232562 3392
rect 233142 3380 233148 3392
rect 232556 3352 233148 3380
rect 232556 3340 232562 3352
rect 233142 3340 233148 3352
rect 233200 3340 233206 3392
rect 275278 3340 275284 3392
rect 275336 3380 275342 3392
rect 277596 3380 277624 3420
rect 419721 3417 419733 3420
rect 419767 3417 419779 3451
rect 419721 3411 419779 3417
rect 432322 3408 432328 3460
rect 432380 3448 432386 3460
rect 473357 3451 473415 3457
rect 473357 3448 473369 3451
rect 432380 3420 473369 3448
rect 432380 3408 432386 3420
rect 473357 3417 473369 3420
rect 473403 3417 473415 3451
rect 473357 3411 473415 3417
rect 473541 3451 473599 3457
rect 473541 3417 473553 3451
rect 473587 3448 473599 3451
rect 509878 3448 509884 3460
rect 473587 3420 509884 3448
rect 473587 3417 473599 3420
rect 473541 3411 473599 3417
rect 509878 3408 509884 3420
rect 509936 3408 509942 3460
rect 510798 3408 510804 3460
rect 510856 3448 510862 3460
rect 520918 3448 520924 3460
rect 510856 3420 520924 3448
rect 510856 3408 510862 3420
rect 520918 3408 520924 3420
rect 520976 3408 520982 3460
rect 522666 3408 522672 3460
rect 522724 3448 522730 3460
rect 526548 3448 526576 3488
rect 522724 3420 526576 3448
rect 522724 3408 522730 3420
rect 527450 3408 527456 3460
rect 527508 3448 527514 3460
rect 528462 3448 528468 3460
rect 527508 3420 528468 3448
rect 527508 3408 527514 3420
rect 528462 3408 528468 3420
rect 528520 3408 528526 3460
rect 275336 3352 277624 3380
rect 275336 3340 275342 3352
rect 277670 3340 277676 3392
rect 277728 3380 277734 3392
rect 278682 3380 278688 3392
rect 277728 3352 278688 3380
rect 277728 3340 277734 3352
rect 278682 3340 278688 3352
rect 278740 3340 278746 3392
rect 284754 3340 284760 3392
rect 284812 3380 284818 3392
rect 285582 3380 285588 3392
rect 284812 3352 285588 3380
rect 284812 3340 284818 3352
rect 285582 3340 285588 3352
rect 285640 3340 285646 3392
rect 300302 3340 300308 3392
rect 300360 3380 300366 3392
rect 303617 3383 303675 3389
rect 303617 3380 303629 3383
rect 300360 3352 303629 3380
rect 300360 3340 300366 3352
rect 303617 3349 303629 3352
rect 303663 3349 303675 3383
rect 303617 3343 303675 3349
rect 309778 3340 309784 3392
rect 309836 3380 309842 3392
rect 310422 3380 310428 3392
rect 309836 3352 310428 3380
rect 309836 3340 309842 3352
rect 310422 3340 310428 3352
rect 310480 3340 310486 3392
rect 310974 3340 310980 3392
rect 311032 3380 311038 3392
rect 311802 3380 311808 3392
rect 311032 3352 311808 3380
rect 311032 3340 311038 3352
rect 311802 3340 311808 3352
rect 311860 3340 311866 3392
rect 313366 3340 313372 3392
rect 313424 3380 313430 3392
rect 314562 3380 314568 3392
rect 313424 3352 314568 3380
rect 313424 3340 313430 3352
rect 314562 3340 314568 3352
rect 314620 3340 314626 3392
rect 318058 3340 318064 3392
rect 318116 3380 318122 3392
rect 318702 3380 318708 3392
rect 318116 3352 318708 3380
rect 318116 3340 318122 3352
rect 318702 3340 318708 3352
rect 318760 3340 318766 3392
rect 320450 3340 320456 3392
rect 320508 3380 320514 3392
rect 321462 3380 321468 3392
rect 320508 3352 321468 3380
rect 320508 3340 320514 3352
rect 321462 3340 321468 3352
rect 321520 3340 321526 3392
rect 334710 3340 334716 3392
rect 334768 3380 334774 3392
rect 335262 3380 335268 3392
rect 334768 3352 335268 3380
rect 334768 3340 334774 3352
rect 335262 3340 335268 3352
rect 335320 3340 335326 3392
rect 338298 3340 338304 3392
rect 338356 3380 338362 3392
rect 339402 3380 339408 3392
rect 338356 3352 339408 3380
rect 338356 3340 338362 3352
rect 339402 3340 339408 3352
rect 339460 3340 339466 3392
rect 339494 3340 339500 3392
rect 339552 3380 339558 3392
rect 340782 3380 340788 3392
rect 339552 3352 340788 3380
rect 339552 3340 339558 3352
rect 340782 3340 340788 3352
rect 340840 3340 340846 3392
rect 345474 3340 345480 3392
rect 345532 3380 345538 3392
rect 346302 3380 346308 3392
rect 345532 3352 346308 3380
rect 345532 3340 345538 3352
rect 346302 3340 346308 3352
rect 346360 3340 346366 3392
rect 347866 3340 347872 3392
rect 347924 3380 347930 3392
rect 349062 3380 349068 3392
rect 347924 3352 349068 3380
rect 347924 3340 347930 3352
rect 349062 3340 349068 3352
rect 349120 3340 349126 3392
rect 351362 3340 351368 3392
rect 351420 3380 351426 3392
rect 351822 3380 351828 3392
rect 351420 3352 351828 3380
rect 351420 3340 351426 3352
rect 351822 3340 351828 3352
rect 351880 3340 351886 3392
rect 352558 3340 352564 3392
rect 352616 3380 352622 3392
rect 353202 3380 353208 3392
rect 352616 3352 353208 3380
rect 352616 3340 352622 3352
rect 353202 3340 353208 3352
rect 353260 3340 353266 3392
rect 353754 3340 353760 3392
rect 353812 3380 353818 3392
rect 354582 3380 354588 3392
rect 353812 3352 354588 3380
rect 353812 3340 353818 3352
rect 354582 3340 354588 3352
rect 354640 3340 354646 3392
rect 356146 3340 356152 3392
rect 356204 3380 356210 3392
rect 357342 3380 357348 3392
rect 356204 3352 357348 3380
rect 356204 3340 356210 3352
rect 357342 3340 357348 3352
rect 357400 3340 357406 3392
rect 360197 3383 360255 3389
rect 360197 3349 360209 3383
rect 360243 3380 360255 3383
rect 452746 3380 452752 3392
rect 360243 3352 452752 3380
rect 360243 3349 360255 3352
rect 360197 3343 360255 3349
rect 452746 3340 452752 3352
rect 452804 3340 452810 3392
rect 453666 3340 453672 3392
rect 453724 3380 453730 3392
rect 457438 3380 457444 3392
rect 453724 3352 457444 3380
rect 453724 3340 453730 3352
rect 457438 3340 457444 3352
rect 457496 3340 457502 3392
rect 467926 3340 467932 3392
rect 467984 3380 467990 3392
rect 469030 3380 469036 3392
rect 467984 3352 469036 3380
rect 467984 3340 467990 3352
rect 469030 3340 469036 3352
rect 469088 3340 469094 3392
rect 475102 3340 475108 3392
rect 475160 3380 475166 3392
rect 476022 3380 476028 3392
rect 475160 3352 476028 3380
rect 475160 3340 475166 3352
rect 476022 3340 476028 3352
rect 476080 3340 476086 3392
rect 477494 3340 477500 3392
rect 477552 3380 477558 3392
rect 478782 3380 478788 3392
rect 477552 3352 478788 3380
rect 477552 3340 477558 3352
rect 478782 3340 478788 3352
rect 478840 3340 478846 3392
rect 481082 3340 481088 3392
rect 481140 3380 481146 3392
rect 481542 3380 481548 3392
rect 481140 3352 481548 3380
rect 481140 3340 481146 3352
rect 481542 3340 481548 3352
rect 481600 3340 481606 3392
rect 482278 3340 482284 3392
rect 482336 3380 482342 3392
rect 482922 3380 482928 3392
rect 482336 3352 482928 3380
rect 482336 3340 482342 3352
rect 482922 3340 482928 3352
rect 482980 3340 482986 3392
rect 485774 3340 485780 3392
rect 485832 3380 485838 3392
rect 487062 3380 487068 3392
rect 485832 3352 487068 3380
rect 485832 3340 485838 3352
rect 487062 3340 487068 3352
rect 487120 3340 487126 3392
rect 489362 3340 489368 3392
rect 489420 3380 489426 3392
rect 489822 3380 489828 3392
rect 489420 3352 489828 3380
rect 489420 3340 489426 3352
rect 489822 3340 489828 3352
rect 489880 3340 489886 3392
rect 490558 3340 490564 3392
rect 490616 3380 490622 3392
rect 491202 3380 491208 3392
rect 490616 3352 491208 3380
rect 490616 3340 490622 3352
rect 491202 3340 491208 3352
rect 491260 3340 491266 3392
rect 498930 3340 498936 3392
rect 498988 3380 498994 3392
rect 499482 3380 499488 3392
rect 498988 3352 499488 3380
rect 498988 3340 498994 3352
rect 499482 3340 499488 3352
rect 499540 3340 499546 3392
rect 501141 3383 501199 3389
rect 501141 3349 501153 3383
rect 501187 3380 501199 3383
rect 511258 3380 511264 3392
rect 501187 3352 511264 3380
rect 501187 3349 501199 3352
rect 501141 3343 501199 3349
rect 511258 3340 511264 3352
rect 511316 3340 511322 3392
rect 514386 3340 514392 3392
rect 514444 3380 514450 3392
rect 522298 3380 522304 3392
rect 514444 3352 522304 3380
rect 514444 3340 514450 3352
rect 522298 3340 522304 3352
rect 522356 3340 522362 3392
rect 201543 3284 203104 3312
rect 201543 3281 201555 3284
rect 201497 3275 201555 3281
rect 282454 3272 282460 3324
rect 282512 3312 282518 3324
rect 364978 3312 364984 3324
rect 282512 3284 364984 3312
rect 282512 3272 282518 3284
rect 364978 3272 364984 3284
rect 365036 3272 365042 3324
rect 377582 3272 377588 3324
rect 377640 3312 377646 3324
rect 378042 3312 378048 3324
rect 377640 3284 378048 3312
rect 377640 3272 377646 3284
rect 378042 3272 378048 3284
rect 378100 3272 378106 3324
rect 381170 3272 381176 3324
rect 381228 3312 381234 3324
rect 382182 3312 382188 3324
rect 381228 3284 382188 3312
rect 381228 3272 381234 3284
rect 382182 3272 382188 3284
rect 382240 3272 382246 3324
rect 382366 3272 382372 3324
rect 382424 3312 382430 3324
rect 383286 3312 383292 3324
rect 382424 3284 383292 3312
rect 382424 3272 382430 3284
rect 383286 3272 383292 3284
rect 383344 3272 383350 3324
rect 383381 3315 383439 3321
rect 383381 3281 383393 3315
rect 383427 3312 383439 3315
rect 471882 3312 471888 3324
rect 383427 3284 471888 3312
rect 383427 3281 383439 3284
rect 383381 3275 383439 3281
rect 471882 3272 471888 3284
rect 471940 3272 471946 3324
rect 492677 3315 492735 3321
rect 492677 3281 492689 3315
rect 492723 3312 492735 3315
rect 502245 3315 502303 3321
rect 502245 3312 502257 3315
rect 492723 3284 502257 3312
rect 492723 3281 492735 3284
rect 492677 3275 492735 3281
rect 502245 3281 502257 3284
rect 502291 3281 502303 3315
rect 502245 3275 502303 3281
rect 521470 3272 521476 3324
rect 521528 3312 521534 3324
rect 524966 3312 524972 3324
rect 521528 3284 524972 3312
rect 521528 3272 521534 3284
rect 524966 3272 524972 3284
rect 525024 3272 525030 3324
rect 528572 3312 528600 3488
rect 528646 3476 528652 3528
rect 528704 3516 528710 3528
rect 529842 3516 529848 3528
rect 528704 3488 529848 3516
rect 528704 3476 528710 3488
rect 529842 3476 529848 3488
rect 529900 3476 529906 3528
rect 533430 3476 533436 3528
rect 533488 3516 533494 3528
rect 533982 3516 533988 3528
rect 533488 3488 533988 3516
rect 533488 3476 533494 3488
rect 533982 3476 533988 3488
rect 534040 3476 534046 3528
rect 534534 3476 534540 3528
rect 534592 3516 534598 3528
rect 535362 3516 535368 3528
rect 534592 3488 535368 3516
rect 534592 3476 534598 3488
rect 535362 3476 535368 3488
rect 535420 3476 535426 3528
rect 543918 3516 543924 3528
rect 538600 3488 543924 3516
rect 538600 3448 538628 3488
rect 543918 3476 543924 3488
rect 543976 3476 543982 3528
rect 563054 3476 563060 3528
rect 563112 3516 563118 3528
rect 564342 3516 564348 3528
rect 563112 3488 564348 3516
rect 563112 3476 563118 3488
rect 564342 3476 564348 3488
rect 564400 3476 564406 3528
rect 580994 3516 581000 3528
rect 564452 3488 581000 3516
rect 529860 3420 538628 3448
rect 529860 3392 529888 3420
rect 542906 3408 542912 3460
rect 542964 3448 542970 3460
rect 543642 3448 543648 3460
rect 542964 3420 543648 3448
rect 542964 3408 542970 3420
rect 543642 3408 543648 3420
rect 543700 3408 543706 3460
rect 561490 3408 561496 3460
rect 561548 3448 561554 3460
rect 564452 3448 564480 3488
rect 580994 3476 581000 3488
rect 581052 3476 581058 3528
rect 579798 3448 579804 3460
rect 561548 3420 564480 3448
rect 564544 3420 579804 3448
rect 561548 3408 561554 3420
rect 529842 3340 529848 3392
rect 529900 3340 529906 3392
rect 539318 3340 539324 3392
rect 539376 3380 539382 3392
rect 545758 3380 545764 3392
rect 539376 3352 545764 3380
rect 539376 3340 539382 3352
rect 545758 3340 545764 3352
rect 545816 3340 545822 3392
rect 546494 3340 546500 3392
rect 546552 3380 546558 3392
rect 547690 3380 547696 3392
rect 546552 3352 547696 3380
rect 546552 3340 546558 3352
rect 547690 3340 547696 3352
rect 547748 3340 547754 3392
rect 560018 3340 560024 3392
rect 560076 3380 560082 3392
rect 564544 3380 564572 3420
rect 579798 3408 579804 3420
rect 579856 3408 579862 3460
rect 560076 3352 564572 3380
rect 564621 3383 564679 3389
rect 560076 3340 560082 3352
rect 564621 3349 564633 3383
rect 564667 3380 564679 3383
rect 571426 3380 571432 3392
rect 564667 3352 571432 3380
rect 564667 3349 564679 3352
rect 564621 3343 564679 3349
rect 571426 3340 571432 3352
rect 571484 3340 571490 3392
rect 534718 3312 534724 3324
rect 528572 3284 534724 3312
rect 534718 3272 534724 3284
rect 534776 3272 534782 3324
rect 535730 3272 535736 3324
rect 535788 3312 535794 3324
rect 536742 3312 536748 3324
rect 535788 3284 536748 3312
rect 535788 3272 535794 3284
rect 536742 3272 536748 3284
rect 536800 3272 536806 3324
rect 557442 3272 557448 3324
rect 557500 3312 557506 3324
rect 569034 3312 569040 3324
rect 557500 3284 569040 3312
rect 557500 3272 557506 3284
rect 569034 3272 569040 3284
rect 569092 3272 569098 3324
rect 60093 3247 60151 3253
rect 60093 3244 60105 3247
rect 58728 3216 60105 3244
rect 57977 3207 58035 3213
rect 60093 3213 60105 3216
rect 60139 3213 60151 3247
rect 60093 3207 60151 3213
rect 68278 3204 68284 3256
rect 68336 3244 68342 3256
rect 162118 3244 162124 3256
rect 68336 3216 162124 3244
rect 68336 3204 68342 3216
rect 162118 3204 162124 3216
rect 162176 3204 162182 3256
rect 162857 3247 162915 3253
rect 162857 3213 162869 3247
rect 162903 3244 162915 3247
rect 171137 3247 171195 3253
rect 171137 3244 171149 3247
rect 162903 3216 171149 3244
rect 162903 3213 162915 3216
rect 162857 3207 162915 3213
rect 171137 3213 171149 3216
rect 171183 3213 171195 3247
rect 171137 3207 171195 3213
rect 181346 3204 181352 3256
rect 181404 3244 181410 3256
rect 186225 3247 186283 3253
rect 186225 3244 186237 3247
rect 181404 3216 186237 3244
rect 181404 3204 181410 3216
rect 186225 3213 186237 3216
rect 186271 3213 186283 3247
rect 186225 3207 186283 3213
rect 357342 3204 357348 3256
rect 357400 3244 357406 3256
rect 360197 3247 360255 3253
rect 360197 3244 360209 3247
rect 357400 3216 360209 3244
rect 357400 3204 357406 3216
rect 360197 3213 360209 3216
rect 360243 3213 360255 3247
rect 360197 3207 360255 3213
rect 387058 3204 387064 3256
rect 387116 3244 387122 3256
rect 387702 3244 387708 3256
rect 387116 3216 387708 3244
rect 387116 3204 387122 3216
rect 387702 3204 387708 3216
rect 387760 3204 387766 3256
rect 388254 3204 388260 3256
rect 388312 3244 388318 3256
rect 389082 3244 389088 3256
rect 388312 3216 389088 3244
rect 388312 3204 388318 3216
rect 389082 3204 389088 3216
rect 389140 3204 389146 3256
rect 389450 3204 389456 3256
rect 389508 3244 389514 3256
rect 390462 3244 390468 3256
rect 389508 3216 390468 3244
rect 389508 3204 389514 3216
rect 390462 3204 390468 3216
rect 390520 3204 390526 3256
rect 390557 3247 390615 3253
rect 390557 3213 390569 3247
rect 390603 3244 390615 3247
rect 476114 3244 476120 3256
rect 390603 3216 476120 3244
rect 390603 3213 390615 3216
rect 390557 3207 390615 3213
rect 476114 3204 476120 3216
rect 476172 3204 476178 3256
rect 541710 3204 541716 3256
rect 541768 3244 541774 3256
rect 548058 3244 548064 3256
rect 541768 3216 548064 3244
rect 541768 3204 541774 3216
rect 548058 3204 548064 3216
rect 548116 3204 548122 3256
rect 557350 3204 557356 3256
rect 557408 3244 557414 3256
rect 567838 3244 567844 3256
rect 557408 3216 567844 3244
rect 557408 3204 557414 3216
rect 567838 3204 567844 3216
rect 567896 3204 567902 3256
rect 5258 3136 5264 3188
rect 5316 3176 5322 3188
rect 68094 3176 68100 3188
rect 5316 3148 68100 3176
rect 5316 3136 5322 3148
rect 68094 3136 68100 3148
rect 68152 3136 68158 3188
rect 81434 3136 81440 3188
rect 81492 3176 81498 3188
rect 82722 3176 82728 3188
rect 81492 3148 82728 3176
rect 81492 3136 81498 3148
rect 82722 3136 82728 3148
rect 82780 3136 82786 3188
rect 163406 3176 163412 3188
rect 82832 3148 163412 3176
rect 39758 3068 39764 3120
rect 39816 3108 39822 3120
rect 53098 3108 53104 3120
rect 39816 3080 53104 3108
rect 39816 3068 39822 3080
rect 53098 3068 53104 3080
rect 53156 3068 53162 3120
rect 55214 3068 55220 3120
rect 55272 3108 55278 3120
rect 56502 3108 56508 3120
rect 55272 3080 56508 3108
rect 55272 3068 55278 3080
rect 56502 3068 56508 3080
rect 56560 3068 56566 3120
rect 57977 3111 58035 3117
rect 57977 3077 57989 3111
rect 58023 3108 58035 3111
rect 61378 3108 61384 3120
rect 58023 3080 61384 3108
rect 58023 3077 58035 3080
rect 57977 3071 58035 3077
rect 61378 3068 61384 3080
rect 61436 3068 61442 3120
rect 79042 3068 79048 3120
rect 79100 3108 79106 3120
rect 82078 3108 82084 3120
rect 79100 3080 82084 3108
rect 79100 3068 79106 3080
rect 82078 3068 82084 3080
rect 82136 3068 82142 3120
rect 82832 3108 82860 3148
rect 163406 3136 163412 3148
rect 163464 3136 163470 3188
rect 182177 3179 182235 3185
rect 182177 3145 182189 3179
rect 182223 3176 182235 3179
rect 193125 3179 193183 3185
rect 193125 3176 193137 3179
rect 182223 3148 193137 3176
rect 182223 3145 182235 3148
rect 182177 3139 182235 3145
rect 193125 3145 193137 3148
rect 193171 3145 193183 3179
rect 193125 3139 193183 3145
rect 327626 3136 327632 3188
rect 327684 3176 327690 3188
rect 328362 3176 328368 3188
rect 327684 3148 328368 3176
rect 327684 3136 327690 3148
rect 328362 3136 328368 3148
rect 328420 3136 328426 3188
rect 371602 3136 371608 3188
rect 371660 3176 371666 3188
rect 458542 3176 458548 3188
rect 371660 3148 458548 3176
rect 371660 3136 371666 3148
rect 458542 3136 458548 3148
rect 458600 3136 458606 3188
rect 556062 3136 556068 3188
rect 556120 3176 556126 3188
rect 566734 3176 566740 3188
rect 556120 3148 566740 3176
rect 556120 3136 556126 3148
rect 566734 3136 566740 3148
rect 566792 3136 566798 3188
rect 82280 3080 82860 3108
rect 50341 3043 50399 3049
rect 50341 3009 50353 3043
rect 50387 3040 50399 3043
rect 57238 3040 57244 3052
rect 50387 3012 57244 3040
rect 50387 3009 50399 3012
rect 50341 3003 50399 3009
rect 57238 3000 57244 3012
rect 57296 3000 57302 3052
rect 74537 3043 74595 3049
rect 74537 3009 74549 3043
rect 74583 3040 74595 3043
rect 74583 3012 75316 3040
rect 74583 3009 74595 3012
rect 74537 3003 74595 3009
rect 55217 2975 55275 2981
rect 55217 2941 55229 2975
rect 55263 2972 55275 2975
rect 62301 2975 62359 2981
rect 62301 2972 62313 2975
rect 55263 2944 62313 2972
rect 55263 2941 55275 2944
rect 55217 2935 55275 2941
rect 62301 2941 62313 2944
rect 62347 2941 62359 2975
rect 62301 2935 62359 2941
rect 62390 2932 62396 2984
rect 62448 2972 62454 2984
rect 63402 2972 63408 2984
rect 62448 2944 63408 2972
rect 62448 2932 62454 2944
rect 63402 2932 63408 2944
rect 63460 2932 63466 2984
rect 71866 2932 71872 2984
rect 71924 2972 71930 2984
rect 75178 2972 75184 2984
rect 71924 2944 75184 2972
rect 71924 2932 71930 2944
rect 75178 2932 75184 2944
rect 75236 2932 75242 2984
rect 75288 2972 75316 3012
rect 75454 3000 75460 3052
rect 75512 3040 75518 3052
rect 82280 3040 82308 3080
rect 84930 3068 84936 3120
rect 84988 3108 84994 3120
rect 85482 3108 85488 3120
rect 84988 3080 85488 3108
rect 84988 3068 84994 3080
rect 85482 3068 85488 3080
rect 85540 3068 85546 3120
rect 88518 3068 88524 3120
rect 88576 3108 88582 3120
rect 89622 3108 89628 3120
rect 88576 3080 89628 3108
rect 88576 3068 88582 3080
rect 89622 3068 89628 3080
rect 89680 3068 89686 3120
rect 164878 3108 164884 3120
rect 89732 3080 164884 3108
rect 75512 3012 82308 3040
rect 75512 3000 75518 3012
rect 82630 3000 82636 3052
rect 82688 3040 82694 3052
rect 89732 3040 89760 3080
rect 164878 3068 164884 3080
rect 164936 3068 164942 3120
rect 171137 3111 171195 3117
rect 171137 3077 171149 3111
rect 171183 3108 171195 3111
rect 180705 3111 180763 3117
rect 180705 3108 180717 3111
rect 171183 3080 180717 3108
rect 171183 3077 171195 3080
rect 171137 3071 171195 3077
rect 180705 3077 180717 3080
rect 180751 3077 180763 3111
rect 180705 3071 180763 3077
rect 193214 3068 193220 3120
rect 193272 3108 193278 3120
rect 194502 3108 194508 3120
rect 193272 3080 194508 3108
rect 193272 3068 193278 3080
rect 194502 3068 194508 3080
rect 194560 3068 194566 3120
rect 303798 3068 303804 3120
rect 303856 3108 303862 3120
rect 385770 3108 385776 3120
rect 303856 3080 385776 3108
rect 303856 3068 303862 3080
rect 385770 3068 385776 3080
rect 385828 3068 385834 3120
rect 395430 3068 395436 3120
rect 395488 3108 395494 3120
rect 395982 3108 395988 3120
rect 395488 3080 395988 3108
rect 395488 3068 395494 3080
rect 395982 3068 395988 3080
rect 396040 3068 396046 3120
rect 396626 3068 396632 3120
rect 396684 3108 396690 3120
rect 397362 3108 397368 3120
rect 396684 3080 397368 3108
rect 396684 3068 396690 3080
rect 397362 3068 397368 3080
rect 397420 3068 397426 3120
rect 399018 3068 399024 3120
rect 399076 3108 399082 3120
rect 400122 3108 400128 3120
rect 399076 3080 400128 3108
rect 399076 3068 399082 3080
rect 400122 3068 400128 3080
rect 400180 3068 400186 3120
rect 400214 3068 400220 3120
rect 400272 3108 400278 3120
rect 403618 3108 403624 3120
rect 400272 3080 403624 3108
rect 400272 3068 400278 3080
rect 403618 3068 403624 3080
rect 403676 3068 403682 3120
rect 403710 3068 403716 3120
rect 403768 3108 403774 3120
rect 477586 3108 477592 3120
rect 403768 3080 477592 3108
rect 403768 3068 403774 3080
rect 477586 3068 477592 3080
rect 477644 3068 477650 3120
rect 555970 3068 555976 3120
rect 556028 3108 556034 3120
rect 565538 3108 565544 3120
rect 556028 3080 565544 3108
rect 556028 3068 556034 3080
rect 565538 3068 565544 3080
rect 565596 3068 565602 3120
rect 166258 3040 166264 3052
rect 82688 3012 89760 3040
rect 89824 3012 166264 3040
rect 82688 3000 82694 3012
rect 84105 2975 84163 2981
rect 84105 2972 84117 2975
rect 75288 2944 84117 2972
rect 84105 2941 84117 2944
rect 84151 2941 84163 2975
rect 84105 2935 84163 2941
rect 86126 2932 86132 2984
rect 86184 2972 86190 2984
rect 89824 2972 89852 3012
rect 166258 3000 166264 3012
rect 166316 3000 166322 3052
rect 378778 3000 378784 3052
rect 378836 3040 378842 3052
rect 383381 3043 383439 3049
rect 383381 3040 383393 3043
rect 378836 3012 383393 3040
rect 378836 3000 378842 3012
rect 383381 3009 383393 3012
rect 383427 3009 383439 3043
rect 383381 3003 383439 3009
rect 385862 3000 385868 3052
rect 385920 3040 385926 3052
rect 390557 3043 390615 3049
rect 390557 3040 390569 3043
rect 385920 3012 390569 3040
rect 385920 3000 385926 3012
rect 390557 3009 390569 3012
rect 390603 3009 390615 3043
rect 390557 3003 390615 3009
rect 406013 3043 406071 3049
rect 406013 3009 406025 3043
rect 406059 3040 406071 3043
rect 410518 3040 410524 3052
rect 406059 3012 410524 3040
rect 406059 3009 406071 3012
rect 406013 3003 406071 3009
rect 410518 3000 410524 3012
rect 410576 3000 410582 3052
rect 414474 3000 414480 3052
rect 414532 3040 414538 3052
rect 418065 3043 418123 3049
rect 418065 3040 418077 3043
rect 414532 3012 418077 3040
rect 414532 3000 414538 3012
rect 418065 3009 418077 3012
rect 418111 3009 418123 3043
rect 418065 3003 418123 3009
rect 419629 3043 419687 3049
rect 419629 3009 419641 3043
rect 419675 3040 419687 3043
rect 421469 3043 421527 3049
rect 421469 3040 421481 3043
rect 419675 3012 421481 3040
rect 419675 3009 419687 3012
rect 419629 3003 419687 3009
rect 421469 3009 421481 3012
rect 421515 3009 421527 3043
rect 421469 3003 421527 3009
rect 421558 3000 421564 3052
rect 421616 3040 421622 3052
rect 480714 3040 480720 3052
rect 421616 3012 480720 3040
rect 421616 3000 421622 3012
rect 480714 3000 480720 3012
rect 480772 3000 480778 3052
rect 558822 3000 558828 3052
rect 558880 3040 558886 3052
rect 564621 3043 564679 3049
rect 564621 3040 564633 3043
rect 558880 3012 564633 3040
rect 558880 3000 558886 3012
rect 564621 3009 564633 3012
rect 564667 3009 564679 3043
rect 564621 3003 564679 3009
rect 86184 2944 89852 2972
rect 86184 2932 86190 2944
rect 93302 2932 93308 2984
rect 93360 2972 93366 2984
rect 169110 2972 169116 2984
rect 93360 2944 169116 2972
rect 93360 2932 93366 2944
rect 169110 2932 169116 2944
rect 169168 2932 169174 2984
rect 393038 2932 393044 2984
rect 393096 2972 393102 2984
rect 464246 2972 464252 2984
rect 393096 2944 464252 2972
rect 393096 2932 393102 2944
rect 464246 2932 464252 2944
rect 464304 2932 464310 2984
rect 466822 2932 466828 2984
rect 466880 2972 466886 2984
rect 467742 2972 467748 2984
rect 466880 2944 467748 2972
rect 466880 2932 466886 2944
rect 467742 2932 467748 2944
rect 467800 2932 467806 2984
rect 55309 2907 55367 2913
rect 55309 2873 55321 2907
rect 55355 2904 55367 2907
rect 66993 2907 67051 2913
rect 66993 2904 67005 2907
rect 55355 2876 67005 2904
rect 55355 2873 55367 2876
rect 55309 2867 55367 2873
rect 66993 2873 67005 2876
rect 67039 2873 67051 2907
rect 66993 2867 67051 2873
rect 74629 2907 74687 2913
rect 74629 2873 74641 2907
rect 74675 2904 74687 2907
rect 84013 2907 84071 2913
rect 84013 2904 84025 2907
rect 74675 2876 84025 2904
rect 74675 2873 74687 2876
rect 74629 2867 74687 2873
rect 84013 2873 84025 2876
rect 84059 2873 84071 2907
rect 84013 2867 84071 2873
rect 93857 2907 93915 2913
rect 93857 2873 93869 2907
rect 93903 2904 93915 2907
rect 93903 2876 95648 2904
rect 93903 2873 93915 2876
rect 93857 2867 93915 2873
rect 89714 2796 89720 2848
rect 89772 2836 89778 2848
rect 95418 2836 95424 2848
rect 89772 2808 95424 2836
rect 89772 2796 89778 2808
rect 95418 2796 95424 2808
rect 95476 2796 95482 2848
rect 95620 2768 95648 2876
rect 95694 2864 95700 2916
rect 95752 2904 95758 2916
rect 96522 2904 96528 2916
rect 95752 2876 96528 2904
rect 95752 2864 95758 2876
rect 96522 2864 96528 2876
rect 96580 2864 96586 2916
rect 96890 2864 96896 2916
rect 96948 2904 96954 2916
rect 102686 2904 102692 2916
rect 96948 2876 102692 2904
rect 96948 2864 96954 2876
rect 102686 2864 102692 2876
rect 102744 2864 102750 2916
rect 102778 2864 102784 2916
rect 102836 2904 102842 2916
rect 103422 2904 103428 2916
rect 102836 2876 103428 2904
rect 102836 2864 102842 2876
rect 103422 2864 103428 2876
rect 103480 2864 103486 2916
rect 103974 2864 103980 2916
rect 104032 2904 104038 2916
rect 105538 2904 105544 2916
rect 104032 2876 105544 2904
rect 104032 2864 104038 2876
rect 105538 2864 105544 2876
rect 105596 2864 105602 2916
rect 106366 2864 106372 2916
rect 106424 2904 106430 2916
rect 107562 2904 107568 2916
rect 106424 2876 107568 2904
rect 106424 2864 106430 2876
rect 107562 2864 107568 2876
rect 107620 2864 107626 2916
rect 107654 2864 107660 2916
rect 107712 2904 107718 2916
rect 107712 2876 111104 2904
rect 107712 2864 107718 2876
rect 95988 2808 100432 2836
rect 95988 2768 96016 2808
rect 95620 2740 96016 2768
rect 100404 2768 100432 2808
rect 100478 2796 100484 2848
rect 100536 2836 100542 2848
rect 110969 2839 111027 2845
rect 110969 2836 110981 2839
rect 100536 2808 110981 2836
rect 100536 2796 100542 2808
rect 110969 2805 110981 2808
rect 111015 2805 111027 2839
rect 110969 2799 111027 2805
rect 103425 2771 103483 2777
rect 103425 2768 103437 2771
rect 100404 2740 103437 2768
rect 103425 2737 103437 2740
rect 103471 2737 103483 2771
rect 111076 2768 111104 2876
rect 111150 2864 111156 2916
rect 111208 2904 111214 2916
rect 111702 2904 111708 2916
rect 111208 2876 111708 2904
rect 111208 2864 111214 2876
rect 111702 2864 111708 2876
rect 111760 2864 111766 2916
rect 169018 2904 169024 2916
rect 111812 2876 169024 2904
rect 111245 2839 111303 2845
rect 111245 2805 111257 2839
rect 111291 2836 111303 2839
rect 111812 2836 111840 2876
rect 169018 2864 169024 2876
rect 169076 2864 169082 2916
rect 253842 2864 253848 2916
rect 253900 2904 253906 2916
rect 292574 2904 292580 2916
rect 253900 2876 292580 2904
rect 253900 2864 253906 2876
rect 292574 2864 292580 2876
rect 292632 2864 292638 2916
rect 410886 2864 410892 2916
rect 410944 2904 410950 2916
rect 479518 2904 479524 2916
rect 410944 2876 479524 2904
rect 410944 2864 410950 2876
rect 479518 2864 479524 2876
rect 479576 2864 479582 2916
rect 540514 2864 540520 2916
rect 540572 2904 540578 2916
rect 547322 2904 547328 2916
rect 540572 2876 547328 2904
rect 540572 2864 540578 2876
rect 547322 2864 547328 2876
rect 547380 2864 547386 2916
rect 171594 2836 171600 2848
rect 111291 2808 111840 2836
rect 111904 2808 171600 2836
rect 111291 2805 111303 2808
rect 111245 2799 111303 2805
rect 111904 2768 111932 2808
rect 171594 2796 171600 2808
rect 171652 2796 171658 2848
rect 261018 2796 261024 2848
rect 261076 2836 261082 2848
rect 311158 2836 311164 2848
rect 261076 2808 311164 2836
rect 261076 2796 261082 2808
rect 311158 2796 311164 2808
rect 311216 2796 311222 2848
rect 346670 2796 346676 2848
rect 346728 2836 346734 2848
rect 419629 2839 419687 2845
rect 419629 2836 419641 2839
rect 346728 2808 419641 2836
rect 346728 2796 346734 2808
rect 419629 2805 419641 2808
rect 419675 2805 419687 2839
rect 419629 2799 419687 2805
rect 419721 2839 419779 2845
rect 419721 2805 419733 2839
rect 419767 2836 419779 2839
rect 425054 2836 425060 2848
rect 419767 2808 425060 2836
rect 419767 2805 419779 2808
rect 419721 2799 419779 2805
rect 425054 2796 425060 2808
rect 425112 2796 425118 2848
rect 425146 2796 425152 2848
rect 425204 2836 425210 2848
rect 485038 2836 485044 2848
rect 425204 2808 485044 2836
rect 425204 2796 425210 2808
rect 485038 2796 485044 2808
rect 485096 2796 485102 2848
rect 550818 2796 550824 2848
rect 550876 2836 550882 2848
rect 550876 2808 551232 2836
rect 550876 2796 550882 2808
rect 551204 2780 551232 2808
rect 553394 2796 553400 2848
rect 553452 2836 553458 2848
rect 553452 2808 553624 2836
rect 553452 2796 553458 2808
rect 553596 2780 553624 2808
rect 111076 2740 111932 2768
rect 103425 2731 103483 2737
rect 274082 2728 274088 2780
rect 274140 2768 274146 2780
rect 461026 2768 461032 2780
rect 274140 2740 461032 2768
rect 274140 2728 274146 2740
rect 461026 2728 461032 2740
rect 461084 2728 461090 2780
rect 551186 2728 551192 2780
rect 551244 2728 551250 2780
rect 553578 2728 553584 2780
rect 553636 2728 553642 2780
rect 269298 2660 269304 2712
rect 269356 2700 269362 2712
rect 459830 2700 459836 2712
rect 269356 2672 459836 2700
rect 269356 2660 269362 2672
rect 459830 2660 459836 2672
rect 459888 2660 459894 2712
rect 262214 2592 262220 2644
rect 262272 2632 262278 2644
rect 456886 2632 456892 2644
rect 262272 2604 456892 2632
rect 262272 2592 262278 2604
rect 456886 2592 456892 2604
rect 456944 2592 456950 2644
rect 243170 2524 243176 2576
rect 243228 2564 243234 2576
rect 451550 2564 451556 2576
rect 243228 2536 451556 2564
rect 243228 2524 243234 2536
rect 451550 2524 451556 2536
rect 451608 2524 451614 2576
rect 183738 2456 183744 2508
rect 183796 2496 183802 2508
rect 184842 2496 184848 2508
rect 183796 2468 184848 2496
rect 183796 2456 183802 2468
rect 184842 2456 184848 2468
rect 184900 2456 184906 2508
rect 235994 2456 236000 2508
rect 236052 2496 236058 2508
rect 448974 2496 448980 2508
rect 236052 2468 446812 2496
rect 448935 2468 448980 2496
rect 236052 2456 236058 2468
rect 228910 2388 228916 2440
rect 228968 2428 228974 2440
rect 415394 2428 415400 2440
rect 228968 2400 415400 2428
rect 228968 2388 228974 2400
rect 415394 2388 415400 2400
rect 415452 2388 415458 2440
rect 424962 2388 424968 2440
rect 425020 2428 425026 2440
rect 434714 2428 434720 2440
rect 425020 2400 434720 2428
rect 425020 2388 425026 2400
rect 434714 2388 434720 2400
rect 434772 2388 434778 2440
rect 446784 2428 446812 2468
rect 448974 2456 448980 2468
rect 449032 2456 449038 2508
rect 449066 2428 449072 2440
rect 446784 2400 449072 2428
rect 449066 2388 449072 2400
rect 449124 2388 449130 2440
rect 214650 2320 214656 2372
rect 214708 2360 214714 2372
rect 342898 2360 342904 2372
rect 214708 2332 342904 2360
rect 214708 2320 214714 2332
rect 342898 2320 342904 2332
rect 342956 2320 342962 2372
rect 347682 2320 347688 2372
rect 347740 2360 347746 2372
rect 441982 2360 441988 2372
rect 347740 2332 441988 2360
rect 347740 2320 347746 2332
rect 441982 2320 441988 2332
rect 442040 2320 442046 2372
rect 442074 2320 442080 2372
rect 442132 2360 442138 2372
rect 447226 2360 447232 2372
rect 442132 2332 447232 2360
rect 442132 2320 442138 2332
rect 447226 2320 447232 2332
rect 447284 2320 447290 2372
rect 200390 2252 200396 2304
rect 200448 2292 200454 2304
rect 347317 2295 347375 2301
rect 347317 2292 347329 2295
rect 200448 2264 347329 2292
rect 200448 2252 200454 2264
rect 347317 2261 347329 2264
rect 347363 2261 347375 2295
rect 347317 2255 347375 2261
rect 347406 2252 347412 2304
rect 347464 2252 347470 2304
rect 347593 2295 347651 2301
rect 347593 2261 347605 2295
rect 347639 2292 347651 2295
rect 437566 2292 437572 2304
rect 347639 2264 437572 2292
rect 347639 2261 347651 2264
rect 347593 2255 347651 2261
rect 437566 2252 437572 2264
rect 437624 2252 437630 2304
rect 199194 2184 199200 2236
rect 199252 2224 199258 2236
rect 328089 2227 328147 2233
rect 328089 2224 328101 2227
rect 199252 2196 328101 2224
rect 199252 2184 199258 2196
rect 328089 2193 328101 2196
rect 328135 2193 328147 2227
rect 328089 2187 328147 2193
rect 328181 2227 328239 2233
rect 328181 2193 328193 2227
rect 328227 2224 328239 2227
rect 347424 2224 347452 2252
rect 328227 2196 347452 2224
rect 328227 2193 328239 2196
rect 328181 2187 328239 2193
rect 347682 2184 347688 2236
rect 347740 2224 347746 2236
rect 386049 2227 386107 2233
rect 386049 2224 386061 2227
rect 347740 2196 386061 2224
rect 347740 2184 347746 2196
rect 386049 2193 386061 2196
rect 386095 2193 386107 2227
rect 386049 2187 386107 2193
rect 386141 2227 386199 2233
rect 386141 2193 386153 2227
rect 386187 2224 386199 2227
rect 437750 2224 437756 2236
rect 386187 2196 437756 2224
rect 386187 2193 386199 2196
rect 386141 2187 386199 2193
rect 437750 2184 437756 2196
rect 437808 2184 437814 2236
rect 192018 2116 192024 2168
rect 192076 2156 192082 2168
rect 347409 2159 347467 2165
rect 347409 2156 347421 2159
rect 192076 2128 347421 2156
rect 192076 2116 192082 2128
rect 347409 2125 347421 2128
rect 347455 2125 347467 2159
rect 347409 2119 347467 2125
rect 347593 2159 347651 2165
rect 347593 2125 347605 2159
rect 347639 2156 347651 2159
rect 385957 2159 386015 2165
rect 385957 2156 385969 2159
rect 347639 2128 385969 2156
rect 347639 2125 347651 2128
rect 347593 2119 347651 2125
rect 385957 2125 385969 2128
rect 386003 2125 386015 2159
rect 385957 2119 386015 2125
rect 386233 2159 386291 2165
rect 386233 2125 386245 2159
rect 386279 2156 386291 2159
rect 434898 2156 434904 2168
rect 386279 2128 434904 2156
rect 386279 2125 386291 2128
rect 386233 2119 386291 2125
rect 434898 2116 434904 2128
rect 434956 2116 434962 2168
rect 133782 2048 133788 2100
rect 133840 2088 133846 2100
rect 327997 2091 328055 2097
rect 327997 2088 328009 2091
rect 133840 2060 328009 2088
rect 133840 2048 133846 2060
rect 327997 2057 328009 2060
rect 328043 2057 328055 2091
rect 327997 2051 328055 2057
rect 328273 2091 328331 2097
rect 328273 2057 328285 2091
rect 328319 2088 328331 2091
rect 347317 2091 347375 2097
rect 347317 2088 347329 2091
rect 328319 2060 347329 2088
rect 328319 2057 328331 2060
rect 328273 2051 328331 2057
rect 347317 2057 347329 2060
rect 347363 2057 347375 2091
rect 347317 2051 347375 2057
rect 347685 2091 347743 2097
rect 347685 2057 347697 2091
rect 347731 2088 347743 2091
rect 381538 2088 381544 2100
rect 347731 2060 381544 2088
rect 347731 2057 347743 2060
rect 347685 2051 347743 2057
rect 381538 2048 381544 2060
rect 381596 2048 381602 2100
rect 386322 2048 386328 2100
rect 386380 2088 386386 2100
rect 415486 2088 415492 2100
rect 386380 2060 415492 2088
rect 386380 2048 386386 2060
rect 415486 2048 415492 2060
rect 415544 2048 415550 2100
rect 450170 2048 450176 2100
rect 450228 2088 450234 2100
rect 453945 2091 454003 2097
rect 453945 2088 453957 2091
rect 450228 2060 453957 2088
rect 450228 2048 450234 2060
rect 453945 2057 453957 2060
rect 453991 2057 454003 2091
rect 453945 2051 454003 2057
rect 276474 1980 276480 2032
rect 276532 2020 276538 2032
rect 462406 2020 462412 2032
rect 276532 1992 462412 2020
rect 276532 1980 276538 1992
rect 462406 1980 462412 1992
rect 462464 1980 462470 2032
rect 281258 1912 281264 1964
rect 281316 1952 281322 1964
rect 328089 1955 328147 1961
rect 328089 1952 328101 1955
rect 281316 1924 328101 1952
rect 281316 1912 281322 1924
rect 328089 1921 328101 1924
rect 328135 1921 328147 1955
rect 328089 1915 328147 1921
rect 328365 1955 328423 1961
rect 328365 1921 328377 1955
rect 328411 1952 328423 1955
rect 463878 1952 463884 1964
rect 328411 1924 463884 1952
rect 328411 1921 328423 1924
rect 328365 1915 328423 1921
rect 463878 1912 463884 1924
rect 463936 1912 463942 1964
rect 288342 1844 288348 1896
rect 288400 1884 288406 1896
rect 327997 1887 328055 1893
rect 327997 1884 328009 1887
rect 288400 1856 328009 1884
rect 288400 1844 288406 1856
rect 327997 1853 328009 1856
rect 328043 1853 328055 1887
rect 327997 1847 328055 1853
rect 328181 1887 328239 1893
rect 328181 1853 328193 1887
rect 328227 1884 328239 1887
rect 347409 1887 347467 1893
rect 347409 1884 347421 1887
rect 328227 1856 347421 1884
rect 328227 1853 328239 1856
rect 328181 1847 328239 1853
rect 347409 1853 347421 1856
rect 347455 1853 347467 1887
rect 347409 1847 347467 1853
rect 347685 1887 347743 1893
rect 347685 1853 347697 1887
rect 347731 1884 347743 1887
rect 386141 1887 386199 1893
rect 386141 1884 386153 1887
rect 347731 1856 386153 1884
rect 347731 1853 347743 1856
rect 347685 1847 347743 1853
rect 386141 1853 386153 1856
rect 386187 1853 386199 1887
rect 386141 1847 386199 1853
rect 386233 1887 386291 1893
rect 386233 1853 386245 1887
rect 386279 1884 386291 1887
rect 465350 1884 465356 1896
rect 386279 1856 465356 1884
rect 386279 1853 386291 1856
rect 386233 1847 386291 1853
rect 465350 1844 465356 1856
rect 465408 1844 465414 1896
rect 299106 1776 299112 1828
rect 299164 1816 299170 1828
rect 385954 1816 385960 1828
rect 299164 1788 385960 1816
rect 299164 1776 299170 1788
rect 385954 1776 385960 1788
rect 386012 1776 386018 1828
rect 386322 1776 386328 1828
rect 386380 1816 386386 1828
rect 469490 1816 469496 1828
rect 386380 1788 469496 1816
rect 386380 1776 386386 1788
rect 469490 1776 469496 1788
rect 469548 1776 469554 1828
rect 292574 1708 292580 1760
rect 292632 1748 292638 1760
rect 454218 1748 454224 1760
rect 292632 1720 454224 1748
rect 292632 1708 292638 1720
rect 454218 1708 454224 1720
rect 454276 1708 454282 1760
rect 311158 1640 311164 1692
rect 311216 1680 311222 1692
rect 456978 1680 456984 1692
rect 311216 1652 456984 1680
rect 311216 1640 311222 1652
rect 456978 1640 456984 1652
rect 457036 1640 457042 1692
rect 362126 1572 362132 1624
rect 362184 1612 362190 1624
rect 490098 1612 490104 1624
rect 362184 1584 490104 1612
rect 362184 1572 362190 1584
rect 490098 1572 490104 1584
rect 490156 1572 490162 1624
rect 165890 960 165896 1012
rect 165948 1000 165954 1012
rect 168009 1003 168067 1009
rect 168009 1000 168021 1003
rect 165948 972 168021 1000
rect 165948 960 165954 972
rect 168009 969 168021 972
rect 168055 969 168067 1003
rect 168009 963 168067 969
rect 65886 552 65892 604
rect 65944 592 65950 604
rect 65978 592 65984 604
rect 65944 564 65984 592
rect 65944 552 65950 564
rect 65978 552 65984 564
rect 66036 552 66042 604
rect 126606 592 126612 604
rect 126567 564 126612 592
rect 126606 552 126612 564
rect 126664 552 126670 604
rect 161106 552 161112 604
rect 161164 592 161170 604
rect 161382 592 161388 604
rect 161164 564 161388 592
rect 161164 552 161170 564
rect 161382 552 161388 564
rect 161440 552 161446 604
rect 178954 552 178960 604
rect 179012 592 179018 604
rect 179322 592 179328 604
rect 179012 564 179328 592
rect 179012 552 179018 564
rect 179322 552 179328 564
rect 179380 552 179386 604
rect 202690 552 202696 604
rect 202748 592 202754 604
rect 202785 595 202843 601
rect 202785 592 202797 595
rect 202748 564 202797 592
rect 202748 552 202754 564
rect 202785 561 202797 564
rect 202831 561 202843 595
rect 202785 555 202843 561
rect 445386 552 445392 604
rect 445444 592 445450 604
rect 445662 592 445668 604
rect 445444 564 445668 592
rect 445444 552 445450 564
rect 445662 552 445668 564
rect 445720 552 445726 604
rect 496538 552 496544 604
rect 496596 592 496602 604
rect 496722 592 496728 604
rect 496596 564 496728 592
rect 496596 552 496602 564
rect 496722 552 496728 564
rect 496780 552 496786 604
rect 554774 552 554780 604
rect 554832 592 554838 604
rect 554958 592 554964 604
rect 554832 564 554964 592
rect 554832 552 554838 564
rect 554958 552 554964 564
rect 555016 552 555022 604
<< via1 >>
rect 305644 700544 305696 700596
rect 332508 700544 332560 700596
rect 138664 700476 138716 700528
rect 154120 700476 154172 700528
rect 202788 700476 202840 700528
rect 250628 700476 250680 700528
rect 267648 700476 267700 700528
rect 282184 700476 282236 700528
rect 301504 700476 301556 700528
rect 397460 700476 397512 700528
rect 51724 700408 51776 700460
rect 72976 700408 73028 700460
rect 89168 700408 89220 700460
rect 138756 700408 138808 700460
rect 218980 700408 219032 700460
rect 282460 700408 282512 700460
rect 313924 700408 313976 700460
rect 413652 700408 413704 700460
rect 40500 700340 40552 700392
rect 282368 700340 282420 700392
rect 312544 700340 312596 700392
rect 462320 700340 462372 700392
rect 8116 700272 8168 700324
rect 8944 700272 8996 700324
rect 24308 700272 24360 700324
rect 282276 700272 282328 700324
rect 315304 700272 315356 700324
rect 527180 700272 527232 700324
rect 250628 698640 250680 698692
rect 252560 698640 252612 698692
rect 283288 698232 283340 698284
rect 283932 698232 283984 698284
rect 136640 697552 136692 697604
rect 137836 697552 137888 697604
rect 576124 696940 576176 696992
rect 580172 696940 580224 696992
rect 252560 696872 252612 696924
rect 260012 696872 260064 696924
rect 260012 694764 260064 694816
rect 267004 694764 267056 694816
rect 283104 694084 283156 694136
rect 283288 694084 283340 694136
rect 283104 692724 283156 692776
rect 283288 692724 283340 692776
rect 48504 691364 48556 691416
rect 51724 691364 51776 691416
rect 46940 685176 46992 685228
rect 48504 685176 48556 685228
rect 282920 683068 282972 683120
rect 3516 681708 3568 681760
rect 453304 681708 453356 681760
rect 42064 680212 42116 680264
rect 46940 680348 46992 680400
rect 133880 674772 133932 674824
rect 136640 674772 136692 674824
rect 40040 672052 40092 672104
rect 42064 672052 42116 672104
rect 131764 670692 131816 670744
rect 133880 670692 133932 670744
rect 267004 670624 267056 670676
rect 269764 670624 269816 670676
rect 3424 667904 3476 667956
rect 287704 667904 287756 667956
rect 37924 666476 37976 666528
rect 40040 666544 40092 666596
rect 283380 666544 283432 666596
rect 269764 659404 269816 659456
rect 271144 659404 271196 659456
rect 3056 652740 3108 652792
rect 10324 652740 10376 652792
rect 271144 651516 271196 651568
rect 271972 651516 272024 651568
rect 36544 650020 36596 650072
rect 37924 650020 37976 650072
rect 577504 650020 577556 650072
rect 579620 650020 579672 650072
rect 271972 648592 272024 648644
rect 274640 648524 274692 648576
rect 129004 648320 129056 648372
rect 131764 648320 131816 648372
rect 283104 647232 283156 647284
rect 283196 647232 283248 647284
rect 274640 645804 274692 645856
rect 276664 645804 276716 645856
rect 283104 640364 283156 640416
rect 283196 640364 283248 640416
rect 126244 640296 126296 640348
rect 129004 640296 129056 640348
rect 35256 634788 35308 634840
rect 36544 634788 36596 634840
rect 276664 633156 276716 633208
rect 278320 633156 278372 633208
rect 283012 630640 283064 630692
rect 283196 630640 283248 630692
rect 116584 629892 116636 629944
rect 126244 629892 126296 629944
rect 33784 629484 33836 629536
rect 35256 629484 35308 629536
rect 278320 627852 278372 627904
rect 279148 627852 279200 627904
rect 551376 627308 551428 627360
rect 551652 627308 551704 627360
rect 23388 619624 23440 619676
rect 84108 619624 84160 619676
rect 551192 618672 551244 618724
rect 551560 618672 551612 618724
rect 29736 618536 29788 618588
rect 33784 618536 33836 618588
rect 453304 616768 453356 616820
rect 456800 616768 456852 616820
rect 282368 614048 282420 614100
rect 313280 614048 313332 614100
rect 283012 611328 283064 611380
rect 283196 611328 283248 611380
rect 551376 611260 551428 611312
rect 551836 611260 551888 611312
rect 3332 609968 3384 610020
rect 13084 609968 13136 610020
rect 551836 606636 551888 606688
rect 551192 606500 551244 606552
rect 551836 606500 551888 606552
rect 551284 606432 551336 606484
rect 551928 606432 551980 606484
rect 551284 606339 551336 606348
rect 551284 606305 551293 606339
rect 551293 606305 551327 606339
rect 551327 606305 551336 606339
rect 551284 606296 551336 606305
rect 551376 601443 551428 601452
rect 551376 601409 551385 601443
rect 551385 601409 551419 601443
rect 551419 601409 551428 601443
rect 551376 601400 551428 601409
rect 283196 598884 283248 598936
rect 28908 598451 28960 598460
rect 28908 598417 28917 598451
rect 28917 598417 28951 598451
rect 28951 598417 28960 598451
rect 28908 598408 28960 598417
rect 28908 598136 28960 598188
rect 551192 598000 551244 598052
rect 551836 598000 551888 598052
rect 26148 597932 26200 597984
rect 28908 597932 28960 597984
rect 551284 596980 551336 597032
rect 551284 596844 551336 596896
rect 551928 596844 551980 596896
rect 551928 596708 551980 596760
rect 551376 596572 551428 596624
rect 551376 596479 551428 596488
rect 551376 596445 551385 596479
rect 551385 596445 551419 596479
rect 551419 596445 551428 596479
rect 551376 596436 551428 596445
rect 28908 595119 28960 595128
rect 28908 595085 28917 595119
rect 28917 595085 28951 595119
rect 28951 595085 28960 595119
rect 28908 595076 28960 595085
rect 551376 595076 551428 595128
rect 3516 594804 3568 594856
rect 9036 594804 9088 594856
rect 139216 594668 139268 594720
rect 139584 594668 139636 594720
rect 551376 592288 551428 592340
rect 551376 592195 551428 592204
rect 551376 592161 551385 592195
rect 551385 592161 551419 592195
rect 551419 592161 551428 592195
rect 551376 592152 551428 592161
rect 551376 592016 551428 592068
rect 551928 592016 551980 592068
rect 554596 590155 554648 590164
rect 554596 590121 554605 590155
rect 554605 590121 554639 590155
rect 554639 590121 554648 590155
rect 554596 590112 554648 590121
rect 28908 589908 28960 589960
rect 28264 589364 28316 589416
rect 28908 589364 28960 589416
rect 283012 589339 283064 589348
rect 283012 589305 283021 589339
rect 283021 589305 283055 589339
rect 283055 589305 283064 589339
rect 283012 589296 283064 589305
rect 554596 589296 554648 589348
rect 556160 589296 556212 589348
rect 28448 589228 28500 589280
rect 28908 589228 28960 589280
rect 554596 588752 554648 588804
rect 557632 588752 557684 588804
rect 28356 588548 28408 588600
rect 28908 588548 28960 588600
rect 551284 587188 551336 587240
rect 551928 587188 551980 587240
rect 554596 587052 554648 587104
rect 556804 587052 556856 587104
rect 551376 586916 551428 586968
rect 554596 586959 554648 586968
rect 554596 586925 554605 586959
rect 554605 586925 554639 586959
rect 554639 586925 554648 586959
rect 554596 586916 554648 586925
rect 554872 586304 554924 586356
rect 558184 586304 558236 586356
rect 551376 586279 551428 586288
rect 551376 586245 551385 586279
rect 551385 586245 551419 586279
rect 551419 586245 551428 586279
rect 551376 586236 551428 586245
rect 24124 586032 24176 586084
rect 26148 586032 26200 586084
rect 554872 585148 554924 585200
rect 560300 585148 560352 585200
rect 554872 583720 554924 583772
rect 561772 583720 561824 583772
rect 551192 582403 551244 582412
rect 551192 582369 551201 582403
rect 551201 582369 551235 582403
rect 551235 582369 551244 582403
rect 551192 582360 551244 582369
rect 554872 581000 554924 581052
rect 563060 581000 563112 581052
rect 28908 580252 28960 580304
rect 283012 579640 283064 579692
rect 283104 579640 283156 579692
rect 554872 579640 554924 579692
rect 564440 579640 564492 579692
rect 576216 579640 576268 579692
rect 580172 579640 580224 579692
rect 554872 578212 554924 578264
rect 565820 578212 565872 578264
rect 551192 576895 551244 576904
rect 551192 576861 551201 576895
rect 551201 576861 551235 576895
rect 551235 576861 551244 576895
rect 551192 576852 551244 576861
rect 551284 576852 551336 576904
rect 551928 576852 551980 576904
rect 553308 576895 553360 576904
rect 553308 576861 553317 576895
rect 553317 576861 553351 576895
rect 553351 576861 553360 576895
rect 553308 576852 553360 576861
rect 554872 576852 554924 576904
rect 567292 576852 567344 576904
rect 28632 576104 28684 576156
rect 28908 576147 28960 576156
rect 28908 576113 28917 576147
rect 28917 576113 28951 576147
rect 28951 576113 28960 576147
rect 28908 576104 28960 576113
rect 28908 575832 28960 575884
rect 553308 575492 553360 575544
rect 560944 575492 560996 575544
rect 28632 575263 28684 575272
rect 28632 575229 28641 575263
rect 28641 575229 28675 575263
rect 28675 575229 28684 575263
rect 28632 575220 28684 575229
rect 28632 575084 28684 575136
rect 28908 575084 28960 575136
rect 28816 575016 28868 575068
rect 28632 574948 28684 575000
rect 28632 574812 28684 574864
rect 28816 574744 28868 574796
rect 553308 574200 553360 574252
rect 568580 574200 568632 574252
rect 553308 574064 553360 574116
rect 569960 574064 570012 574116
rect 29368 573452 29420 573504
rect 30012 573427 30064 573436
rect 30012 573393 30021 573427
rect 30021 573393 30055 573427
rect 30055 573393 30064 573427
rect 30012 573384 30064 573393
rect 29092 572772 29144 572824
rect 30104 572772 30156 572824
rect 26424 572704 26476 572756
rect 29276 572704 29328 572756
rect 553308 572704 553360 572756
rect 571432 572704 571484 572756
rect 29920 572679 29972 572688
rect 29920 572645 29929 572679
rect 29929 572645 29963 572679
rect 29963 572645 29972 572679
rect 29920 572636 29972 572645
rect 26424 572568 26476 572620
rect 551928 572568 551980 572620
rect 199292 572432 199344 572484
rect 204260 572432 204312 572484
rect 189540 572296 189592 572348
rect 195980 572296 196032 572348
rect 198096 572296 198148 572348
rect 202880 572296 202932 572348
rect 188344 572160 188396 572212
rect 194600 572160 194652 572212
rect 196808 572160 196860 572212
rect 202972 572160 203024 572212
rect 209044 572160 209096 572212
rect 213920 572160 213972 572212
rect 206652 572092 206704 572144
rect 211160 572092 211212 572144
rect 218888 572092 218940 572144
rect 222200 572092 222252 572144
rect 190276 572024 190328 572076
rect 197360 572024 197412 572076
rect 207848 572024 207900 572076
rect 212540 572024 212592 572076
rect 194416 571888 194468 571940
rect 200120 571888 200172 571940
rect 205364 571888 205416 571940
rect 209780 571888 209832 571940
rect 227444 571888 227496 571940
rect 229100 571888 229152 571940
rect 195612 571820 195664 571872
rect 201500 571820 201552 571872
rect 23296 571752 23348 571804
rect 24676 571752 24728 571804
rect 267648 571752 267700 571804
rect 268292 571752 268344 571804
rect 217600 571684 217652 571736
rect 220820 571684 220872 571736
rect 216404 571616 216456 571668
rect 219440 571616 219492 571668
rect 228640 571616 228692 571668
rect 230480 571616 230532 571668
rect 553308 571616 553360 571668
rect 558276 571616 558328 571668
rect 202788 571548 202840 571600
rect 208400 571548 208452 571600
rect 213828 571548 213880 571600
rect 218060 571548 218112 571600
rect 220084 571548 220136 571600
rect 223672 571548 223724 571600
rect 224868 571548 224920 571600
rect 227812 571548 227864 571600
rect 201408 571480 201460 571532
rect 207020 571480 207072 571532
rect 212448 571480 212500 571532
rect 216680 571480 216732 571532
rect 223488 571480 223540 571532
rect 226340 571480 226392 571532
rect 231032 571480 231084 571532
rect 233332 571480 233384 571532
rect 273076 571480 273128 571532
rect 275652 571480 275704 571532
rect 278688 571480 278740 571532
rect 281724 571480 281776 571532
rect 191748 571412 191800 571464
rect 198832 571412 198884 571464
rect 200488 571412 200540 571464
rect 205640 571412 205692 571464
rect 211528 571412 211580 571464
rect 215300 571412 215352 571464
rect 222108 571412 222160 571464
rect 224960 571412 225012 571464
rect 233148 571412 233200 571464
rect 234620 571412 234672 571464
rect 235908 571412 235960 571464
rect 237472 571412 237524 571464
rect 269028 571412 269080 571464
rect 270776 571412 270828 571464
rect 271788 571412 271840 571464
rect 273260 571412 273312 571464
rect 274548 571412 274600 571464
rect 276848 571412 276900 571464
rect 277308 571412 277360 571464
rect 279332 571412 279384 571464
rect 193128 571344 193180 571396
rect 198740 571344 198792 571396
rect 204168 571344 204220 571396
rect 208492 571344 208544 571396
rect 210332 571344 210384 571396
rect 214012 571344 214064 571396
rect 215208 571344 215260 571396
rect 218152 571344 218204 571396
rect 221280 571344 221332 571396
rect 223580 571344 223632 571396
rect 226156 571344 226208 571396
rect 227720 571344 227772 571396
rect 229836 571344 229888 571396
rect 231860 571344 231912 571396
rect 232320 571344 232372 571396
rect 233240 571344 233292 571396
rect 234528 571344 234580 571396
rect 236000 571344 236052 571396
rect 239588 571344 239640 571396
rect 240140 571344 240192 571396
rect 240876 571344 240928 571396
rect 241520 571344 241572 571396
rect 242072 571344 242124 571396
rect 242900 571344 242952 571396
rect 254860 571344 254912 571396
rect 255320 571344 255372 571396
rect 256056 571344 256108 571396
rect 256700 571344 256752 571396
rect 257344 571344 257396 571396
rect 263416 571344 263468 571396
rect 264612 571344 264664 571396
rect 264888 571344 264940 571396
rect 265900 571344 265952 571396
rect 266268 571344 266320 571396
rect 267096 571344 267148 571396
rect 268936 571344 268988 571396
rect 269488 571344 269540 571396
rect 270408 571344 270460 571396
rect 271972 571344 272024 571396
rect 273168 571344 273220 571396
rect 274640 571344 274692 571396
rect 275928 571344 275980 571396
rect 278044 571344 278096 571396
rect 278596 571344 278648 571396
rect 280528 571344 280580 571396
rect 29000 571276 29052 571328
rect 31852 571276 31904 571328
rect 253940 571276 253992 571328
rect 30288 570596 30340 570648
rect 74540 570596 74592 570648
rect 30288 570460 30340 570512
rect 31760 570120 31812 570172
rect 29000 569984 29052 570036
rect 29644 569984 29696 570036
rect 318524 569916 318576 569968
rect 318708 569916 318760 569968
rect 354404 569916 354456 569968
rect 354588 569916 354640 569968
rect 553308 569916 553360 569968
rect 572720 569916 572772 569968
rect 112536 569848 112588 569900
rect 138664 569848 138716 569900
rect 282276 569848 282328 569900
rect 284300 569848 284352 569900
rect 30196 569236 30248 569288
rect 78680 569236 78732 569288
rect 56416 569168 56468 569220
rect 281540 569168 281592 569220
rect 282276 569168 282328 569220
rect 286324 569168 286376 569220
rect 580448 569168 580500 569220
rect 327540 568488 327592 568540
rect 328276 568488 328328 568540
rect 338304 568488 338356 568540
rect 339316 568488 339368 568540
rect 346124 568488 346176 568540
rect 408224 568488 408276 568540
rect 456064 568488 456116 568540
rect 483020 568488 483072 568540
rect 529020 568488 529072 568540
rect 529848 568488 529900 568540
rect 329380 568420 329432 568472
rect 392032 568420 392084 568472
rect 343548 568352 343600 568404
rect 411812 568352 411864 568404
rect 325792 568284 325844 568336
rect 394884 568284 394936 568336
rect 341984 568216 342036 568268
rect 415400 568216 415452 568268
rect 339408 568148 339460 568200
rect 418988 568148 419040 568200
rect 336556 568080 336608 568132
rect 422576 568080 422628 568132
rect 335268 568012 335320 568064
rect 426164 568012 426216 568064
rect 332416 567944 332468 567996
rect 429752 567944 429804 567996
rect 29276 567876 29328 567928
rect 56600 567876 56652 567928
rect 331128 567876 331180 567928
rect 433340 567876 433392 567928
rect 29460 567808 29512 567860
rect 66352 567808 66404 567860
rect 328368 567808 328420 567860
rect 436928 567808 436980 567860
rect 347688 567740 347740 567792
rect 404636 567740 404688 567792
rect 332968 567672 333020 567724
rect 389180 567672 389232 567724
rect 336464 567604 336516 567656
rect 387800 567604 387852 567656
rect 350448 567536 350500 567588
rect 401048 567536 401100 567588
rect 351736 567468 351788 567520
rect 397460 567468 397512 567520
rect 340144 567400 340196 567452
rect 385040 567400 385092 567452
rect 343732 567332 343784 567384
rect 383660 567332 383712 567384
rect 347320 567264 347372 567316
rect 380992 567264 381044 567316
rect 3516 567196 3568 567248
rect 9128 567196 9180 567248
rect 29092 567196 29144 567248
rect 320364 567196 320416 567248
rect 321468 567196 321520 567248
rect 350908 567196 350960 567248
rect 356244 567196 356296 567248
rect 357348 567196 357400 567248
rect 358820 567196 358872 567248
rect 359832 567196 359884 567248
rect 379520 567196 379572 567248
rect 29368 566448 29420 566500
rect 60832 566448 60884 566500
rect 361580 566448 361632 566500
rect 372620 566448 372672 566500
rect 368388 565836 368440 565888
rect 369860 565836 369912 565888
rect 29092 565156 29144 565208
rect 49700 565156 49752 565208
rect 358084 565156 358136 565208
rect 29552 565088 29604 565140
rect 63500 565088 63552 565140
rect 375564 565088 375616 565140
rect 29920 563660 29972 563712
rect 67640 563660 67692 563712
rect 355876 563660 355928 563712
rect 389272 563660 389324 563712
rect 29184 563524 29236 563576
rect 29920 563524 29972 563576
rect 364340 563048 364392 563100
rect 369860 563048 369912 563100
rect 30288 562300 30340 562352
rect 71780 562300 71832 562352
rect 362960 562300 363012 562352
rect 364248 562300 364300 562352
rect 365720 562300 365772 562352
rect 367008 562300 367060 562352
rect 365628 562232 365680 562284
rect 375380 562300 375432 562352
rect 29828 560940 29880 560992
rect 86960 560940 87012 560992
rect 362868 560940 362920 560992
rect 379612 560940 379664 560992
rect 283196 560260 283248 560312
rect 283288 560260 283340 560312
rect 358820 558152 358872 558204
rect 360108 558152 360160 558204
rect 304264 556180 304316 556232
rect 580172 556180 580224 556232
rect 364248 554004 364300 554056
rect 371240 554004 371292 554056
rect 317328 552644 317380 552696
rect 400312 552644 400364 552696
rect 3148 552032 3200 552084
rect 279516 552032 279568 552084
rect 29552 551284 29604 551336
rect 95240 551284 95292 551336
rect 543648 547204 543700 547256
rect 553124 547204 553176 547256
rect 540888 547136 540940 547188
rect 553032 547136 553084 547188
rect 545028 547068 545080 547120
rect 553216 547068 553268 547120
rect 366916 546456 366968 546508
rect 371332 546456 371384 546508
rect 354496 542988 354548 543040
rect 393320 542988 393372 543040
rect 322848 541628 322900 541680
rect 396080 541628 396132 541680
rect 282920 540948 282972 541000
rect 283196 540948 283248 541000
rect 358728 540200 358780 540252
rect 386420 540200 386472 540252
rect 366824 538840 366876 538892
rect 374000 538840 374052 538892
rect 3516 538228 3568 538280
rect 10416 538228 10468 538280
rect 360108 537480 360160 537532
rect 374092 537480 374144 537532
rect 357164 536120 357216 536172
rect 376116 536120 376168 536172
rect 360568 536052 360620 536104
rect 382280 536052 382332 536104
rect 26608 535619 26660 535628
rect 26608 535585 26617 535619
rect 26617 535585 26651 535619
rect 26651 535585 26660 535619
rect 26608 535576 26660 535585
rect 26792 535440 26844 535492
rect 26792 535236 26844 535288
rect 367008 535236 367060 535288
rect 369860 535236 369912 535288
rect 353208 535168 353260 535220
rect 378232 535168 378284 535220
rect 152464 535100 152516 535152
rect 436008 535100 436060 535152
rect 156328 535032 156380 535084
rect 446128 535032 446180 535084
rect 27068 534964 27120 535016
rect 148140 534964 148192 535016
rect 442908 534964 442960 535016
rect 147956 534896 148008 534948
rect 450452 534896 450504 534948
rect 143816 534828 143868 534880
rect 452568 534828 452620 534880
rect 167000 534760 167052 534812
rect 483848 534760 483900 534812
rect 139492 534692 139544 534744
rect 456984 534692 457036 534744
rect 137376 534624 137428 534676
rect 459100 534624 459152 534676
rect 135260 534556 135312 534608
rect 461216 534556 461268 534608
rect 131948 534488 132000 534540
rect 464528 534488 464580 534540
rect 129832 534420 129884 534472
rect 466644 534420 466696 534472
rect 127716 534352 127768 534404
rect 468760 534352 468812 534404
rect 125508 534284 125560 534336
rect 470968 534284 471020 534336
rect 123392 534216 123444 534268
rect 473452 534216 473504 534268
rect 121184 534148 121236 534200
rect 475292 534148 475344 534200
rect 111064 534080 111116 534132
rect 487160 534080 487212 534132
rect 339316 534012 339368 534064
rect 386880 534012 386932 534064
rect 335176 533944 335228 533996
rect 389180 533944 389232 533996
rect 26148 533876 26200 533928
rect 34980 533876 35032 533928
rect 331036 533876 331088 533928
rect 391204 533876 391256 533928
rect 25044 533808 25096 533860
rect 37188 533808 37240 533860
rect 328276 533808 328328 533860
rect 393320 533808 393372 533860
rect 25136 533740 25188 533792
rect 39304 533740 39356 533792
rect 318708 533740 318760 533792
rect 398932 533740 398984 533792
rect 25228 533672 25280 533724
rect 41420 533672 41472 533724
rect 323952 533672 324004 533724
rect 443000 533672 443052 533724
rect 25320 533604 25372 533656
rect 43628 533604 43680 533656
rect 322848 533604 322900 533656
rect 445760 533604 445812 533656
rect 530860 533604 530912 533656
rect 551468 533604 551520 533656
rect 27160 533536 27212 533588
rect 29736 533536 29788 533588
rect 56508 533536 56560 533588
rect 321284 533536 321336 533588
rect 447140 533536 447192 533588
rect 514668 533536 514720 533588
rect 552296 533536 552348 533588
rect 27252 533468 27304 533520
rect 84568 533468 84620 533520
rect 320732 533468 320784 533520
rect 448520 533468 448572 533520
rect 512552 533468 512604 533520
rect 552204 533468 552256 533520
rect 86684 533400 86736 533452
rect 319628 533400 319680 533452
rect 451280 533400 451332 533452
rect 510436 533400 510488 533452
rect 552020 533400 552072 533452
rect 26240 533332 26292 533384
rect 27068 533332 27120 533384
rect 27712 533332 27764 533384
rect 91008 533332 91060 533384
rect 266728 533332 266780 533384
rect 267648 533332 267700 533384
rect 318524 533332 318576 533384
rect 452660 533332 452712 533384
rect 529848 533332 529900 533384
rect 574376 533332 574428 533384
rect 342076 533264 342128 533316
rect 385132 533264 385184 533316
rect 346216 533196 346268 533248
rect 382556 533196 382608 533248
rect 349068 533128 349120 533180
rect 380440 533128 380492 533180
rect 354588 533060 354640 533112
rect 377220 533060 377272 533112
rect 193404 532992 193456 533044
rect 403072 532992 403124 533044
rect 192392 532924 192444 532976
rect 404452 532924 404504 532976
rect 189080 532856 189132 532908
rect 407396 532856 407448 532908
rect 183744 532788 183796 532840
rect 412732 532788 412784 532840
rect 177304 532720 177356 532772
rect 419632 532720 419684 532772
rect 28724 532652 28776 532704
rect 33876 532652 33928 532704
rect 42524 532652 42576 532704
rect 344376 532652 344428 532704
rect 409880 532652 409932 532704
rect 554320 532652 554372 532704
rect 25504 532584 25556 532636
rect 45744 532584 45796 532636
rect 342168 532584 342220 532636
rect 412640 532584 412692 532636
rect 547052 532584 547104 532636
rect 551744 532584 551796 532636
rect 25688 532516 25740 532568
rect 47952 532516 48004 532568
rect 324136 532516 324188 532568
rect 395528 532516 395580 532568
rect 536288 532516 536340 532568
rect 551560 532516 551612 532568
rect 21364 532448 21416 532500
rect 24124 532448 24176 532500
rect 25780 532448 25832 532500
rect 52276 532448 52328 532500
rect 340144 532448 340196 532500
rect 416780 532448 416832 532500
rect 538128 532448 538180 532500
rect 28448 532380 28500 532432
rect 54392 532380 54444 532432
rect 321468 532380 321520 532432
rect 397644 532380 397696 532432
rect 401508 532380 401560 532432
rect 455420 532380 455472 532432
rect 531964 532380 532016 532432
rect 554136 532448 554188 532500
rect 553952 532380 554004 532432
rect 25872 532312 25924 532364
rect 58716 532312 58768 532364
rect 337936 532312 337988 532364
rect 419540 532312 419592 532364
rect 527640 532312 527692 532364
rect 551376 532312 551428 532364
rect 26056 532244 26108 532296
rect 60832 532244 60884 532296
rect 335820 532244 335872 532296
rect 423680 532244 423732 532296
rect 529756 532244 529808 532296
rect 24952 532176 25004 532228
rect 63040 532176 63092 532228
rect 333612 532176 333664 532228
rect 427820 532176 427872 532228
rect 525524 532176 525576 532228
rect 553860 532244 553912 532296
rect 26516 532108 26568 532160
rect 67364 532108 67416 532160
rect 331496 532108 331548 532160
rect 430580 532108 430632 532160
rect 523316 532108 523368 532160
rect 553768 532176 553820 532228
rect 549168 532108 549220 532160
rect 551836 532108 551888 532160
rect 28172 532040 28224 532092
rect 69480 532040 69532 532092
rect 329288 532040 329340 532092
rect 434720 532040 434772 532092
rect 521200 532040 521252 532092
rect 553584 532040 553636 532092
rect 26976 531972 27028 532024
rect 75920 531972 75972 532024
rect 326988 531972 327040 532024
rect 437480 531972 437532 532024
rect 518716 531972 518768 532024
rect 551100 531972 551152 532024
rect 25412 531904 25464 531956
rect 40408 531904 40460 531956
rect 346308 531904 346360 531956
rect 405740 531904 405792 531956
rect 26792 531836 26844 531888
rect 36084 531836 36136 531888
rect 348700 531836 348752 531888
rect 401600 531836 401652 531888
rect 28632 531768 28684 531820
rect 38200 531768 38252 531820
rect 350908 531768 350960 531820
rect 398840 531768 398892 531820
rect 353024 531700 353076 531752
rect 394792 531700 394844 531752
rect 26424 531632 26476 531684
rect 355232 531632 355284 531684
rect 391940 531632 391992 531684
rect 167552 531564 167604 531616
rect 339500 531564 339552 531616
rect 357348 531564 357400 531616
rect 387892 531564 387944 531616
rect 163228 531496 163280 531548
rect 344928 531496 344980 531548
rect 359464 531496 359516 531548
rect 383752 531496 383804 531548
rect 161112 531428 161164 531480
rect 347780 531428 347832 531480
rect 361488 531428 361540 531480
rect 380900 531428 380952 531480
rect 158904 531360 158956 531412
rect 353208 531360 353260 531412
rect 363788 531360 363840 531412
rect 376760 531360 376812 531412
rect 26608 531224 26660 531276
rect 29920 531224 29972 531276
rect 30656 531224 30708 531276
rect 156788 531292 156840 531344
rect 59820 531224 59872 531276
rect 353208 531224 353260 531276
rect 27988 531156 28040 531208
rect 70584 531156 70636 531208
rect 22100 531088 22152 531140
rect 23388 531088 23440 531140
rect 26700 531088 26752 531140
rect 65156 531088 65208 531140
rect 150348 531088 150400 531140
rect 156328 531088 156380 531140
rect 26884 531020 26936 531072
rect 71596 531020 71648 531072
rect 184848 531020 184900 531072
rect 198740 531020 198792 531072
rect 199660 531020 199712 531072
rect 202880 531020 202932 531072
rect 203892 531020 203944 531072
rect 223580 531088 223632 531140
rect 224316 531088 224368 531140
rect 227720 531088 227772 531140
rect 228732 531088 228784 531140
rect 233240 531088 233292 531140
rect 234068 531088 234120 531140
rect 237380 531088 237432 531140
rect 238300 531088 238352 531140
rect 339500 531156 339552 531208
rect 261300 531088 261352 531140
rect 262128 531088 262180 531140
rect 262404 531088 262456 531140
rect 263508 531088 263560 531140
rect 267832 531088 267884 531140
rect 268936 531088 268988 531140
rect 271052 531088 271104 531140
rect 271788 531088 271840 531140
rect 272064 531088 272116 531140
rect 273168 531088 273220 531140
rect 276388 531088 276440 531140
rect 277308 531088 277360 531140
rect 277492 531088 277544 531140
rect 278596 531088 278648 531140
rect 28080 530952 28132 531004
rect 77024 530952 77076 531004
rect 298192 531020 298244 531072
rect 326068 531088 326120 531140
rect 326896 531088 326948 531140
rect 330392 531088 330444 531140
rect 331128 531088 331180 531140
rect 334716 531088 334768 531140
rect 335268 531088 335320 531140
rect 341156 531088 341208 531140
rect 341984 531088 342036 531140
rect 347780 531156 347832 531208
rect 439688 531224 439740 531276
rect 442908 531224 442960 531276
rect 448520 531224 448572 531276
rect 535184 531224 535236 531276
rect 345480 531088 345532 531140
rect 346124 531088 346176 531140
rect 349804 531088 349856 531140
rect 350448 531088 350500 531140
rect 354036 531088 354088 531140
rect 354496 531088 354548 531140
rect 437664 531156 437716 531208
rect 533988 531156 534040 531208
rect 551376 531224 551428 531276
rect 551928 531224 551980 531276
rect 552388 531224 552440 531276
rect 552940 531224 552992 531276
rect 552572 531156 552624 531208
rect 435364 531088 435416 531140
rect 533068 531088 533120 531140
rect 552480 531088 552532 531140
rect 429292 531020 429344 531072
rect 528468 531020 528520 531072
rect 551284 531020 551336 531072
rect 298100 530952 298152 531004
rect 344928 530952 344980 531004
rect 433340 530952 433392 531004
rect 526536 530952 526588 531004
rect 27896 530884 27948 530936
rect 78128 530884 78180 530936
rect 186964 530884 187016 530936
rect 409880 530884 409932 530936
rect 522212 530884 522264 530936
rect 551192 530952 551244 531004
rect 548156 530884 548208 530936
rect 552756 530884 552808 530936
rect 27344 530816 27396 530868
rect 81348 530816 81400 530868
rect 146024 530816 146076 530868
rect 147956 530816 148008 530868
rect 411628 530816 411680 530868
rect 524328 530816 524380 530868
rect 554044 530816 554096 530868
rect 27804 530748 27856 530800
rect 83464 530748 83516 530800
rect 182640 530748 182692 530800
rect 414020 530748 414072 530800
rect 520096 530748 520148 530800
rect 552296 530748 552348 530800
rect 27436 530680 27488 530732
rect 85672 530680 85724 530732
rect 180524 530680 180576 530732
rect 415952 530680 416004 530732
rect 517980 530680 518032 530732
rect 550272 530680 550324 530732
rect 552848 530680 552900 530732
rect 27620 530612 27672 530664
rect 88892 530612 88944 530664
rect 90364 530612 90416 530664
rect 99656 530612 99708 530664
rect 178316 530612 178368 530664
rect 418252 530612 418304 530664
rect 513656 530612 513708 530664
rect 552112 530612 552164 530664
rect 555424 530612 555476 530664
rect 562600 530612 562652 530664
rect 27528 530544 27580 530596
rect 89996 530544 90048 530596
rect 90548 530544 90600 530596
rect 105084 530544 105136 530596
rect 112628 530544 112680 530596
rect 167000 530544 167052 530596
rect 176200 530544 176252 530596
rect 420276 530544 420328 530596
rect 436008 530544 436060 530596
rect 444380 530544 444432 530596
rect 511448 530544 511500 530596
rect 553492 530544 553544 530596
rect 558276 530544 558328 530596
rect 572260 530544 572312 530596
rect 25964 530476 26016 530528
rect 55496 530476 55548 530528
rect 173992 530476 174044 530528
rect 422484 530476 422536 530528
rect 542728 530476 542780 530528
rect 543648 530476 543700 530528
rect 553676 530476 553728 530528
rect 28264 530408 28316 530460
rect 53288 530408 53340 530460
rect 171876 530408 171928 530460
rect 424600 530408 424652 530460
rect 537300 530408 537352 530460
rect 551652 530408 551704 530460
rect 553308 530408 553360 530460
rect 554596 530408 554648 530460
rect 28356 530340 28408 530392
rect 51172 530340 51224 530392
rect 169760 530340 169812 530392
rect 426716 530340 426768 530392
rect 541624 530340 541676 530392
rect 553400 530340 553452 530392
rect 28540 530272 28592 530324
rect 48964 530272 49016 530324
rect 133052 530272 133104 530324
rect 463792 530272 463844 530324
rect 543648 530272 543700 530324
rect 552664 530272 552716 530324
rect 558184 530272 558236 530324
rect 559288 530272 559340 530324
rect 27160 530204 27212 530256
rect 46848 530204 46900 530256
rect 109316 530204 109368 530256
rect 111064 530204 111116 530256
rect 130936 530204 130988 530256
rect 465540 530204 465592 530256
rect 471704 530204 471756 530256
rect 481732 530204 481784 530256
rect 539508 530204 539560 530256
rect 554228 530204 554280 530256
rect 25596 530136 25648 530188
rect 44732 530136 44784 530188
rect 128728 530136 128780 530188
rect 467840 530136 467892 530188
rect 478880 530136 478932 530188
rect 493140 530136 493192 530188
rect 493968 530136 494020 530188
rect 554412 530136 554464 530188
rect 126612 530068 126664 530120
rect 469864 530068 469916 530120
rect 554504 530068 554556 530120
rect 124404 530000 124456 530052
rect 472072 530000 472124 530052
rect 482928 530000 482980 530052
rect 488540 530000 488592 530052
rect 556804 530000 556856 530052
rect 558276 530000 558328 530052
rect 122288 529932 122340 529984
rect 474188 529932 474240 529984
rect 481548 529932 481600 529984
rect 484952 529932 485004 529984
rect 560944 529932 560996 529984
rect 567936 529932 567988 529984
rect 431040 529864 431092 529916
rect 191288 529796 191340 529848
rect 405188 529796 405240 529848
rect 165436 529728 165488 529780
rect 179420 529728 179472 529780
rect 417056 529728 417108 529780
rect 160008 529660 160060 529712
rect 436468 529660 436520 529712
rect 157892 529592 157944 529644
rect 438952 529592 439004 529644
rect 151360 529524 151412 529576
rect 445116 529524 445168 529576
rect 149244 529456 149296 529508
rect 447324 529456 447376 529508
rect 147036 529388 147088 529440
rect 449440 529388 449492 529440
rect 144920 529320 144972 529372
rect 451556 529320 451608 529372
rect 111524 529252 111576 529304
rect 481548 529252 481600 529304
rect 108304 529184 108356 529236
rect 482928 529184 482980 529236
rect 142804 529116 142856 529168
rect 454040 529116 454092 529168
rect 140596 529048 140648 529100
rect 456202 529048 456254 529100
rect 138480 528980 138532 529032
rect 458318 528980 458370 529032
rect 136548 528912 136600 528964
rect 460204 528912 460256 528964
rect 134432 528844 134484 528896
rect 462320 528844 462372 528896
rect 120448 528776 120500 528828
rect 476304 528776 476356 528828
rect 117136 528708 117188 528760
rect 479616 528708 479668 528760
rect 114008 528640 114060 528692
rect 483020 528640 483072 528692
rect 110696 528572 110748 528624
rect 486056 528572 486108 528624
rect 315948 528504 316000 528556
rect 456064 528504 456116 528556
rect 194600 528436 194652 528488
rect 401968 528436 402020 528488
rect 190368 528368 190420 528420
rect 406292 528368 406344 528420
rect 186136 528300 186188 528352
rect 410616 528300 410668 528352
rect 115940 528232 115992 528284
rect 125324 528232 125376 528284
rect 181904 528232 181956 528284
rect 414940 528232 414992 528284
rect 118240 528164 118292 528216
rect 164516 528164 164568 528216
rect 169024 528164 169076 528216
rect 173256 528164 173308 528216
rect 423680 528164 423732 528216
rect 427820 528164 427872 528216
rect 432144 528164 432196 528216
rect 298100 527416 298152 527468
rect 302976 527416 303028 527468
rect 288532 527212 288584 527264
rect 296628 527212 296680 527264
rect 282920 514700 282972 514752
rect 283104 514700 283156 514752
rect 577596 509600 577648 509652
rect 579620 509600 579672 509652
rect 2872 509260 2924 509312
rect 14556 509260 14608 509312
rect 283104 509192 283156 509244
rect 416596 503004 416648 503056
rect 418160 503004 418212 503056
rect 418804 503004 418856 503056
rect 420276 503004 420328 503056
rect 413284 502936 413336 502988
rect 580356 502936 580408 502988
rect 481272 502868 481324 502920
rect 484308 502868 484360 502920
rect 487160 502868 487212 502920
rect 459468 502664 459520 502716
rect 461216 502664 461268 502716
rect 114560 502596 114612 502648
rect 115572 502596 115624 502648
rect 158720 501168 158772 501220
rect 159732 501168 159784 501220
rect 164240 501168 164292 501220
rect 165068 501168 165120 501220
rect 173900 501168 173952 501220
rect 174820 501168 174872 501220
rect 183652 501168 183704 501220
rect 184572 501168 184624 501220
rect 24216 500896 24268 500948
rect 25320 500896 25372 500948
rect 27528 500896 27580 500948
rect 29644 500896 29696 500948
rect 50068 500896 50120 500948
rect 50988 500896 51040 500948
rect 59820 500896 59872 500948
rect 60648 500896 60700 500948
rect 60832 500896 60884 500948
rect 61936 500896 61988 500948
rect 64052 500896 64104 500948
rect 64788 500896 64840 500948
rect 69480 500896 69532 500948
rect 70308 500896 70360 500948
rect 99656 500896 99708 500948
rect 100668 500896 100720 500948
rect 100760 500896 100812 500948
rect 102048 500896 102100 500948
rect 105084 500896 105136 500948
rect 106188 500896 106240 500948
rect 121460 500896 121512 500948
rect 153476 500896 153528 500948
rect 195244 500896 195296 500948
rect 197728 500896 197780 500948
rect 201684 500896 201736 500948
rect 203156 500896 203208 500948
rect 204628 500896 204680 500948
rect 208492 500896 208544 500948
rect 214656 500896 214708 500948
rect 217140 500896 217192 500948
rect 224868 500896 224920 500948
rect 225788 500896 225840 500948
rect 229100 500896 229152 500948
rect 230112 500896 230164 500948
rect 230572 500896 230624 500948
rect 232228 500896 232280 500948
rect 234528 500896 234580 500948
rect 235448 500896 235500 500948
rect 235908 500896 235960 500948
rect 236552 500896 236604 500948
rect 255320 500896 255372 500948
rect 256976 500896 257028 500948
rect 259460 500896 259512 500948
rect 261300 500896 261352 500948
rect 262312 500896 262364 500948
rect 263508 500896 263560 500948
rect 267924 500896 267976 500948
rect 268844 500896 268896 500948
rect 269120 500896 269172 500948
rect 269948 500896 270000 500948
rect 340144 500896 340196 500948
rect 340788 500896 340840 500948
rect 341156 500896 341208 500948
rect 342076 500896 342128 500948
rect 343180 500896 343232 500948
rect 343732 500896 343784 500948
rect 345480 500896 345532 500948
rect 346216 500896 346268 500948
rect 354128 500896 354180 500948
rect 354588 500896 354640 500948
rect 359464 500896 359516 500948
rect 360108 500896 360160 500948
rect 364892 500896 364944 500948
rect 365628 500896 365680 500948
rect 365996 500896 366048 500948
rect 367008 500896 367060 500948
rect 370320 500896 370372 500948
rect 371148 500896 371200 500948
rect 375656 500896 375708 500948
rect 376576 500896 376628 500948
rect 384304 500896 384356 500948
rect 384948 500896 385000 500948
rect 385408 500896 385460 500948
rect 386328 500896 386380 500948
rect 395068 500896 395120 500948
rect 395988 500896 396040 500948
rect 400496 500896 400548 500948
rect 401416 500896 401468 500948
rect 404728 500896 404780 500948
rect 411628 500896 411680 500948
rect 420828 500896 420880 500948
rect 423128 500896 423180 500948
rect 424968 500896 425020 500948
rect 427084 500896 427136 500948
rect 429292 500896 429344 500948
rect 431408 500896 431460 500948
rect 433432 500896 433484 500948
rect 435548 500896 435600 500948
rect 437572 500896 437624 500948
rect 439688 500896 439740 500948
rect 441988 500896 442040 500948
rect 444380 500896 444432 500948
rect 446312 500896 446364 500948
rect 448520 500896 448572 500948
rect 450452 500896 450504 500948
rect 453304 500896 453356 500948
rect 455328 500896 455380 500948
rect 457352 500896 457404 500948
rect 461860 500896 461912 500948
rect 464068 500896 464120 500948
rect 465908 500896 465960 500948
rect 468116 500896 468168 500948
rect 470232 500896 470284 500948
rect 472716 500896 472768 500948
rect 474648 500896 474700 500948
rect 477776 500896 477828 500948
rect 480812 500896 480864 500948
rect 492036 500896 492088 500948
rect 492588 500896 492640 500948
rect 498384 500896 498436 500948
rect 498936 500896 498988 500948
rect 502432 500896 502484 500948
rect 503260 500896 503312 500948
rect 509240 500896 509292 500948
rect 509792 500896 509844 500948
rect 511448 500896 511500 500948
rect 511908 500896 511960 500948
rect 522212 500896 522264 500948
rect 522948 500896 523000 500948
rect 527640 500896 527692 500948
rect 528376 500896 528428 500948
rect 531964 500896 532016 500948
rect 532608 500896 532660 500948
rect 533068 500896 533120 500948
rect 533988 500896 534040 500948
rect 536288 500896 536340 500948
rect 536748 500896 536800 500948
rect 541624 500896 541676 500948
rect 542268 500896 542320 500948
rect 545948 500896 546000 500948
rect 546408 500896 546460 500948
rect 547052 500896 547104 500948
rect 547788 500896 547840 500948
rect 553308 500896 553360 500948
rect 554044 500896 554096 500948
rect 558184 500896 558236 500948
rect 559288 500896 559340 500948
rect 31668 500828 31720 500880
rect 31760 500828 31812 500880
rect 45744 500828 45796 500880
rect 53932 500828 53984 500880
rect 126612 500828 126664 500880
rect 153384 500828 153436 500880
rect 195336 500828 195388 500880
rect 198832 500828 198884 500880
rect 200212 500828 200264 500880
rect 205272 500828 205324 500880
rect 205640 500828 205692 500880
rect 209596 500828 209648 500880
rect 213460 500828 213512 500880
rect 216036 500828 216088 500880
rect 251180 500828 251232 500880
rect 253756 500828 253808 500880
rect 253940 500828 253992 500880
rect 255964 500828 256016 500880
rect 260840 500828 260892 500880
rect 262404 500828 262456 500880
rect 403716 500828 403768 500880
rect 409880 500828 409932 500880
rect 129832 500760 129884 500812
rect 153292 500760 153344 500812
rect 214932 500760 214984 500812
rect 218244 500760 218296 500812
rect 355232 500760 355284 500812
rect 355968 500760 356020 500812
rect 554136 500760 554188 500812
rect 41420 500692 41472 500744
rect 47032 500692 47084 500744
rect 128728 500692 128780 500744
rect 151912 500692 151964 500744
rect 197176 500692 197228 500744
rect 202052 500692 202104 500744
rect 211344 500692 211396 500744
rect 215024 500692 215076 500744
rect 542728 500692 542780 500744
rect 551376 500692 551428 500744
rect 130936 500624 130988 500676
rect 154764 500624 154816 500676
rect 223488 500624 223540 500676
rect 224684 500624 224736 500676
rect 350908 500624 350960 500676
rect 351828 500624 351880 500676
rect 507124 500624 507176 500676
rect 507768 500624 507820 500676
rect 544844 500624 544896 500676
rect 127716 500556 127768 500608
rect 154488 500556 154540 500608
rect 201592 500556 201644 500608
rect 206376 500556 206428 500608
rect 215300 500556 215352 500608
rect 219256 500556 219308 500608
rect 219532 500556 219584 500608
rect 222568 500556 222620 500608
rect 533896 500556 533948 500608
rect 554228 500556 554280 500608
rect 124404 500488 124456 500540
rect 152004 500488 152056 500540
rect 196072 500488 196124 500540
rect 200948 500488 201000 500540
rect 363788 500488 363840 500540
rect 364248 500488 364300 500540
rect 523316 500488 523368 500540
rect 548156 500488 548208 500540
rect 549168 500488 549220 500540
rect 42524 500420 42576 500472
rect 47584 500420 47636 500472
rect 125508 500420 125560 500472
rect 153384 500420 153436 500472
rect 187792 500420 187844 500472
rect 192392 500420 192444 500472
rect 199476 500420 199528 500472
rect 204168 500420 204220 500472
rect 209872 500420 209924 500472
rect 213920 500420 213972 500472
rect 218152 500420 218204 500472
rect 221464 500420 221516 500472
rect 224224 500420 224276 500472
rect 226800 500420 226852 500472
rect 515772 500420 515824 500472
rect 551468 500420 551520 500472
rect 43628 500352 43680 500404
rect 48964 500352 49016 500404
rect 123392 500352 123444 500404
rect 153476 500352 153528 500404
rect 209136 500352 209188 500404
rect 212816 500352 212868 500404
rect 322848 500352 322900 500404
rect 323308 500352 323360 500404
rect 349804 500352 349856 500404
rect 350448 500352 350500 500404
rect 398288 500352 398340 500404
rect 398748 500352 398800 500404
rect 506112 500352 506164 500404
rect 512644 500352 512696 500404
rect 513656 500352 513708 500404
rect 551560 500352 551612 500404
rect 44732 500284 44784 500336
rect 52552 500284 52604 500336
rect 55496 500284 55548 500336
rect 56416 500284 56468 500336
rect 120264 500284 120316 500336
rect 153844 500284 153896 500336
rect 509056 500284 509108 500336
rect 551652 500284 551704 500336
rect 85672 500216 85724 500268
rect 112444 500216 112496 500268
rect 117320 500216 117372 500268
rect 153108 500216 153160 500268
rect 187884 500216 187936 500268
rect 193404 500216 193456 500268
rect 195612 500216 195664 500268
rect 279608 500216 279660 500268
rect 289728 500216 289780 500268
rect 416136 500216 416188 500268
rect 498568 500216 498620 500268
rect 499488 500216 499540 500268
rect 502892 500216 502944 500268
rect 551744 500216 551796 500268
rect 556804 500216 556856 500268
rect 571340 500216 571392 500268
rect 70584 500148 70636 500200
rect 131948 500148 132000 500200
rect 154396 500148 154448 500200
rect 549904 500148 549956 500200
rect 65156 500080 65208 500132
rect 66168 500080 66220 500132
rect 135260 500080 135312 500132
rect 154304 500080 154356 500132
rect 220820 500080 220872 500132
rect 223580 500080 223632 500132
rect 369216 500080 369268 500132
rect 369768 500080 369820 500132
rect 379980 500080 380032 500132
rect 380808 500080 380860 500132
rect 94504 500012 94556 500064
rect 137376 500012 137428 500064
rect 154120 500012 154172 500064
rect 191840 500012 191892 500064
rect 199936 500012 199988 500064
rect 501788 500012 501840 500064
rect 502248 500012 502300 500064
rect 516876 500012 516928 500064
rect 517428 500012 517480 500064
rect 140596 499944 140648 499996
rect 154212 499944 154264 499996
rect 360568 499944 360620 499996
rect 361488 499944 361540 499996
rect 374552 499944 374604 499996
rect 375288 499944 375340 499996
rect 378876 499944 378928 499996
rect 379428 499944 379480 499996
rect 389640 499944 389692 499996
rect 390468 499944 390520 499996
rect 393964 499944 394016 499996
rect 394608 499944 394660 499996
rect 399392 499944 399444 499996
rect 400128 499944 400180 499996
rect 526536 499944 526588 499996
rect 527088 499944 527140 499996
rect 537300 499944 537352 499996
rect 538128 499944 538180 499996
rect 139492 499876 139544 499928
rect 154028 499876 154080 499928
rect 223580 499876 223632 499928
rect 229008 499876 229060 499928
rect 388628 499876 388680 499928
rect 389088 499876 389140 499928
rect 141700 499808 141752 499860
rect 153936 499808 153988 499860
rect 344376 499808 344428 499860
rect 344928 499808 344980 499860
rect 493140 499808 493192 499860
rect 494704 499808 494756 499860
rect 517980 499808 518032 499860
rect 518808 499808 518860 499860
rect 22100 499740 22152 499792
rect 24124 499740 24176 499792
rect 51172 499740 51224 499792
rect 52368 499740 52420 499792
rect 66260 499740 66312 499792
rect 67548 499740 67600 499792
rect 142804 499740 142856 499792
rect 153660 499740 153712 499792
rect 191932 499740 191984 499792
rect 196624 499740 196676 499792
rect 233056 499740 233108 499792
rect 234344 499740 234396 499792
rect 259368 499740 259420 499792
rect 260288 499740 260340 499792
rect 263600 499740 263652 499792
rect 264520 499740 264572 499792
rect 549076 499740 549128 499792
rect 551284 499740 551336 499792
rect 24308 499672 24360 499724
rect 26332 499672 26384 499724
rect 143816 499672 143868 499724
rect 153568 499672 153620 499724
rect 206376 499672 206428 499724
rect 210700 499672 210752 499724
rect 26148 499604 26200 499656
rect 28540 499604 28592 499656
rect 103980 499604 104032 499656
rect 104808 499604 104860 499656
rect 203708 499604 203760 499656
rect 207480 499604 207532 499656
rect 207756 499604 207808 499656
rect 211712 499604 211764 499656
rect 216680 499604 216732 499656
rect 220360 499604 220412 499656
rect 252652 499604 252704 499656
rect 254860 499604 254912 499656
rect 271972 499604 272024 499656
rect 273168 499604 273220 499656
rect 25504 499536 25556 499588
rect 27436 499536 27488 499588
rect 31944 499536 31996 499588
rect 32864 499536 32916 499588
rect 34980 499536 35032 499588
rect 35808 499536 35860 499588
rect 36084 499536 36136 499588
rect 37096 499536 37148 499588
rect 40408 499536 40460 499588
rect 41328 499536 41380 499588
rect 75920 499536 75972 499588
rect 77208 499536 77260 499588
rect 79140 499536 79192 499588
rect 79968 499536 80020 499588
rect 80244 499536 80296 499588
rect 81256 499536 81308 499588
rect 84568 499536 84620 499588
rect 85488 499536 85540 499588
rect 86960 499536 87012 499588
rect 87788 499536 87840 499588
rect 88892 499536 88944 499588
rect 89628 499536 89680 499588
rect 89996 499536 90048 499588
rect 91008 499536 91060 499588
rect 94228 499536 94280 499588
rect 95148 499536 95200 499588
rect 95332 499536 95384 499588
rect 96528 499536 96580 499588
rect 144920 499536 144972 499588
rect 153752 499536 153804 499588
rect 230388 499536 230440 499588
rect 231124 499536 231176 499588
rect 247040 499536 247092 499588
rect 249432 499536 249484 499588
rect 256792 499536 256844 499588
rect 259184 499536 259236 499588
rect 266360 499536 266412 499588
rect 267832 499536 267884 499588
rect 277584 499536 277636 499588
rect 278596 499536 278648 499588
rect 283012 499579 283064 499588
rect 283012 499545 283021 499579
rect 283021 499545 283055 499579
rect 283055 499545 283064 499579
rect 283012 499536 283064 499545
rect 317328 499536 317380 499588
rect 317880 499536 317932 499588
rect 560944 499536 560996 499588
rect 567200 499536 567252 499588
rect 551468 499468 551520 499520
rect 551836 499468 551888 499520
rect 81348 498788 81400 498840
rect 113180 498788 113232 498840
rect 527824 498788 527876 498840
rect 574100 498788 574152 498840
rect 77024 497428 77076 497480
rect 106280 497428 106332 497480
rect 132500 497428 132552 497480
rect 154856 497428 154908 497480
rect 498384 497428 498436 497480
rect 553308 497428 553360 497480
rect 299388 496068 299440 496120
rect 414020 496068 414072 496120
rect 3516 495456 3568 495508
rect 298100 495456 298152 495508
rect 299388 495456 299440 495508
rect 320456 495456 320508 495508
rect 321100 495456 321152 495508
rect 283012 495388 283064 495440
rect 283196 495388 283248 495440
rect 13084 494708 13136 494760
rect 443644 494708 443696 494760
rect 502432 494708 502484 494760
rect 553216 494708 553268 494760
rect 190920 493960 190972 494012
rect 195336 493960 195388 494012
rect 196900 493960 196952 494012
rect 199476 493960 199528 494012
rect 200488 493960 200540 494012
rect 203708 493960 203760 494012
rect 205272 493960 205324 494012
rect 207756 493960 207808 494012
rect 213644 493960 213696 494012
rect 215300 493960 215352 494012
rect 216036 493960 216088 494012
rect 218152 493960 218204 494012
rect 231584 493960 231636 494012
rect 234528 493960 234580 494012
rect 235172 493960 235224 494012
rect 237564 493960 237616 494012
rect 241152 493960 241204 494012
rect 243084 493960 243136 494012
rect 245936 493960 245988 494012
rect 248420 493960 248472 494012
rect 256792 493960 256844 494012
rect 257896 493960 257948 494012
rect 259460 493960 259512 494012
rect 260288 493960 260340 494012
rect 266360 493960 266412 494012
rect 267464 493960 267516 494012
rect 226800 493892 226852 493944
rect 230388 493892 230440 493944
rect 232780 493892 232832 493944
rect 235908 493892 235960 493944
rect 201684 493824 201736 493876
rect 204628 493824 204680 493876
rect 210056 493824 210108 493876
rect 213460 493824 213512 493876
rect 219624 493824 219676 493876
rect 223488 493824 223540 493876
rect 229192 493824 229244 493876
rect 233148 493824 233200 493876
rect 237564 493824 237616 493876
rect 240140 493824 240192 493876
rect 236368 493756 236420 493808
rect 238760 493756 238812 493808
rect 248328 493756 248380 493808
rect 249800 493756 249852 493808
rect 206468 493688 206520 493740
rect 209136 493688 209188 493740
rect 212448 493688 212500 493740
rect 214932 493688 214984 493740
rect 193312 493620 193364 493672
rect 196072 493620 196124 493672
rect 204076 493620 204128 493672
rect 206376 493620 206428 493672
rect 211252 493620 211304 493672
rect 214656 493620 214708 493672
rect 222016 493620 222068 493672
rect 224224 493620 224276 493672
rect 198096 493552 198148 493604
rect 200212 493552 200264 493604
rect 218428 493552 218480 493604
rect 220820 493552 220872 493604
rect 225604 493552 225656 493604
rect 229008 493552 229060 493604
rect 230388 493552 230440 493604
rect 233056 493552 233108 493604
rect 233976 493552 234028 493604
rect 237288 493552 237340 493604
rect 194508 493484 194560 493536
rect 197176 493484 197228 493536
rect 217232 493484 217284 493536
rect 219532 493484 219584 493536
rect 239956 493484 240008 493536
rect 242808 493484 242860 493536
rect 202880 493416 202932 493468
rect 205640 493416 205692 493468
rect 207664 493416 207716 493468
rect 209872 493416 209924 493468
rect 220820 493416 220872 493468
rect 224868 493416 224920 493468
rect 238760 493416 238812 493468
rect 241520 493416 241572 493468
rect 243544 493416 243596 493468
rect 245660 493416 245712 493468
rect 74540 493348 74592 493400
rect 102140 493348 102192 493400
rect 189724 493348 189776 493400
rect 195244 493348 195296 493400
rect 86960 493280 87012 493332
rect 124220 493280 124272 493332
rect 199292 493280 199344 493332
rect 201592 493280 201644 493332
rect 244740 493280 244792 493332
rect 247224 493280 247276 493332
rect 249524 493280 249576 493332
rect 251272 493280 251324 493332
rect 509240 493280 509292 493332
rect 553124 493280 553176 493332
rect 214840 493212 214892 493264
rect 216680 493212 216732 493264
rect 242348 493212 242400 493264
rect 244280 493212 244332 493264
rect 195704 493144 195756 493196
rect 201868 493144 201920 493196
rect 208860 493144 208912 493196
rect 211344 493144 211396 493196
rect 256700 493144 256752 493196
rect 257988 493144 258040 493196
rect 277584 493144 277636 493196
rect 279424 493144 279476 493196
rect 188620 493008 188672 493060
rect 191932 493008 191984 493060
rect 227996 493008 228048 493060
rect 230572 493008 230624 493060
rect 250720 492940 250772 492992
rect 252744 492940 252796 492992
rect 223212 492872 223264 492924
rect 227904 492872 227956 492924
rect 271972 492804 272024 492856
rect 273444 492804 273496 492856
rect 223580 492736 223632 492788
rect 224408 492736 224460 492788
rect 282920 492600 282972 492652
rect 283196 492600 283248 492652
rect 320272 492600 320324 492652
rect 320732 492600 320784 492652
rect 73068 491988 73120 492040
rect 99012 491988 99064 492040
rect 84108 491920 84160 491972
rect 117136 491920 117188 491972
rect 495348 491920 495400 491972
rect 555700 491920 555752 491972
rect 94504 491240 94556 491292
rect 95700 491240 95752 491292
rect 68928 490628 68980 490680
rect 92112 490628 92164 490680
rect 79968 490560 80020 490612
rect 109960 490560 110012 490612
rect 112444 490560 112496 490612
rect 120724 490560 120776 490612
rect 499488 490560 499540 490612
rect 555976 490560 556028 490612
rect 551468 489880 551520 489932
rect 551836 489880 551888 489932
rect 35808 489812 35860 489864
rect 36544 489812 36596 489864
rect 61936 489812 61988 489864
rect 79508 489812 79560 489864
rect 95148 489812 95200 489864
rect 135076 489812 135128 489864
rect 62028 489744 62080 489796
rect 81348 489744 81400 489796
rect 90916 489744 90968 489796
rect 129740 489744 129792 489796
rect 64788 489676 64840 489728
rect 84936 489676 84988 489728
rect 96528 489676 96580 489728
rect 136916 489676 136968 489728
rect 49608 489608 49660 489660
rect 59820 489608 59872 489660
rect 63408 489608 63460 489660
rect 83096 489608 83148 489660
rect 97908 489608 97960 489660
rect 140504 489608 140556 489660
rect 50988 489540 51040 489592
rect 61660 489540 61712 489592
rect 66168 489540 66220 489592
rect 86684 489540 86736 489592
rect 96436 489540 96488 489592
rect 138664 489540 138716 489592
rect 52368 489472 52420 489524
rect 63408 489472 63460 489524
rect 67548 489472 67600 489524
rect 88524 489472 88576 489524
rect 102048 489472 102100 489524
rect 145840 489472 145892 489524
rect 53748 489404 53800 489456
rect 66996 489404 67048 489456
rect 67456 489404 67508 489456
rect 90272 489404 90324 489456
rect 100668 489404 100720 489456
rect 144092 489404 144144 489456
rect 52276 489336 52328 489388
rect 65156 489336 65208 489388
rect 70308 489336 70360 489388
rect 93860 489336 93912 489388
rect 99288 489336 99340 489388
rect 142252 489336 142304 489388
rect 56416 489268 56468 489320
rect 70584 489268 70636 489320
rect 71688 489268 71740 489320
rect 97448 489268 97500 489320
rect 103428 489268 103480 489320
rect 149428 489268 149480 489320
rect 37096 489200 37148 489252
rect 38292 489200 38344 489252
rect 48228 489200 48280 489252
rect 58072 489200 58124 489252
rect 59268 489200 59320 489252
rect 75920 489200 75972 489252
rect 77208 489200 77260 489252
rect 104624 489200 104676 489252
rect 104808 489200 104860 489252
rect 151268 489200 151320 489252
rect 37188 489132 37240 489184
rect 40132 489132 40184 489184
rect 46848 489132 46900 489184
rect 56232 489132 56284 489184
rect 56508 489132 56560 489184
rect 72332 489132 72384 489184
rect 74448 489132 74500 489184
rect 101036 489132 101088 489184
rect 101956 489132 102008 489184
rect 147680 489132 147732 489184
rect 60648 489064 60700 489116
rect 77760 489064 77812 489116
rect 93768 489064 93820 489116
rect 133328 489064 133380 489116
rect 57888 488996 57940 489048
rect 74172 488996 74224 489048
rect 92388 488996 92440 489048
rect 131488 488996 131540 489048
rect 55128 488928 55180 488980
rect 68744 488928 68796 488980
rect 89628 488928 89680 488980
rect 126152 488928 126204 488980
rect 91008 488860 91060 488912
rect 127900 488860 127952 488912
rect 86868 488792 86920 488844
rect 122564 488792 122616 488844
rect 20352 488724 20404 488776
rect 24216 488724 24268 488776
rect 39948 488724 40000 488776
rect 43720 488724 43772 488776
rect 85488 488724 85540 488776
rect 118976 488724 119028 488776
rect 16856 488656 16908 488708
rect 22284 488656 22336 488708
rect 38568 488656 38620 488708
rect 41880 488656 41932 488708
rect 82728 488656 82780 488708
rect 115388 488656 115440 488708
rect 22192 488588 22244 488640
rect 24308 488588 24360 488640
rect 48964 488588 49016 488640
rect 50896 488588 50948 488640
rect 81256 488588 81308 488640
rect 111800 488588 111852 488640
rect 18604 488520 18656 488572
rect 23480 488520 23532 488572
rect 23940 488520 23992 488572
rect 25504 488520 25556 488572
rect 29368 488520 29420 488572
rect 30288 488520 30340 488572
rect 41328 488520 41380 488572
rect 45468 488520 45520 488572
rect 47584 488520 47636 488572
rect 49056 488520 49108 488572
rect 78588 488520 78640 488572
rect 108212 488520 108264 488572
rect 24124 486412 24176 486464
rect 156052 486412 156104 486464
rect 505008 486412 505060 486464
rect 555240 486412 555292 486464
rect 3424 485052 3476 485104
rect 185584 485052 185636 485104
rect 521568 483692 521620 483744
rect 552664 483692 552716 483744
rect 511908 483624 511960 483676
rect 555148 483624 555200 483676
rect 528376 482264 528428 482316
rect 552388 482264 552440 482316
rect 529848 481040 529900 481092
rect 555792 481040 555844 481092
rect 520188 480972 520240 481024
rect 554596 480972 554648 481024
rect 517428 480904 517480 480956
rect 551008 480904 551060 480956
rect 551468 480904 551520 480956
rect 553032 480768 553084 480820
rect 3148 480224 3200 480276
rect 14464 480224 14516 480276
rect 183652 480224 183704 480276
rect 183836 480224 183888 480276
rect 525708 479612 525760 479664
rect 552480 479612 552532 479664
rect 527088 479544 527140 479596
rect 554504 479544 554556 479596
rect 494704 479476 494756 479528
rect 554780 479476 554832 479528
rect 542268 478388 542320 478440
rect 553676 478388 553728 478440
rect 540888 478320 540940 478372
rect 555608 478320 555660 478372
rect 532608 478252 532660 478304
rect 552848 478252 552900 478304
rect 522948 478184 523000 478236
rect 551192 478184 551244 478236
rect 496728 478116 496780 478168
rect 555884 478116 555936 478168
rect 344928 477436 344980 477488
rect 346032 477436 346084 477488
rect 353208 477436 353260 477488
rect 355784 477436 355836 477488
rect 369768 477436 369820 477488
rect 374092 477436 374144 477488
rect 354588 477368 354640 477420
rect 356980 477368 357032 477420
rect 378048 477368 378100 477420
rect 383844 477368 383896 477420
rect 390468 477300 390520 477352
rect 397276 477300 397328 477352
rect 395988 477232 396040 477284
rect 403440 477232 403492 477284
rect 362868 477164 362920 477216
rect 366732 477164 366784 477216
rect 383568 477164 383620 477216
rect 390008 477164 390060 477216
rect 391848 477164 391900 477216
rect 399760 477164 399812 477216
rect 400128 477164 400180 477216
rect 408316 477164 408368 477216
rect 375288 477096 375340 477148
rect 380164 477096 380216 477148
rect 386328 477028 386380 477080
rect 392400 477028 392452 477080
rect 393228 477028 393280 477080
rect 400956 477028 401008 477080
rect 401416 477028 401468 477080
rect 409512 477028 409564 477080
rect 546408 477028 546460 477080
rect 553584 477028 553636 477080
rect 317880 476960 317932 477012
rect 318708 476960 318760 477012
rect 319076 476960 319128 477012
rect 320088 476960 320140 477012
rect 364248 476960 364300 477012
rect 368020 476960 368072 477012
rect 371148 476960 371200 477012
rect 375288 476960 375340 477012
rect 376576 476960 376628 477012
rect 381452 476960 381504 477012
rect 382188 476960 382240 477012
rect 388720 476960 388772 477012
rect 389088 476960 389140 477012
rect 396080 476960 396132 477012
rect 397368 476960 397420 477012
rect 405832 476960 405884 477012
rect 536748 476960 536800 477012
rect 552572 476960 552624 477012
rect 351828 476892 351880 476944
rect 353300 476892 353352 476944
rect 355876 476892 355928 476944
rect 359464 476892 359516 476944
rect 361396 476892 361448 476944
rect 365536 476892 365588 476944
rect 372528 476892 372580 476944
rect 377772 476892 377824 476944
rect 380808 476892 380860 476944
rect 386328 476892 386380 476944
rect 398748 476892 398800 476944
rect 407120 476892 407172 476944
rect 535368 476892 535420 476944
rect 554320 476892 554372 476944
rect 332600 476824 332652 476876
rect 333796 476824 333848 476876
rect 335360 476824 335412 476876
rect 336188 476824 336240 476876
rect 336648 476824 336700 476876
rect 337476 476824 337528 476876
rect 342168 476824 342220 476876
rect 343548 476824 343600 476876
rect 346216 476824 346268 476876
rect 347228 476824 347280 476876
rect 350448 476824 350500 476876
rect 352104 476824 352156 476876
rect 355968 476824 356020 476876
rect 358176 476824 358228 476876
rect 358728 476824 358780 476876
rect 361856 476824 361908 476876
rect 365628 476824 365680 476876
rect 369216 476824 369268 476876
rect 373908 476824 373960 476876
rect 378968 476824 379020 476876
rect 380716 476824 380768 476876
rect 387524 476824 387576 476876
rect 390376 476824 390428 476876
rect 398564 476824 398616 476876
rect 401508 476824 401560 476876
rect 410708 476824 410760 476876
rect 524328 476824 524380 476876
rect 551836 476824 551888 476876
rect 351736 476756 351788 476808
rect 354588 476756 354640 476808
rect 371056 476756 371108 476808
rect 376576 476756 376628 476808
rect 386236 476756 386288 476808
rect 393688 476756 393740 476808
rect 395896 476756 395948 476808
rect 404636 476756 404688 476808
rect 492588 476756 492640 476808
rect 552112 476756 552164 476808
rect 361488 476688 361540 476740
rect 364340 476688 364392 476740
rect 368388 476688 368440 476740
rect 372896 476688 372948 476740
rect 394608 476688 394660 476740
rect 402244 476688 402296 476740
rect 367008 476620 367060 476672
rect 370412 476620 370464 476672
rect 316684 476552 316736 476604
rect 317328 476552 317380 476604
rect 333980 476552 334032 476604
rect 334992 476552 335044 476604
rect 349068 476552 349120 476604
rect 350908 476552 350960 476604
rect 357348 476552 357400 476604
rect 360660 476552 360712 476604
rect 366916 476552 366968 476604
rect 371608 476552 371660 476604
rect 360108 476484 360160 476536
rect 363052 476484 363104 476536
rect 331404 476416 331456 476468
rect 332508 476416 332560 476468
rect 387708 476416 387760 476468
rect 394884 476416 394936 476468
rect 347688 476348 347740 476400
rect 349620 476348 349672 476400
rect 346308 476280 346360 476332
rect 348424 476280 348476 476332
rect 379428 476280 379480 476332
rect 385132 476280 385184 476332
rect 376668 476212 376720 476264
rect 382648 476212 382700 476264
rect 384948 476212 385000 476264
rect 391204 476212 391256 476264
rect 550548 475804 550600 475856
rect 553400 475804 553452 475856
rect 549168 475668 549220 475720
rect 553768 475668 553820 475720
rect 543648 475600 543700 475652
rect 553860 475600 553912 475652
rect 538036 475532 538088 475584
rect 555056 475532 555108 475584
rect 531228 475464 531280 475516
rect 554412 475464 554464 475516
rect 499304 475396 499356 475448
rect 527824 475396 527876 475448
rect 528468 475396 528520 475448
rect 552940 475396 552992 475448
rect 518716 475328 518768 475380
rect 555424 475328 555476 475380
rect 287704 474648 287756 474700
rect 551928 474648 551980 474700
rect 550916 474580 550968 474632
rect 553492 474580 553544 474632
rect 549904 474512 549956 474564
rect 555332 474512 555384 474564
rect 538128 474308 538180 474360
rect 552296 474308 552348 474360
rect 539508 474240 539560 474292
rect 553952 474240 554004 474292
rect 533988 474172 534040 474224
rect 552756 474172 552808 474224
rect 518808 474104 518860 474156
rect 552204 474104 552256 474156
rect 512644 474036 512696 474088
rect 556068 474036 556120 474088
rect 502248 473968 502300 474020
rect 554964 473968 555016 474020
rect 551192 473492 551244 473544
rect 551928 473492 551980 473544
rect 546592 473467 546644 473476
rect 546592 473433 546601 473467
rect 546601 473433 546635 473467
rect 546635 473433 546644 473467
rect 546592 473424 546644 473433
rect 547788 473424 547840 473476
rect 551008 473424 551060 473476
rect 551468 473424 551520 473476
rect 554780 471996 554832 472048
rect 283104 471928 283156 471980
rect 283288 471928 283340 471980
rect 551652 471903 551704 471912
rect 551652 471869 551661 471903
rect 551661 471869 551695 471903
rect 551695 471869 551704 471903
rect 551652 471860 551704 471869
rect 551468 471724 551520 471776
rect 552756 471563 552808 471572
rect 552756 471529 552765 471563
rect 552765 471529 552799 471563
rect 552799 471529 552808 471563
rect 552756 471520 552808 471529
rect 552940 471520 552992 471572
rect 551744 471384 551796 471436
rect 552112 471384 552164 471436
rect 552296 471384 552348 471436
rect 552480 471384 552532 471436
rect 552756 471384 552808 471436
rect 552940 471384 552992 471436
rect 553308 471384 553360 471436
rect 553124 471248 553176 471300
rect 553308 471248 553360 471300
rect 552480 471180 552532 471232
rect 552572 471180 552624 471232
rect 552848 471180 552900 471232
rect 553124 471155 553176 471164
rect 553124 471121 553133 471155
rect 553133 471121 553167 471155
rect 553167 471121 553176 471155
rect 553124 471112 553176 471121
rect 552756 470951 552808 470960
rect 552756 470917 552765 470951
rect 552765 470917 552799 470951
rect 552799 470917 552808 470951
rect 552756 470908 552808 470917
rect 554228 470364 554280 470416
rect 555700 470364 555752 470416
rect 552940 468503 552992 468512
rect 552940 468469 552949 468503
rect 552949 468469 552983 468503
rect 552983 468469 552992 468503
rect 552940 468460 552992 468469
rect 554136 467576 554188 467628
rect 555976 467576 556028 467628
rect 551652 467440 551704 467492
rect 551744 467347 551796 467356
rect 551744 467313 551753 467347
rect 551753 467313 551787 467347
rect 551787 467313 551796 467347
rect 551744 467304 551796 467313
rect 552204 466964 552256 467016
rect 552480 466964 552532 467016
rect 552480 466828 552532 466880
rect 552756 466828 552808 466880
rect 552756 466692 552808 466744
rect 553124 466692 553176 466744
rect 554688 464992 554740 465044
rect 555884 464992 555936 465044
rect 279700 463632 279752 463684
rect 313280 463632 313332 463684
rect 551744 463564 551796 463616
rect 553032 463564 553084 463616
rect 551744 463360 551796 463412
rect 553032 463360 553084 463412
rect 563704 462340 563756 462392
rect 580172 462340 580224 462392
rect 283104 462315 283156 462324
rect 283104 462281 283113 462315
rect 283113 462281 283147 462315
rect 283147 462281 283156 462315
rect 283104 462272 283156 462281
rect 552848 461796 552900 461848
rect 553216 461796 553268 461848
rect 552940 461728 552992 461780
rect 551744 461388 551796 461440
rect 552848 461388 552900 461440
rect 552940 461388 552992 461440
rect 183652 460912 183704 460964
rect 183836 460912 183888 460964
rect 552756 459688 552808 459740
rect 554044 459552 554096 459604
rect 554964 459552 555016 459604
rect 552756 459484 552808 459536
rect 551928 456492 551980 456544
rect 552112 456492 552164 456544
rect 551836 455268 551888 455320
rect 552112 455268 552164 455320
rect 283196 452616 283248 452668
rect 3424 451256 3476 451308
rect 11704 451256 11756 451308
rect 283012 447108 283064 447160
rect 283196 447108 283248 447160
rect 9128 444320 9180 444372
rect 12532 444320 12584 444372
rect 183652 441600 183704 441652
rect 183836 441600 183888 441652
rect 283012 437520 283064 437572
rect 554964 437316 555016 437368
rect 557724 437316 557776 437368
rect 554780 437112 554832 437164
rect 557632 437112 557684 437164
rect 554872 436024 554924 436076
rect 560300 436024 560352 436076
rect 554780 435956 554832 436008
rect 558184 435956 558236 436008
rect 282920 434843 282972 434852
rect 282920 434809 282929 434843
rect 282929 434809 282963 434843
rect 282963 434809 282972 434843
rect 282920 434800 282972 434809
rect 554780 434664 554832 434716
rect 561680 434664 561732 434716
rect 554872 434596 554924 434648
rect 561956 434596 562008 434648
rect 282920 433279 282972 433288
rect 282920 433245 282929 433279
rect 282929 433245 282963 433279
rect 282963 433245 282972 433279
rect 282920 433236 282972 433245
rect 554872 433236 554924 433288
rect 564440 433236 564492 433288
rect 554780 433168 554832 433220
rect 563060 433168 563112 433220
rect 554964 431876 555016 431928
rect 567292 431876 567344 431928
rect 554780 431808 554832 431860
rect 565820 431808 565872 431860
rect 554872 431740 554924 431792
rect 560944 431740 560996 431792
rect 554872 430516 554924 430568
rect 569960 430516 570012 430568
rect 554780 430448 554832 430500
rect 568580 430448 568632 430500
rect 554780 429088 554832 429140
rect 571616 429088 571668 429140
rect 554872 428884 554924 428936
rect 556804 428884 556856 428936
rect 554780 427728 554832 427780
rect 572720 427728 572772 427780
rect 314660 426368 314712 426420
rect 499304 426368 499356 426420
rect 289636 425688 289688 425740
rect 314660 425688 314712 425740
rect 3516 423648 3568 423700
rect 13084 423648 13136 423700
rect 283012 423648 283064 423700
rect 183652 422288 183704 422340
rect 183836 422288 183888 422340
rect 281632 421540 281684 421592
rect 282276 421540 282328 421592
rect 292580 421540 292632 421592
rect 304356 415420 304408 415472
rect 580172 415420 580224 415472
rect 283104 415395 283156 415404
rect 283104 415361 283113 415395
rect 283113 415361 283147 415395
rect 283147 415361 283156 415395
rect 283104 415352 283156 415361
rect 283196 405696 283248 405748
rect 183652 402976 183704 403028
rect 183836 402976 183888 403028
rect 283196 402296 283248 402348
rect 143448 401548 143500 401600
rect 153660 401548 153712 401600
rect 142068 401480 142120 401532
rect 153936 401480 153988 401532
rect 140688 401412 140740 401464
rect 154028 401412 154080 401464
rect 140596 401344 140648 401396
rect 154212 401344 154264 401396
rect 137928 401276 137980 401328
rect 154120 401276 154172 401328
rect 136456 401208 136508 401260
rect 154304 401208 154356 401260
rect 133788 401140 133840 401192
rect 154856 401140 154908 401192
rect 132408 401072 132460 401124
rect 154396 401072 154448 401124
rect 128268 401004 128320 401056
rect 154488 401004 154540 401056
rect 121276 400936 121328 400988
rect 153844 400936 153896 400988
rect 118608 400868 118660 400920
rect 153108 400868 153160 400920
rect 144828 400800 144880 400852
rect 153568 400800 153620 400852
rect 146116 400460 146168 400512
rect 153752 400460 153804 400512
rect 77944 396584 77996 396636
rect 183652 383664 183704 383716
rect 183836 383664 183888 383716
rect 282276 377000 282328 377052
rect 284300 377000 284352 377052
rect 304448 368500 304500 368552
rect 580172 368500 580224 368552
rect 183652 364352 183704 364404
rect 183836 364352 183888 364404
rect 282276 360136 282328 360188
rect 282552 360136 282604 360188
rect 187792 358300 187844 358352
rect 191932 358300 191984 358352
rect 187884 358096 187936 358148
rect 193312 358096 193364 358148
rect 282552 357348 282604 357400
rect 194416 355988 194468 356040
rect 198924 355988 198976 356040
rect 201408 355988 201460 356040
rect 206928 355988 206980 356040
rect 210332 355988 210384 356040
rect 214748 355988 214800 356040
rect 215208 355988 215260 356040
rect 218980 355988 219032 356040
rect 221280 355988 221332 356040
rect 223212 355988 223264 356040
rect 226156 355988 226208 356040
rect 226984 355988 227036 356040
rect 233148 355988 233200 356040
rect 233700 355988 233752 356040
rect 234528 355988 234580 356040
rect 235908 355988 235960 356040
rect 239588 355988 239640 356040
rect 240508 355988 240560 356040
rect 242072 355988 242124 356040
rect 242900 355988 242952 356040
rect 258080 355988 258132 356040
rect 258540 355988 258592 356040
rect 261576 355988 261628 356040
rect 262220 355988 262272 356040
rect 262680 355988 262732 356040
rect 263600 355988 263652 356040
rect 191748 355920 191800 355972
rect 198648 355920 198700 355972
rect 200488 355920 200540 355972
rect 206100 355920 206152 355972
rect 222108 355920 222160 355972
rect 225420 355920 225472 355972
rect 232320 355920 232372 355972
rect 234068 355920 234120 355972
rect 193128 355852 193180 355904
rect 199660 355852 199712 355904
rect 204168 355852 204220 355904
rect 209228 355852 209280 355904
rect 213828 355852 213880 355904
rect 218060 355852 218112 355904
rect 220084 355852 220136 355904
rect 223672 355852 223724 355904
rect 231032 355852 231084 355904
rect 233148 355852 233200 355904
rect 211528 355784 211580 355836
rect 215668 355784 215720 355836
rect 229836 355784 229888 355836
rect 230480 355784 230532 355836
rect 235816 355784 235868 355836
rect 237288 355784 237340 355836
rect 240876 355784 240928 355836
rect 241704 355784 241756 355836
rect 199292 355716 199344 355768
rect 204996 355716 205048 355768
rect 209044 355716 209096 355768
rect 214012 355716 214064 355768
rect 198096 355648 198148 355700
rect 203892 355648 203944 355700
rect 217600 355648 217652 355700
rect 221188 355648 221240 355700
rect 255320 355648 255372 355700
rect 256056 355648 256108 355700
rect 196808 355580 196860 355632
rect 201500 355580 201552 355632
rect 218888 355512 218940 355564
rect 222384 355512 222436 355564
rect 224868 355512 224920 355564
rect 227720 355512 227772 355564
rect 263416 355512 263468 355564
rect 264612 355512 264664 355564
rect 207848 355376 207900 355428
rect 212632 355376 212684 355428
rect 227444 355376 227496 355428
rect 228824 355376 228876 355428
rect 256700 355376 256752 355428
rect 257344 355376 257396 355428
rect 266084 355376 266136 355428
rect 267096 355376 267148 355428
rect 243268 355308 243320 355360
rect 243820 355308 243872 355360
rect 244096 355308 244148 355360
rect 244924 355308 244976 355360
rect 264888 355240 264940 355292
rect 265900 355240 265952 355292
rect 202788 355172 202840 355224
rect 208308 355172 208360 355224
rect 254124 355104 254176 355156
rect 254860 355104 254912 355156
rect 268200 355104 268252 355156
rect 269488 355104 269540 355156
rect 212356 354968 212408 355020
rect 216772 354968 216824 355020
rect 237196 354968 237248 355020
rect 238300 354968 238352 355020
rect 189540 354832 189592 354884
rect 193680 354832 193732 354884
rect 190368 354764 190420 354816
rect 193864 354764 193916 354816
rect 206652 354764 206704 354816
rect 211436 354764 211488 354816
rect 223396 354764 223448 354816
rect 226524 354764 226576 354816
rect 238392 354764 238444 354816
rect 239404 354764 239456 354816
rect 248052 354764 248104 354816
rect 248604 354764 248656 354816
rect 188344 354696 188396 354748
rect 195244 354696 195296 354748
rect 195612 354696 195664 354748
rect 201408 354696 201460 354748
rect 205364 354696 205416 354748
rect 210332 354696 210384 354748
rect 216404 354696 216456 354748
rect 220084 354696 220136 354748
rect 228640 354696 228692 354748
rect 230388 354696 230440 354748
rect 260564 354696 260616 354748
rect 261024 354696 261076 354748
rect 267096 354696 267148 354748
rect 268292 354696 268344 354748
rect 278780 354696 278832 354748
rect 280528 354696 280580 354748
rect 46848 354628 46900 354680
rect 58532 354628 58584 354680
rect 48320 354560 48372 354612
rect 59636 354560 59688 354612
rect 29920 354492 29972 354544
rect 35808 354492 35860 354544
rect 45468 354492 45520 354544
rect 57520 354492 57572 354544
rect 34980 354424 35032 354476
rect 40040 354424 40092 354476
rect 47860 354424 47912 354476
rect 59360 354424 59412 354476
rect 35624 354356 35676 354408
rect 40224 354356 40276 354408
rect 46480 354356 46532 354408
rect 58072 354356 58124 354408
rect 38384 354288 38436 354340
rect 48596 354288 48648 354340
rect 49332 354288 49384 354340
rect 64972 354288 65024 354340
rect 39948 354220 40000 354272
rect 50988 354220 51040 354272
rect 52920 354220 52972 354272
rect 70400 354220 70452 354272
rect 41236 354152 41288 354204
rect 53012 354152 53064 354204
rect 55772 354152 55824 354204
rect 74724 354152 74776 354204
rect 25596 354084 25648 354136
rect 29276 354084 29328 354136
rect 32772 354084 32824 354136
rect 38200 354084 38252 354136
rect 42708 354084 42760 354136
rect 55128 354084 55180 354136
rect 58624 354084 58676 354136
rect 78772 354084 78824 354136
rect 26148 354016 26200 354068
rect 30380 354016 30432 354068
rect 34244 354016 34296 354068
rect 39212 354016 39264 354068
rect 45008 354016 45060 354068
rect 56784 354016 56836 354068
rect 61568 354016 61620 354068
rect 83188 354016 83240 354068
rect 44088 353948 44140 354000
rect 57244 353948 57296 354000
rect 64420 353948 64472 354000
rect 87420 353948 87472 354000
rect 39304 353880 39356 353932
rect 49700 353880 49752 353932
rect 50712 353880 50764 353932
rect 62212 353880 62264 353932
rect 33416 353812 33468 353864
rect 38660 353812 38712 353864
rect 51448 353812 51500 353864
rect 63500 353812 63552 353864
rect 30288 353676 30340 353728
rect 34520 353676 34572 353728
rect 37096 353676 37148 353728
rect 42248 353676 42300 353728
rect 43536 353676 43588 353728
rect 56140 353676 56192 353728
rect 28908 353608 28960 353660
rect 34428 353608 34480 353660
rect 42156 353608 42208 353660
rect 54116 353608 54168 353660
rect 27068 353540 27120 353592
rect 31852 353540 31904 353592
rect 40684 353540 40736 353592
rect 51908 353540 51960 353592
rect 24768 353472 24820 353524
rect 28172 353472 28224 353524
rect 31668 353472 31720 353524
rect 37188 353472 37240 353524
rect 50068 353472 50120 353524
rect 62120 353472 62172 353524
rect 22008 353404 22060 353456
rect 23940 353404 23992 353456
rect 24216 353404 24268 353456
rect 27068 353404 27120 353456
rect 31392 353404 31444 353456
rect 37096 353404 37148 353456
rect 21272 353336 21324 353388
rect 22836 353336 22888 353388
rect 23388 353336 23440 353388
rect 26240 353336 26292 353388
rect 28448 353336 28500 353388
rect 33508 353336 33560 353388
rect 36360 353336 36412 353388
rect 41604 353336 41656 353388
rect 20628 353268 20680 353320
rect 22192 353268 22244 353320
rect 22744 353268 22796 353320
rect 25044 353268 25096 353320
rect 27528 353268 27580 353320
rect 32588 353268 32640 353320
rect 37832 353268 37884 353320
rect 42800 353268 42852 353320
rect 54300 353268 54352 353320
rect 57888 353268 57940 353320
rect 57888 352792 57940 352844
rect 72424 352792 72476 352844
rect 57336 352724 57388 352776
rect 76748 352724 76800 352776
rect 60096 352656 60148 352708
rect 80980 352656 81032 352708
rect 62948 352588 63000 352640
rect 85580 352588 85632 352640
rect 65800 352520 65852 352572
rect 89720 352520 89772 352572
rect 37188 351840 37240 351892
rect 39028 351840 39080 351892
rect 56784 351840 56836 351892
rect 58348 351840 58400 351892
rect 62120 351840 62172 351892
rect 66352 351840 66404 351892
rect 68008 351840 68060 351892
rect 92940 351840 92992 351892
rect 198924 351840 198976 351892
rect 200580 351840 200632 351892
rect 274548 351840 274600 351892
rect 276848 351840 276900 351892
rect 58072 351772 58124 351824
rect 60740 351772 60792 351824
rect 68744 351772 68796 351824
rect 94044 351772 94096 351824
rect 275744 351772 275796 351824
rect 278044 351772 278096 351824
rect 59360 351704 59412 351756
rect 62764 351704 62816 351756
rect 70124 351704 70176 351756
rect 96068 351704 96120 351756
rect 276664 351704 276716 351756
rect 279332 351704 279384 351756
rect 42800 351636 42852 351688
rect 47676 351636 47728 351688
rect 62212 351636 62264 351688
rect 66996 351636 67048 351688
rect 70860 351636 70912 351688
rect 97172 351636 97224 351688
rect 277768 351636 277820 351688
rect 278780 351636 278832 351688
rect 58532 351568 58584 351620
rect 61660 351568 61712 351620
rect 69388 351568 69440 351620
rect 95240 351568 95292 351620
rect 278688 351568 278740 351620
rect 281724 351568 281776 351620
rect 59636 351500 59688 351552
rect 63684 351500 63736 351552
rect 73712 351500 73764 351552
rect 101404 351500 101456 351552
rect 271328 351500 271380 351552
rect 273352 351500 273404 351552
rect 57520 351432 57572 351484
rect 59452 351432 59504 351484
rect 71596 351432 71648 351484
rect 98276 351432 98328 351484
rect 114008 351432 114060 351484
rect 114468 351432 114520 351484
rect 115112 351432 115164 351484
rect 115756 351432 115808 351484
rect 118148 351432 118200 351484
rect 118608 351432 118660 351484
rect 133328 351432 133380 351484
rect 133788 351432 133840 351484
rect 138848 351432 138900 351484
rect 139308 351432 139360 351484
rect 143080 351432 143132 351484
rect 143448 351432 143500 351484
rect 145288 351432 145340 351484
rect 146116 351432 146168 351484
rect 155960 351432 156012 351484
rect 156420 351432 156472 351484
rect 160100 351432 160152 351484
rect 160836 351432 160888 351484
rect 161480 351432 161532 351484
rect 161940 351432 161992 351484
rect 165620 351432 165672 351484
rect 166172 351432 166224 351484
rect 169852 351432 169904 351484
rect 170404 351432 170456 351484
rect 171140 351432 171192 351484
rect 171600 351432 171652 351484
rect 175280 351432 175332 351484
rect 175924 351432 175976 351484
rect 176660 351432 176712 351484
rect 177120 351432 177172 351484
rect 179604 351432 179656 351484
rect 180156 351432 180208 351484
rect 180800 351432 180852 351484
rect 181260 351432 181312 351484
rect 184940 351432 184992 351484
rect 185492 351432 185544 351484
rect 193680 351432 193732 351484
rect 196348 351432 196400 351484
rect 269028 351432 269080 351484
rect 270500 351432 270552 351484
rect 273076 351432 273128 351484
rect 275652 351432 275704 351484
rect 40040 351364 40092 351416
rect 43260 351364 43312 351416
rect 63500 351364 63552 351416
rect 68100 351364 68152 351416
rect 72332 351364 72384 351416
rect 99380 351364 99432 351416
rect 130200 351364 130252 351416
rect 153292 351364 153344 351416
rect 193864 351364 193916 351416
rect 197452 351364 197504 351416
rect 270224 351364 270276 351416
rect 271880 351364 271932 351416
rect 39212 351296 39264 351348
rect 42156 351296 42208 351348
rect 42248 351296 42300 351348
rect 46572 351296 46624 351348
rect 52184 351296 52236 351348
rect 69204 351296 69256 351348
rect 72976 351296 73028 351348
rect 100852 351296 100904 351348
rect 131028 351296 131080 351348
rect 154764 351296 154816 351348
rect 40224 351228 40276 351280
rect 44364 351228 44416 351280
rect 53656 351228 53708 351280
rect 71228 351228 71280 351280
rect 75184 351228 75236 351280
rect 103704 351228 103756 351280
rect 125416 351228 125468 351280
rect 153384 351228 153436 351280
rect 226984 351228 227036 351280
rect 228732 351228 228784 351280
rect 38660 351160 38712 351212
rect 41512 351160 41564 351212
rect 41604 351160 41656 351212
rect 45652 351160 45704 351212
rect 55036 351160 55088 351212
rect 73436 351160 73488 351212
rect 74448 351160 74500 351212
rect 102508 351160 102560 351212
rect 123760 351160 123812 351212
rect 153476 351160 153528 351212
rect 228824 351160 228876 351212
rect 229836 351160 229888 351212
rect 38200 351092 38252 351144
rect 40132 351092 40184 351144
rect 64788 351092 64840 351144
rect 88524 351092 88576 351144
rect 66168 351024 66220 351076
rect 90732 351024 90784 351076
rect 183836 351024 183888 351076
rect 184572 351024 184624 351076
rect 67272 350956 67324 351008
rect 91836 350956 91888 351008
rect 110696 350956 110748 351008
rect 111708 350956 111760 351008
rect 173900 350956 173952 351008
rect 174820 350956 174872 351008
rect 230480 350956 230532 351008
rect 231860 350956 231912 351008
rect 62028 350888 62080 350940
rect 84384 350888 84436 350940
rect 135536 350888 135588 350940
rect 136456 350888 136508 350940
rect 201500 350888 201552 350940
rect 202880 350888 202932 350940
rect 233700 350888 233752 350940
rect 235172 350888 235224 350940
rect 272432 350888 272484 350940
rect 274640 350888 274692 350940
rect 63408 350820 63460 350872
rect 86316 350820 86368 350872
rect 120448 350820 120500 350872
rect 121368 350820 121420 350872
rect 158720 350820 158772 350872
rect 159732 350820 159784 350872
rect 34520 350752 34572 350804
rect 36820 350752 36872 350804
rect 37096 350752 37148 350804
rect 37924 350752 37976 350804
rect 60648 350752 60700 350804
rect 82084 350752 82136 350804
rect 134432 350752 134484 350804
rect 135168 350752 135220 350804
rect 139768 350752 139820 350804
rect 140688 350752 140740 350804
rect 223212 350752 223264 350804
rect 224316 350752 224368 350804
rect 59268 350684 59320 350736
rect 80060 350684 80112 350736
rect 57796 350616 57848 350668
rect 77852 350616 77904 350668
rect 144184 350616 144236 350668
rect 144828 350616 144880 350668
rect 164240 350616 164292 350668
rect 165068 350616 165120 350668
rect 56508 350548 56560 350600
rect 76012 350548 76064 350600
rect 282368 347803 282420 347812
rect 282368 347769 282377 347803
rect 282377 347769 282411 347803
rect 282411 347769 282420 347803
rect 282368 347760 282420 347769
rect 3148 336744 3200 336796
rect 6184 336744 6236 336796
rect 303620 327020 303672 327072
rect 577596 327020 577648 327072
rect 303620 325592 303672 325644
rect 563704 325592 563756 325644
rect 21364 322736 21416 322788
rect 22192 322736 22244 322788
rect 303620 321580 303672 321632
rect 580172 321580 580224 321632
rect 100760 321240 100812 321292
rect 106280 321240 106332 321292
rect 231768 321172 231820 321224
rect 235448 321172 235500 321224
rect 108304 321104 108356 321156
rect 115204 321104 115256 321156
rect 92112 321036 92164 321088
rect 96620 321036 96672 321088
rect 111524 321036 111576 321088
rect 117964 321036 118016 321088
rect 101772 320968 101824 321020
rect 106372 320968 106424 321020
rect 109316 320968 109368 321020
rect 119344 320968 119396 321020
rect 228272 320968 228324 321020
rect 232228 320968 232280 321020
rect 22100 320900 22152 320952
rect 24768 320832 24820 320884
rect 26332 320832 26384 320884
rect 75920 320900 75972 320952
rect 78680 320900 78732 320952
rect 102876 320900 102928 320952
rect 108948 320900 109000 320952
rect 42892 320832 42944 320884
rect 64052 320832 64104 320884
rect 64880 320832 64932 320884
rect 72700 320832 72752 320884
rect 74540 320832 74592 320884
rect 82452 320832 82504 320884
rect 85120 320832 85172 320884
rect 93216 320832 93268 320884
rect 98000 320832 98052 320884
rect 106096 320832 106148 320884
rect 121552 320832 121604 320884
rect 279516 320832 279568 320884
rect 73804 320764 73856 320816
rect 75920 320764 75972 320816
rect 83464 320764 83516 320816
rect 85764 320764 85816 320816
rect 91008 320764 91060 320816
rect 95240 320764 95292 320816
rect 195612 320764 195664 320816
rect 227076 320764 227128 320816
rect 231124 320764 231176 320816
rect 248236 320764 248288 320816
rect 250536 320764 250588 320816
rect 256608 320764 256660 320816
rect 258080 320764 258132 320816
rect 226248 320628 226300 320680
rect 230112 320628 230164 320680
rect 204260 320560 204312 320612
rect 206376 320560 206428 320612
rect 208400 320560 208452 320612
rect 210700 320560 210752 320612
rect 110420 320492 110472 320544
rect 113824 320492 113876 320544
rect 23388 320424 23440 320476
rect 25320 320424 25372 320476
rect 88892 320424 88944 320476
rect 91284 320424 91336 320476
rect 94228 320424 94280 320476
rect 99472 320424 99524 320476
rect 99656 320424 99708 320476
rect 104900 320424 104952 320476
rect 235448 320424 235500 320476
rect 238668 320424 238720 320476
rect 246120 320424 246172 320476
rect 248420 320424 248472 320476
rect 78128 320356 78180 320408
rect 81256 320356 81308 320408
rect 87788 320356 87840 320408
rect 90088 320356 90140 320408
rect 97540 320356 97592 320408
rect 102140 320356 102192 320408
rect 200120 320356 200172 320408
rect 203156 320356 203208 320408
rect 236644 320356 236696 320408
rect 239772 320356 239824 320408
rect 25320 320288 25372 320340
rect 27436 320288 27488 320340
rect 54392 320288 54444 320340
rect 55220 320288 55272 320340
rect 66260 320288 66312 320340
rect 67640 320288 67692 320340
rect 69480 320288 69532 320340
rect 71780 320288 71832 320340
rect 80244 320288 80296 320340
rect 82820 320288 82872 320340
rect 86684 320288 86736 320340
rect 91100 320288 91152 320340
rect 98552 320288 98604 320340
rect 103520 320288 103572 320340
rect 103980 320288 104032 320340
rect 109776 320288 109828 320340
rect 198740 320288 198792 320340
rect 200948 320288 201000 320340
rect 229468 320288 229520 320340
rect 233332 320288 233384 320340
rect 238668 320288 238720 320340
rect 241888 320288 241940 320340
rect 242624 320288 242676 320340
rect 245200 320288 245252 320340
rect 253388 320288 253440 320340
rect 254860 320288 254912 320340
rect 27712 320220 27764 320272
rect 29644 320220 29696 320272
rect 30288 320220 30340 320272
rect 31760 320220 31812 320272
rect 33692 320220 33744 320272
rect 34980 320220 35032 320272
rect 61936 320220 61988 320272
rect 63500 320220 63552 320272
rect 68376 320220 68428 320272
rect 70400 320220 70452 320272
rect 70584 320220 70636 320272
rect 73160 320220 73212 320272
rect 77024 320220 77076 320272
rect 79968 320220 80020 320272
rect 81348 320220 81400 320272
rect 83096 320220 83148 320272
rect 85672 320220 85724 320272
rect 89628 320220 89680 320272
rect 96436 320220 96488 320272
rect 100760 320220 100812 320272
rect 105084 320220 105136 320272
rect 110420 320220 110472 320272
rect 163228 320220 163280 320272
rect 167644 320220 167696 320272
rect 197544 320220 197596 320272
rect 199936 320220 199988 320272
rect 201500 320220 201552 320272
rect 204168 320220 204220 320272
rect 233148 320220 233200 320272
rect 236552 320220 236604 320272
rect 237840 320220 237892 320272
rect 240876 320220 240928 320272
rect 241428 320220 241480 320272
rect 244096 320220 244148 320272
rect 245016 320220 245068 320272
rect 247316 320220 247368 320272
rect 247408 320220 247460 320272
rect 249432 320220 249484 320272
rect 251088 320220 251140 320272
rect 252744 320220 252796 320272
rect 254584 320220 254636 320272
rect 255964 320220 256016 320272
rect 257988 320220 258040 320272
rect 259184 320220 259236 320272
rect 22008 320152 22060 320204
rect 24216 320152 24268 320204
rect 26516 320152 26568 320204
rect 28540 320152 28592 320204
rect 28908 320152 28960 320204
rect 30656 320152 30708 320204
rect 31668 320152 31720 320204
rect 32864 320152 32916 320204
rect 33048 320152 33100 320204
rect 33876 320152 33928 320204
rect 35900 320152 35952 320204
rect 37188 320152 37240 320204
rect 37280 320152 37332 320204
rect 38200 320152 38252 320204
rect 38568 320152 38620 320204
rect 39304 320152 39356 320204
rect 42524 320152 42576 320204
rect 42800 320152 42852 320204
rect 43628 320152 43680 320204
rect 46940 320152 46992 320204
rect 47952 320152 48004 320204
rect 59820 320152 59872 320204
rect 60740 320152 60792 320204
rect 60832 320152 60884 320204
rect 62120 320152 62172 320204
rect 63040 320152 63092 320204
rect 64328 320152 64380 320204
rect 65156 320152 65208 320204
rect 66260 320152 66312 320204
rect 67364 320152 67416 320204
rect 69020 320152 69072 320204
rect 71596 320152 71648 320204
rect 73252 320152 73304 320204
rect 74908 320152 74960 320204
rect 77300 320152 77352 320204
rect 79140 320152 79192 320204
rect 81624 320152 81676 320204
rect 84568 320152 84620 320204
rect 88064 320152 88116 320204
rect 89996 320152 90048 320204
rect 92664 320152 92716 320204
rect 95332 320152 95384 320204
rect 99104 320152 99156 320204
rect 107200 320152 107252 320204
rect 112444 320152 112496 320204
rect 113640 320152 113692 320204
rect 114468 320152 114520 320204
rect 114744 320152 114796 320204
rect 115848 320152 115900 320204
rect 119068 320152 119120 320204
rect 119988 320152 120040 320204
rect 120172 320152 120224 320204
rect 121368 320152 121420 320204
rect 124404 320152 124456 320204
rect 125416 320152 125468 320204
rect 128728 320152 128780 320204
rect 129648 320152 129700 320204
rect 129832 320152 129884 320204
rect 130936 320152 130988 320204
rect 133052 320152 133104 320204
rect 133788 320152 133840 320204
rect 134156 320152 134208 320204
rect 135168 320152 135220 320204
rect 135260 320152 135312 320204
rect 136548 320152 136600 320204
rect 138480 320152 138532 320204
rect 139308 320152 139360 320204
rect 139492 320152 139544 320204
rect 140688 320152 140740 320204
rect 143816 320152 143868 320204
rect 144828 320152 144880 320204
rect 144920 320152 144972 320204
rect 146116 320152 146168 320204
rect 148140 320152 148192 320204
rect 148968 320152 149020 320204
rect 149244 320152 149296 320204
rect 150256 320152 150308 320204
rect 153568 320152 153620 320204
rect 154488 320152 154540 320204
rect 154672 320152 154724 320204
rect 155776 320152 155828 320204
rect 157892 320152 157944 320204
rect 158628 320152 158680 320204
rect 158904 320152 158956 320204
rect 159916 320152 159968 320204
rect 164332 320152 164384 320204
rect 165436 320152 165488 320204
rect 168656 320152 168708 320204
rect 169668 320152 169720 320204
rect 169760 320152 169812 320204
rect 170956 320152 171008 320204
rect 172980 320152 173032 320204
rect 173808 320152 173860 320204
rect 173992 320152 174044 320204
rect 175096 320152 175148 320204
rect 178316 320152 178368 320204
rect 179328 320152 179380 320204
rect 179420 320152 179472 320204
rect 180708 320152 180760 320204
rect 182640 320152 182692 320204
rect 183468 320152 183520 320204
rect 183744 320152 183796 320204
rect 184756 320152 184808 320204
rect 191840 320152 191892 320204
rect 196624 320152 196676 320204
rect 197268 320152 197320 320204
rect 198832 320152 198884 320204
rect 199016 320152 199068 320204
rect 202052 320152 202104 320204
rect 202880 320152 202932 320204
rect 205272 320152 205324 320204
rect 207112 320152 207164 320204
rect 209596 320152 209648 320204
rect 219900 320152 219952 320204
rect 224684 320152 224736 320204
rect 224868 320152 224920 320204
rect 229008 320152 229060 320204
rect 230296 320152 230348 320204
rect 234344 320152 234396 320204
rect 234528 320152 234580 320204
rect 237656 320152 237708 320204
rect 240048 320152 240100 320204
rect 242992 320152 243044 320204
rect 243820 320152 243872 320204
rect 246212 320152 246264 320204
rect 249708 320152 249760 320204
rect 251640 320152 251692 320204
rect 252468 320152 252520 320204
rect 253756 320152 253808 320204
rect 255780 320152 255832 320204
rect 256976 320152 257028 320204
rect 259368 320152 259420 320204
rect 260288 320152 260340 320204
rect 41420 320084 41472 320136
rect 263508 320152 263560 320204
rect 263600 320152 263652 320204
rect 264520 320152 264572 320204
rect 267740 320152 267792 320204
rect 268844 320152 268896 320204
rect 269120 320152 269172 320204
rect 269948 320152 270000 320204
rect 276020 320152 276072 320204
rect 276664 320152 276716 320204
rect 277400 320152 277452 320204
rect 277860 320152 277912 320204
rect 278688 320152 278740 320204
rect 279056 320152 279108 320204
rect 262220 320016 262272 320068
rect 22192 319404 22244 319456
rect 36544 319404 36596 319456
rect 20628 318724 20680 318776
rect 23112 318724 23164 318776
rect 91284 318724 91336 318776
rect 93492 318724 93544 318776
rect 99104 318724 99156 318776
rect 100668 318724 100720 318776
rect 191196 318724 191248 318776
rect 197268 318724 197320 318776
rect 200764 318724 200816 318776
rect 206928 318724 206980 318776
rect 211528 318724 211580 318776
rect 217140 318724 217192 318776
rect 223488 318724 223540 318776
rect 227904 318724 227956 318776
rect 201960 318656 202012 318708
rect 208308 318656 208360 318708
rect 220636 318656 220688 318708
rect 225788 318656 225840 318708
rect 106372 318520 106424 318572
rect 107844 318520 107896 318572
rect 192392 318520 192444 318572
rect 197544 318520 197596 318572
rect 193588 318452 193640 318504
rect 198740 318452 198792 318504
rect 34888 318384 34940 318436
rect 35808 318384 35860 318436
rect 85120 318384 85172 318436
rect 86316 318384 86368 318436
rect 88064 318384 88116 318436
rect 88708 318384 88760 318436
rect 194508 318384 194560 318436
rect 199016 318384 199068 318436
rect 209136 318384 209188 318436
rect 215024 318384 215076 318436
rect 85764 318316 85816 318368
rect 87512 318316 87564 318368
rect 195796 318248 195848 318300
rect 200120 318248 200172 318300
rect 204168 318248 204220 318300
rect 208400 318248 208452 318300
rect 217508 318248 217560 318300
rect 222568 318248 222620 318300
rect 198372 318180 198424 318232
rect 202880 318180 202932 318232
rect 218704 318180 218756 318232
rect 223580 318180 223632 318232
rect 202788 318112 202840 318164
rect 207112 318112 207164 318164
rect 207940 318112 207992 318164
rect 213828 318112 213880 318164
rect 42892 318044 42944 318096
rect 113364 318044 113416 318096
rect 190000 318044 190052 318096
rect 197176 318044 197228 318096
rect 90088 317976 90140 318028
rect 92296 317976 92348 318028
rect 197176 317908 197228 317960
rect 201500 317908 201552 317960
rect 213828 317908 213880 317960
rect 219256 317908 219308 317960
rect 222016 317908 222068 317960
rect 226800 317908 226852 317960
rect 199568 317704 199620 317756
rect 204260 317704 204312 317756
rect 210332 317704 210384 317756
rect 216036 317704 216088 317756
rect 206744 317568 206796 317620
rect 212448 317568 212500 317620
rect 216312 317568 216364 317620
rect 221464 317568 221516 317620
rect 83096 317500 83148 317552
rect 85120 317500 85172 317552
rect 188896 317500 188948 317552
rect 191840 317500 191892 317552
rect 205364 317500 205416 317552
rect 211068 317500 211120 317552
rect 217968 317500 218020 317552
rect 92664 317432 92716 317484
rect 94688 317432 94740 317484
rect 212448 317432 212500 317484
rect 215116 317432 215168 317484
rect 220360 317432 220412 317484
rect 2780 316684 2832 316736
rect 3516 316684 3568 316736
rect 288900 316684 288952 316736
rect 36544 315324 36596 315376
rect 111800 315324 111852 315376
rect 14556 315256 14608 315308
rect 185584 315256 185636 315308
rect 111800 313216 111852 313268
rect 114376 313216 114428 313268
rect 303620 311856 303672 311908
rect 336004 311856 336056 311908
rect 114376 310768 114428 310820
rect 116584 310768 116636 310820
rect 303620 310496 303672 310548
rect 341524 310496 341576 310548
rect 303620 309136 303672 309188
rect 340144 309136 340196 309188
rect 282092 309111 282144 309120
rect 282092 309077 282101 309111
rect 282101 309077 282135 309111
rect 282135 309077 282144 309111
rect 282092 309068 282144 309077
rect 113180 306348 113232 306400
rect 113364 306348 113416 306400
rect 303620 306348 303672 306400
rect 560944 306348 560996 306400
rect 300860 305600 300912 305652
rect 296168 303560 296220 303612
rect 580356 303560 580408 303612
rect 282552 299480 282604 299532
rect 282368 292544 282420 292596
rect 282552 292544 282604 292596
rect 282276 278740 282328 278792
rect 282368 278740 282420 278792
rect 11704 275952 11756 276004
rect 17132 275952 17184 276004
rect 304356 275952 304408 276004
rect 580172 275952 580224 276004
rect 282184 263576 282236 263628
rect 282368 263576 282420 263628
rect 146024 254124 146076 254176
rect 149520 254124 149572 254176
rect 214564 233860 214616 233912
rect 315304 233860 315356 233912
rect 67180 230392 67232 230444
rect 72424 230392 72476 230444
rect 214748 229712 214800 229764
rect 305644 229712 305696 229764
rect 245568 229100 245620 229152
rect 250444 229100 250496 229152
rect 304264 229032 304316 229084
rect 579988 229032 580040 229084
rect 214932 228352 214984 228404
rect 301504 228352 301556 228404
rect 72424 227060 72476 227112
rect 79324 227060 79376 227112
rect 13084 226992 13136 227044
rect 411904 226992 411956 227044
rect 214656 225632 214708 225684
rect 312544 225632 312596 225684
rect 9128 225564 9180 225616
rect 299480 225564 299532 225616
rect 125508 224952 125560 225004
rect 214472 224995 214524 225004
rect 114468 224884 114520 224936
rect 214472 224961 214481 224995
rect 214481 224961 214515 224995
rect 214515 224961 214524 224995
rect 214472 224952 214524 224961
rect 119344 224816 119396 224868
rect 125416 224816 125468 224868
rect 130936 224884 130988 224936
rect 145748 224884 145800 224936
rect 155776 224884 155828 224936
rect 170312 224884 170364 224936
rect 179328 224884 179380 224936
rect 193864 224884 193916 224936
rect 128268 224816 128320 224868
rect 143540 224816 143592 224868
rect 150256 224816 150308 224868
rect 164976 224816 165028 224868
rect 167644 224816 167696 224868
rect 178868 224816 178920 224868
rect 180708 224816 180760 224868
rect 194876 224816 194928 224868
rect 115204 224748 115256 224800
rect 124312 224748 124364 224800
rect 132868 224748 132920 224800
rect 146116 224748 146168 224800
rect 160652 224748 160704 224800
rect 161388 224748 161440 224800
rect 176752 224748 176804 224800
rect 183468 224748 183520 224800
rect 198096 224748 198148 224800
rect 122748 224680 122800 224732
rect 138204 224680 138256 224732
rect 151728 224680 151780 224732
rect 167092 224680 167144 224732
rect 170956 224680 171008 224732
rect 185308 224680 185360 224732
rect 187608 224680 187660 224732
rect 202420 224680 202472 224732
rect 115848 224612 115900 224664
rect 113088 224544 113140 224596
rect 130752 224612 130804 224664
rect 131028 224612 131080 224664
rect 146760 224612 146812 224664
rect 147588 224612 147640 224664
rect 162860 224612 162912 224664
rect 165436 224612 165488 224664
rect 179972 224612 180024 224664
rect 186228 224612 186280 224664
rect 201316 224612 201368 224664
rect 117228 224476 117280 224528
rect 113824 224408 113876 224460
rect 126428 224408 126480 224460
rect 129372 224544 129424 224596
rect 132408 224544 132460 224596
rect 147864 224544 147916 224596
rect 150348 224544 150400 224596
rect 166080 224544 166132 224596
rect 175096 224544 175148 224596
rect 189540 224544 189592 224596
rect 133972 224476 134024 224528
rect 137928 224476 137980 224528
rect 153200 224476 153252 224528
rect 155868 224476 155920 224528
rect 171416 224476 171468 224528
rect 184756 224476 184808 224528
rect 199200 224476 199252 224528
rect 128636 224408 128688 224460
rect 112444 224340 112496 224392
rect 123208 224340 123260 224392
rect 126888 224340 126940 224392
rect 142528 224408 142580 224460
rect 146208 224408 146260 224460
rect 161756 224408 161808 224460
rect 175188 224408 175240 224460
rect 190644 224408 190696 224460
rect 141424 224340 141476 224392
rect 142068 224340 142120 224392
rect 157432 224340 157484 224392
rect 171048 224340 171100 224392
rect 186320 224340 186372 224392
rect 188436 224340 188488 224392
rect 203432 224340 203484 224392
rect 79324 224272 79376 224324
rect 100300 224272 100352 224324
rect 115756 224272 115808 224324
rect 131764 224272 131816 224324
rect 136456 224272 136508 224324
rect 152096 224272 152148 224324
rect 165528 224272 165580 224324
rect 180984 224272 181036 224324
rect 184848 224272 184900 224324
rect 200304 224272 200356 224324
rect 3608 224204 3660 224256
rect 120080 224204 120132 224256
rect 121276 224204 121328 224256
rect 137192 224204 137244 224256
rect 140596 224204 140648 224256
rect 156420 224204 156472 224256
rect 160008 224204 160060 224256
rect 175648 224204 175700 224256
rect 180616 224204 180668 224256
rect 195980 224204 196032 224256
rect 210976 224204 211028 224256
rect 286324 224204 286376 224256
rect 118608 224136 118660 224188
rect 125232 224068 125284 224120
rect 140320 224136 140372 224188
rect 144828 224136 144880 224188
rect 159640 224136 159692 224188
rect 159916 224136 159968 224188
rect 174636 224136 174688 224188
rect 177948 224136 178000 224188
rect 192760 224136 192812 224188
rect 139308 224068 139360 224120
rect 140688 224068 140740 224120
rect 155316 224068 155368 224120
rect 166908 224068 166960 224120
rect 182088 224068 182140 224120
rect 182180 224068 182232 224120
rect 197084 224068 197136 224120
rect 119988 224000 120040 224052
rect 134984 224000 135036 224052
rect 136548 224000 136600 224052
rect 151084 224000 151136 224052
rect 153108 224000 153160 224052
rect 168196 224000 168248 224052
rect 169668 224000 169720 224052
rect 184204 224000 184256 224052
rect 121368 223932 121420 223984
rect 136088 223932 136140 223984
rect 143448 223932 143500 223984
rect 158536 223932 158588 223984
rect 158628 223932 158680 223984
rect 173532 223932 173584 223984
rect 173808 223932 173860 223984
rect 188528 223932 188580 223984
rect 117964 223864 118016 223916
rect 127532 223864 127584 223916
rect 139400 223864 139452 223916
rect 154304 223864 154356 223916
rect 162768 223864 162820 223916
rect 177764 223864 177816 223916
rect 124128 223796 124180 223848
rect 135168 223796 135220 223848
rect 149980 223796 150032 223848
rect 154488 223796 154540 223848
rect 169208 223796 169260 223848
rect 176568 223796 176620 223848
rect 191748 223796 191800 223848
rect 133788 223728 133840 223780
rect 148876 223728 148928 223780
rect 148968 223728 149020 223780
rect 163872 223728 163924 223780
rect 168288 223728 168340 223780
rect 183192 223728 183244 223780
rect 129648 223660 129700 223712
rect 144644 223660 144696 223712
rect 157248 223660 157300 223712
rect 172428 223660 172480 223712
rect 172520 223660 172572 223712
rect 187424 223660 187476 223712
rect 3516 223592 3568 223644
rect 121092 223592 121144 223644
rect 229744 223592 229796 223644
rect 283380 223592 283432 223644
rect 231124 222912 231176 222964
rect 245568 222912 245620 222964
rect 229008 222844 229060 222896
rect 313924 222844 313976 222896
rect 214472 222207 214524 222216
rect 214472 222173 214481 222207
rect 214481 222173 214515 222207
rect 214515 222173 214524 222207
rect 214472 222164 214524 222173
rect 214472 222071 214524 222080
rect 214472 222037 214481 222071
rect 214481 222037 214515 222071
rect 214515 222037 214524 222071
rect 214472 222028 214524 222037
rect 55220 220804 55272 220856
rect 116400 220804 116452 220856
rect 213920 220804 213972 220856
rect 226340 220804 226392 220856
rect 214012 220124 214064 220176
rect 226340 220124 226392 220176
rect 14464 220056 14516 220108
rect 116676 220056 116728 220108
rect 213920 220056 213972 220108
rect 226432 220056 226484 220108
rect 104808 219376 104860 219428
rect 116124 219444 116176 219496
rect 213920 218764 213972 218816
rect 226340 218764 226392 218816
rect 214012 218696 214064 218748
rect 226432 218696 226484 218748
rect 104808 217948 104860 218000
rect 116400 218016 116452 218068
rect 213920 217268 213972 217320
rect 226340 217268 226392 217320
rect 104808 216588 104860 216640
rect 116400 216588 116452 216640
rect 213920 216588 213972 216640
rect 226432 216588 226484 216640
rect 104808 215908 104860 215960
rect 115940 215908 115992 215960
rect 213920 215908 213972 215960
rect 226340 215908 226392 215960
rect 104808 215228 104860 215280
rect 116400 215296 116452 215348
rect 213920 215228 213972 215280
rect 226432 215228 226484 215280
rect 214012 215160 214064 215212
rect 226340 215160 226392 215212
rect 104808 213868 104860 213920
rect 116400 213936 116452 213988
rect 213920 213868 213972 213920
rect 226432 213868 226484 213920
rect 214012 213800 214064 213852
rect 226340 213800 226392 213852
rect 104440 212440 104492 212492
rect 115940 212508 115992 212560
rect 214564 212508 214616 212560
rect 213920 212440 213972 212492
rect 226432 212440 226484 212492
rect 214012 212372 214064 212424
rect 226340 212372 226392 212424
rect 104808 211080 104860 211132
rect 116308 211148 116360 211200
rect 213920 211080 213972 211132
rect 226524 211080 226576 211132
rect 104808 209720 104860 209772
rect 116308 209788 116360 209840
rect 214012 209720 214064 209772
rect 226248 209720 226300 209772
rect 213920 209652 213972 209704
rect 226064 209652 226116 209704
rect 104808 208292 104860 208344
rect 116032 208360 116084 208412
rect 214012 208292 214064 208344
rect 226156 208292 226208 208344
rect 213920 208224 213972 208276
rect 225972 208224 226024 208276
rect 113824 207068 113876 207120
rect 116400 207068 116452 207120
rect 104716 206932 104768 206984
rect 116308 207000 116360 207052
rect 213920 206932 213972 206984
rect 226064 206932 226116 206984
rect 104808 206864 104860 206916
rect 113824 206864 113876 206916
rect 214012 206864 214064 206916
rect 226248 206864 226300 206916
rect 104808 205572 104860 205624
rect 115940 205640 115992 205692
rect 214472 205683 214524 205692
rect 214472 205649 214481 205683
rect 214481 205649 214515 205683
rect 214515 205649 214524 205683
rect 214472 205640 214524 205649
rect 213920 205572 213972 205624
rect 226156 205572 226208 205624
rect 104808 204212 104860 204264
rect 116400 204280 116452 204332
rect 214012 204212 214064 204264
rect 225972 204212 226024 204264
rect 213920 204144 213972 204196
rect 225788 204144 225840 204196
rect 104808 202784 104860 202836
rect 116308 202852 116360 202904
rect 214472 202895 214524 202904
rect 214472 202861 214481 202895
rect 214481 202861 214515 202895
rect 214515 202861 214524 202895
rect 214472 202852 214524 202861
rect 213920 202784 213972 202836
rect 225880 202784 225932 202836
rect 214012 202716 214064 202768
rect 226156 202716 226208 202768
rect 104808 201424 104860 201476
rect 116124 201492 116176 201544
rect 213920 201424 213972 201476
rect 225604 201424 225656 201476
rect 214012 201356 214064 201408
rect 225696 201356 225748 201408
rect 214472 200540 214524 200592
rect 214840 200540 214892 200592
rect 104808 200064 104860 200116
rect 116124 200200 116176 200252
rect 113272 200132 113324 200184
rect 115940 200132 115992 200184
rect 213920 200064 213972 200116
rect 226248 200064 226300 200116
rect 224132 198772 224184 198824
rect 226432 198772 226484 198824
rect 114468 198704 114520 198756
rect 115940 198704 115992 198756
rect 223948 198704 224000 198756
rect 226340 198704 226392 198756
rect 104808 198636 104860 198688
rect 113272 198636 113324 198688
rect 214012 198636 214064 198688
rect 225972 198636 226024 198688
rect 213920 198568 213972 198620
rect 226064 198568 226116 198620
rect 224500 197412 224552 197464
rect 226432 197412 226484 197464
rect 104716 197276 104768 197328
rect 116124 197344 116176 197396
rect 224040 197344 224092 197396
rect 226340 197344 226392 197396
rect 214012 197276 214064 197328
rect 226156 197276 226208 197328
rect 104808 197208 104860 197260
rect 114468 197208 114520 197260
rect 213920 197208 213972 197260
rect 225788 197208 225840 197260
rect 224316 196052 224368 196104
rect 226340 196052 226392 196104
rect 104808 195916 104860 195968
rect 116400 195984 116452 196036
rect 224408 195984 224460 196036
rect 226708 195984 226760 196036
rect 213920 195916 213972 195968
rect 226248 195916 226300 195968
rect 214012 195848 214064 195900
rect 225880 195848 225932 195900
rect 224224 194692 224276 194744
rect 226524 194692 226576 194744
rect 221464 194624 221516 194676
rect 226432 194624 226484 194676
rect 104808 194488 104860 194540
rect 115940 194556 115992 194608
rect 214196 194556 214248 194608
rect 226340 194556 226392 194608
rect 213920 194488 213972 194540
rect 225696 194488 225748 194540
rect 220084 193264 220136 193316
rect 226432 193264 226484 193316
rect 104440 193128 104492 193180
rect 116124 193196 116176 193248
rect 214472 193196 214524 193248
rect 226340 193196 226392 193248
rect 213920 193128 213972 193180
rect 224132 193128 224184 193180
rect 214012 193060 214064 193112
rect 223948 193060 224000 193112
rect 113916 191972 113968 192024
rect 116400 191972 116452 192024
rect 113180 191904 113232 191956
rect 116032 191904 116084 191956
rect 215300 191904 215352 191956
rect 226340 191904 226392 191956
rect 214104 191836 214156 191888
rect 226432 191836 226484 191888
rect 104440 191768 104492 191820
rect 113916 191768 113968 191820
rect 214012 191768 214064 191820
rect 224040 191768 224092 191820
rect 213920 191700 213972 191752
rect 224500 191700 224552 191752
rect 113272 190612 113324 190664
rect 116492 190612 116544 190664
rect 214288 190544 214340 190596
rect 226340 190544 226392 190596
rect 215024 190476 215076 190528
rect 226432 190476 226484 190528
rect 104716 190408 104768 190460
rect 113180 190408 113232 190460
rect 214012 190408 214064 190460
rect 224408 190408 224460 190460
rect 213920 190340 213972 190392
rect 224316 190340 224368 190392
rect 218704 189116 218756 189168
rect 226432 189116 226484 189168
rect 114468 189048 114520 189100
rect 116400 189048 116452 189100
rect 214380 189048 214432 189100
rect 226340 189048 226392 189100
rect 104808 188980 104860 189032
rect 113272 188980 113324 189032
rect 213920 188980 213972 189032
rect 224224 188980 224276 189032
rect 222936 187756 222988 187808
rect 226432 187756 226484 187808
rect 114100 187688 114152 187740
rect 116400 187688 116452 187740
rect 215944 187688 215996 187740
rect 226340 187688 226392 187740
rect 104808 187620 104860 187672
rect 114468 187620 114520 187672
rect 213920 186532 213972 186584
rect 221464 186532 221516 186584
rect 224408 186396 224460 186448
rect 226432 186396 226484 186448
rect 104716 186260 104768 186312
rect 115940 186328 115992 186380
rect 214196 186328 214248 186380
rect 226340 186328 226392 186380
rect 104808 186192 104860 186244
rect 114100 186192 114152 186244
rect 213920 185036 213972 185088
rect 220084 185036 220136 185088
rect 114468 184968 114520 185020
rect 116400 184968 116452 185020
rect 220176 184968 220228 185020
rect 226432 184968 226484 185020
rect 104808 184832 104860 184884
rect 116032 184900 116084 184952
rect 214012 184900 214064 184952
rect 226340 184900 226392 184952
rect 215300 184152 215352 184204
rect 226524 184152 226576 184204
rect 114376 183540 114428 183592
rect 116400 183540 116452 183592
rect 213920 183540 213972 183592
rect 226340 183540 226392 183592
rect 104808 183472 104860 183524
rect 114468 183472 114520 183524
rect 214472 182316 214524 182368
rect 226432 182316 226484 182368
rect 215024 182248 215076 182300
rect 226340 182248 226392 182300
rect 113180 182180 113232 182232
rect 115940 182180 115992 182232
rect 104808 182112 104860 182164
rect 114376 182112 114428 182164
rect 336004 182112 336056 182164
rect 579988 182112 580040 182164
rect 221464 181228 221516 181280
rect 226340 181228 226392 181280
rect 113272 181092 113324 181144
rect 115940 181092 115992 181144
rect 215116 180820 215168 180872
rect 226340 180820 226392 180872
rect 227720 180820 227772 180872
rect 230848 180820 230900 180872
rect 104808 180752 104860 180804
rect 113180 180752 113232 180804
rect 213920 180548 213972 180600
rect 218704 180548 218756 180600
rect 214840 179528 214892 179580
rect 222844 179460 222896 179512
rect 226432 179460 226484 179512
rect 113916 179392 113968 179444
rect 116400 179392 116452 179444
rect 214840 179392 214892 179444
rect 226340 179392 226392 179444
rect 104808 179324 104860 179376
rect 113272 179324 113324 179376
rect 214012 179324 214064 179376
rect 222936 179324 222988 179376
rect 213920 179052 213972 179104
rect 215944 179052 215996 179104
rect 221556 178100 221608 178152
rect 226432 178100 226484 178152
rect 114192 178032 114244 178084
rect 115940 178032 115992 178084
rect 224316 178032 224368 178084
rect 226340 178032 226392 178084
rect 104164 177964 104216 178016
rect 113916 177964 113968 178016
rect 213920 177964 213972 178016
rect 227076 177964 227128 178016
rect 114100 176740 114152 176792
rect 115940 176740 115992 176792
rect 114468 176672 114520 176724
rect 116400 176672 116452 176724
rect 218704 176672 218756 176724
rect 226340 176672 226392 176724
rect 104164 176604 104216 176656
rect 114192 176604 114244 176656
rect 214012 176604 214064 176656
rect 224408 176604 224460 176656
rect 114284 175244 114336 175296
rect 116400 175244 116452 175296
rect 224224 175244 224276 175296
rect 226892 175244 226944 175296
rect 104808 175176 104860 175228
rect 114100 175176 114152 175228
rect 104532 175108 104584 175160
rect 114468 175108 114520 175160
rect 213920 174156 213972 174208
rect 220176 174156 220228 174208
rect 223580 174088 223632 174140
rect 227720 174088 227772 174140
rect 220084 174020 220136 174072
rect 226432 174020 226484 174072
rect 114376 173884 114428 173936
rect 115940 173884 115992 173936
rect 214472 173927 214524 173936
rect 214472 173893 214481 173927
rect 214481 173893 214515 173927
rect 214515 173893 214524 173927
rect 214472 173884 214524 173893
rect 104808 173816 104860 173868
rect 114284 173816 114336 173868
rect 213920 173816 213972 173868
rect 226984 173816 227036 173868
rect 113180 172524 113232 172576
rect 116400 172524 116452 172576
rect 104440 172456 104492 172508
rect 114376 172456 114428 172508
rect 213920 172456 213972 172508
rect 225696 172456 225748 172508
rect 218796 171776 218848 171828
rect 223580 171776 223632 171828
rect 113272 171572 113324 171624
rect 116124 171572 116176 171624
rect 104808 171028 104860 171080
rect 113180 171028 113232 171080
rect 218060 170348 218112 170400
rect 227444 170348 227496 170400
rect 113916 169804 113968 169856
rect 116308 169804 116360 169856
rect 104256 169736 104308 169788
rect 116400 169736 116452 169788
rect 104808 169668 104860 169720
rect 113272 169668 113324 169720
rect 213920 169056 213972 169108
rect 221464 169056 221516 169108
rect 104808 168376 104860 168428
rect 116400 168376 116452 168428
rect 104164 168308 104216 168360
rect 113916 168308 113968 168360
rect 213920 168308 213972 168360
rect 222844 168308 222896 168360
rect 114468 167016 114520 167068
rect 115940 167016 115992 167068
rect 213920 166948 213972 167000
rect 224316 166948 224368 167000
rect 232228 166948 232280 167000
rect 232596 166948 232648 167000
rect 214196 166880 214248 166932
rect 214472 166880 214524 166932
rect 214012 166540 214064 166592
rect 221556 166540 221608 166592
rect 113824 165588 113876 165640
rect 115940 165588 115992 165640
rect 104624 165520 104676 165572
rect 114468 165520 114520 165572
rect 213920 165520 213972 165572
rect 225604 165520 225656 165572
rect 114468 164228 114520 164280
rect 116124 164228 116176 164280
rect 104808 164160 104860 164212
rect 113824 164160 113876 164212
rect 232320 164160 232372 164212
rect 232596 164160 232648 164212
rect 213920 164092 213972 164144
rect 218704 164092 218756 164144
rect 213920 163548 213972 163600
rect 220084 163548 220136 163600
rect 113180 162868 113232 162920
rect 116400 162868 116452 162920
rect 104808 162800 104860 162852
rect 114468 162800 114520 162852
rect 213920 162800 213972 162852
rect 224224 162800 224276 162852
rect 213920 162256 213972 162308
rect 218060 162256 218112 162308
rect 113272 161984 113324 162036
rect 116216 161984 116268 162036
rect 103704 161440 103756 161492
rect 116400 161440 116452 161492
rect 104808 161372 104860 161424
rect 113180 161372 113232 161424
rect 213920 161372 213972 161424
rect 229744 161372 229796 161424
rect 213920 160828 213972 160880
rect 218796 160828 218848 160880
rect 104256 160080 104308 160132
rect 116400 160080 116452 160132
rect 104808 160012 104860 160064
rect 113272 160012 113324 160064
rect 104808 158720 104860 158772
rect 116400 158720 116452 158772
rect 104348 157360 104400 157412
rect 116400 157360 116452 157412
rect 114284 155932 114336 155984
rect 116032 155932 116084 155984
rect 213920 155932 213972 155984
rect 224684 155932 224736 155984
rect 113456 154640 113508 154692
rect 116032 154640 116084 154692
rect 104256 154572 104308 154624
rect 116400 154572 116452 154624
rect 213920 154572 213972 154624
rect 224776 154572 224828 154624
rect 104624 154504 104676 154556
rect 114284 154504 114336 154556
rect 213920 153280 213972 153332
rect 224592 153280 224644 153332
rect 103796 153212 103848 153264
rect 115940 153212 115992 153264
rect 214012 153212 214064 153264
rect 224868 153212 224920 153264
rect 104808 153144 104860 153196
rect 113456 153144 113508 153196
rect 213920 151852 213972 151904
rect 224500 151852 224552 151904
rect 103704 151784 103756 151836
rect 116400 151784 116452 151836
rect 215944 151784 215996 151836
rect 286140 151784 286192 151836
rect 213920 150832 213972 150884
rect 216680 150832 216732 150884
rect 104348 150424 104400 150476
rect 116400 150424 116452 150476
rect 213920 150424 213972 150476
rect 224224 150424 224276 150476
rect 224684 150356 224736 150408
rect 227444 150356 227496 150408
rect 232136 149676 232188 149728
rect 232504 149676 232556 149728
rect 213920 149336 213972 149388
rect 216772 149336 216824 149388
rect 104808 149064 104860 149116
rect 116400 149064 116452 149116
rect 213920 149064 213972 149116
rect 224132 149064 224184 149116
rect 214104 148996 214156 149048
rect 227444 148996 227496 149048
rect 224776 148928 224828 148980
rect 227536 148928 227588 148980
rect 214564 148316 214616 148368
rect 214748 148316 214800 148368
rect 213920 147976 213972 148028
rect 216864 147976 216916 148028
rect 104716 147636 104768 147688
rect 116400 147636 116452 147688
rect 214932 147568 214984 147620
rect 227444 147568 227496 147620
rect 224868 147500 224920 147552
rect 226984 147500 227036 147552
rect 224592 147432 224644 147484
rect 227536 147432 227588 147484
rect 113640 146344 113692 146396
rect 115940 146344 115992 146396
rect 213920 146344 213972 146396
rect 217600 146344 217652 146396
rect 104532 146276 104584 146328
rect 116400 146276 116452 146328
rect 214012 146276 214064 146328
rect 227628 146276 227680 146328
rect 216680 146208 216732 146260
rect 226708 146208 226760 146260
rect 224500 146140 224552 146192
rect 227444 146140 227496 146192
rect 213920 144984 213972 145036
rect 217324 144984 217376 145036
rect 104164 144916 104216 144968
rect 116032 144916 116084 144968
rect 214012 144916 214064 144968
rect 227260 144916 227312 144968
rect 104624 144848 104676 144900
rect 113640 144848 113692 144900
rect 216772 144848 216824 144900
rect 226524 144848 226576 144900
rect 224224 144780 224276 144832
rect 227444 144780 227496 144832
rect 213920 143624 213972 143676
rect 216772 143624 216824 143676
rect 103520 143556 103572 143608
rect 116400 143556 116452 143608
rect 214012 143556 214064 143608
rect 227536 143556 227588 143608
rect 216864 143488 216916 143540
rect 226892 143488 226944 143540
rect 214380 143420 214432 143472
rect 214564 143420 214616 143472
rect 224132 143420 224184 143472
rect 227444 143420 227496 143472
rect 213920 142196 213972 142248
rect 216680 142196 216732 142248
rect 103704 142128 103756 142180
rect 116400 142128 116452 142180
rect 214012 142128 214064 142180
rect 227352 142128 227404 142180
rect 217600 142060 217652 142112
rect 226708 142060 226760 142112
rect 104348 140768 104400 140820
rect 116400 140768 116452 140820
rect 213920 140768 213972 140820
rect 226708 140768 226760 140820
rect 217324 140700 217376 140752
rect 227076 140700 227128 140752
rect 113548 139476 113600 139528
rect 116308 139476 116360 139528
rect 213920 139476 213972 139528
rect 226616 139476 226668 139528
rect 104808 139408 104860 139460
rect 116400 139408 116452 139460
rect 214012 139408 214064 139460
rect 226524 139408 226576 139460
rect 216772 139340 216824 139392
rect 227444 139340 227496 139392
rect 214012 138048 214064 138100
rect 226432 138048 226484 138100
rect 213920 137980 213972 138032
rect 226800 137980 226852 138032
rect 216680 137912 216732 137964
rect 227444 137912 227496 137964
rect 213920 136688 213972 136740
rect 227076 136688 227128 136740
rect 104716 136620 104768 136672
rect 116400 136620 116452 136672
rect 214012 136620 214064 136672
rect 227444 136620 227496 136672
rect 104348 135260 104400 135312
rect 115940 135260 115992 135312
rect 213920 135260 213972 135312
rect 227628 135260 227680 135312
rect 104808 135192 104860 135244
rect 113548 135192 113600 135244
rect 341524 135192 341576 135244
rect 580172 135192 580224 135244
rect 214012 133968 214064 134020
rect 227536 133968 227588 134020
rect 100484 133900 100536 133952
rect 103612 133900 103664 133952
rect 109868 133900 109920 133952
rect 116400 133900 116452 133952
rect 213920 133900 213972 133952
rect 227352 133900 227404 133952
rect 104808 133832 104860 133884
rect 115848 133832 115900 133884
rect 114560 132880 114612 132932
rect 117136 132880 117188 132932
rect 213920 132540 213972 132592
rect 226708 132540 226760 132592
rect 214012 132472 214064 132524
rect 227444 132472 227496 132524
rect 113916 131180 113968 131232
rect 116400 131180 116452 131232
rect 213920 131180 213972 131232
rect 226524 131180 226576 131232
rect 100392 131112 100444 131164
rect 115940 131112 115992 131164
rect 214012 131112 214064 131164
rect 227076 131112 227128 131164
rect 103980 130704 104032 130756
rect 109868 130704 109920 130756
rect 213920 129752 213972 129804
rect 227536 129752 227588 129804
rect 104808 129684 104860 129736
rect 114560 129684 114612 129736
rect 116400 129276 116452 129328
rect 10416 129208 10468 129260
rect 213920 129004 213972 129056
rect 227444 129004 227496 129056
rect 213920 128324 213972 128376
rect 226340 128324 226392 128376
rect 9036 128256 9088 128308
rect 116400 128256 116452 128308
rect 104808 128188 104860 128240
rect 113916 128188 113968 128240
rect 103612 127576 103664 127628
rect 116308 127576 116360 127628
rect 213920 127576 213972 127628
rect 227444 127576 227496 127628
rect 213920 126964 213972 127016
rect 227444 126964 227496 127016
rect 10324 126896 10376 126948
rect 116400 126896 116452 126948
rect 213920 126216 213972 126268
rect 227444 126216 227496 126268
rect 213920 125604 213972 125656
rect 227444 125604 227496 125656
rect 8944 125536 8996 125588
rect 116400 125536 116452 125588
rect 214380 125536 214432 125588
rect 214472 125536 214524 125588
rect 78220 125468 78272 125520
rect 100392 125468 100444 125520
rect 213920 124856 213972 124908
rect 227260 124856 227312 124908
rect 213920 124108 213972 124160
rect 227260 124108 227312 124160
rect 213920 123428 213972 123480
rect 227260 123428 227312 123480
rect 213920 122748 213972 122800
rect 227444 122748 227496 122800
rect 213920 122068 213972 122120
rect 227444 122068 227496 122120
rect 50988 121456 51040 121508
rect 116400 121456 116452 121508
rect 213920 121388 213972 121440
rect 227444 121388 227496 121440
rect 213920 120708 213972 120760
rect 227444 120708 227496 120760
rect 94504 120096 94556 120148
rect 116400 120096 116452 120148
rect 213920 120028 213972 120080
rect 227444 120028 227496 120080
rect 94688 118668 94740 118720
rect 116400 118668 116452 118720
rect 213920 118600 213972 118652
rect 226432 118600 226484 118652
rect 214012 118532 214064 118584
rect 226340 118532 226392 118584
rect 94596 117308 94648 117360
rect 116400 117308 116452 117360
rect 214012 117240 214064 117292
rect 227444 117240 227496 117292
rect 213920 117172 213972 117224
rect 226248 117172 226300 117224
rect 94964 116016 95016 116068
rect 116124 116016 116176 116068
rect 94780 115948 94832 116000
rect 116400 115948 116452 116000
rect 214012 115880 214064 115932
rect 227444 115880 227496 115932
rect 213920 115812 213972 115864
rect 226156 115812 226208 115864
rect 94872 114520 94924 114572
rect 116400 114520 116452 114572
rect 214012 114452 214064 114504
rect 227076 114452 227128 114504
rect 213920 114384 213972 114436
rect 226248 114384 226300 114436
rect 97264 113160 97316 113212
rect 116400 113160 116452 113212
rect 213920 113092 213972 113144
rect 226156 113092 226208 113144
rect 94412 111800 94464 111852
rect 116400 111800 116452 111852
rect 214012 111732 214064 111784
rect 226248 111732 226300 111784
rect 213920 111664 213972 111716
rect 226064 111664 226116 111716
rect 95884 110440 95936 110492
rect 116400 110440 116452 110492
rect 214012 110372 214064 110424
rect 226156 110372 226208 110424
rect 213920 110304 213972 110356
rect 225972 110304 226024 110356
rect 95148 109012 95200 109064
rect 116400 109012 116452 109064
rect 214012 108944 214064 108996
rect 226248 108944 226300 108996
rect 213920 108876 213972 108928
rect 225880 108876 225932 108928
rect 102784 107720 102836 107772
rect 116308 107720 116360 107772
rect 95056 107652 95108 107704
rect 116400 107652 116452 107704
rect 213920 107584 213972 107636
rect 226064 107584 226116 107636
rect 98644 106292 98696 106344
rect 116400 106292 116452 106344
rect 213920 106224 213972 106276
rect 225788 106224 225840 106276
rect 214012 106156 214064 106208
rect 226248 106156 226300 106208
rect 94320 104864 94372 104916
rect 116400 104864 116452 104916
rect 224776 104864 224828 104916
rect 227444 104864 227496 104916
rect 214012 104796 214064 104848
rect 226156 104796 226208 104848
rect 213920 104728 213972 104780
rect 225604 104728 225656 104780
rect 224868 103640 224920 103692
rect 227444 103640 227496 103692
rect 101404 103504 101456 103556
rect 116400 103504 116452 103556
rect 214012 103436 214064 103488
rect 225972 103436 226024 103488
rect 213920 103368 213972 103420
rect 225696 103368 225748 103420
rect 94228 102144 94280 102196
rect 116308 102144 116360 102196
rect 213920 102076 213972 102128
rect 225880 102076 225932 102128
rect 314200 102076 314252 102128
rect 338396 102076 338448 102128
rect 105544 100784 105596 100836
rect 116400 100784 116452 100836
rect 104164 100716 104216 100768
rect 116308 100716 116360 100768
rect 213920 100648 213972 100700
rect 226156 100648 226208 100700
rect 232136 100648 232188 100700
rect 258080 100648 258132 100700
rect 214012 100580 214064 100632
rect 226064 100580 226116 100632
rect 97356 99356 97408 99408
rect 116400 99356 116452 99408
rect 214656 99288 214708 99340
rect 226248 99288 226300 99340
rect 232136 99288 232188 99340
rect 232504 99288 232556 99340
rect 215116 99220 215168 99272
rect 224776 99220 224828 99272
rect 94136 97996 94188 98048
rect 116400 97996 116452 98048
rect 214104 97928 214156 97980
rect 224868 97928 224920 97980
rect 213920 97588 213972 97640
rect 215944 97588 215996 97640
rect 100024 96636 100076 96688
rect 116400 96636 116452 96688
rect 94688 95208 94740 95260
rect 116308 95208 116360 95260
rect 215116 95140 215168 95192
rect 576124 95140 576176 95192
rect 94504 93848 94556 93900
rect 116400 93848 116452 93900
rect 215208 93780 215260 93832
rect 578884 93780 578936 93832
rect 215116 93712 215168 93764
rect 577504 93712 577556 93764
rect 95148 93508 95200 93560
rect 97264 93508 97316 93560
rect 95976 92488 96028 92540
rect 116400 92488 116452 92540
rect 94596 91808 94648 91860
rect 95884 91808 95936 91860
rect 94596 91060 94648 91112
rect 116400 91060 116452 91112
rect 94780 90992 94832 91044
rect 102784 90992 102836 91044
rect 98736 90312 98788 90364
rect 116492 90312 116544 90364
rect 102876 89700 102928 89752
rect 116400 89700 116452 89752
rect 94964 88340 95016 88392
rect 115940 88340 115992 88392
rect 340144 88272 340196 88324
rect 580172 88272 580224 88324
rect 95148 88204 95200 88256
rect 98644 88204 98696 88256
rect 97264 86980 97316 87032
rect 116400 86980 116452 87032
rect 94412 86572 94464 86624
rect 101404 86572 101456 86624
rect 101496 85620 101548 85672
rect 116400 85620 116452 85672
rect 94780 85552 94832 85604
rect 116308 85552 116360 85604
rect 215116 85552 215168 85604
rect 224224 85552 224276 85604
rect 95148 85484 95200 85536
rect 104164 85484 104216 85536
rect 94872 84192 94924 84244
rect 116400 84192 116452 84244
rect 215116 84192 215168 84244
rect 225604 84192 225656 84244
rect 95148 84124 95200 84176
rect 105544 84124 105596 84176
rect 214012 83512 214064 83564
rect 214380 83512 214432 83564
rect 284484 83512 284536 83564
rect 413284 83512 413336 83564
rect 320824 83444 320876 83496
rect 580264 83444 580316 83496
rect 94228 83376 94280 83428
rect 97356 83376 97408 83428
rect 95884 82832 95936 82884
rect 116400 82832 116452 82884
rect 215944 82832 215996 82884
rect 248144 82832 248196 82884
rect 95056 81404 95108 81456
rect 115940 81404 115992 81456
rect 214196 81404 214248 81456
rect 226984 81404 227036 81456
rect 215024 81336 215076 81388
rect 227352 81336 227404 81388
rect 94412 81268 94464 81320
rect 100024 81268 100076 81320
rect 214840 81268 214892 81320
rect 227444 81268 227496 81320
rect 215116 80112 215168 80164
rect 220176 80112 220228 80164
rect 98644 80044 98696 80096
rect 116400 80044 116452 80096
rect 232412 80112 232464 80164
rect 94412 79976 94464 80028
rect 98736 79976 98788 80028
rect 214288 79976 214340 80028
rect 227536 79976 227588 80028
rect 232320 79976 232372 80028
rect 214564 79908 214616 79960
rect 227444 79908 227496 79960
rect 100024 78752 100076 78804
rect 116400 78752 116452 78804
rect 213920 78752 213972 78804
rect 220820 78752 220872 78804
rect 95148 78684 95200 78736
rect 116216 78684 116268 78736
rect 214012 78616 214064 78668
rect 227536 78616 227588 78668
rect 214748 78548 214800 78600
rect 227444 78548 227496 78600
rect 94228 78208 94280 78260
rect 95976 78208 96028 78260
rect 94688 77256 94740 77308
rect 116400 77256 116452 77308
rect 213920 77256 213972 77308
rect 218796 77256 218848 77308
rect 214656 77188 214708 77240
rect 227444 77188 227496 77240
rect 214472 77120 214524 77172
rect 227536 77120 227588 77172
rect 213920 76032 213972 76084
rect 219440 76032 219492 76084
rect 97356 75896 97408 75948
rect 116400 75896 116452 75948
rect 224224 75828 224276 75880
rect 227444 75828 227496 75880
rect 94596 75692 94648 75744
rect 102876 75692 102928 75744
rect 214196 75692 214248 75744
rect 227444 75692 227496 75744
rect 213920 74604 213972 74656
rect 216036 74604 216088 74656
rect 94504 74536 94556 74588
rect 116400 74536 116452 74588
rect 214380 74400 214432 74452
rect 227444 74468 227496 74520
rect 94596 74264 94648 74316
rect 97264 74264 97316 74316
rect 95976 73176 96028 73228
rect 116400 73176 116452 73228
rect 213920 73176 213972 73228
rect 218060 73176 218112 73228
rect 215208 73108 215260 73160
rect 227444 73108 227496 73160
rect 220176 73040 220228 73092
rect 227536 73040 227588 73092
rect 94412 72904 94464 72956
rect 101496 72904 101548 72956
rect 94964 71748 95016 71800
rect 116400 71748 116452 71800
rect 214932 71680 214984 71732
rect 227444 71680 227496 71732
rect 220820 71612 220872 71664
rect 227536 71612 227588 71664
rect 214012 70456 214064 70508
rect 224500 70456 224552 70508
rect 94596 70388 94648 70440
rect 116400 70388 116452 70440
rect 213920 70388 213972 70440
rect 224408 70388 224460 70440
rect 214840 70320 214892 70372
rect 227444 70320 227496 70372
rect 94872 70252 94924 70304
rect 95884 70252 95936 70304
rect 218796 70252 218848 70304
rect 226524 70252 226576 70304
rect 215116 69096 215168 69148
rect 224224 69096 224276 69148
rect 94412 69028 94464 69080
rect 116400 69028 116452 69080
rect 214656 69028 214708 69080
rect 224132 69028 224184 69080
rect 215024 68960 215076 69012
rect 227444 68960 227496 69012
rect 219440 68892 219492 68944
rect 227536 68892 227588 68944
rect 93860 68484 93912 68536
rect 98644 68484 98696 68536
rect 214472 67668 214524 67720
rect 224684 67668 224736 67720
rect 94872 67600 94924 67652
rect 116400 67600 116452 67652
rect 215116 67600 215168 67652
rect 224868 67600 224920 67652
rect 214748 67532 214800 67584
rect 227444 67532 227496 67584
rect 216036 67464 216088 67516
rect 227536 67464 227588 67516
rect 95148 66852 95200 66904
rect 100024 66852 100076 66904
rect 94780 66240 94832 66292
rect 116400 66240 116452 66292
rect 215116 66240 215168 66292
rect 224316 66240 224368 66292
rect 214104 66172 214156 66224
rect 227444 66172 227496 66224
rect 218060 66104 218112 66156
rect 227536 66104 227588 66156
rect 214380 65492 214432 65544
rect 216772 65492 216824 65544
rect 94688 65288 94740 65340
rect 97356 65288 97408 65340
rect 94320 64880 94372 64932
rect 116400 64880 116452 64932
rect 214012 64880 214064 64932
rect 224592 64880 224644 64932
rect 214564 64812 214616 64864
rect 227444 64812 227496 64864
rect 224500 64472 224552 64524
rect 227444 64472 227496 64524
rect 224408 64268 224460 64320
rect 227536 64268 227588 64320
rect 94228 63656 94280 63708
rect 94780 63656 94832 63708
rect 214564 63588 214616 63640
rect 216956 63588 217008 63640
rect 95148 63520 95200 63572
rect 115940 63520 115992 63572
rect 215116 63520 215168 63572
rect 224040 63520 224092 63572
rect 94872 63452 94924 63504
rect 95976 63452 96028 63504
rect 224132 63452 224184 63504
rect 227444 63452 227496 63504
rect 224224 63384 224276 63436
rect 227536 63384 227588 63436
rect 487620 62772 487672 62824
rect 576216 62772 576268 62824
rect 94688 62160 94740 62212
rect 116216 62160 116268 62212
rect 214656 62160 214708 62212
rect 216680 62160 216732 62212
rect 94504 62092 94556 62144
rect 116400 62092 116452 62144
rect 215116 62092 215168 62144
rect 224132 62092 224184 62144
rect 93952 62024 94004 62076
rect 116584 62024 116636 62076
rect 224684 62024 224736 62076
rect 227536 62024 227588 62076
rect 224868 61956 224920 62008
rect 226708 61956 226760 62008
rect 214564 61208 214616 61260
rect 216864 61208 216916 61260
rect 94964 60732 95016 60784
rect 116400 60732 116452 60784
rect 215116 60732 215168 60784
rect 224224 60732 224276 60784
rect 216772 60664 216824 60716
rect 227444 60664 227496 60716
rect 224316 60596 224368 60648
rect 227076 60596 227128 60648
rect 95056 59372 95108 59424
rect 116400 59372 116452 59424
rect 214564 59372 214616 59424
rect 217600 59372 217652 59424
rect 216956 59304 217008 59356
rect 227536 59304 227588 59356
rect 224592 59236 224644 59288
rect 227444 59236 227496 59288
rect 214104 58012 214156 58064
rect 217508 58012 217560 58064
rect 94412 57944 94464 57996
rect 116400 57944 116452 57996
rect 214196 57944 214248 57996
rect 217416 57944 217468 57996
rect 216680 57876 216732 57928
rect 227444 57876 227496 57928
rect 224040 57808 224092 57860
rect 227260 57808 227312 57860
rect 213920 56652 213972 56704
rect 216772 56652 216824 56704
rect 93860 56584 93912 56636
rect 116308 56584 116360 56636
rect 214012 56584 214064 56636
rect 216680 56584 216732 56636
rect 216864 56516 216916 56568
rect 227444 56516 227496 56568
rect 224132 56448 224184 56500
rect 227260 56448 227312 56500
rect 94044 55292 94096 55344
rect 116400 55292 116452 55344
rect 93952 55224 94004 55276
rect 116308 55224 116360 55276
rect 215116 55224 215168 55276
rect 227536 55224 227588 55276
rect 217600 55156 217652 55208
rect 224224 55156 224276 55208
rect 227444 55156 227496 55208
rect 226524 55020 226576 55072
rect 215116 53864 215168 53916
rect 226984 53864 227036 53916
rect 94780 53796 94832 53848
rect 116400 53796 116452 53848
rect 214748 53796 214800 53848
rect 226616 53796 226668 53848
rect 217508 53728 217560 53780
rect 227444 53728 227496 53780
rect 217416 53660 217468 53712
rect 226524 53660 226576 53712
rect 215116 52504 215168 52556
rect 226800 52504 226852 52556
rect 95148 52436 95200 52488
rect 116400 52436 116452 52488
rect 214748 52436 214800 52488
rect 226708 52436 226760 52488
rect 216680 52368 216732 52420
rect 227444 52368 227496 52420
rect 216772 52300 216824 52352
rect 227260 52300 227312 52352
rect 215116 51144 215168 51196
rect 226340 51144 226392 51196
rect 94228 51076 94280 51128
rect 115940 51076 115992 51128
rect 214104 51076 214156 51128
rect 226524 51076 226576 51128
rect 215116 49784 215168 49836
rect 227628 49784 227680 49836
rect 95056 49716 95108 49768
rect 116400 49716 116452 49768
rect 215208 49716 215260 49768
rect 227536 49716 227588 49768
rect 94504 48356 94556 48408
rect 116124 48356 116176 48408
rect 94412 48288 94464 48340
rect 116400 48288 116452 48340
rect 215116 48288 215168 48340
rect 227352 48288 227404 48340
rect 214748 46996 214800 47048
rect 227444 46996 227496 47048
rect 94136 46928 94188 46980
rect 116400 46928 116452 46980
rect 214012 46928 214064 46980
rect 226708 46928 226760 46980
rect 215116 45636 215168 45688
rect 227260 45636 227312 45688
rect 93952 45568 94004 45620
rect 116400 45568 116452 45620
rect 215208 45568 215260 45620
rect 227076 45568 227128 45620
rect 215208 44208 215260 44260
rect 227444 44208 227496 44260
rect 94780 44140 94832 44192
rect 116400 44140 116452 44192
rect 215116 44140 215168 44192
rect 227536 44140 227588 44192
rect 94596 42780 94648 42832
rect 115940 42780 115992 42832
rect 214380 42780 214432 42832
rect 226432 42780 226484 42832
rect 215116 41488 215168 41540
rect 226616 41488 226668 41540
rect 95148 41420 95200 41472
rect 116400 41420 116452 41472
rect 214104 41420 214156 41472
rect 226340 41420 226392 41472
rect 560944 41352 560996 41404
rect 580172 41352 580224 41404
rect 94504 40128 94556 40180
rect 116308 40128 116360 40180
rect 215116 40128 215168 40180
rect 227444 40128 227496 40180
rect 95056 40060 95108 40112
rect 116400 40060 116452 40112
rect 214656 40060 214708 40112
rect 227076 40060 227128 40112
rect 215116 38700 215168 38752
rect 227536 38700 227588 38752
rect 94596 38632 94648 38684
rect 116400 38632 116452 38684
rect 214564 38632 214616 38684
rect 226708 38632 226760 38684
rect 93860 37272 93912 37324
rect 116400 37272 116452 37324
rect 215116 37272 215168 37324
rect 227444 37272 227496 37324
rect 214104 35980 214156 36032
rect 226708 35980 226760 36032
rect 93952 35912 94004 35964
rect 116400 35912 116452 35964
rect 215116 35912 215168 35964
rect 227444 35912 227496 35964
rect 215116 34552 215168 34604
rect 227352 34552 227404 34604
rect 95148 34484 95200 34536
rect 116400 34484 116452 34536
rect 214656 34484 214708 34536
rect 227444 34484 227496 34536
rect 214564 33192 214616 33244
rect 227444 33192 227496 33244
rect 95148 33124 95200 33176
rect 116308 33124 116360 33176
rect 215116 33124 215168 33176
rect 227536 33124 227588 33176
rect 213920 32512 213972 32564
rect 215944 32512 215996 32564
rect 95148 32376 95200 32428
rect 116400 32376 116452 32428
rect 215116 32376 215168 32428
rect 227444 32376 227496 32428
rect 71688 31764 71740 31816
rect 116400 31764 116452 31816
rect 29920 31288 29972 31340
rect 32312 31288 32364 31340
rect 105544 30268 105596 30320
rect 195428 30268 195480 30320
rect 95884 30200 95936 30252
rect 185032 30200 185084 30252
rect 50344 30132 50396 30184
rect 163504 30132 163556 30184
rect 174636 30132 174688 30184
rect 82084 30064 82136 30116
rect 177212 30064 177264 30116
rect 53104 29996 53156 30048
rect 148600 29996 148652 30048
rect 164884 29996 164936 30048
rect 179788 29996 179840 30048
rect 75184 29928 75236 29980
rect 172060 29928 172112 29980
rect 31024 29860 31076 29912
rect 127716 29860 127768 29912
rect 143356 29860 143408 29912
rect 166264 29860 166316 29912
rect 182456 29860 182508 29912
rect 66904 29792 66956 29844
rect 166816 29792 166868 29844
rect 169116 29792 169168 29844
rect 187608 29792 187660 29844
rect 25504 29724 25556 29776
rect 126888 29724 126940 29776
rect 169024 29724 169076 29776
rect 192852 29724 192904 29776
rect 60004 29656 60056 29708
rect 161572 29656 161624 29708
rect 171784 29656 171836 29708
rect 198096 29656 198148 29708
rect 28264 29588 28316 29640
rect 130384 29588 130436 29640
rect 173164 29588 173216 29640
rect 205824 29588 205876 29640
rect 111708 29520 111760 29572
rect 200672 29520 200724 29572
rect 46204 29384 46256 29436
rect 115848 29452 115900 29504
rect 203248 29452 203300 29504
rect 133788 29384 133840 29436
rect 102784 29316 102836 29368
rect 190276 29316 190328 29368
rect 117964 29248 118016 29300
rect 122748 29248 122800 29300
rect 208492 29248 208544 29300
rect 68008 29180 68060 29232
rect 123392 29180 123444 29232
rect 125508 29180 125560 29232
rect 211068 29180 211120 29232
rect 57244 29112 57296 29164
rect 131212 29112 131264 29164
rect 61384 29044 61436 29096
rect 134708 29044 134760 29096
rect 162124 29044 162176 29096
rect 119988 28976 120040 29028
rect 124312 28976 124364 29028
rect 152464 28976 152516 29028
rect 156420 28976 156472 29028
rect 156604 28976 156656 29028
rect 158996 28976 159048 29028
rect 159364 28976 159416 29028
rect 164240 28976 164292 29028
rect 169392 28976 169444 29028
rect 68008 28951 68060 28960
rect 68008 28917 68017 28951
rect 68017 28917 68051 28951
rect 68051 28917 68060 28951
rect 68008 28908 68060 28917
rect 103428 28364 103480 28416
rect 194600 28364 194652 28416
rect 60648 28296 60700 28348
rect 163320 28296 163372 28348
rect 10324 28228 10376 28280
rect 121644 28228 121696 28280
rect 3424 27548 3476 27600
rect 411260 27548 411312 27600
rect 110328 26868 110380 26920
rect 199752 26868 199804 26920
rect 138112 26732 138164 26784
rect 138756 26732 138808 26784
rect 144920 26732 144972 26784
rect 145748 26732 145800 26784
rect 149060 26732 149112 26784
rect 149980 26732 150032 26784
rect 154580 26732 154632 26784
rect 155132 26732 155184 26784
rect 197176 26188 197228 26240
rect 67548 25576 67600 25628
rect 168564 25576 168616 25628
rect 11704 25508 11756 25560
rect 125140 25508 125192 25560
rect 114468 24216 114520 24268
rect 202420 24216 202472 24268
rect 74448 24148 74500 24200
rect 173716 24148 173768 24200
rect 52368 24080 52420 24132
rect 157248 24080 157300 24132
rect 125416 22856 125468 22908
rect 210240 22856 210292 22908
rect 85488 22788 85540 22840
rect 181536 22788 181588 22840
rect 63408 22720 63460 22772
rect 165068 22720 165120 22772
rect 121460 22448 121512 22500
rect 122196 22448 122248 22500
rect 203064 22108 203116 22160
rect 203892 22108 203944 22160
rect 121460 22040 121512 22092
rect 121644 22040 121696 22092
rect 96528 21428 96580 21480
rect 189172 21428 189224 21480
rect 59268 21360 59320 21412
rect 161572 21360 161624 21412
rect 107568 20680 107620 20732
rect 99196 20000 99248 20052
rect 191932 20000 191984 20052
rect 66168 19932 66220 19984
rect 167000 19932 167052 19984
rect 68100 19320 68152 19372
rect 66168 19252 66220 19304
rect 121644 19295 121696 19304
rect 121644 19261 121653 19295
rect 121653 19261 121687 19295
rect 121687 19261 121696 19295
rect 121644 19252 121696 19261
rect 182272 19252 182324 19304
rect 184572 19252 184624 19304
rect 185032 19252 185084 19304
rect 117136 18708 117188 18760
rect 204260 18708 204312 18760
rect 89628 18640 89680 18692
rect 183560 18640 183612 18692
rect 53748 18572 53800 18624
rect 157340 18572 157392 18624
rect 121368 17348 121420 17400
rect 207020 17348 207072 17400
rect 92388 17280 92440 17332
rect 186412 17280 186464 17332
rect 56508 17212 56560 17264
rect 158812 17212 158864 17264
rect 492864 16396 492916 16448
rect 493600 16396 493652 16448
rect 378048 16328 378100 16380
rect 494796 16328 494848 16380
rect 318064 16260 318116 16312
rect 458364 16260 458416 16312
rect 300124 16192 300176 16244
rect 456340 16192 456392 16244
rect 286324 16124 286376 16176
rect 452844 16124 452896 16176
rect 296628 16056 296680 16108
rect 468576 16056 468628 16108
rect 285588 15988 285640 16040
rect 465172 15988 465224 16040
rect 82728 15920 82780 15972
rect 178132 15920 178184 15972
rect 280068 15920 280120 15972
rect 463608 15920 463660 15972
rect 48228 15852 48280 15904
rect 154672 15852 154724 15904
rect 278688 15852 278740 15904
rect 462872 15852 462924 15904
rect 273168 15784 273220 15836
rect 461308 15784 461360 15836
rect 266268 15716 266320 15768
rect 459008 15716 459060 15768
rect 259368 15648 259420 15700
rect 456708 15648 456760 15700
rect 240048 15580 240100 15632
rect 450544 15580 450596 15632
rect 233148 15512 233200 15564
rect 448244 15512 448296 15564
rect 222108 15444 222160 15496
rect 444840 15444 444892 15496
rect 202788 15376 202840 15428
rect 438676 15376 438728 15428
rect 204168 15308 204220 15360
rect 439044 15308 439096 15360
rect 195888 15240 195940 15292
rect 436376 15240 436428 15292
rect 188988 15172 189040 15224
rect 434076 15172 434128 15224
rect 456984 15172 457036 15224
rect 457444 15172 457496 15224
rect 354588 15104 354640 15156
rect 487344 15104 487396 15156
rect 503628 15104 503680 15156
rect 535644 15104 535696 15156
rect 538128 15104 538180 15156
rect 546776 15104 546828 15156
rect 340788 15036 340840 15088
rect 482744 15036 482796 15088
rect 489828 15036 489880 15088
rect 531044 15036 531096 15088
rect 535368 15036 535420 15088
rect 545672 15036 545724 15088
rect 332508 14968 332560 15020
rect 480444 14968 480496 15020
rect 496728 14968 496780 15020
rect 533344 14968 533396 15020
rect 533988 14968 534040 15020
rect 545304 14968 545356 15020
rect 325608 14900 325660 14952
rect 478144 14900 478196 14952
rect 487068 14900 487120 14952
rect 529940 14900 529992 14952
rect 531228 14900 531280 14952
rect 544476 14900 544528 14952
rect 555240 14900 555292 14952
rect 563060 14900 563112 14952
rect 318708 14832 318760 14884
rect 475844 14832 475896 14884
rect 482928 14832 482980 14884
rect 528744 14832 528796 14884
rect 532608 14832 532660 14884
rect 544844 14832 544896 14884
rect 311808 14764 311860 14816
rect 473544 14764 473596 14816
rect 478788 14764 478840 14816
rect 527272 14764 527324 14816
rect 529848 14764 529900 14816
rect 543740 14764 543792 14816
rect 305000 14696 305052 14748
rect 468944 14696 468996 14748
rect 476028 14696 476080 14748
rect 526444 14696 526496 14748
rect 526628 14696 526680 14748
rect 542544 14696 542596 14748
rect 302240 14628 302292 14680
rect 466644 14628 466696 14680
rect 469036 14628 469088 14680
rect 214564 14560 214616 14612
rect 424140 14560 424192 14612
rect 447784 14560 447836 14612
rect 517244 14560 517296 14612
rect 523684 14628 523736 14680
rect 540244 14628 540296 14680
rect 524144 14560 524196 14612
rect 524328 14560 524380 14612
rect 542176 14560 542228 14612
rect 204904 14492 204956 14544
rect 422944 14492 422996 14544
rect 443828 14492 443880 14544
rect 514944 14492 514996 14544
rect 521568 14492 521620 14544
rect 541072 14492 541124 14544
rect 546316 14492 546368 14544
rect 549076 14492 549128 14544
rect 554872 14492 554924 14544
rect 563152 14492 563204 14544
rect 13728 14424 13780 14476
rect 128544 14424 128596 14476
rect 174176 14424 174228 14476
rect 421840 14424 421892 14476
rect 511540 14424 511592 14476
rect 513564 14424 513616 14476
rect 514024 14424 514076 14476
rect 517428 14424 517480 14476
rect 539876 14424 539928 14476
rect 547788 14424 547840 14476
rect 549904 14424 549956 14476
rect 361488 14356 361540 14408
rect 489644 14356 489696 14408
rect 502524 14356 502576 14408
rect 503168 14356 503220 14408
rect 507768 14356 507820 14408
rect 536840 14356 536892 14408
rect 544384 14356 544436 14408
rect 546408 14356 546460 14408
rect 547696 14356 547748 14408
rect 549444 14356 549496 14408
rect 551376 14356 551428 14408
rect 551928 14356 551980 14408
rect 368388 14288 368440 14340
rect 491944 14288 491996 14340
rect 514024 14288 514076 14340
rect 521844 14288 521896 14340
rect 522304 14288 522356 14340
rect 539140 14288 539192 14340
rect 548340 14288 548392 14340
rect 375196 14220 375248 14272
rect 494244 14220 494296 14272
rect 520924 14220 520976 14272
rect 537944 14220 537996 14272
rect 383568 14152 383620 14204
rect 496544 14152 496596 14204
rect 525156 14152 525208 14204
rect 541440 14152 541492 14204
rect 390468 14084 390520 14136
rect 498844 14084 498896 14136
rect 519728 14084 519780 14136
rect 534540 14084 534592 14136
rect 536748 14084 536800 14136
rect 546040 14220 546092 14272
rect 553676 14220 553728 14272
rect 556988 14220 557040 14272
rect 543648 14152 543700 14204
rect 545764 14152 545816 14204
rect 547144 14152 547196 14204
rect 554044 14152 554096 14204
rect 556896 14152 556948 14204
rect 552572 14084 552624 14136
rect 555240 14084 555292 14136
rect 313280 14016 313332 14068
rect 420644 14016 420696 14068
rect 420828 14016 420880 14068
rect 508044 14016 508096 14068
rect 528468 14016 528520 14068
rect 543372 14016 543424 14068
rect 545028 14016 545080 14068
rect 548708 14016 548760 14068
rect 552940 14016 552992 14068
rect 555424 14016 555476 14068
rect 397368 13948 397420 14000
rect 501144 13948 501196 14000
rect 509884 13948 509936 14000
rect 512644 13948 512696 14000
rect 518348 13948 518400 14000
rect 532240 13948 532292 14000
rect 553308 13948 553360 14000
rect 555516 13948 555568 14000
rect 408408 13880 408460 13932
rect 504640 13880 504692 13932
rect 511264 13880 511316 13932
rect 513840 13880 513892 13932
rect 555608 13880 555660 13932
rect 555976 13880 556028 13932
rect 556344 13880 556396 13932
rect 557356 13880 557408 13932
rect 557540 13880 557592 13932
rect 558828 13880 558880 13932
rect 559104 13880 559156 13932
rect 560116 13880 560168 13932
rect 330300 13812 330352 13864
rect 425244 13812 425296 13864
rect 425428 13812 425480 13864
rect 268384 13744 268436 13796
rect 422300 13744 422352 13796
rect 457444 13812 457496 13864
rect 519544 13812 519596 13864
rect 551744 13812 551796 13864
rect 553400 13812 553452 13864
rect 554504 13812 554556 13864
rect 556712 13812 556764 13864
rect 556804 13812 556856 13864
rect 557448 13812 557500 13864
rect 557908 13812 557960 13864
rect 558644 13812 558696 13864
rect 559840 13812 559892 13864
rect 560208 13812 560260 13864
rect 560576 13812 560628 13864
rect 561496 13812 561548 13864
rect 463240 13744 463292 13796
rect 261484 13676 261536 13728
rect 433708 13676 433760 13728
rect 433984 13676 434036 13728
rect 470140 13676 470192 13728
rect 257344 13608 257396 13660
rect 431408 13608 431460 13660
rect 436008 13608 436060 13660
rect 438860 13608 438912 13660
rect 439320 13608 439372 13660
rect 211068 13540 211120 13592
rect 441344 13540 441396 13592
rect 219256 13472 219308 13524
rect 443644 13472 443696 13524
rect 208308 13404 208360 13456
rect 440240 13404 440292 13456
rect 191748 13336 191800 13388
rect 434904 13336 434956 13388
rect 435364 13336 435416 13388
rect 474740 13608 474792 13660
rect 464252 13472 464304 13524
rect 500040 13472 500092 13524
rect 445668 13404 445720 13456
rect 461584 13404 461636 13456
rect 490840 13404 490892 13456
rect 491208 13404 491260 13456
rect 531504 13404 531556 13456
rect 461032 13336 461084 13388
rect 461676 13336 461728 13388
rect 467748 13336 467800 13388
rect 523776 13336 523828 13388
rect 432604 13268 432656 13320
rect 439320 13268 439372 13320
rect 506940 13268 506992 13320
rect 131028 13200 131080 13252
rect 415308 13200 415360 13252
rect 419448 13200 419500 13252
rect 508504 13200 508556 13252
rect 516048 13200 516100 13252
rect 539508 13200 539560 13252
rect 46848 13132 46900 13184
rect 152096 13132 152148 13184
rect 173808 13132 173860 13184
rect 429108 13132 429160 13184
rect 429200 13132 429252 13184
rect 437572 13132 437624 13184
rect 437940 13132 437992 13184
rect 516876 13132 516928 13184
rect 126888 13064 126940 13116
rect 414204 13064 414256 13116
rect 416688 13064 416740 13116
rect 507308 13064 507360 13116
rect 510528 13064 510580 13116
rect 537576 13064 537628 13116
rect 304264 12996 304316 13048
rect 454040 12996 454092 13048
rect 349068 12928 349120 12980
rect 485504 12928 485556 12980
rect 351828 12860 351880 12912
rect 393228 12860 393280 12912
rect 402980 12860 403032 12912
rect 412548 12860 412600 12912
rect 422300 12860 422352 12912
rect 431868 12860 431920 12912
rect 486608 12860 486660 12912
rect 488908 12792 488960 12844
rect 358728 12656 358780 12708
rect 387708 12724 387760 12776
rect 498108 12724 498160 12776
rect 364984 12656 365036 12708
rect 464344 12656 464396 12708
rect 409788 12588 409840 12640
rect 505008 12588 505060 12640
rect 423588 12520 423640 12572
rect 509608 12520 509660 12572
rect 528836 12520 528888 12572
rect 529296 12520 529348 12572
rect 67548 12452 67600 12504
rect 179512 12452 179564 12504
rect 393228 12452 393280 12504
rect 403072 12452 403124 12504
rect 410432 12452 410484 12504
rect 410524 12452 410576 12504
rect 460940 12452 460992 12504
rect 121644 12427 121696 12436
rect 121644 12393 121653 12427
rect 121653 12393 121687 12427
rect 121687 12393 121696 12427
rect 121644 12384 121696 12393
rect 275284 12384 275336 12436
rect 445944 12384 445996 12436
rect 497096 12384 497148 12436
rect 497740 12384 497792 12436
rect 555240 12384 555292 12436
rect 555884 12384 555936 12436
rect 225604 12316 225656 12368
rect 427544 12316 427596 12368
rect 428924 12359 428976 12368
rect 428924 12325 428933 12359
rect 428933 12325 428967 12359
rect 428967 12325 428976 12359
rect 428924 12316 428976 12325
rect 431684 12316 431736 12368
rect 467840 12316 467892 12368
rect 196808 12248 196860 12300
rect 436744 12248 436796 12300
rect 194508 12180 194560 12232
rect 435640 12180 435692 12232
rect 190368 12112 190420 12164
rect 229100 12112 229152 12164
rect 238668 12112 238720 12164
rect 248420 12112 248472 12164
rect 257988 12112 258040 12164
rect 267740 12112 267792 12164
rect 277308 12112 277360 12164
rect 287060 12112 287112 12164
rect 306380 12112 306432 12164
rect 315948 12112 316000 12164
rect 325700 12112 325752 12164
rect 335268 12112 335320 12164
rect 186228 12044 186280 12096
rect 433340 12112 433392 12164
rect 182548 11976 182600 12028
rect 432144 12044 432196 12096
rect 433432 12044 433484 12096
rect 441712 12044 441764 12096
rect 442632 12044 442684 12096
rect 456892 12044 456944 12096
rect 457628 12044 457680 12096
rect 179328 11908 179380 11960
rect 431040 11976 431092 12028
rect 465540 12112 465592 12164
rect 175464 11840 175516 11892
rect 429568 11908 429620 11960
rect 430488 11908 430540 11960
rect 463792 11976 463844 12028
rect 464436 11976 464488 12028
rect 469404 11976 469456 12028
rect 470232 11976 470284 12028
rect 479340 11976 479392 12028
rect 436100 11908 436152 11960
rect 38568 11772 38620 11824
rect 147772 11772 147824 11824
rect 160008 11772 160060 11824
rect 434444 11840 434496 11892
rect 437480 11840 437532 11892
rect 438032 11840 438084 11892
rect 472440 11908 472492 11960
rect 470692 11840 470744 11892
rect 471428 11840 471480 11892
rect 426440 11772 426492 11824
rect 485044 11908 485096 11960
rect 503536 11840 503588 11892
rect 535276 11840 535328 11892
rect 483112 11772 483164 11824
rect 484032 11772 484084 11824
rect 502248 11772 502300 11824
rect 534908 11772 534960 11824
rect 132500 11704 132552 11756
rect 416044 11704 416096 11756
rect 417976 11704 418028 11756
rect 507676 11704 507728 11756
rect 524420 11704 524472 11756
rect 524696 11704 524748 11756
rect 534724 11704 534776 11756
rect 541808 11704 541860 11756
rect 382188 11636 382240 11688
rect 496176 11636 496228 11688
rect 507860 11636 507912 11688
rect 508688 11636 508740 11688
rect 510712 11636 510764 11688
rect 511632 11636 511684 11688
rect 524604 11636 524656 11688
rect 525432 11636 525484 11688
rect 527272 11636 527324 11688
rect 527732 11636 527784 11688
rect 384948 11568 385000 11620
rect 497372 11568 497424 11620
rect 229100 11500 229152 11552
rect 238668 11500 238720 11552
rect 248420 11500 248472 11552
rect 257988 11500 258040 11552
rect 267740 11500 267792 11552
rect 277308 11500 277360 11552
rect 287060 11500 287112 11552
rect 306380 11500 306432 11552
rect 315948 11500 316000 11552
rect 325700 11500 325752 11552
rect 335268 11500 335320 11552
rect 389088 11500 389140 11552
rect 498476 11500 498528 11552
rect 391848 11432 391900 11484
rect 499672 11432 499724 11484
rect 395988 11364 396040 11416
rect 500776 11364 500828 11416
rect 400128 11296 400180 11348
rect 501972 11296 502024 11348
rect 552204 11296 552256 11348
rect 554964 11296 555016 11348
rect 407028 11228 407080 11280
rect 504272 11228 504324 11280
rect 409696 11160 409748 11212
rect 505376 11160 505428 11212
rect 413928 11092 413980 11144
rect 506572 11092 506624 11144
rect 415492 11024 415544 11076
rect 416320 11024 416372 11076
rect 424876 11024 424928 11076
rect 425060 11024 425112 11076
rect 462044 11024 462096 11076
rect 465356 11024 465408 11076
rect 466184 11024 466236 11076
rect 339408 10956 339460 11008
rect 482376 10956 482428 11008
rect 335268 10888 335320 10940
rect 481272 10888 481324 10940
rect 328368 10820 328420 10872
rect 478972 10820 479024 10872
rect 324228 10752 324280 10804
rect 477776 10752 477828 10804
rect 321468 10684 321520 10736
rect 476672 10684 476724 10736
rect 298008 10616 298060 10668
rect 305000 10616 305052 10668
rect 317328 10616 317380 10668
rect 475476 10616 475528 10668
rect 485044 10616 485096 10668
rect 510344 10616 510396 10668
rect 310428 10548 310480 10600
rect 473176 10548 473228 10600
rect 479524 10548 479576 10600
rect 505744 10548 505796 10600
rect 306288 10480 306340 10532
rect 472072 10480 472124 10532
rect 499488 10480 499540 10532
rect 534172 10480 534224 10532
rect 146852 10412 146904 10464
rect 313280 10412 313332 10464
rect 314568 10412 314620 10464
rect 474372 10412 474424 10464
rect 498108 10412 498160 10464
rect 533804 10412 533856 10464
rect 289728 10344 289780 10396
rect 302240 10344 302292 10396
rect 303528 10344 303580 10396
rect 470876 10344 470928 10396
rect 486976 10344 487028 10396
rect 530308 10344 530360 10396
rect 10416 10276 10468 10328
rect 120080 10276 120132 10328
rect 161388 10276 161440 10328
rect 330300 10276 330352 10328
rect 332416 10276 332468 10328
rect 480076 10276 480128 10328
rect 481548 10276 481600 10328
rect 528376 10276 528428 10328
rect 342168 10208 342220 10260
rect 483572 10208 483624 10260
rect 346308 10140 346360 10192
rect 484676 10140 484728 10192
rect 348976 10072 349028 10124
rect 485872 10072 485924 10124
rect 353208 10004 353260 10056
rect 486700 10004 486752 10056
rect 357348 9936 357400 9988
rect 488172 9936 488224 9988
rect 360108 9868 360160 9920
rect 489276 9868 489328 9920
rect 363328 9800 363380 9852
rect 490472 9800 490524 9852
rect 367008 9732 367060 9784
rect 491576 9732 491628 9784
rect 65984 9707 66036 9716
rect 65984 9673 65993 9707
rect 65993 9673 66027 9707
rect 66027 9673 66036 9707
rect 65984 9664 66036 9673
rect 67180 9707 67232 9716
rect 67180 9673 67189 9707
rect 67189 9673 67223 9707
rect 67223 9673 67232 9707
rect 67180 9664 67232 9673
rect 179420 9707 179472 9716
rect 179420 9673 179429 9707
rect 179429 9673 179463 9707
rect 179463 9673 179472 9707
rect 179420 9664 179472 9673
rect 182180 9707 182232 9716
rect 182180 9673 182189 9707
rect 182189 9673 182223 9707
rect 182223 9673 182232 9707
rect 182180 9664 182232 9673
rect 184848 9707 184900 9716
rect 184848 9673 184857 9707
rect 184857 9673 184891 9707
rect 184891 9673 184900 9707
rect 184848 9664 184900 9673
rect 205732 9664 205784 9716
rect 206008 9664 206060 9716
rect 208492 9664 208544 9716
rect 208860 9664 208912 9716
rect 403624 9664 403676 9716
rect 502340 9664 502392 9716
rect 530124 9664 530176 9716
rect 530676 9664 530728 9716
rect 548892 9664 548944 9716
rect 550272 9664 550324 9716
rect 126888 9596 126940 9648
rect 202788 9639 202840 9648
rect 202788 9605 202797 9639
rect 202797 9605 202831 9639
rect 202831 9605 202840 9639
rect 202788 9596 202840 9605
rect 245568 9596 245620 9648
rect 241980 9528 242032 9580
rect 451280 9528 451332 9580
rect 477040 9596 477092 9648
rect 452476 9528 452528 9580
rect 452660 9528 452712 9580
rect 486240 9528 486292 9580
rect 238392 9460 238444 9512
rect 234804 9392 234856 9444
rect 448796 9460 448848 9512
rect 451188 9460 451240 9512
rect 483940 9460 483992 9512
rect 231308 9324 231360 9376
rect 447876 9392 447928 9444
rect 458548 9392 458600 9444
rect 493140 9392 493192 9444
rect 494244 9392 494296 9444
rect 532332 9392 532384 9444
rect 227720 9256 227772 9308
rect 446772 9324 446824 9376
rect 452752 9324 452804 9376
rect 488540 9324 488592 9376
rect 495348 9324 495400 9376
rect 532976 9324 533028 9376
rect 224132 9188 224184 9240
rect 445576 9256 445628 9308
rect 446220 9256 446272 9308
rect 481640 9256 481692 9308
rect 483480 9256 483532 9308
rect 529204 9256 529256 9308
rect 445300 9188 445352 9240
rect 463240 9188 463292 9240
rect 522672 9188 522724 9240
rect 220544 9120 220596 9172
rect 444472 9120 444524 9172
rect 459744 9120 459796 9172
rect 521476 9120 521528 9172
rect 217048 9052 217100 9104
rect 443000 9052 443052 9104
rect 450176 9052 450228 9104
rect 456064 9052 456116 9104
rect 520280 9052 520332 9104
rect 150624 8984 150676 9036
rect 174176 8984 174228 9036
rect 213460 8984 213512 9036
rect 442172 8984 442224 9036
rect 452476 8984 452528 9036
rect 518992 8984 519044 9036
rect 18328 8916 18380 8968
rect 132592 8916 132644 8968
rect 153936 8916 153988 8968
rect 204904 8916 204956 8968
rect 209872 8916 209924 8968
rect 440976 8916 441028 8968
rect 518072 8916 518124 8968
rect 533252 8916 533304 8968
rect 543004 8916 543056 8968
rect 249156 8848 249208 8900
rect 453672 8848 453724 8900
rect 252652 8780 252704 8832
rect 454776 8780 454828 8832
rect 256240 8712 256292 8764
rect 455972 8712 456024 8764
rect 259828 8644 259880 8696
rect 457076 8644 457128 8696
rect 263416 8576 263468 8628
rect 458272 8576 458324 8628
rect 267004 8508 267056 8560
rect 459376 8508 459428 8560
rect 270500 8440 270552 8492
rect 460572 8440 460624 8492
rect 370412 8372 370464 8424
rect 492772 8372 492824 8424
rect 402520 8304 402572 8356
rect 503076 8304 503128 8356
rect 372804 8236 372856 8288
rect 493508 8236 493560 8288
rect 369216 8168 369268 8220
rect 492404 8168 492456 8220
rect 365720 8100 365772 8152
rect 490932 8100 490984 8152
rect 292304 8032 292356 8084
rect 459560 8032 459612 8084
rect 220820 7964 220872 8016
rect 432972 7964 433024 8016
rect 195520 7896 195572 7948
rect 431776 7896 431828 7948
rect 428372 7828 428424 7880
rect 441896 7828 441948 7880
rect 515772 7828 515824 7880
rect 177764 7760 177816 7812
rect 430672 7760 430724 7812
rect 438216 7760 438268 7812
rect 514576 7760 514628 7812
rect 174176 7692 174228 7744
rect 429476 7692 429528 7744
rect 434628 7692 434680 7744
rect 513472 7692 513524 7744
rect 167092 7624 167144 7676
rect 427176 7624 427228 7676
rect 431132 7624 431184 7676
rect 512276 7624 512328 7676
rect 513196 7624 513248 7676
rect 538772 7624 538824 7676
rect 31484 7556 31536 7608
rect 142252 7556 142304 7608
rect 143264 7556 143316 7608
rect 144184 7556 144236 7608
rect 163504 7556 163556 7608
rect 426072 7556 426124 7608
rect 427544 7556 427596 7608
rect 511172 7556 511224 7608
rect 512000 7556 512052 7608
rect 538404 7556 538456 7608
rect 376392 7488 376444 7540
rect 494704 7488 494756 7540
rect 379980 7420 380032 7472
rect 495808 7420 495860 7472
rect 383476 7352 383528 7404
rect 497004 7352 497056 7404
rect 390652 7284 390704 7336
rect 499304 7284 499356 7336
rect 394240 7216 394292 7268
rect 500408 7216 500460 7268
rect 397828 7148 397880 7200
rect 501604 7148 501656 7200
rect 401324 7080 401376 7132
rect 502708 7080 502760 7132
rect 404912 7012 404964 7064
rect 503904 7012 503956 7064
rect 412088 6944 412140 6996
rect 506204 6944 506256 6996
rect 539600 6876 539652 6928
rect 540520 6876 540572 6928
rect 77852 6808 77904 6860
rect 175372 6808 175424 6860
rect 315764 6808 315816 6860
rect 474924 6808 474976 6860
rect 70676 6740 70728 6792
rect 171232 6740 171284 6792
rect 312176 6740 312228 6792
rect 473452 6740 473504 6792
rect 63592 6672 63644 6724
rect 165712 6672 165764 6724
rect 308588 6672 308640 6724
rect 472164 6672 472216 6724
rect 56416 6604 56468 6656
rect 160100 6604 160152 6656
rect 305000 6604 305052 6656
rect 470692 6604 470744 6656
rect 476120 6604 476172 6656
rect 496912 6604 496964 6656
rect 49332 6536 49384 6588
rect 154580 6536 154632 6588
rect 301412 6536 301464 6588
rect 469404 6536 469456 6588
rect 480720 6536 480772 6588
rect 509332 6536 509384 6588
rect 44548 6468 44600 6520
rect 151820 6468 151872 6520
rect 297916 6468 297968 6520
rect 469312 6468 469364 6520
rect 471888 6468 471940 6520
rect 495624 6468 495676 6520
rect 506020 6468 506072 6520
rect 535644 6468 535696 6520
rect 40960 6400 41012 6452
rect 149152 6400 149204 6452
rect 294328 6400 294380 6452
rect 468024 6400 468076 6452
rect 477592 6400 477644 6452
rect 502524 6400 502576 6452
rect 504824 6400 504876 6452
rect 535552 6400 535604 6452
rect 37372 6332 37424 6384
rect 146300 6332 146352 6384
rect 290740 6332 290792 6384
rect 466552 6332 466604 6384
rect 473912 6332 473964 6384
rect 525892 6332 525944 6384
rect 33876 6264 33928 6316
rect 143540 6264 143592 6316
rect 287152 6264 287204 6316
rect 465172 6264 465224 6316
rect 470324 6264 470376 6316
rect 524420 6264 524472 6316
rect 8852 6196 8904 6248
rect 125692 6196 125744 6248
rect 149244 6196 149296 6248
rect 421196 6196 421248 6248
rect 423956 6196 424008 6248
rect 509516 6196 509568 6248
rect 4068 6128 4120 6180
rect 121644 6128 121696 6180
rect 144460 6128 144512 6180
rect 419724 6128 419776 6180
rect 420368 6128 420420 6180
rect 507860 6128 507912 6180
rect 519084 6128 519136 6180
rect 539600 6128 539652 6180
rect 319260 6060 319312 6112
rect 476212 6060 476264 6112
rect 322848 5992 322900 6044
rect 476304 5992 476356 6044
rect 326436 5924 326488 5976
rect 477500 5924 477552 5976
rect 330024 5856 330076 5908
rect 479064 5856 479116 5908
rect 333612 5788 333664 5840
rect 480352 5788 480404 5840
rect 337108 5720 337160 5772
rect 481824 5720 481876 5772
rect 340696 5652 340748 5704
rect 483296 5652 483348 5704
rect 344284 5584 344336 5636
rect 483112 5584 483164 5636
rect 385776 5516 385828 5568
rect 470876 5516 470928 5568
rect 90916 5448 90968 5500
rect 184756 5448 184808 5500
rect 240784 5448 240836 5500
rect 450636 5448 450688 5500
rect 469128 5448 469180 5500
rect 524512 5448 524564 5500
rect 87328 5380 87380 5432
rect 182180 5380 182232 5432
rect 237196 5380 237248 5432
rect 449532 5380 449584 5432
rect 465632 5380 465684 5432
rect 523316 5380 523368 5432
rect 83832 5312 83884 5364
rect 179420 5312 179472 5364
rect 233700 5312 233752 5364
rect 448704 5312 448756 5364
rect 462044 5312 462096 5364
rect 521936 5312 521988 5364
rect 80244 5244 80296 5296
rect 178040 5244 178092 5296
rect 230112 5244 230164 5296
rect 447324 5244 447376 5296
rect 458456 5244 458508 5296
rect 520832 5244 520884 5296
rect 76656 5176 76708 5228
rect 175280 5176 175332 5228
rect 226524 5176 226576 5228
rect 445852 5176 445904 5228
rect 454868 5176 454920 5228
rect 519636 5176 519688 5228
rect 69480 5108 69532 5160
rect 169760 5108 169812 5160
rect 222936 5108 222988 5160
rect 444472 5108 444524 5160
rect 451280 5108 451332 5160
rect 518532 5108 518584 5160
rect 73068 5040 73120 5092
rect 172520 5040 172572 5092
rect 219348 5040 219400 5092
rect 443184 5040 443236 5092
rect 447876 5040 447928 5092
rect 517704 5040 517756 5092
rect 30288 4972 30340 5024
rect 140872 4972 140924 5024
rect 215852 4972 215904 5024
rect 441712 4972 441764 5024
rect 444196 4972 444248 5024
rect 516324 4972 516376 5024
rect 26700 4904 26752 4956
rect 138112 4904 138164 4956
rect 416780 4904 416832 4956
rect 426348 4904 426400 4956
rect 510896 4904 510948 4956
rect 17224 4836 17276 4888
rect 131212 4836 131264 4888
rect 208676 4836 208728 4888
rect 440424 4836 440476 4888
rect 440608 4836 440660 4888
rect 515128 4836 515180 4888
rect 21916 4768 21968 4820
rect 135352 4768 135404 4820
rect 198004 4768 198056 4820
rect 436836 4768 436888 4820
rect 437020 4768 437072 4820
rect 513564 4768 513616 4820
rect 94504 4700 94556 4752
rect 187700 4700 187752 4752
rect 244372 4700 244424 4752
rect 451832 4700 451884 4752
rect 472716 4700 472768 4752
rect 524604 4700 524656 4752
rect 98092 4632 98144 4684
rect 190460 4632 190512 4684
rect 247960 4632 248012 4684
rect 452936 4632 452988 4684
rect 476304 4632 476356 4684
rect 525984 4632 526036 4684
rect 101588 4564 101640 4616
rect 193220 4564 193272 4616
rect 251456 4564 251508 4616
rect 454132 4564 454184 4616
rect 479892 4564 479944 4616
rect 527272 4564 527324 4616
rect 108764 4496 108816 4548
rect 198740 4496 198792 4548
rect 255044 4496 255096 4548
rect 455420 4496 455472 4548
rect 484584 4496 484636 4548
rect 528744 4496 528796 4548
rect 105176 4428 105228 4480
rect 195980 4428 196032 4480
rect 291936 4428 291988 4480
rect 466736 4428 466788 4480
rect 488172 4428 488224 4480
rect 530124 4428 530176 4480
rect 112352 4360 112404 4412
rect 201408 4360 201460 4412
rect 354956 4360 355008 4412
rect 487252 4360 487304 4412
rect 491760 4360 491812 4412
rect 531504 4360 531556 4412
rect 119436 4292 119488 4344
rect 122932 4292 122984 4344
rect 123024 4292 123076 4344
rect 125692 4292 125744 4344
rect 206008 4292 206060 4344
rect 374000 4292 374052 4344
rect 492864 4292 492916 4344
rect 508412 4292 508464 4344
rect 537024 4292 537076 4344
rect 115940 4224 115992 4276
rect 203064 4224 203116 4276
rect 429936 4224 429988 4276
rect 510712 4224 510764 4276
rect 208860 4156 208912 4208
rect 383292 4156 383344 4208
rect 383568 4156 383620 4208
rect 418068 4156 418120 4208
rect 420828 4156 420880 4208
rect 433524 4156 433576 4208
rect 512092 4156 512144 4208
rect 45468 4088 45520 4140
rect 50344 4088 50396 4140
rect 57612 4088 57664 4140
rect 60004 4088 60056 4140
rect 19524 4020 19576 4072
rect 46204 4020 46256 4072
rect 46940 4020 46992 4072
rect 139676 4088 139728 4140
rect 140688 4088 140740 4140
rect 152464 4020 152516 4072
rect 43352 3952 43404 4004
rect 150440 3952 150492 4004
rect 172980 4088 173032 4140
rect 173808 4088 173860 4140
rect 220820 4088 220872 4140
rect 360936 4088 360988 4140
rect 361488 4088 361540 4140
rect 364524 4088 364576 4140
rect 461584 4088 461636 4140
rect 500132 4088 500184 4140
rect 502340 4088 502392 4140
rect 502524 4088 502576 4140
rect 515588 4088 515640 4140
rect 516048 4088 516100 4140
rect 516784 4088 516836 4140
rect 517428 4088 517480 4140
rect 157524 4020 157576 4072
rect 207480 4020 207532 4072
rect 208308 4020 208360 4072
rect 225328 4020 225380 4072
rect 275284 4020 275336 4072
rect 350264 4020 350316 4072
rect 492956 4020 493008 4072
rect 518348 4088 518400 4140
rect 520280 4088 520332 4140
rect 521568 4088 521620 4140
rect 523868 4088 523920 4140
rect 524328 4088 524380 4140
rect 550088 4088 550140 4140
rect 550548 4088 550600 4140
rect 551928 4088 551980 4140
rect 552388 4088 552440 4140
rect 555424 4088 555476 4140
rect 557172 4088 557224 4140
rect 558644 4088 558696 4140
rect 572628 4088 572680 4140
rect 517888 4020 517940 4072
rect 523684 4020 523736 4072
rect 556988 4020 557040 4072
rect 559564 4020 559616 4072
rect 168196 3952 168248 4004
rect 225604 3952 225656 4004
rect 246764 3952 246816 4004
rect 286324 3952 286376 4004
rect 343088 3952 343140 4004
rect 451188 3952 451240 4004
rect 42156 3884 42208 3936
rect 149060 3884 149112 3936
rect 232504 3884 232556 3936
rect 257436 3884 257488 3936
rect 300124 3884 300176 3936
rect 328828 3884 328880 3936
rect 436100 3884 436152 3936
rect 439412 3884 439464 3936
rect 443552 3884 443604 3936
rect 36176 3816 36228 3868
rect 64788 3816 64840 3868
rect 66904 3816 66956 3868
rect 113180 3816 113232 3868
rect 118700 3816 118752 3868
rect 130200 3816 130252 3868
rect 131028 3816 131080 3868
rect 11244 3748 11296 3800
rect 31024 3748 31076 3800
rect 34980 3748 35032 3800
rect 139400 3748 139452 3800
rect 153200 3748 153252 3800
rect 184756 3816 184808 3868
rect 268384 3816 268436 3868
rect 331220 3816 331272 3868
rect 332416 3816 332468 3868
rect 335912 3816 335964 3868
rect 446220 3816 446272 3868
rect 478696 3952 478748 4004
rect 527364 3952 527416 4004
rect 555516 3952 555568 4004
rect 558368 3952 558420 4004
rect 471520 3884 471572 3936
rect 524696 3884 524748 3936
rect 557264 3884 557316 3936
rect 570236 4020 570288 4072
rect 573824 3952 573876 4004
rect 560116 3884 560168 3936
rect 576216 3884 576268 3936
rect 460848 3816 460900 3868
rect 514024 3816 514076 3868
rect 519728 3816 519780 3868
rect 545304 3816 545356 3868
rect 546316 3816 546368 3868
rect 558736 3816 558788 3868
rect 575020 3816 575072 3868
rect 187240 3748 187292 3800
rect 261484 3748 261536 3800
rect 314476 3748 314528 3800
rect 435364 3748 435416 3800
rect 452660 3748 452712 3800
rect 464436 3748 464488 3800
rect 523224 3748 523276 3800
rect 559748 3748 559800 3800
rect 577412 3748 577464 3800
rect 2872 3680 2924 3732
rect 10324 3680 10376 3732
rect 14832 3680 14884 3732
rect 28264 3680 28316 3732
rect 29092 3680 29144 3732
rect 45468 3680 45520 3732
rect 120632 3680 120684 3732
rect 121368 3680 121420 3732
rect 121828 3680 121880 3732
rect 122748 3680 122800 3732
rect 124220 3680 124272 3732
rect 125416 3680 125468 3732
rect 144920 3680 144972 3732
rect 176476 3680 176528 3732
rect 250444 3680 250496 3732
rect 264612 3680 264664 3732
rect 318064 3680 318116 3732
rect 321652 3680 321704 3732
rect 445300 3680 445352 3732
rect 457260 3680 457312 3732
rect 10048 3612 10100 3664
rect 25504 3612 25556 3664
rect 27896 3612 27948 3664
rect 133236 3612 133288 3664
rect 136640 3612 136692 3664
rect 137284 3612 137336 3664
rect 169392 3612 169444 3664
rect 243544 3612 243596 3664
rect 250352 3612 250404 3664
rect 304264 3612 304316 3664
rect 307392 3612 307444 3664
rect 6460 3544 6512 3596
rect 113456 3544 113508 3596
rect 113548 3544 113600 3596
rect 114468 3544 114520 3596
rect 114744 3544 114796 3596
rect 115848 3544 115900 3596
rect 116032 3544 116084 3596
rect 117964 3544 118016 3596
rect 118240 3544 118292 3596
rect 173164 3544 173216 3596
rect 180156 3544 180208 3596
rect 182180 3544 182232 3596
rect 182640 3544 182692 3596
rect 257344 3544 257396 3596
rect 268108 3544 268160 3596
rect 292304 3544 292356 3596
rect 295524 3544 295576 3596
rect 296628 3544 296680 3596
rect 296720 3544 296772 3596
rect 298008 3544 298060 3596
rect 302608 3544 302660 3596
rect 303528 3544 303580 3596
rect 433984 3612 434036 3664
rect 443000 3612 443052 3664
rect 1676 3476 1728 3528
rect 10416 3476 10468 3528
rect 24308 3476 24360 3528
rect 129832 3476 129884 3528
rect 572 3408 624 3460
rect 9128 3408 9180 3460
rect 23112 3408 23164 3460
rect 135444 3476 135496 3528
rect 145012 3476 145064 3528
rect 152740 3476 152792 3528
rect 140780 3408 140832 3460
rect 7656 3340 7708 3392
rect 11704 3340 11756 3392
rect 32680 3340 32732 3392
rect 45744 3340 45796 3392
rect 46848 3340 46900 3392
rect 51632 3340 51684 3392
rect 52368 3340 52420 3392
rect 52828 3340 52880 3392
rect 53748 3340 53800 3392
rect 54024 3340 54076 3392
rect 156604 3340 156656 3392
rect 162308 3476 162360 3528
rect 239404 3476 239456 3528
rect 239588 3476 239640 3528
rect 240048 3476 240100 3528
rect 258632 3476 258684 3528
rect 259368 3476 259420 3528
rect 265808 3476 265860 3528
rect 266268 3476 266320 3528
rect 271696 3476 271748 3528
rect 406108 3476 406160 3528
rect 407028 3476 407080 3528
rect 407304 3476 407356 3528
rect 408408 3476 408460 3528
rect 408500 3476 408552 3528
rect 409788 3476 409840 3528
rect 413284 3476 413336 3528
rect 413928 3476 413980 3528
rect 415676 3476 415728 3528
rect 416688 3476 416740 3528
rect 416872 3476 416924 3528
rect 417976 3476 418028 3528
rect 421380 3476 421432 3528
rect 422760 3476 422812 3528
rect 423588 3476 423640 3528
rect 426440 3476 426492 3528
rect 426532 3476 426584 3528
rect 439320 3544 439372 3596
rect 446588 3544 446640 3596
rect 447784 3544 447836 3596
rect 520556 3680 520608 3732
rect 544108 3680 544160 3732
rect 545028 3680 545080 3732
rect 558552 3680 558604 3732
rect 560208 3680 560260 3732
rect 578608 3680 578660 3732
rect 518164 3612 518216 3664
rect 556896 3612 556948 3664
rect 560760 3612 560812 3664
rect 561588 3612 561640 3664
rect 582196 3612 582248 3664
rect 473360 3544 473412 3596
rect 473452 3544 473504 3596
rect 516232 3544 516284 3596
rect 526260 3544 526312 3596
rect 533252 3544 533304 3596
rect 536932 3544 536984 3596
rect 544384 3544 544436 3596
rect 556712 3544 556764 3596
rect 561956 3544 562008 3596
rect 563704 3544 563756 3596
rect 583392 3544 583444 3596
rect 433432 3476 433484 3528
rect 435824 3476 435876 3528
rect 501236 3476 501288 3528
rect 502248 3476 502300 3528
rect 502432 3476 502484 3528
rect 503536 3476 503588 3528
rect 507216 3476 507268 3528
rect 507768 3476 507820 3528
rect 509608 3476 509660 3528
rect 510528 3476 510580 3528
rect 525064 3476 525116 3528
rect 526352 3476 526404 3528
rect 170588 3340 170640 3392
rect 16028 3272 16080 3324
rect 50528 3272 50580 3324
rect 20720 3204 20772 3256
rect 58808 3272 58860 3324
rect 59268 3272 59320 3324
rect 60004 3272 60056 3324
rect 60648 3272 60700 3324
rect 61200 3272 61252 3324
rect 159364 3272 159416 3324
rect 188436 3272 188488 3324
rect 188988 3272 189040 3324
rect 189632 3340 189684 3392
rect 190368 3340 190420 3392
rect 190828 3340 190880 3392
rect 191748 3340 191800 3392
rect 194416 3340 194468 3392
rect 195520 3272 195572 3324
rect 246304 3408 246356 3460
rect 214564 3340 214616 3392
rect 218152 3340 218204 3392
rect 219256 3340 219308 3392
rect 232504 3340 232556 3392
rect 233148 3340 233200 3392
rect 275284 3340 275336 3392
rect 432328 3408 432380 3460
rect 509884 3408 509936 3460
rect 510804 3408 510856 3460
rect 520924 3408 520976 3460
rect 522672 3408 522724 3460
rect 527456 3408 527508 3460
rect 528468 3408 528520 3460
rect 277676 3340 277728 3392
rect 278688 3340 278740 3392
rect 284760 3340 284812 3392
rect 285588 3340 285640 3392
rect 300308 3340 300360 3392
rect 309784 3340 309836 3392
rect 310428 3340 310480 3392
rect 310980 3340 311032 3392
rect 311808 3340 311860 3392
rect 313372 3340 313424 3392
rect 314568 3340 314620 3392
rect 318064 3340 318116 3392
rect 318708 3340 318760 3392
rect 320456 3340 320508 3392
rect 321468 3340 321520 3392
rect 334716 3340 334768 3392
rect 335268 3340 335320 3392
rect 338304 3340 338356 3392
rect 339408 3340 339460 3392
rect 339500 3340 339552 3392
rect 340788 3340 340840 3392
rect 345480 3340 345532 3392
rect 346308 3340 346360 3392
rect 347872 3340 347924 3392
rect 349068 3340 349120 3392
rect 351368 3340 351420 3392
rect 351828 3340 351880 3392
rect 352564 3340 352616 3392
rect 353208 3340 353260 3392
rect 353760 3340 353812 3392
rect 354588 3340 354640 3392
rect 356152 3340 356204 3392
rect 357348 3340 357400 3392
rect 452752 3340 452804 3392
rect 453672 3340 453724 3392
rect 457444 3340 457496 3392
rect 467932 3340 467984 3392
rect 469036 3340 469088 3392
rect 475108 3340 475160 3392
rect 476028 3340 476080 3392
rect 477500 3340 477552 3392
rect 478788 3340 478840 3392
rect 481088 3340 481140 3392
rect 481548 3340 481600 3392
rect 482284 3340 482336 3392
rect 482928 3340 482980 3392
rect 485780 3340 485832 3392
rect 487068 3340 487120 3392
rect 489368 3340 489420 3392
rect 489828 3340 489880 3392
rect 490564 3340 490616 3392
rect 491208 3340 491260 3392
rect 498936 3340 498988 3392
rect 499488 3340 499540 3392
rect 511264 3340 511316 3392
rect 514392 3340 514444 3392
rect 522304 3340 522356 3392
rect 282460 3272 282512 3324
rect 364984 3272 365036 3324
rect 377588 3272 377640 3324
rect 378048 3272 378100 3324
rect 381176 3272 381228 3324
rect 382188 3272 382240 3324
rect 382372 3272 382424 3324
rect 383292 3272 383344 3324
rect 471888 3272 471940 3324
rect 521476 3272 521528 3324
rect 524972 3272 525024 3324
rect 528652 3476 528704 3528
rect 529848 3476 529900 3528
rect 533436 3476 533488 3528
rect 533988 3476 534040 3528
rect 534540 3476 534592 3528
rect 535368 3476 535420 3528
rect 543924 3476 543976 3528
rect 563060 3476 563112 3528
rect 564348 3476 564400 3528
rect 542912 3408 542964 3460
rect 543648 3408 543700 3460
rect 561496 3408 561548 3460
rect 581000 3476 581052 3528
rect 529848 3340 529900 3392
rect 539324 3340 539376 3392
rect 545764 3340 545816 3392
rect 546500 3340 546552 3392
rect 547696 3340 547748 3392
rect 560024 3340 560076 3392
rect 579804 3408 579856 3460
rect 571432 3340 571484 3392
rect 534724 3272 534776 3324
rect 535736 3272 535788 3324
rect 536748 3272 536800 3324
rect 557448 3272 557500 3324
rect 569040 3272 569092 3324
rect 68284 3204 68336 3256
rect 162124 3204 162176 3256
rect 181352 3204 181404 3256
rect 357348 3204 357400 3256
rect 387064 3204 387116 3256
rect 387708 3204 387760 3256
rect 388260 3204 388312 3256
rect 389088 3204 389140 3256
rect 389456 3204 389508 3256
rect 390468 3204 390520 3256
rect 476120 3204 476172 3256
rect 541716 3204 541768 3256
rect 548064 3204 548116 3256
rect 557356 3204 557408 3256
rect 567844 3204 567896 3256
rect 5264 3136 5316 3188
rect 68100 3136 68152 3188
rect 81440 3136 81492 3188
rect 82728 3136 82780 3188
rect 39764 3068 39816 3120
rect 53104 3068 53156 3120
rect 55220 3068 55272 3120
rect 56508 3068 56560 3120
rect 61384 3068 61436 3120
rect 79048 3068 79100 3120
rect 82084 3068 82136 3120
rect 163412 3136 163464 3188
rect 327632 3136 327684 3188
rect 328368 3136 328420 3188
rect 371608 3136 371660 3188
rect 458548 3136 458600 3188
rect 556068 3136 556120 3188
rect 566740 3136 566792 3188
rect 57244 3000 57296 3052
rect 62396 2932 62448 2984
rect 63408 2932 63460 2984
rect 71872 2932 71924 2984
rect 75184 2932 75236 2984
rect 75460 3000 75512 3052
rect 84936 3068 84988 3120
rect 85488 3068 85540 3120
rect 88524 3068 88576 3120
rect 89628 3068 89680 3120
rect 82636 3000 82688 3052
rect 164884 3068 164936 3120
rect 193220 3068 193272 3120
rect 194508 3068 194560 3120
rect 303804 3068 303856 3120
rect 385776 3068 385828 3120
rect 395436 3068 395488 3120
rect 395988 3068 396040 3120
rect 396632 3068 396684 3120
rect 397368 3068 397420 3120
rect 399024 3068 399076 3120
rect 400128 3068 400180 3120
rect 400220 3068 400272 3120
rect 403624 3068 403676 3120
rect 403716 3068 403768 3120
rect 477592 3068 477644 3120
rect 555976 3068 556028 3120
rect 565544 3068 565596 3120
rect 86132 2932 86184 2984
rect 166264 3000 166316 3052
rect 378784 3000 378836 3052
rect 385868 3000 385920 3052
rect 410524 3000 410576 3052
rect 414480 3000 414532 3052
rect 421564 3000 421616 3052
rect 480720 3000 480772 3052
rect 558828 3000 558880 3052
rect 93308 2932 93360 2984
rect 169116 2932 169168 2984
rect 393044 2932 393096 2984
rect 464252 2932 464304 2984
rect 466828 2932 466880 2984
rect 467748 2932 467800 2984
rect 89720 2796 89772 2848
rect 95424 2796 95476 2848
rect 95700 2864 95752 2916
rect 96528 2864 96580 2916
rect 96896 2864 96948 2916
rect 102692 2864 102744 2916
rect 102784 2864 102836 2916
rect 103428 2864 103480 2916
rect 103980 2864 104032 2916
rect 105544 2864 105596 2916
rect 106372 2864 106424 2916
rect 107568 2864 107620 2916
rect 107660 2864 107712 2916
rect 100484 2796 100536 2848
rect 111156 2864 111208 2916
rect 111708 2864 111760 2916
rect 169024 2864 169076 2916
rect 253848 2864 253900 2916
rect 292580 2864 292632 2916
rect 410892 2864 410944 2916
rect 479524 2864 479576 2916
rect 540520 2864 540572 2916
rect 547328 2864 547380 2916
rect 171600 2796 171652 2848
rect 261024 2796 261076 2848
rect 311164 2796 311216 2848
rect 346676 2796 346728 2848
rect 425060 2796 425112 2848
rect 425152 2796 425204 2848
rect 485044 2796 485096 2848
rect 550824 2796 550876 2848
rect 553400 2796 553452 2848
rect 274088 2728 274140 2780
rect 461032 2728 461084 2780
rect 551192 2728 551244 2780
rect 553584 2728 553636 2780
rect 269304 2660 269356 2712
rect 459836 2660 459888 2712
rect 262220 2592 262272 2644
rect 456892 2592 456944 2644
rect 243176 2524 243228 2576
rect 451556 2524 451608 2576
rect 183744 2456 183796 2508
rect 184848 2456 184900 2508
rect 236000 2456 236052 2508
rect 448980 2499 449032 2508
rect 228916 2388 228968 2440
rect 415400 2388 415452 2440
rect 424968 2388 425020 2440
rect 434720 2388 434772 2440
rect 448980 2465 448989 2499
rect 448989 2465 449023 2499
rect 449023 2465 449032 2499
rect 448980 2456 449032 2465
rect 449072 2388 449124 2440
rect 214656 2320 214708 2372
rect 342904 2320 342956 2372
rect 347688 2320 347740 2372
rect 441988 2320 442040 2372
rect 442080 2320 442132 2372
rect 447232 2320 447284 2372
rect 200396 2252 200448 2304
rect 347412 2252 347464 2304
rect 437572 2252 437624 2304
rect 199200 2184 199252 2236
rect 347688 2184 347740 2236
rect 437756 2184 437808 2236
rect 192024 2116 192076 2168
rect 434904 2116 434956 2168
rect 133788 2048 133840 2100
rect 381544 2048 381596 2100
rect 386328 2048 386380 2100
rect 415492 2048 415544 2100
rect 450176 2048 450228 2100
rect 276480 1980 276532 2032
rect 462412 1980 462464 2032
rect 281264 1912 281316 1964
rect 463884 1912 463936 1964
rect 288348 1844 288400 1896
rect 465356 1844 465408 1896
rect 299112 1776 299164 1828
rect 385960 1776 386012 1828
rect 386328 1776 386380 1828
rect 469496 1776 469548 1828
rect 292580 1708 292632 1760
rect 454224 1708 454276 1760
rect 311164 1640 311216 1692
rect 456984 1640 457036 1692
rect 362132 1572 362184 1624
rect 490104 1572 490156 1624
rect 165896 960 165948 1012
rect 65892 552 65944 604
rect 65984 552 66036 604
rect 126612 595 126664 604
rect 126612 561 126621 595
rect 126621 561 126655 595
rect 126655 561 126664 595
rect 126612 552 126664 561
rect 161112 552 161164 604
rect 161388 552 161440 604
rect 178960 552 179012 604
rect 179328 552 179380 604
rect 202696 552 202748 604
rect 445392 552 445444 604
rect 445668 552 445720 604
rect 496544 552 496596 604
rect 496728 552 496780 604
rect 554780 552 554832 604
rect 554964 552 555016 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700330 8156 703520
rect 24320 700330 24348 703520
rect 40512 700398 40540 703520
rect 72988 700466 73016 703520
rect 89180 700466 89208 703520
rect 51724 700460 51776 700466
rect 51724 700402 51776 700408
rect 72976 700460 73028 700466
rect 72976 700402 73028 700408
rect 89168 700460 89220 700466
rect 89168 700402 89220 700408
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 8944 700324 8996 700330
rect 8944 700266 8996 700272
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3528 681766 3556 682207
rect 3516 681760 3568 681766
rect 3516 681702 3568 681708
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 3422 624880 3478 624889
rect 3422 624815 3478 624824
rect 3330 610464 3386 610473
rect 3330 610399 3386 610408
rect 3344 610026 3372 610399
rect 3332 610020 3384 610026
rect 3332 609962 3384 609968
rect 3146 553072 3202 553081
rect 3146 553007 3202 553016
rect 3160 552090 3188 553007
rect 3148 552084 3200 552090
rect 3148 552026 3200 552032
rect 2870 509960 2926 509969
rect 2870 509895 2926 509904
rect 2884 509318 2912 509895
rect 2872 509312 2924 509318
rect 2872 509254 2924 509260
rect 3436 485110 3464 624815
rect 3514 596048 3570 596057
rect 3514 595983 3570 595992
rect 3528 594862 3556 595983
rect 3516 594856 3568 594862
rect 3516 594798 3568 594804
rect 3514 567352 3570 567361
rect 3514 567287 3570 567296
rect 3528 567254 3556 567287
rect 3516 567248 3568 567254
rect 3516 567190 3568 567196
rect 3514 538656 3570 538665
rect 3514 538591 3570 538600
rect 3528 538286 3556 538591
rect 3516 538280 3568 538286
rect 3516 538222 3568 538228
rect 3514 495544 3570 495553
rect 3514 495479 3516 495488
rect 3568 495479 3570 495488
rect 3516 495450 3568 495456
rect 3424 485104 3476 485110
rect 3424 485046 3476 485052
rect 3146 481128 3202 481137
rect 3146 481063 3202 481072
rect 3160 480282 3188 481063
rect 3148 480276 3200 480282
rect 3148 480218 3200 480224
rect 3422 452432 3478 452441
rect 3422 452367 3478 452376
rect 3436 451314 3464 452367
rect 3424 451308 3476 451314
rect 3424 451250 3476 451256
rect 3422 438016 3478 438025
rect 3422 437951 3478 437960
rect 2778 380624 2834 380633
rect 2778 380559 2834 380568
rect 2792 366217 2820 380559
rect 2778 366208 2834 366217
rect 2778 366143 2834 366152
rect 2792 323105 2820 366143
rect 3146 337512 3202 337521
rect 3146 337447 3202 337456
rect 3160 336802 3188 337447
rect 3148 336796 3200 336802
rect 3148 336738 3200 336744
rect 2778 323096 2834 323105
rect 2778 323031 2834 323040
rect 2792 316742 2820 323031
rect 2780 316736 2832 316742
rect 2780 316678 2832 316684
rect 2778 309088 2834 309097
rect 2778 309023 2834 309032
rect 2792 308825 2820 309023
rect 2778 308816 2834 308825
rect 2778 308751 2834 308760
rect 2792 280129 2820 308751
rect 2778 280120 2834 280129
rect 2778 280055 2834 280064
rect 2792 265713 2820 280055
rect 2778 265704 2834 265713
rect 2778 265639 2834 265648
rect 2792 237017 2820 265639
rect 2778 237008 2834 237017
rect 2778 236943 2834 236952
rect 2792 222601 2820 236943
rect 2778 222592 2834 222601
rect 2778 222527 2834 222536
rect 2792 193905 2820 222527
rect 2778 193896 2834 193905
rect 2778 193831 2834 193840
rect 2792 179489 2820 193831
rect 2778 179480 2834 179489
rect 2778 179415 2834 179424
rect 2792 150793 2820 179415
rect 2778 150784 2834 150793
rect 2778 150719 2834 150728
rect 2792 136377 2820 150719
rect 2778 136368 2834 136377
rect 2778 136303 2834 136312
rect 2792 107681 2820 136303
rect 2778 107672 2834 107681
rect 2778 107607 2834 107616
rect 2792 93265 2820 107607
rect 2778 93256 2834 93265
rect 2778 93191 2834 93200
rect 2792 64569 2820 93191
rect 2778 64560 2834 64569
rect 2778 64495 2834 64504
rect 2792 50153 2820 64495
rect 2778 50144 2834 50153
rect 2778 50079 2834 50088
rect 2792 21457 2820 50079
rect 3436 27606 3464 437951
rect 3514 423736 3570 423745
rect 3514 423671 3516 423680
rect 3568 423671 3570 423680
rect 3516 423642 3568 423648
rect 4802 395040 4858 395049
rect 4802 394975 4858 394984
rect 3516 316736 3568 316742
rect 3516 316678 3568 316684
rect 3528 309097 3556 316678
rect 3514 309088 3570 309097
rect 3514 309023 3570 309032
rect 3606 294400 3662 294409
rect 3606 294335 3662 294344
rect 3620 224262 3648 294335
rect 3608 224256 3660 224262
rect 3608 224198 3660 224204
rect 3516 223644 3568 223650
rect 3516 223586 3568 223592
rect 3528 35873 3556 223586
rect 4816 173777 4844 394975
rect 6184 336796 6236 336802
rect 6184 336738 6236 336744
rect 4802 173768 4858 173777
rect 4802 173703 4858 173712
rect 6196 65521 6224 336738
rect 8956 125594 8984 700266
rect 51736 691422 51764 700402
rect 137848 697610 137876 703520
rect 154132 700534 154160 703520
rect 202800 700534 202828 703520
rect 138664 700528 138716 700534
rect 138664 700470 138716 700476
rect 154120 700528 154172 700534
rect 154120 700470 154172 700476
rect 202788 700528 202840 700534
rect 202788 700470 202840 700476
rect 136640 697604 136692 697610
rect 136640 697546 136692 697552
rect 137836 697604 137888 697610
rect 137836 697546 137888 697552
rect 48504 691416 48556 691422
rect 48504 691358 48556 691364
rect 51724 691416 51776 691422
rect 51724 691358 51776 691364
rect 48516 685234 48544 691358
rect 46940 685228 46992 685234
rect 46940 685170 46992 685176
rect 48504 685228 48556 685234
rect 48504 685170 48556 685176
rect 46952 680406 46980 685170
rect 46940 680400 46992 680406
rect 46940 680342 46992 680348
rect 42064 680264 42116 680270
rect 42064 680206 42116 680212
rect 42076 672110 42104 680206
rect 136652 674830 136680 697546
rect 133880 674824 133932 674830
rect 133880 674766 133932 674772
rect 136640 674824 136692 674830
rect 136640 674766 136692 674772
rect 40040 672104 40092 672110
rect 40040 672046 40092 672052
rect 42064 672104 42116 672110
rect 42064 672046 42116 672052
rect 40052 666602 40080 672046
rect 133892 670750 133920 674766
rect 131764 670744 131816 670750
rect 131764 670686 131816 670692
rect 133880 670744 133932 670750
rect 133880 670686 133932 670692
rect 40040 666596 40092 666602
rect 40040 666538 40092 666544
rect 37924 666528 37976 666534
rect 37924 666470 37976 666476
rect 10324 652792 10376 652798
rect 10324 652734 10376 652740
rect 9036 594856 9088 594862
rect 9036 594798 9088 594804
rect 9048 128314 9076 594798
rect 9128 567248 9180 567254
rect 9128 567190 9180 567196
rect 9140 444378 9168 567190
rect 9128 444372 9180 444378
rect 9128 444314 9180 444320
rect 9128 225616 9180 225622
rect 9128 225558 9180 225564
rect 9036 128308 9088 128314
rect 9036 128250 9088 128256
rect 8944 125588 8996 125594
rect 8944 125530 8996 125536
rect 6182 65512 6238 65521
rect 6182 65447 6238 65456
rect 3514 35864 3570 35873
rect 3514 35799 3570 35808
rect 3424 27600 3476 27606
rect 3424 27542 3476 27548
rect 2778 21448 2834 21457
rect 2778 21383 2834 21392
rect 2792 7177 2820 21383
rect 2778 7168 2834 7177
rect 2778 7103 2834 7112
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3470
rect 2884 480 2912 3674
rect 4080 480 4108 6122
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5276 480 5304 3130
rect 6472 480 6500 3538
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 7668 480 7696 3334
rect 8864 480 8892 6190
rect 9140 3466 9168 225558
rect 10336 126954 10364 652734
rect 37936 650078 37964 666470
rect 36544 650072 36596 650078
rect 36544 650014 36596 650020
rect 37924 650072 37976 650078
rect 37924 650014 37976 650020
rect 36556 634846 36584 650014
rect 131776 648378 131804 670686
rect 129004 648372 129056 648378
rect 129004 648314 129056 648320
rect 131764 648372 131816 648378
rect 131764 648314 131816 648320
rect 129016 640354 129044 648314
rect 126244 640348 126296 640354
rect 126244 640290 126296 640296
rect 129004 640348 129056 640354
rect 129004 640290 129056 640296
rect 35256 634840 35308 634846
rect 35256 634782 35308 634788
rect 36544 634840 36596 634846
rect 36544 634782 36596 634788
rect 35268 629542 35296 634782
rect 126256 629950 126284 640290
rect 116584 629944 116636 629950
rect 116584 629886 116636 629892
rect 126244 629944 126296 629950
rect 126244 629886 126296 629892
rect 33784 629536 33836 629542
rect 33784 629478 33836 629484
rect 35256 629536 35308 629542
rect 35256 629478 35308 629484
rect 23388 619676 23440 619682
rect 23388 619618 23440 619624
rect 13084 610020 13136 610026
rect 13084 609962 13136 609968
rect 10416 538280 10468 538286
rect 10416 538222 10468 538228
rect 10428 129266 10456 538222
rect 13096 494766 13124 609962
rect 23296 571804 23348 571810
rect 23296 571746 23348 571752
rect 21364 532500 21416 532506
rect 21364 532442 21416 532448
rect 14556 509312 14608 509318
rect 14556 509254 14608 509260
rect 13084 494760 13136 494766
rect 13084 494702 13136 494708
rect 14464 480276 14516 480282
rect 14464 480218 14516 480224
rect 11704 451308 11756 451314
rect 11704 451250 11756 451256
rect 11716 276010 11744 451250
rect 12532 444372 12584 444378
rect 12532 444314 12584 444320
rect 12544 443601 12572 444314
rect 12530 443592 12586 443601
rect 12530 443527 12586 443536
rect 13084 423700 13136 423706
rect 13084 423642 13136 423648
rect 11704 276004 11756 276010
rect 11704 275946 11756 275952
rect 13096 227050 13124 423642
rect 13084 227044 13136 227050
rect 13084 226986 13136 226992
rect 14476 220114 14504 480218
rect 14568 315314 14596 509254
rect 21376 492561 21404 532442
rect 22100 531140 22152 531146
rect 22100 531082 22152 531088
rect 22112 528836 22140 531082
rect 23308 528850 23336 571746
rect 23400 531146 23428 619618
rect 33796 618594 33824 629478
rect 116596 622441 116624 629886
rect 116582 622432 116638 622441
rect 116582 622367 116638 622376
rect 84108 619676 84160 619682
rect 84108 619618 84160 619624
rect 29736 618588 29788 618594
rect 29736 618530 29788 618536
rect 33784 618588 33836 618594
rect 33784 618530 33836 618536
rect 28630 611552 28686 611561
rect 28686 611510 29132 611538
rect 28630 611487 28686 611496
rect 27710 609648 27766 609657
rect 29104 609634 29132 611510
rect 29748 610722 29776 618530
rect 84120 617658 84148 619618
rect 84120 617630 84180 617658
rect 29748 610694 30144 610722
rect 29104 609606 29408 609634
rect 27710 609583 27766 609592
rect 27526 608968 27582 608977
rect 27526 608903 27582 608912
rect 27158 607200 27214 607209
rect 27158 607135 27214 607144
rect 27066 601216 27122 601225
rect 27066 601151 27122 601160
rect 26974 598768 27030 598777
rect 26974 598703 27030 598712
rect 26148 597984 26200 597990
rect 26148 597926 26200 597932
rect 24950 594008 25006 594017
rect 24950 593943 25006 593952
rect 24124 586084 24176 586090
rect 24124 586026 24176 586032
rect 24136 532506 24164 586026
rect 24858 572928 24914 572937
rect 24858 572863 24914 572872
rect 24766 572384 24822 572393
rect 24766 572319 24822 572328
rect 24674 571840 24730 571849
rect 24674 571775 24676 571784
rect 24728 571775 24730 571784
rect 24676 571746 24728 571752
rect 24124 532500 24176 532506
rect 24124 532442 24176 532448
rect 23388 531140 23440 531146
rect 23388 531082 23440 531088
rect 23138 528822 23336 528850
rect 24780 528714 24808 572319
rect 24872 528850 24900 572863
rect 24964 532234 24992 593943
rect 26054 592784 26110 592793
rect 26054 592719 26110 592728
rect 25870 591560 25926 591569
rect 25870 591495 25926 591504
rect 25778 588024 25834 588033
rect 25778 587959 25834 587968
rect 25686 585576 25742 585585
rect 25686 585511 25742 585520
rect 25502 584352 25558 584361
rect 25502 584287 25558 584296
rect 25318 583128 25374 583137
rect 25318 583063 25374 583072
rect 25226 582040 25282 582049
rect 25226 581975 25282 581984
rect 25134 580816 25190 580825
rect 25134 580751 25190 580760
rect 25042 579592 25098 579601
rect 25042 579527 25098 579536
rect 25056 533866 25084 579527
rect 25044 533860 25096 533866
rect 25044 533802 25096 533808
rect 25148 533798 25176 580751
rect 25136 533792 25188 533798
rect 25136 533734 25188 533740
rect 25240 533730 25268 581975
rect 25228 533724 25280 533730
rect 25228 533666 25280 533672
rect 25332 533662 25360 583063
rect 25410 581360 25466 581369
rect 25410 581295 25466 581304
rect 25320 533656 25372 533662
rect 25320 533598 25372 533604
rect 24952 532228 25004 532234
rect 24952 532170 25004 532176
rect 25424 531962 25452 581295
rect 25516 532642 25544 584287
rect 25594 583808 25650 583817
rect 25594 583743 25650 583752
rect 25504 532636 25556 532642
rect 25504 532578 25556 532584
rect 25412 531956 25464 531962
rect 25412 531898 25464 531904
rect 25608 530194 25636 583743
rect 25700 532574 25728 585511
rect 25688 532568 25740 532574
rect 25688 532510 25740 532516
rect 25792 532506 25820 587959
rect 25780 532500 25832 532506
rect 25780 532442 25832 532448
rect 25884 532370 25912 591495
rect 25962 589792 26018 589801
rect 25962 589727 26018 589736
rect 25872 532364 25924 532370
rect 25872 532306 25924 532312
rect 25976 530534 26004 589727
rect 26068 532302 26096 592719
rect 26160 586090 26188 597926
rect 26790 596456 26846 596465
rect 26790 596391 26846 596400
rect 26698 592240 26754 592249
rect 26698 592175 26754 592184
rect 26148 586084 26200 586090
rect 26148 586026 26200 586032
rect 26606 585032 26662 585041
rect 26606 584967 26662 584976
rect 26514 582584 26570 582593
rect 26514 582519 26570 582528
rect 26422 578912 26478 578921
rect 26422 578847 26478 578856
rect 26146 578368 26202 578377
rect 26146 578303 26202 578312
rect 26160 533934 26188 578303
rect 26238 574152 26294 574161
rect 26238 574087 26294 574096
rect 26148 533928 26200 533934
rect 26148 533870 26200 533876
rect 26252 533390 26280 574087
rect 26330 573608 26386 573617
rect 26330 573543 26386 573552
rect 26240 533384 26292 533390
rect 26240 533326 26292 533332
rect 26056 532296 26108 532302
rect 26056 532238 26108 532244
rect 25964 530528 26016 530534
rect 25964 530470 26016 530476
rect 25596 530188 25648 530194
rect 25596 530130 25648 530136
rect 24872 528822 25346 528850
rect 26344 528836 26372 573543
rect 26436 572762 26464 578847
rect 26424 572756 26476 572762
rect 26424 572698 26476 572704
rect 26424 572620 26476 572626
rect 26424 572562 26476 572568
rect 26436 531690 26464 572562
rect 26528 532166 26556 582519
rect 26620 535634 26648 584967
rect 26608 535628 26660 535634
rect 26608 535570 26660 535576
rect 26712 535514 26740 592175
rect 26620 535486 26740 535514
rect 26804 535498 26832 596391
rect 26882 595232 26938 595241
rect 26882 595167 26938 595176
rect 26792 535492 26844 535498
rect 26516 532160 26568 532166
rect 26516 532102 26568 532108
rect 26424 531684 26476 531690
rect 26424 531626 26476 531632
rect 26620 531282 26648 535486
rect 26792 535434 26844 535440
rect 26896 535378 26924 595167
rect 26712 535350 26924 535378
rect 26608 531276 26660 531282
rect 26608 531218 26660 531224
rect 26712 531146 26740 535350
rect 26792 535288 26844 535294
rect 26988 535242 27016 598703
rect 26792 535230 26844 535236
rect 26804 531894 26832 535230
rect 26896 535214 27016 535242
rect 26792 531888 26844 531894
rect 26792 531830 26844 531836
rect 26700 531140 26752 531146
rect 26700 531082 26752 531088
rect 26896 531078 26924 535214
rect 27080 535106 27108 601151
rect 26988 535078 27108 535106
rect 26988 532030 27016 535078
rect 27068 535016 27120 535022
rect 27068 534958 27120 534964
rect 27080 533474 27108 534958
rect 27172 533594 27200 607135
rect 27434 606656 27490 606665
rect 27434 606591 27490 606600
rect 27250 605976 27306 605985
rect 27250 605911 27306 605920
rect 27160 533588 27212 533594
rect 27160 533530 27212 533536
rect 27264 533526 27292 605911
rect 27342 604208 27398 604217
rect 27342 604143 27398 604152
rect 27252 533520 27304 533526
rect 27080 533446 27200 533474
rect 27252 533462 27304 533468
rect 27068 533384 27120 533390
rect 27068 533326 27120 533332
rect 26976 532024 27028 532030
rect 26976 531966 27028 531972
rect 26884 531072 26936 531078
rect 26884 531014 26936 531020
rect 27080 528850 27108 533326
rect 27172 530262 27200 533446
rect 27356 530874 27384 604143
rect 27344 530868 27396 530874
rect 27344 530810 27396 530816
rect 27448 530738 27476 606591
rect 27436 530732 27488 530738
rect 27436 530674 27488 530680
rect 27540 530602 27568 608903
rect 27618 608424 27674 608433
rect 27618 608359 27674 608368
rect 27632 530670 27660 608359
rect 27724 533390 27752 609583
rect 28630 607336 28686 607345
rect 28686 607294 29132 607322
rect 28630 607271 28686 607280
rect 29104 605826 29132 607294
rect 28920 605798 29132 605826
rect 27802 605432 27858 605441
rect 27802 605367 27858 605376
rect 27712 533384 27764 533390
rect 27712 533326 27764 533332
rect 27816 530806 27844 605367
rect 28538 602576 28594 602585
rect 28538 602511 28594 602520
rect 27894 602032 27950 602041
rect 27894 601967 27950 601976
rect 27908 530942 27936 601967
rect 28078 601896 28134 601905
rect 28078 601831 28134 601840
rect 27986 597680 28042 597689
rect 27986 597615 28042 597624
rect 28000 531214 28028 597615
rect 27988 531208 28040 531214
rect 27988 531150 28040 531156
rect 28092 531010 28120 601831
rect 28552 599026 28580 602511
rect 28630 600264 28686 600273
rect 28686 600222 28764 600250
rect 28630 600199 28686 600208
rect 28552 598998 28672 599026
rect 28538 598904 28594 598913
rect 28538 598839 28594 598848
rect 28170 597136 28226 597145
rect 28170 597071 28226 597080
rect 28184 532098 28212 597071
rect 28552 595490 28580 598839
rect 28644 597666 28672 598998
rect 28736 597802 28764 600222
rect 28920 598466 28948 605798
rect 28908 598460 28960 598466
rect 28908 598402 28960 598408
rect 29380 598210 29408 609606
rect 30116 598210 30144 610694
rect 28920 598194 29408 598210
rect 28908 598188 29408 598194
rect 28960 598182 29408 598188
rect 29472 598182 30144 598210
rect 28908 598130 28960 598136
rect 28908 597984 28960 597990
rect 29472 597972 29500 598182
rect 28960 597944 29500 597972
rect 28908 597926 28960 597932
rect 28736 597774 30328 597802
rect 28644 597638 30236 597666
rect 28630 597136 28686 597145
rect 28686 597094 29868 597122
rect 28630 597071 28686 597080
rect 29840 596850 29868 597094
rect 29840 596822 30144 596850
rect 28552 595462 30052 595490
rect 28446 595368 28502 595377
rect 28446 595303 28502 595312
rect 28262 594144 28318 594153
rect 28262 594079 28318 594088
rect 28276 589422 28304 594079
rect 28354 592920 28410 592929
rect 28354 592855 28410 592864
rect 28264 589416 28316 589422
rect 28264 589358 28316 589364
rect 28368 588606 28396 592855
rect 28460 589286 28488 595303
rect 28908 595128 28960 595134
rect 28960 595088 29868 595116
rect 28908 595070 28960 595076
rect 28538 590472 28594 590481
rect 28538 590407 28594 590416
rect 28448 589280 28500 589286
rect 28448 589222 28500 589228
rect 28446 588704 28502 588713
rect 28552 588690 28580 590407
rect 29288 590294 29776 590322
rect 28630 590064 28686 590073
rect 29288 590050 29316 590294
rect 28686 590022 29316 590050
rect 28630 589999 28686 590008
rect 28908 589960 28960 589966
rect 28960 589908 29684 589914
rect 28908 589902 29684 589908
rect 28920 589886 29684 589902
rect 28908 589416 28960 589422
rect 28960 589364 29592 589370
rect 28908 589358 29592 589364
rect 28920 589342 29592 589358
rect 28908 589280 28960 589286
rect 28960 589228 29500 589234
rect 28908 589222 29500 589228
rect 28920 589206 29500 589222
rect 28552 588662 29316 588690
rect 28446 588639 28502 588648
rect 28356 588600 28408 588606
rect 28356 588542 28408 588548
rect 28262 588160 28318 588169
rect 28262 588095 28318 588104
rect 28172 532092 28224 532098
rect 28172 532034 28224 532040
rect 28080 531004 28132 531010
rect 28080 530946 28132 530952
rect 27896 530936 27948 530942
rect 27896 530878 27948 530884
rect 27804 530800 27856 530806
rect 27804 530742 27856 530748
rect 27620 530664 27672 530670
rect 27620 530606 27672 530612
rect 27528 530596 27580 530602
rect 27528 530538 27580 530544
rect 28276 530466 28304 588095
rect 28354 586936 28410 586945
rect 28354 586871 28410 586880
rect 28264 530460 28316 530466
rect 28264 530402 28316 530408
rect 28368 530398 28396 586871
rect 28460 532438 28488 588639
rect 28908 588600 28960 588606
rect 28960 588548 29224 588554
rect 28908 588542 29224 588548
rect 28920 588526 29224 588542
rect 28630 586936 28686 586945
rect 28686 586894 29040 586922
rect 28630 586871 28686 586880
rect 28630 585712 28686 585721
rect 28686 585670 28856 585698
rect 28630 585647 28686 585656
rect 28828 579850 28856 585670
rect 29012 582298 29040 586894
rect 28920 582270 29040 582298
rect 28920 580310 28948 582270
rect 28908 580304 28960 580310
rect 28908 580246 28960 580252
rect 28552 579822 28856 579850
rect 28448 532432 28500 532438
rect 28448 532374 28500 532380
rect 28356 530392 28408 530398
rect 28356 530334 28408 530340
rect 28552 530330 28580 579822
rect 28630 579728 28686 579737
rect 28686 579686 28856 579714
rect 28630 579663 28686 579672
rect 28630 577280 28686 577289
rect 28686 577238 28764 577266
rect 28630 577215 28686 577224
rect 28630 576736 28686 576745
rect 28630 576671 28686 576680
rect 28644 576162 28672 576671
rect 28632 576156 28684 576162
rect 28632 576098 28684 576104
rect 28630 576056 28686 576065
rect 28630 575991 28686 576000
rect 28644 575278 28672 575991
rect 28632 575272 28684 575278
rect 28632 575214 28684 575220
rect 28632 575136 28684 575142
rect 28630 575104 28632 575113
rect 28684 575104 28686 575113
rect 28630 575039 28686 575048
rect 28632 575000 28684 575006
rect 28630 574968 28632 574977
rect 28684 574968 28686 574977
rect 28630 574903 28686 574912
rect 28632 574864 28684 574870
rect 28632 574806 28684 574812
rect 28644 531826 28672 574806
rect 28736 532710 28764 577238
rect 28828 575074 28856 579686
rect 28908 576156 28960 576162
rect 29196 576144 29224 588526
rect 29288 586378 29316 588662
rect 29288 586350 29408 586378
rect 28960 576116 29224 576144
rect 28908 576098 28960 576104
rect 28908 575884 28960 575890
rect 28960 575844 29040 575872
rect 28908 575826 28960 575832
rect 28908 575136 28960 575142
rect 28908 575078 28960 575084
rect 28816 575068 28868 575074
rect 28816 575010 28868 575016
rect 28816 574796 28868 574802
rect 28816 574738 28868 574744
rect 28724 532704 28776 532710
rect 28724 532646 28776 532652
rect 28632 531820 28684 531826
rect 28632 531762 28684 531768
rect 28540 530324 28592 530330
rect 28540 530266 28592 530272
rect 27160 530256 27212 530262
rect 27160 530198 27212 530204
rect 28828 528850 28856 574738
rect 28920 529938 28948 575078
rect 29012 571334 29040 575844
rect 29380 573730 29408 586350
rect 29104 573702 29408 573730
rect 29104 572830 29132 573702
rect 29368 573504 29420 573510
rect 29368 573446 29420 573452
rect 29092 572824 29144 572830
rect 29092 572766 29144 572772
rect 29276 572756 29328 572762
rect 29276 572698 29328 572704
rect 29182 571568 29238 571577
rect 29182 571503 29238 571512
rect 29000 571328 29052 571334
rect 29000 571270 29052 571276
rect 29000 570036 29052 570042
rect 29000 569978 29052 569984
rect 29012 563394 29040 569978
rect 29092 567248 29144 567254
rect 29092 567190 29144 567196
rect 29104 565214 29132 567190
rect 29092 565208 29144 565214
rect 29092 565150 29144 565156
rect 29196 563582 29224 571503
rect 29288 567934 29316 572698
rect 29276 567928 29328 567934
rect 29276 567870 29328 567876
rect 29380 566506 29408 573446
rect 29472 567866 29500 589206
rect 29460 567860 29512 567866
rect 29460 567802 29512 567808
rect 29368 566500 29420 566506
rect 29368 566442 29420 566448
rect 29564 565146 29592 589342
rect 29656 570042 29684 589886
rect 29644 570036 29696 570042
rect 29644 569978 29696 569984
rect 29552 565140 29604 565146
rect 29552 565082 29604 565088
rect 29184 563576 29236 563582
rect 29184 563518 29236 563524
rect 29012 563366 29500 563394
rect 29472 562986 29500 563366
rect 29472 562958 29592 562986
rect 29564 551342 29592 562958
rect 29552 551336 29604 551342
rect 29552 551278 29604 551284
rect 29748 533594 29776 590294
rect 29840 560998 29868 595088
rect 30024 573442 30052 595462
rect 30012 573436 30064 573442
rect 30012 573378 30064 573384
rect 30116 572830 30144 596822
rect 30104 572824 30156 572830
rect 30104 572766 30156 572772
rect 29920 572688 29972 572694
rect 29920 572630 29972 572636
rect 29932 563718 29960 572630
rect 30208 569294 30236 597638
rect 30300 570654 30328 597774
rect 56120 571526 56456 571554
rect 112240 571526 112576 571554
rect 31852 571328 31904 571334
rect 31852 571270 31904 571276
rect 30288 570648 30340 570654
rect 30288 570590 30340 570596
rect 30288 570512 30340 570518
rect 30288 570454 30340 570460
rect 30196 569288 30248 569294
rect 30196 569230 30248 569236
rect 29920 563712 29972 563718
rect 29920 563654 29972 563660
rect 29920 563576 29972 563582
rect 29920 563518 29972 563524
rect 29828 560992 29880 560998
rect 29828 560934 29880 560940
rect 29736 533588 29788 533594
rect 29736 533530 29788 533536
rect 29932 531282 29960 563518
rect 30300 562358 30328 570454
rect 31760 570172 31812 570178
rect 31760 570114 31812 570120
rect 30288 562352 30340 562358
rect 30288 562294 30340 562300
rect 29920 531276 29972 531282
rect 29920 531218 29972 531224
rect 30656 531276 30708 531282
rect 30656 531218 30708 531224
rect 28920 529910 29224 529938
rect 27080 528822 27462 528850
rect 28566 528822 28856 528850
rect 29196 528850 29224 529910
rect 29196 528822 29670 528850
rect 30668 528836 30696 531218
rect 31772 528836 31800 570114
rect 24242 528686 24808 528714
rect 31864 528714 31892 571270
rect 56428 569226 56456 571526
rect 74540 570648 74592 570654
rect 74540 570590 74592 570596
rect 56416 569220 56468 569226
rect 56416 569162 56468 569168
rect 56600 567928 56652 567934
rect 56600 567870 56652 567876
rect 49700 565208 49752 565214
rect 49700 565150 49752 565156
rect 34980 533928 35032 533934
rect 34980 533870 35032 533876
rect 33876 532704 33928 532710
rect 33876 532646 33928 532652
rect 33888 528836 33916 532646
rect 34992 528836 35020 533870
rect 37188 533860 37240 533866
rect 37188 533802 37240 533808
rect 36084 531888 36136 531894
rect 36084 531830 36136 531836
rect 36096 528836 36124 531830
rect 37200 528836 37228 533802
rect 39304 533792 39356 533798
rect 39304 533734 39356 533740
rect 38200 531820 38252 531826
rect 38200 531762 38252 531768
rect 38212 528836 38240 531762
rect 39316 528836 39344 533734
rect 41420 533724 41472 533730
rect 41420 533666 41472 533672
rect 40408 531956 40460 531962
rect 40408 531898 40460 531904
rect 40420 528836 40448 531898
rect 41432 528836 41460 533666
rect 43628 533656 43680 533662
rect 43628 533598 43680 533604
rect 42524 532704 42576 532710
rect 42524 532646 42576 532652
rect 42536 528836 42564 532646
rect 43640 528836 43668 533598
rect 45744 532636 45796 532642
rect 45744 532578 45796 532584
rect 44732 530188 44784 530194
rect 44732 530130 44784 530136
rect 44744 528836 44772 530130
rect 45756 528836 45784 532578
rect 47952 532568 48004 532574
rect 47952 532510 48004 532516
rect 46848 530256 46900 530262
rect 46848 530198 46900 530204
rect 46860 528836 46888 530198
rect 47964 528836 47992 532510
rect 48964 530324 49016 530330
rect 48964 530266 49016 530272
rect 48976 528836 49004 530266
rect 49712 528850 49740 565150
rect 56508 533588 56560 533594
rect 56508 533530 56560 533536
rect 52276 532500 52328 532506
rect 52276 532442 52328 532448
rect 51172 530392 51224 530398
rect 51172 530334 51224 530340
rect 49712 528822 50094 528850
rect 51184 528836 51212 530334
rect 52288 528836 52316 532442
rect 54392 532432 54444 532438
rect 54392 532374 54444 532380
rect 53288 530460 53340 530466
rect 53288 530402 53340 530408
rect 53300 528836 53328 530402
rect 54404 528836 54432 532374
rect 55496 530528 55548 530534
rect 55496 530470 55548 530476
rect 55508 528836 55536 530470
rect 56520 528836 56548 533530
rect 56612 528986 56640 567870
rect 66352 567860 66404 567866
rect 66352 567802 66404 567808
rect 60832 566500 60884 566506
rect 60832 566442 60884 566448
rect 60844 532386 60872 566442
rect 63500 565140 63552 565146
rect 63500 565082 63552 565088
rect 58716 532364 58768 532370
rect 60844 532358 61700 532386
rect 58716 532306 58768 532312
rect 56612 528958 57284 528986
rect 57256 528850 57284 528958
rect 57256 528822 57638 528850
rect 58728 528836 58756 532306
rect 60832 532296 60884 532302
rect 60832 532238 60884 532244
rect 59820 531276 59872 531282
rect 59820 531218 59872 531224
rect 59832 528836 59860 531218
rect 60844 528836 60872 532238
rect 61672 528850 61700 532358
rect 63040 532228 63092 532234
rect 63040 532170 63092 532176
rect 61672 528822 61962 528850
rect 63052 528836 63080 532170
rect 63512 528986 63540 565082
rect 65156 531140 65208 531146
rect 65156 531082 65208 531088
rect 63512 528958 63724 528986
rect 63696 528850 63724 528958
rect 63696 528822 64078 528850
rect 65168 528836 65196 531082
rect 66364 528850 66392 567802
rect 67640 563712 67692 563718
rect 67640 563654 67692 563660
rect 67364 532160 67416 532166
rect 67364 532102 67416 532108
rect 66286 528822 66392 528850
rect 67376 528836 67404 532102
rect 67652 528986 67680 563654
rect 71780 562352 71832 562358
rect 71780 562294 71832 562300
rect 69480 532092 69532 532098
rect 69480 532034 69532 532040
rect 67652 528958 68140 528986
rect 68112 528850 68140 528958
rect 68112 528822 68402 528850
rect 69492 528836 69520 532034
rect 70584 531208 70636 531214
rect 70584 531150 70636 531156
rect 70596 528836 70624 531150
rect 71596 531072 71648 531078
rect 71596 531014 71648 531020
rect 71608 528836 71636 531014
rect 71792 529258 71820 562294
rect 73802 532672 73858 532681
rect 73802 532607 73858 532616
rect 71792 529230 72372 529258
rect 72344 528850 72372 529230
rect 72344 528822 72726 528850
rect 73816 528836 73844 532607
rect 74552 528850 74580 570590
rect 112548 569906 112576 571526
rect 138676 569906 138704 700470
rect 218992 700466 219020 703520
rect 267660 700534 267688 703520
rect 283852 703474 283880 703520
rect 283852 703446 283972 703474
rect 250628 700528 250680 700534
rect 250628 700470 250680 700476
rect 267648 700528 267700 700534
rect 267648 700470 267700 700476
rect 282184 700528 282236 700534
rect 282184 700470 282236 700476
rect 138756 700460 138808 700466
rect 138756 700402 138808 700408
rect 218980 700460 219032 700466
rect 218980 700402 219032 700408
rect 138768 605826 138796 700402
rect 250640 698698 250668 700470
rect 250628 698692 250680 698698
rect 250628 698634 250680 698640
rect 252560 698692 252612 698698
rect 252560 698634 252612 698640
rect 252572 696930 252600 698634
rect 252560 696924 252612 696930
rect 252560 696866 252612 696872
rect 260012 696924 260064 696930
rect 260012 696866 260064 696872
rect 260024 694822 260052 696866
rect 260012 694816 260064 694822
rect 260012 694758 260064 694764
rect 267004 694816 267056 694822
rect 267004 694758 267056 694764
rect 267016 670682 267044 694758
rect 267004 670676 267056 670682
rect 267004 670618 267056 670624
rect 269764 670676 269816 670682
rect 269764 670618 269816 670624
rect 269776 659462 269804 670618
rect 269764 659456 269816 659462
rect 269764 659398 269816 659404
rect 271144 659456 271196 659462
rect 271144 659398 271196 659404
rect 271156 651574 271184 659398
rect 271144 651568 271196 651574
rect 271144 651510 271196 651516
rect 271972 651568 272024 651574
rect 271972 651510 272024 651516
rect 271984 648650 272012 651510
rect 271972 648644 272024 648650
rect 271972 648586 272024 648592
rect 274640 648576 274692 648582
rect 274640 648518 274692 648524
rect 274652 645862 274680 648518
rect 274640 645856 274692 645862
rect 274640 645798 274692 645804
rect 276664 645856 276716 645862
rect 276664 645798 276716 645804
rect 276676 633214 276704 645798
rect 276664 633208 276716 633214
rect 276664 633150 276716 633156
rect 278320 633208 278372 633214
rect 278320 633150 278372 633156
rect 278332 627910 278360 633150
rect 278320 627904 278372 627910
rect 278320 627846 278372 627852
rect 279148 627904 279200 627910
rect 279148 627846 279200 627852
rect 279160 618361 279188 627846
rect 279146 618352 279202 618361
rect 279146 618287 279202 618296
rect 138768 605798 138888 605826
rect 138860 605418 138888 605798
rect 138860 605390 139164 605418
rect 139136 594674 139164 605390
rect 139582 594824 139638 594833
rect 139582 594759 139638 594768
rect 139596 594726 139624 594759
rect 139216 594720 139268 594726
rect 139136 594668 139216 594674
rect 139136 594662 139268 594668
rect 139584 594720 139636 594726
rect 139584 594662 139636 594668
rect 139136 594646 139256 594662
rect 188048 574110 188384 574138
rect 189244 574110 189580 574138
rect 188356 572218 188384 574110
rect 189552 572354 189580 574110
rect 190288 574110 190440 574138
rect 191636 574110 191788 574138
rect 192924 574110 193168 574138
rect 194120 574110 194456 574138
rect 195316 574110 195652 574138
rect 196512 574110 196848 574138
rect 197800 574110 198136 574138
rect 198996 574110 199332 574138
rect 200192 574110 200528 574138
rect 189540 572348 189592 572354
rect 189540 572290 189592 572296
rect 188344 572212 188396 572218
rect 188344 572154 188396 572160
rect 190288 572082 190316 574110
rect 190276 572076 190328 572082
rect 190276 572018 190328 572024
rect 191760 571470 191788 574110
rect 191748 571464 191800 571470
rect 191748 571406 191800 571412
rect 193140 571402 193168 574110
rect 194428 571946 194456 574110
rect 194600 572212 194652 572218
rect 194600 572154 194652 572160
rect 194416 571940 194468 571946
rect 194416 571882 194468 571888
rect 193128 571396 193180 571402
rect 193128 571338 193180 571344
rect 112536 569900 112588 569906
rect 112536 569842 112588 569848
rect 138664 569900 138716 569906
rect 138664 569842 138716 569848
rect 78680 569288 78732 569294
rect 78680 569230 78732 569236
rect 75920 532024 75972 532030
rect 75920 531966 75972 531972
rect 74552 528822 74934 528850
rect 75932 528836 75960 531966
rect 77024 531004 77076 531010
rect 77024 530946 77076 530952
rect 77036 528836 77064 530946
rect 78128 530936 78180 530942
rect 78128 530878 78180 530884
rect 78140 528836 78168 530878
rect 78692 528850 78720 569230
rect 86960 560992 87012 560998
rect 86960 560934 87012 560940
rect 80242 533624 80298 533633
rect 80242 533559 80298 533568
rect 78692 528822 79166 528850
rect 80256 528836 80284 533559
rect 84568 533520 84620 533526
rect 82450 533488 82506 533497
rect 84568 533462 84620 533468
rect 82450 533423 82506 533432
rect 81348 530868 81400 530874
rect 81348 530810 81400 530816
rect 81360 528836 81388 530810
rect 82464 528836 82492 533423
rect 83464 530800 83516 530806
rect 83464 530742 83516 530748
rect 83476 528836 83504 530742
rect 84580 528836 84608 533462
rect 86684 533452 86736 533458
rect 86684 533394 86736 533400
rect 85672 530732 85724 530738
rect 85672 530674 85724 530680
rect 85684 528836 85712 530674
rect 86696 528836 86724 533394
rect 86972 528986 87000 560934
rect 100758 559600 100814 559609
rect 100758 559535 100814 559544
rect 90546 554160 90602 554169
rect 90546 554095 90602 554104
rect 90362 554024 90418 554033
rect 90362 553959 90418 553968
rect 90376 530670 90404 553959
rect 88892 530664 88944 530670
rect 88892 530606 88944 530612
rect 90364 530664 90416 530670
rect 90364 530606 90416 530612
rect 86972 528958 87184 528986
rect 87156 528850 87184 528958
rect 87156 528822 87814 528850
rect 88904 528836 88932 530606
rect 90560 530602 90588 554095
rect 95240 551336 95292 551342
rect 95240 551278 95292 551284
rect 91008 533384 91060 533390
rect 91008 533326 91060 533332
rect 89996 530596 90048 530602
rect 89996 530538 90048 530544
rect 90548 530596 90600 530602
rect 90548 530538 90600 530544
rect 90008 528836 90036 530538
rect 91020 528836 91048 533326
rect 92110 530904 92166 530913
rect 92110 530839 92166 530848
rect 92124 528836 92152 530839
rect 93214 530768 93270 530777
rect 93214 530703 93270 530712
rect 93228 528836 93256 530703
rect 94226 530632 94282 530641
rect 94226 530567 94282 530576
rect 94240 528836 94268 530567
rect 95252 528850 95280 551278
rect 97538 533352 97594 533361
rect 97538 533287 97594 533296
rect 96434 532536 96490 532545
rect 96434 532471 96490 532480
rect 95252 528822 95358 528850
rect 96448 528836 96476 532471
rect 97552 528836 97580 533287
rect 98550 532400 98606 532409
rect 100772 532386 100800 559535
rect 152464 535152 152516 535158
rect 152464 535094 152516 535100
rect 148140 535016 148192 535022
rect 148140 534958 148192 534964
rect 147956 534948 148008 534954
rect 147956 534890 148008 534896
rect 143816 534880 143868 534886
rect 143816 534822 143868 534828
rect 139492 534744 139544 534750
rect 139492 534686 139544 534692
rect 137376 534676 137428 534682
rect 137376 534618 137428 534624
rect 135260 534608 135312 534614
rect 135260 534550 135312 534556
rect 131948 534540 132000 534546
rect 131948 534482 132000 534488
rect 129832 534472 129884 534478
rect 129832 534414 129884 534420
rect 127716 534404 127768 534410
rect 127716 534346 127768 534352
rect 125508 534336 125560 534342
rect 125508 534278 125560 534284
rect 123392 534268 123444 534274
rect 123392 534210 123444 534216
rect 121184 534200 121236 534206
rect 121184 534142 121236 534148
rect 111064 534132 111116 534138
rect 111064 534074 111116 534080
rect 100772 532358 101260 532386
rect 98550 532335 98606 532344
rect 98564 528836 98592 532335
rect 100758 532264 100814 532273
rect 100758 532199 100814 532208
rect 99656 530664 99708 530670
rect 99656 530606 99708 530612
rect 99668 528836 99696 530606
rect 100772 528836 100800 532199
rect 101232 528714 101260 532358
rect 102874 532128 102930 532137
rect 102874 532063 102930 532072
rect 102888 528836 102916 532063
rect 103978 531992 104034 532001
rect 103978 531927 104034 531936
rect 103992 528836 104020 531927
rect 105084 530596 105136 530602
rect 105084 530538 105136 530544
rect 105096 528836 105124 530538
rect 111076 530262 111104 534074
rect 112628 530596 112680 530602
rect 112628 530538 112680 530544
rect 109316 530256 109368 530262
rect 109316 530198 109368 530204
rect 111064 530256 111116 530262
rect 111064 530198 111116 530204
rect 106094 529952 106150 529961
rect 106094 529887 106150 529896
rect 106108 528836 106136 529887
rect 108304 529236 108356 529242
rect 108304 529178 108356 529184
rect 108316 528836 108344 529178
rect 109328 528836 109356 530198
rect 111524 529304 111576 529310
rect 111524 529246 111576 529252
rect 111536 528836 111564 529246
rect 112640 528836 112668 530538
rect 119066 530224 119122 530233
rect 119066 530159 119122 530168
rect 115846 530088 115902 530097
rect 115846 530023 115902 530032
rect 115860 528836 115888 530023
rect 119080 528836 119108 530159
rect 120198 528834 120488 528850
rect 121196 528836 121224 534142
rect 122288 529984 122340 529990
rect 122288 529926 122340 529932
rect 122300 528836 122328 529926
rect 123404 528836 123432 534210
rect 124404 530052 124456 530058
rect 124404 529994 124456 530000
rect 124416 528836 124444 529994
rect 125520 528836 125548 534278
rect 126612 530120 126664 530126
rect 126612 530062 126664 530068
rect 126624 528836 126652 530062
rect 127728 528836 127756 534346
rect 128728 530188 128780 530194
rect 128728 530130 128780 530136
rect 128740 528836 128768 530130
rect 129844 528836 129872 534414
rect 130936 530256 130988 530262
rect 130936 530198 130988 530204
rect 130948 528836 130976 530198
rect 131960 528836 131988 534482
rect 133052 530324 133104 530330
rect 133052 530266 133104 530272
rect 133064 528836 133092 530266
rect 134432 528896 134484 528902
rect 134182 528844 134432 528850
rect 134182 528838 134484 528844
rect 120198 528828 120500 528834
rect 120198 528822 120448 528828
rect 134182 528822 134472 528838
rect 135272 528836 135300 534550
rect 136548 528964 136600 528970
rect 136548 528906 136600 528912
rect 136560 528850 136588 528906
rect 136298 528822 136588 528850
rect 137388 528836 137416 534618
rect 138480 529032 138532 529038
rect 138480 528974 138532 528980
rect 138492 528836 138520 528974
rect 139504 528836 139532 534686
rect 141698 531448 141754 531457
rect 141698 531383 141754 531392
rect 140596 529100 140648 529106
rect 140596 529042 140648 529048
rect 140608 528836 140636 529042
rect 141712 528836 141740 531383
rect 142804 529168 142856 529174
rect 142804 529110 142856 529116
rect 142816 528836 142844 529110
rect 143828 528836 143856 534822
rect 147968 530874 147996 534890
rect 146024 530868 146076 530874
rect 146024 530810 146076 530816
rect 147956 530868 148008 530874
rect 147956 530810 148008 530816
rect 144920 529372 144972 529378
rect 144920 529314 144972 529320
rect 144932 528836 144960 529314
rect 146036 528836 146064 530810
rect 147036 529440 147088 529446
rect 147036 529382 147088 529388
rect 147048 528836 147076 529382
rect 148152 528836 148180 534958
rect 150348 531140 150400 531146
rect 150348 531082 150400 531088
rect 149244 529508 149296 529514
rect 149244 529450 149296 529456
rect 149256 528836 149284 529450
rect 150360 528836 150388 531082
rect 151360 529576 151412 529582
rect 151360 529518 151412 529524
rect 151372 528836 151400 529518
rect 152476 528836 152504 535094
rect 156328 535084 156380 535090
rect 156328 535026 156380 535032
rect 154670 532808 154726 532817
rect 154670 532743 154726 532752
rect 153566 531584 153622 531593
rect 153566 531519 153622 531528
rect 153580 528836 153608 531519
rect 154684 528836 154712 532743
rect 155682 531720 155738 531729
rect 155682 531655 155738 531664
rect 155696 528836 155724 531655
rect 156340 531146 156368 535026
rect 167000 534812 167052 534818
rect 167000 534754 167052 534760
rect 166446 532944 166502 532953
rect 166446 532879 166502 532888
rect 162214 531856 162270 531865
rect 162214 531791 162270 531800
rect 161112 531480 161164 531486
rect 161112 531422 161164 531428
rect 158904 531412 158956 531418
rect 158904 531354 158956 531360
rect 156788 531344 156840 531350
rect 156788 531286 156840 531292
rect 156328 531140 156380 531146
rect 156328 531082 156380 531088
rect 156800 528836 156828 531286
rect 157892 529644 157944 529650
rect 157892 529586 157944 529592
rect 157904 528836 157932 529586
rect 158916 528836 158944 531354
rect 160008 529712 160060 529718
rect 160008 529654 160060 529660
rect 160020 528836 160048 529654
rect 161124 528836 161152 531422
rect 162228 528836 162256 531791
rect 163228 531548 163280 531554
rect 163228 531490 163280 531496
rect 163240 528836 163268 531490
rect 165436 529780 165488 529786
rect 165436 529722 165488 529728
rect 165448 528836 165476 529722
rect 166460 528836 166488 532879
rect 167012 530602 167040 534754
rect 175094 533216 175150 533225
rect 175094 533151 175150 533160
rect 170770 533080 170826 533089
rect 170770 533015 170826 533024
rect 167552 531616 167604 531622
rect 167552 531558 167604 531564
rect 167000 530596 167052 530602
rect 167000 530538 167052 530544
rect 167564 528836 167592 531558
rect 169760 530392 169812 530398
rect 169760 530334 169812 530340
rect 169772 528836 169800 530334
rect 170784 528836 170812 533015
rect 173992 530528 174044 530534
rect 173992 530470 174044 530476
rect 171876 530460 171928 530466
rect 171876 530402 171928 530408
rect 171888 528836 171916 530402
rect 174004 528836 174032 530470
rect 175108 528836 175136 533151
rect 193404 533044 193456 533050
rect 193404 532986 193456 532992
rect 192392 532976 192444 532982
rect 192392 532918 192444 532924
rect 189080 532908 189132 532914
rect 189080 532850 189132 532856
rect 183744 532840 183796 532846
rect 183744 532782 183796 532788
rect 177304 532772 177356 532778
rect 177304 532714 177356 532720
rect 176200 530596 176252 530602
rect 176200 530538 176252 530544
rect 176212 528836 176240 530538
rect 177316 528836 177344 532714
rect 182640 530800 182692 530806
rect 182640 530742 182692 530748
rect 180524 530732 180576 530738
rect 180524 530674 180576 530680
rect 178316 530664 178368 530670
rect 178316 530606 178368 530612
rect 178328 528836 178356 530606
rect 179420 529780 179472 529786
rect 179420 529722 179472 529728
rect 179432 528836 179460 529722
rect 180536 528836 180564 530674
rect 182652 528836 182680 530742
rect 183756 528836 183784 532782
rect 188066 531992 188122 532001
rect 188066 531927 188122 531936
rect 184848 531072 184900 531078
rect 184848 531014 184900 531020
rect 184860 528836 184888 531014
rect 186964 530936 187016 530942
rect 186964 530878 187016 530884
rect 186976 528836 187004 530878
rect 188080 528836 188108 531927
rect 189092 528836 189120 532850
rect 191288 529848 191340 529854
rect 191288 529790 191340 529796
rect 191300 528836 191328 529790
rect 192404 528836 192432 532918
rect 193416 528836 193444 532986
rect 194612 528986 194640 572154
rect 195624 571878 195652 574110
rect 195980 572348 196032 572354
rect 195980 572290 196032 572296
rect 195612 571872 195664 571878
rect 195612 571814 195664 571820
rect 194612 528958 195100 528986
rect 120448 528770 120500 528776
rect 117136 528760 117188 528766
rect 31864 528686 32890 528714
rect 101232 528686 101798 528714
rect 113666 528698 114048 528714
rect 116886 528708 117136 528714
rect 116886 528702 117188 528708
rect 195072 528714 195100 528958
rect 195992 528714 196020 572290
rect 196820 572218 196848 574110
rect 198108 572354 198136 574110
rect 199304 572490 199332 574110
rect 199292 572484 199344 572490
rect 199292 572426 199344 572432
rect 198096 572348 198148 572354
rect 198096 572290 198148 572296
rect 196808 572212 196860 572218
rect 196808 572154 196860 572160
rect 197360 572076 197412 572082
rect 197360 572018 197412 572024
rect 197372 528850 197400 572018
rect 200120 571940 200172 571946
rect 200120 571882 200172 571888
rect 198832 571464 198884 571470
rect 198832 571406 198884 571412
rect 198740 571396 198792 571402
rect 198740 571338 198792 571344
rect 198752 531078 198780 571338
rect 198740 531072 198792 531078
rect 198740 531014 198792 531020
rect 197372 528822 197754 528850
rect 198844 528836 198872 571406
rect 199660 531072 199712 531078
rect 199660 531014 199712 531020
rect 199672 528850 199700 531014
rect 199672 528822 199962 528850
rect 200132 528714 200160 571882
rect 200500 571470 200528 574110
rect 201420 574110 201480 574138
rect 202676 574110 202828 574138
rect 203872 574110 204208 574138
rect 205068 574110 205404 574138
rect 206356 574110 206692 574138
rect 207552 574110 207888 574138
rect 208748 574110 209084 574138
rect 210036 574110 210372 574138
rect 211232 574110 211568 574138
rect 212428 574110 212488 574138
rect 213624 574110 213868 574138
rect 214912 574110 215248 574138
rect 216108 574110 216444 574138
rect 217304 574110 217640 574138
rect 218592 574110 218928 574138
rect 219788 574110 220124 574138
rect 220984 574110 221320 574138
rect 201420 571538 201448 574110
rect 201500 571872 201552 571878
rect 201500 571814 201552 571820
rect 201408 571532 201460 571538
rect 201408 571474 201460 571480
rect 200488 571464 200540 571470
rect 200488 571406 200540 571412
rect 201512 528714 201540 571814
rect 202800 571606 202828 574110
rect 202880 572348 202932 572354
rect 202880 572290 202932 572296
rect 202788 571600 202840 571606
rect 202788 571542 202840 571548
rect 202892 531078 202920 572290
rect 202972 572212 203024 572218
rect 202972 572154 203024 572160
rect 202880 531072 202932 531078
rect 202880 531014 202932 531020
rect 202984 528850 203012 572154
rect 204180 571402 204208 574110
rect 204260 572484 204312 572490
rect 204260 572426 204312 572432
rect 204168 571396 204220 571402
rect 204168 571338 204220 571344
rect 203892 531072 203944 531078
rect 203892 531014 203944 531020
rect 203904 528850 203932 531014
rect 204272 528986 204300 572426
rect 205376 571946 205404 574110
rect 206664 572150 206692 574110
rect 206652 572144 206704 572150
rect 206652 572086 206704 572092
rect 207860 572082 207888 574110
rect 209056 572218 209084 574110
rect 209044 572212 209096 572218
rect 209044 572154 209096 572160
rect 207848 572076 207900 572082
rect 207848 572018 207900 572024
rect 205364 571940 205416 571946
rect 205364 571882 205416 571888
rect 209780 571940 209832 571946
rect 209780 571882 209832 571888
rect 208400 571600 208452 571606
rect 208400 571542 208452 571548
rect 207020 571532 207072 571538
rect 207020 571474 207072 571480
rect 205640 571464 205692 571470
rect 205640 571406 205692 571412
rect 205652 528986 205680 571406
rect 207032 528986 207060 571474
rect 204272 528958 204852 528986
rect 205652 528958 206140 528986
rect 207032 528958 207244 528986
rect 202984 528822 203182 528850
rect 203904 528822 204194 528850
rect 204824 528714 204852 528958
rect 206112 528850 206140 528958
rect 207216 528850 207244 528958
rect 208412 528850 208440 571542
rect 208492 571396 208544 571402
rect 208492 571338 208544 571344
rect 208504 529258 208532 571338
rect 208504 529230 209268 529258
rect 209240 528850 209268 529230
rect 209792 528986 209820 571882
rect 210344 571402 210372 574110
rect 211160 572144 211212 572150
rect 211160 572086 211212 572092
rect 210332 571396 210384 571402
rect 210332 571338 210384 571344
rect 211172 528986 211200 572086
rect 211540 571470 211568 574110
rect 212460 571538 212488 574110
rect 212540 572076 212592 572082
rect 212540 572018 212592 572024
rect 212448 571532 212500 571538
rect 212448 571474 212500 571480
rect 211528 571464 211580 571470
rect 211528 571406 211580 571412
rect 209792 528958 210372 528986
rect 211172 528958 211476 528986
rect 210344 528850 210372 528958
rect 211448 528850 211476 528958
rect 212552 528850 212580 572018
rect 213840 571606 213868 574110
rect 213920 572212 213972 572218
rect 213920 572154 213972 572160
rect 213828 571600 213880 571606
rect 213828 571542 213880 571548
rect 206112 528822 206402 528850
rect 207216 528822 207506 528850
rect 208412 528822 208518 528850
rect 209240 528822 209622 528850
rect 210344 528822 210726 528850
rect 211448 528822 211738 528850
rect 212552 528822 212842 528850
rect 213932 528836 213960 572154
rect 215220 571402 215248 574110
rect 216416 571674 216444 574110
rect 217612 571742 217640 574110
rect 218900 572150 218928 574110
rect 218888 572144 218940 572150
rect 218888 572086 218940 572092
rect 217600 571736 217652 571742
rect 217600 571678 217652 571684
rect 216404 571668 216456 571674
rect 216404 571610 216456 571616
rect 219440 571668 219492 571674
rect 219440 571610 219492 571616
rect 218060 571600 218112 571606
rect 218060 571542 218112 571548
rect 216680 571532 216732 571538
rect 216680 571474 216732 571480
rect 215300 571464 215352 571470
rect 215300 571406 215352 571412
rect 214012 571396 214064 571402
rect 214012 571338 214064 571344
rect 215208 571396 215260 571402
rect 215208 571338 215260 571344
rect 214024 528986 214052 571338
rect 214024 528958 214788 528986
rect 214760 528850 214788 528958
rect 214760 528822 215050 528850
rect 215312 528714 215340 571406
rect 216692 528850 216720 571474
rect 218072 528850 218100 571542
rect 218152 571396 218204 571402
rect 218152 571338 218204 571344
rect 218164 528986 218192 571338
rect 218164 528958 218836 528986
rect 216692 528822 217166 528850
rect 218072 528822 218270 528850
rect 218808 528714 218836 528958
rect 219452 528714 219480 571610
rect 220096 571606 220124 574110
rect 220820 571736 220872 571742
rect 220820 571678 220872 571684
rect 220084 571600 220136 571606
rect 220084 571542 220136 571548
rect 220832 528714 220860 571678
rect 221292 571402 221320 574110
rect 222120 574110 222180 574138
rect 223468 574110 223528 574138
rect 224664 574110 224908 574138
rect 225860 574110 226196 574138
rect 227148 574110 227484 574138
rect 228344 574110 228680 574138
rect 229540 574110 229876 574138
rect 230736 574110 231072 574138
rect 232024 574110 232360 574138
rect 222120 571470 222148 574110
rect 222200 572144 222252 572150
rect 222200 572086 222252 572092
rect 222108 571464 222160 571470
rect 222108 571406 222160 571412
rect 221280 571396 221332 571402
rect 221280 571338 221332 571344
rect 222212 528850 222240 572086
rect 223500 571538 223528 574110
rect 224880 571606 224908 574110
rect 223672 571600 223724 571606
rect 223672 571542 223724 571548
rect 224868 571600 224920 571606
rect 224868 571542 224920 571548
rect 223488 571532 223540 571538
rect 223488 571474 223540 571480
rect 223580 571396 223632 571402
rect 223580 571338 223632 571344
rect 223592 531146 223620 571338
rect 223580 531140 223632 531146
rect 223580 531082 223632 531088
rect 223684 528850 223712 571542
rect 224960 571464 225012 571470
rect 224960 571406 225012 571412
rect 224316 531140 224368 531146
rect 224316 531082 224368 531088
rect 222212 528822 222594 528850
rect 223606 528822 223712 528850
rect 224328 528850 224356 531082
rect 224972 528986 225000 571406
rect 226168 571402 226196 574110
rect 227456 571946 227484 574110
rect 227444 571940 227496 571946
rect 227444 571882 227496 571888
rect 228652 571674 228680 574110
rect 229100 571940 229152 571946
rect 229100 571882 229152 571888
rect 228640 571668 228692 571674
rect 228640 571610 228692 571616
rect 227812 571600 227864 571606
rect 227812 571542 227864 571548
rect 226340 571532 226392 571538
rect 226340 571474 226392 571480
rect 226156 571396 226208 571402
rect 226156 571338 226208 571344
rect 224972 528958 225276 528986
rect 224328 528822 224710 528850
rect 225248 528714 225276 528958
rect 226352 528714 226380 571474
rect 227720 571396 227772 571402
rect 227720 571338 227772 571344
rect 227732 531146 227760 571338
rect 227720 531140 227772 531146
rect 227720 531082 227772 531088
rect 227824 528850 227852 571542
rect 228732 531140 228784 531146
rect 228732 531082 228784 531088
rect 228744 528850 228772 531082
rect 229112 528986 229140 571882
rect 229848 571402 229876 574110
rect 230480 571668 230532 571674
rect 230480 571610 230532 571616
rect 229836 571396 229888 571402
rect 229836 571338 229888 571344
rect 229112 528958 229692 528986
rect 227824 528822 227930 528850
rect 228744 528822 229034 528850
rect 229664 528714 229692 528958
rect 230492 528714 230520 571610
rect 231044 571538 231072 574110
rect 231032 571532 231084 571538
rect 231032 571474 231084 571480
rect 232332 571402 232360 574110
rect 233160 574110 233220 574138
rect 234416 574110 234568 574138
rect 235704 574110 235948 574138
rect 236900 574110 237328 574138
rect 238096 574110 238616 574138
rect 239292 574110 239628 574138
rect 240580 574110 240916 574138
rect 241776 574110 242112 574138
rect 242972 574110 243032 574138
rect 244168 574110 244228 574138
rect 245456 574110 245608 574138
rect 246652 574110 246988 574138
rect 247848 574110 248368 574138
rect 233160 571470 233188 574110
rect 233332 571532 233384 571538
rect 233332 571474 233384 571480
rect 233148 571464 233200 571470
rect 233148 571406 233200 571412
rect 231860 571396 231912 571402
rect 231860 571338 231912 571344
rect 232320 571396 232372 571402
rect 232320 571338 232372 571344
rect 233240 571396 233292 571402
rect 233240 571338 233292 571344
rect 231872 528850 231900 571338
rect 233252 531146 233280 571338
rect 233240 531140 233292 531146
rect 233240 531082 233292 531088
rect 231872 528822 232254 528850
rect 233344 528836 233372 571474
rect 234540 571402 234568 574110
rect 235920 571470 235948 574110
rect 234620 571464 234672 571470
rect 234620 571406 234672 571412
rect 235908 571464 235960 571470
rect 235908 571406 235960 571412
rect 237300 571418 237328 574110
rect 238588 572098 238616 574110
rect 238588 572070 238800 572098
rect 237472 571464 237524 571470
rect 234528 571396 234580 571402
rect 234528 571338 234580 571344
rect 234068 531140 234120 531146
rect 234068 531082 234120 531088
rect 234080 528850 234108 531082
rect 234080 528822 234370 528850
rect 234632 528714 234660 571406
rect 236000 571396 236052 571402
rect 237300 571390 237420 571418
rect 237472 571406 237524 571412
rect 236000 571338 236052 571344
rect 236012 528714 236040 571338
rect 237392 531146 237420 571390
rect 237380 531140 237432 531146
rect 237380 531082 237432 531088
rect 237484 528850 237512 571406
rect 238300 531140 238352 531146
rect 238300 531082 238352 531088
rect 238312 528850 238340 531082
rect 237484 528822 237682 528850
rect 238312 528822 238694 528850
rect 238772 528714 238800 572070
rect 239600 571402 239628 574110
rect 240888 571402 240916 574110
rect 242084 571402 242112 574110
rect 239588 571396 239640 571402
rect 239588 571338 239640 571344
rect 240140 571396 240192 571402
rect 240140 571338 240192 571344
rect 240876 571396 240928 571402
rect 240876 571338 240928 571344
rect 241520 571396 241572 571402
rect 241520 571338 241572 571344
rect 242072 571396 242124 571402
rect 242072 571338 242124 571344
rect 242900 571396 242952 571402
rect 242900 571338 242952 571344
rect 240152 528714 240180 571338
rect 241532 528850 241560 571338
rect 242912 528850 242940 571338
rect 243004 529258 243032 574110
rect 244200 571418 244228 574110
rect 245580 571418 245608 574110
rect 246960 571418 246988 574110
rect 248340 572098 248368 574110
rect 248524 574110 249136 574138
rect 249812 574110 250332 574138
rect 251192 574110 251528 574138
rect 252664 574110 252724 574138
rect 253952 574110 254012 574138
rect 254872 574110 255208 574138
rect 256068 574110 256404 574138
rect 257356 574110 257692 574138
rect 258184 574110 258888 574138
rect 259472 574110 260084 574138
rect 260852 574110 261280 574138
rect 262232 574110 262568 574138
rect 263612 574110 263764 574138
rect 264624 574110 264960 574138
rect 265912 574110 266248 574138
rect 267108 574110 267444 574138
rect 268304 574110 268640 574138
rect 269500 574110 269836 574138
rect 270788 574110 271124 574138
rect 271984 574110 272320 574138
rect 273272 574110 273516 574138
rect 274652 574110 274804 574138
rect 275664 574110 276000 574138
rect 276860 574110 277196 574138
rect 278056 574110 278392 574138
rect 279344 574110 279680 574138
rect 280540 574110 280876 574138
rect 281736 574110 282072 574138
rect 248340 572070 248460 572098
rect 244200 571390 244320 571418
rect 245580 571390 245700 571418
rect 246960 571390 247080 571418
rect 243004 529230 243676 529258
rect 241532 528822 241914 528850
rect 242912 528822 243018 528850
rect 243648 528714 243676 529230
rect 244292 528986 244320 571390
rect 244292 528958 244780 528986
rect 244752 528714 244780 528958
rect 245672 528714 245700 571390
rect 247052 528850 247080 571390
rect 247052 528822 247342 528850
rect 248432 528836 248460 572070
rect 248524 528714 248552 574110
rect 249812 528714 249840 574110
rect 251192 528714 251220 574110
rect 252664 528850 252692 574110
rect 253952 571418 253980 574110
rect 253860 571390 253980 571418
rect 254872 571402 254900 574110
rect 256068 571402 256096 574110
rect 257356 571402 257384 574110
rect 254860 571396 254912 571402
rect 253860 528850 253888 571390
rect 254860 571338 254912 571344
rect 255320 571396 255372 571402
rect 255320 571338 255372 571344
rect 256056 571396 256108 571402
rect 256056 571338 256108 571344
rect 256700 571396 256752 571402
rect 256700 571338 256752 571344
rect 257344 571396 257396 571402
rect 257344 571338 257396 571344
rect 253940 571328 253992 571334
rect 253940 571270 253992 571276
rect 252664 528822 252770 528850
rect 253782 528822 253888 528850
rect 253952 528714 253980 571270
rect 255332 528714 255360 571338
rect 256712 528850 256740 571338
rect 258184 528850 258212 574110
rect 259472 571418 259500 574110
rect 260852 571418 260880 574110
rect 262232 571418 262260 574110
rect 263612 571418 263640 574110
rect 259380 571390 259500 571418
rect 260760 571390 260880 571418
rect 262140 571390 262260 571418
rect 263416 571396 263468 571402
rect 259380 528850 259408 571390
rect 260760 528850 260788 571390
rect 262140 531146 262168 571390
rect 263416 571338 263468 571344
rect 263520 571390 263640 571418
rect 264624 571402 264652 574110
rect 265912 571402 265940 574110
rect 267108 571402 267136 574110
rect 268304 571810 268332 574110
rect 267648 571804 267700 571810
rect 267648 571746 267700 571752
rect 268292 571804 268344 571810
rect 268292 571746 268344 571752
rect 264612 571396 264664 571402
rect 261300 531140 261352 531146
rect 261300 531082 261352 531088
rect 262128 531140 262180 531146
rect 262128 531082 262180 531088
rect 262404 531140 262456 531146
rect 262404 531082 262456 531088
rect 256712 528822 257002 528850
rect 258106 528822 258212 528850
rect 259210 528822 259408 528850
rect 260314 528822 260788 528850
rect 261312 528836 261340 531082
rect 262416 528836 262444 531082
rect 263428 528850 263456 571338
rect 263520 531146 263548 571390
rect 264612 571338 264664 571344
rect 264888 571396 264940 571402
rect 264888 571338 264940 571344
rect 265900 571396 265952 571402
rect 265900 571338 265952 571344
rect 266268 571396 266320 571402
rect 266268 571338 266320 571344
rect 267096 571396 267148 571402
rect 267096 571338 267148 571344
rect 263508 531140 263560 531146
rect 263508 531082 263560 531088
rect 264900 528850 264928 571338
rect 263428 528822 263534 528850
rect 264546 528822 264928 528850
rect 266280 528714 266308 571338
rect 267660 533390 267688 571746
rect 269028 571464 269080 571470
rect 269028 571406 269080 571412
rect 268936 571396 268988 571402
rect 268936 571338 268988 571344
rect 266728 533384 266780 533390
rect 266728 533326 266780 533332
rect 267648 533384 267700 533390
rect 267648 533326 267700 533332
rect 266740 528836 266768 533326
rect 268948 531146 268976 571338
rect 267832 531140 267884 531146
rect 267832 531082 267884 531088
rect 268936 531140 268988 531146
rect 268936 531082 268988 531088
rect 267844 528836 267872 531082
rect 269040 528850 269068 571406
rect 269500 571402 269528 574110
rect 270788 571470 270816 574110
rect 270776 571464 270828 571470
rect 270776 571406 270828 571412
rect 271788 571464 271840 571470
rect 271788 571406 271840 571412
rect 269488 571396 269540 571402
rect 269488 571338 269540 571344
rect 270408 571396 270460 571402
rect 270408 571338 270460 571344
rect 268870 528822 269068 528850
rect 270420 528714 270448 571338
rect 271800 531146 271828 571406
rect 271984 571402 272012 574110
rect 273076 571532 273128 571538
rect 273076 571474 273128 571480
rect 271972 571396 272024 571402
rect 271972 571338 272024 571344
rect 271052 531140 271104 531146
rect 271052 531082 271104 531088
rect 271788 531140 271840 531146
rect 271788 531082 271840 531088
rect 272064 531140 272116 531146
rect 272064 531082 272116 531088
rect 271064 528836 271092 531082
rect 272076 528836 272104 531082
rect 273088 528850 273116 571474
rect 273272 571470 273300 574110
rect 273260 571464 273312 571470
rect 273260 571406 273312 571412
rect 274548 571464 274600 571470
rect 274548 571406 274600 571412
rect 273168 571396 273220 571402
rect 273168 571338 273220 571344
rect 273180 531146 273208 571338
rect 273168 531140 273220 531146
rect 273168 531082 273220 531088
rect 274560 528850 274588 571406
rect 274652 571402 274680 574110
rect 275664 571538 275692 574110
rect 275652 571532 275704 571538
rect 275652 571474 275704 571480
rect 276860 571470 276888 574110
rect 276848 571464 276900 571470
rect 276848 571406 276900 571412
rect 277308 571464 277360 571470
rect 277308 571406 277360 571412
rect 274640 571396 274692 571402
rect 274640 571338 274692 571344
rect 275928 571396 275980 571402
rect 275928 571338 275980 571344
rect 273088 528822 273194 528850
rect 274298 528822 274588 528850
rect 275940 528714 275968 571338
rect 277320 531146 277348 571406
rect 278056 571402 278084 574110
rect 278688 571532 278740 571538
rect 278688 571474 278740 571480
rect 278044 571396 278096 571402
rect 278044 571338 278096 571344
rect 278596 571396 278648 571402
rect 278596 571338 278648 571344
rect 278608 531146 278636 571338
rect 276388 531140 276440 531146
rect 276388 531082 276440 531088
rect 277308 531140 277360 531146
rect 277308 531082 277360 531088
rect 277492 531140 277544 531146
rect 277492 531082 277544 531088
rect 278596 531140 278648 531146
rect 278596 531082 278648 531088
rect 276400 528836 276428 531082
rect 277504 528836 277532 531082
rect 278700 528850 278728 571474
rect 279344 571470 279372 574110
rect 279332 571464 279384 571470
rect 279332 571406 279384 571412
rect 280540 571402 280568 574110
rect 281736 571538 281764 574110
rect 281724 571532 281776 571538
rect 281724 571474 281776 571480
rect 280528 571396 280580 571402
rect 280528 571338 280580 571344
rect 281540 569220 281592 569226
rect 281540 569162 281592 569168
rect 280158 563816 280214 563825
rect 280158 563751 280214 563760
rect 280172 553217 280200 563751
rect 280158 553208 280214 553217
rect 280158 553143 280214 553152
rect 279516 552084 279568 552090
rect 279516 552026 279568 552032
rect 278622 528822 278728 528850
rect 113666 528692 114060 528698
rect 113666 528686 114008 528692
rect 116886 528686 117176 528702
rect 195072 528686 195638 528714
rect 195992 528686 196650 528714
rect 200132 528686 200974 528714
rect 201512 528686 202078 528714
rect 204824 528686 205298 528714
rect 215312 528686 216062 528714
rect 218808 528686 219282 528714
rect 219452 528686 220386 528714
rect 220832 528686 221490 528714
rect 225248 528686 225814 528714
rect 226352 528686 226826 528714
rect 229664 528686 230138 528714
rect 230492 528686 231150 528714
rect 234632 528686 235474 528714
rect 236012 528686 236578 528714
rect 238772 528686 239798 528714
rect 240152 528686 240902 528714
rect 243648 528686 244122 528714
rect 244752 528686 245226 528714
rect 245672 528686 246238 528714
rect 248524 528686 249458 528714
rect 249812 528686 250562 528714
rect 251192 528686 251666 528714
rect 253952 528686 254886 528714
rect 255332 528686 255990 528714
rect 265650 528686 266308 528714
rect 269974 528686 270448 528714
rect 275402 528686 275968 528714
rect 114008 528634 114060 528640
rect 110696 528624 110748 528630
rect 107566 528592 107622 528601
rect 107226 528550 107566 528578
rect 110446 528572 110696 528578
rect 110446 528566 110748 528572
rect 110446 528550 110736 528566
rect 107566 528527 107622 528536
rect 194600 528488 194652 528494
rect 190210 528426 190408 528442
rect 194534 528436 194600 528442
rect 194534 528430 194652 528436
rect 190210 528420 190420 528426
rect 190210 528414 190368 528420
rect 194534 528414 194640 528430
rect 190368 528362 190420 528368
rect 186136 528352 186188 528358
rect 115110 528320 115166 528329
rect 114770 528278 115110 528306
rect 115110 528255 115166 528264
rect 115938 528320 115994 528329
rect 181562 528290 181944 528306
rect 185886 528300 186136 528306
rect 185886 528294 186188 528300
rect 115938 528255 115940 528264
rect 115992 528255 115994 528264
rect 125324 528284 125376 528290
rect 115940 528226 115992 528232
rect 181562 528284 181956 528290
rect 181562 528278 181904 528284
rect 125324 528227 125376 528232
rect 185886 528278 186176 528294
rect 118240 528216 118292 528222
rect 117990 528164 118240 528170
rect 117990 528158 118292 528164
rect 125322 528218 125378 528227
rect 181904 528226 181956 528232
rect 164516 528216 164568 528222
rect 117990 528142 118280 528158
rect 125322 528153 125378 528162
rect 164358 528164 164516 528170
rect 169024 528216 169076 528222
rect 164358 528158 164568 528164
rect 168682 528164 169024 528170
rect 173256 528216 173308 528222
rect 168682 528158 169076 528164
rect 173006 528164 173256 528170
rect 173006 528158 173308 528164
rect 164358 528142 164556 528158
rect 168682 528142 169064 528158
rect 173006 528142 173296 528158
rect 105188 502982 106122 503010
rect 22112 499798 22140 502860
rect 22296 502846 23138 502874
rect 23492 502846 24242 502874
rect 22100 499792 22152 499798
rect 22100 499734 22152 499740
rect 21362 492552 21418 492561
rect 21362 492487 21418 492496
rect 20352 488776 20404 488782
rect 20352 488718 20404 488724
rect 16856 488708 16908 488714
rect 16856 488650 16908 488656
rect 16868 486948 16896 488650
rect 18604 488572 18656 488578
rect 18604 488514 18656 488520
rect 18616 486948 18644 488514
rect 20364 486948 20392 488718
rect 22296 488714 22324 502846
rect 22284 488708 22336 488714
rect 22284 488650 22336 488656
rect 22192 488640 22244 488646
rect 22192 488582 22244 488588
rect 22204 486948 22232 488582
rect 23492 488578 23520 502846
rect 25332 500954 25360 502860
rect 24216 500948 24268 500954
rect 24216 500890 24268 500896
rect 25320 500948 25372 500954
rect 25320 500890 25372 500896
rect 24124 499792 24176 499798
rect 24124 499734 24176 499740
rect 23480 488572 23532 488578
rect 23480 488514 23532 488520
rect 23940 488572 23992 488578
rect 23940 488514 23992 488520
rect 23952 486948 23980 488514
rect 24136 486470 24164 499734
rect 24228 488782 24256 500890
rect 26344 499730 26372 502860
rect 24308 499724 24360 499730
rect 24308 499666 24360 499672
rect 26332 499724 26384 499730
rect 26332 499666 26384 499672
rect 24216 488776 24268 488782
rect 24216 488718 24268 488724
rect 24320 488646 24348 499666
rect 26148 499656 26200 499662
rect 26148 499598 26200 499604
rect 25504 499588 25556 499594
rect 25504 499530 25556 499536
rect 24308 488640 24360 488646
rect 24308 488582 24360 488588
rect 25516 488578 25544 499530
rect 25504 488572 25556 488578
rect 25504 488514 25556 488520
rect 26160 486962 26188 499598
rect 27448 499594 27476 502860
rect 27528 500948 27580 500954
rect 27528 500890 27580 500896
rect 27436 499588 27488 499594
rect 27436 499530 27488 499536
rect 25806 486934 26188 486962
rect 27540 486948 27568 500890
rect 28552 499662 28580 502860
rect 29656 500954 29684 502860
rect 30484 502846 30682 502874
rect 29644 500948 29696 500954
rect 29644 500890 29696 500896
rect 30484 500834 30512 502846
rect 31772 500886 31800 502860
rect 30300 500806 30512 500834
rect 31668 500880 31720 500886
rect 31668 500822 31720 500828
rect 31760 500880 31812 500886
rect 31760 500822 31812 500828
rect 28540 499656 28592 499662
rect 28540 499598 28592 499604
rect 30300 488578 30328 500806
rect 29368 488572 29420 488578
rect 29368 488514 29420 488520
rect 30288 488572 30340 488578
rect 30288 488514 30340 488520
rect 29380 486948 29408 488514
rect 31680 486826 31708 500822
rect 32876 499594 32904 502860
rect 33902 502846 34468 502874
rect 31944 499588 31996 499594
rect 31944 499530 31996 499536
rect 32864 499588 32916 499594
rect 32864 499530 32916 499536
rect 31956 487098 31984 499530
rect 34440 488594 34468 502846
rect 34992 499594 35020 502860
rect 36096 499594 36124 502860
rect 34980 499588 35032 499594
rect 34980 499530 35032 499536
rect 35808 499588 35860 499594
rect 35808 499530 35860 499536
rect 36084 499588 36136 499594
rect 36084 499530 36136 499536
rect 37096 499588 37148 499594
rect 37096 499530 37148 499536
rect 35820 489870 35848 499530
rect 35808 489864 35860 489870
rect 35808 489806 35860 489812
rect 36544 489864 36596 489870
rect 36544 489806 36596 489812
rect 34440 488566 34560 488594
rect 31956 487070 32628 487098
rect 32600 486962 32628 487070
rect 34532 486962 34560 488566
rect 32600 486934 32982 486962
rect 34532 486934 34730 486962
rect 36556 486948 36584 489806
rect 37108 489258 37136 499530
rect 37096 489252 37148 489258
rect 37096 489194 37148 489200
rect 37200 489190 37228 502860
rect 38226 502846 38608 502874
rect 39330 502846 39988 502874
rect 38292 489252 38344 489258
rect 38292 489194 38344 489200
rect 37188 489184 37240 489190
rect 37188 489126 37240 489132
rect 38304 486948 38332 489194
rect 38580 488714 38608 502846
rect 39960 488782 39988 502846
rect 40420 499594 40448 502860
rect 41432 500750 41460 502860
rect 41420 500744 41472 500750
rect 41420 500686 41472 500692
rect 42536 500478 42564 502860
rect 42524 500472 42576 500478
rect 42524 500414 42576 500420
rect 43640 500410 43668 502860
rect 43628 500404 43680 500410
rect 43628 500346 43680 500352
rect 44744 500342 44772 502860
rect 45756 500886 45784 502860
rect 45744 500880 45796 500886
rect 45744 500822 45796 500828
rect 44732 500336 44784 500342
rect 44732 500278 44784 500284
rect 40408 499588 40460 499594
rect 40408 499530 40460 499536
rect 41328 499588 41380 499594
rect 41328 499530 41380 499536
rect 40132 489184 40184 489190
rect 40132 489126 40184 489132
rect 39948 488776 40000 488782
rect 39948 488718 40000 488724
rect 38568 488708 38620 488714
rect 38568 488650 38620 488656
rect 40144 486948 40172 489126
rect 41340 488578 41368 499530
rect 46860 489190 46888 502860
rect 47978 502846 48268 502874
rect 48990 502846 49648 502874
rect 47032 500744 47084 500750
rect 47032 500686 47084 500692
rect 46848 489184 46900 489190
rect 46848 489126 46900 489132
rect 43720 488776 43772 488782
rect 43720 488718 43772 488724
rect 41880 488708 41932 488714
rect 41880 488650 41932 488656
rect 41328 488572 41380 488578
rect 41328 488514 41380 488520
rect 41892 486948 41920 488650
rect 43732 486948 43760 488718
rect 45468 488572 45520 488578
rect 45468 488514 45520 488520
rect 45480 486948 45508 488514
rect 47044 486962 47072 500686
rect 47584 500472 47636 500478
rect 47584 500414 47636 500420
rect 47596 488578 47624 500414
rect 48240 489258 48268 502846
rect 48964 500404 49016 500410
rect 48964 500346 49016 500352
rect 48228 489252 48280 489258
rect 48228 489194 48280 489200
rect 48976 488646 49004 500346
rect 49620 489666 49648 502846
rect 50080 500954 50108 502860
rect 50068 500948 50120 500954
rect 50068 500890 50120 500896
rect 50988 500948 51040 500954
rect 50988 500890 51040 500896
rect 49608 489660 49660 489666
rect 49608 489602 49660 489608
rect 51000 489598 51028 500890
rect 51184 499798 51212 502860
rect 51172 499792 51224 499798
rect 51172 499734 51224 499740
rect 50988 489592 51040 489598
rect 50988 489534 51040 489540
rect 52288 489394 52316 502860
rect 53314 502846 53788 502874
rect 54418 502846 55168 502874
rect 52552 500336 52604 500342
rect 52552 500278 52604 500284
rect 52368 499792 52420 499798
rect 52368 499734 52420 499740
rect 52380 489530 52408 499734
rect 52368 489524 52420 489530
rect 52368 489466 52420 489472
rect 52276 489388 52328 489394
rect 52276 489330 52328 489336
rect 48964 488640 49016 488646
rect 48964 488582 49016 488588
rect 50896 488640 50948 488646
rect 50896 488582 50948 488588
rect 47584 488572 47636 488578
rect 47584 488514 47636 488520
rect 49056 488572 49108 488578
rect 49056 488514 49108 488520
rect 47044 486934 47334 486962
rect 49068 486948 49096 488514
rect 50908 486948 50936 488582
rect 52564 486962 52592 500278
rect 53760 489462 53788 502846
rect 53932 500880 53984 500886
rect 53932 500822 53984 500828
rect 53748 489456 53800 489462
rect 53748 489398 53800 489404
rect 53944 486962 53972 500822
rect 55140 488986 55168 502846
rect 55508 500342 55536 502860
rect 55496 500336 55548 500342
rect 55496 500278 55548 500284
rect 56416 500336 56468 500342
rect 56416 500278 56468 500284
rect 56428 489326 56456 500278
rect 56416 489320 56468 489326
rect 56416 489262 56468 489268
rect 56520 489190 56548 502860
rect 57638 502846 57928 502874
rect 58742 502846 59308 502874
rect 56232 489184 56284 489190
rect 56232 489126 56284 489132
rect 56508 489184 56560 489190
rect 56508 489126 56560 489132
rect 55128 488980 55180 488986
rect 55128 488922 55180 488928
rect 52564 486934 52670 486962
rect 53944 486934 54510 486962
rect 56244 486948 56272 489126
rect 57900 489054 57928 502846
rect 59280 489258 59308 502846
rect 59832 500954 59860 502860
rect 60844 500954 60872 502860
rect 61962 502846 62068 502874
rect 63066 502846 63448 502874
rect 59820 500948 59872 500954
rect 59820 500890 59872 500896
rect 60648 500948 60700 500954
rect 60648 500890 60700 500896
rect 60832 500948 60884 500954
rect 60832 500890 60884 500896
rect 61936 500948 61988 500954
rect 61936 500890 61988 500896
rect 59820 489660 59872 489666
rect 59820 489602 59872 489608
rect 58072 489252 58124 489258
rect 58072 489194 58124 489200
rect 59268 489252 59320 489258
rect 59268 489194 59320 489200
rect 57888 489048 57940 489054
rect 57888 488990 57940 488996
rect 58084 486948 58112 489194
rect 59832 486948 59860 489602
rect 60660 489122 60688 500890
rect 61948 489870 61976 500890
rect 61936 489864 61988 489870
rect 61936 489806 61988 489812
rect 62040 489802 62068 502846
rect 62028 489796 62080 489802
rect 62028 489738 62080 489744
rect 63420 489666 63448 502846
rect 64064 500954 64092 502860
rect 64052 500948 64104 500954
rect 64052 500890 64104 500896
rect 64788 500948 64840 500954
rect 64788 500890 64840 500896
rect 64800 489734 64828 500890
rect 65168 500138 65196 502860
rect 65156 500132 65208 500138
rect 65156 500074 65208 500080
rect 66168 500132 66220 500138
rect 66168 500074 66220 500080
rect 64788 489728 64840 489734
rect 64788 489670 64840 489676
rect 63408 489660 63460 489666
rect 63408 489602 63460 489608
rect 66180 489598 66208 500074
rect 66272 499798 66300 502860
rect 67390 502846 67496 502874
rect 68402 502846 68968 502874
rect 66260 499792 66312 499798
rect 66260 499734 66312 499740
rect 61660 489592 61712 489598
rect 61660 489534 61712 489540
rect 66168 489592 66220 489598
rect 66168 489534 66220 489540
rect 60648 489116 60700 489122
rect 60648 489058 60700 489064
rect 61672 486948 61700 489534
rect 63408 489524 63460 489530
rect 63408 489466 63460 489472
rect 63420 486948 63448 489466
rect 67468 489462 67496 502846
rect 67548 499792 67600 499798
rect 67548 499734 67600 499740
rect 67560 489530 67588 499734
rect 68940 490686 68968 502846
rect 69492 500954 69520 502860
rect 69480 500948 69532 500954
rect 69480 500890 69532 500896
rect 70308 500948 70360 500954
rect 70308 500890 70360 500896
rect 68928 490680 68980 490686
rect 68928 490622 68980 490628
rect 67548 489524 67600 489530
rect 67548 489466 67600 489472
rect 66996 489456 67048 489462
rect 66996 489398 67048 489404
rect 67456 489456 67508 489462
rect 67456 489398 67508 489404
rect 65156 489388 65208 489394
rect 65156 489330 65208 489336
rect 65168 486948 65196 489330
rect 67008 486948 67036 489398
rect 70320 489394 70348 500890
rect 70596 500206 70624 502860
rect 71622 502846 71728 502874
rect 72726 502846 73108 502874
rect 73830 502846 74488 502874
rect 70584 500200 70636 500206
rect 70584 500142 70636 500148
rect 70308 489388 70360 489394
rect 70308 489330 70360 489336
rect 71700 489326 71728 502846
rect 73080 492046 73108 502846
rect 73068 492040 73120 492046
rect 73068 491982 73120 491988
rect 70584 489320 70636 489326
rect 70584 489262 70636 489268
rect 71688 489320 71740 489326
rect 71688 489262 71740 489268
rect 68744 488980 68796 488986
rect 68744 488922 68796 488928
rect 68756 486948 68784 488922
rect 70596 486948 70624 489262
rect 74460 489190 74488 502846
rect 74552 502846 74934 502874
rect 74552 493406 74580 502846
rect 75932 499594 75960 502860
rect 75920 499588 75972 499594
rect 75920 499530 75972 499536
rect 77036 497486 77064 502860
rect 78154 502846 78628 502874
rect 77208 499588 77260 499594
rect 77208 499530 77260 499536
rect 77024 497480 77076 497486
rect 77024 497422 77076 497428
rect 74540 493400 74592 493406
rect 74540 493342 74592 493348
rect 77220 489258 77248 499530
rect 75920 489252 75972 489258
rect 75920 489194 75972 489200
rect 77208 489252 77260 489258
rect 77208 489194 77260 489200
rect 72332 489184 72384 489190
rect 72332 489126 72384 489132
rect 74448 489184 74500 489190
rect 74448 489126 74500 489132
rect 72344 486948 72372 489126
rect 74172 489048 74224 489054
rect 74172 488990 74224 488996
rect 74184 486948 74212 488990
rect 75932 486948 75960 489194
rect 77760 489116 77812 489122
rect 77760 489058 77812 489064
rect 77772 486948 77800 489058
rect 78600 488578 78628 502846
rect 79152 499594 79180 502860
rect 80256 499594 80284 502860
rect 79140 499588 79192 499594
rect 79140 499530 79192 499536
rect 79968 499588 80020 499594
rect 79968 499530 80020 499536
rect 80244 499588 80296 499594
rect 80244 499530 80296 499536
rect 81256 499588 81308 499594
rect 81256 499530 81308 499536
rect 79980 490618 80008 499530
rect 79968 490612 80020 490618
rect 79968 490554 80020 490560
rect 79508 489864 79560 489870
rect 79508 489806 79560 489812
rect 78588 488572 78640 488578
rect 78588 488514 78640 488520
rect 79520 486948 79548 489806
rect 81268 488646 81296 499530
rect 81360 498846 81388 502860
rect 82478 502846 82768 502874
rect 83490 502846 84148 502874
rect 81348 498840 81400 498846
rect 81348 498782 81400 498788
rect 81348 489796 81400 489802
rect 81348 489738 81400 489744
rect 81256 488640 81308 488646
rect 81256 488582 81308 488588
rect 81360 486948 81388 489738
rect 82740 488714 82768 502846
rect 84120 491978 84148 502846
rect 84580 499594 84608 502860
rect 85684 500274 85712 502860
rect 86710 502846 86908 502874
rect 85672 500268 85724 500274
rect 85672 500210 85724 500216
rect 84568 499588 84620 499594
rect 84568 499530 84620 499536
rect 85488 499588 85540 499594
rect 85488 499530 85540 499536
rect 84108 491972 84160 491978
rect 84108 491914 84160 491920
rect 84936 489728 84988 489734
rect 84936 489670 84988 489676
rect 83096 489660 83148 489666
rect 83096 489602 83148 489608
rect 82728 488708 82780 488714
rect 82728 488650 82780 488656
rect 83108 486948 83136 489602
rect 84948 486948 84976 489670
rect 85500 488782 85528 499530
rect 86684 489592 86736 489598
rect 86684 489534 86736 489540
rect 85488 488776 85540 488782
rect 85488 488718 85540 488724
rect 86696 486948 86724 489534
rect 86880 488850 86908 502846
rect 87800 499594 87828 502860
rect 88904 499594 88932 502860
rect 90008 499594 90036 502860
rect 90928 502846 91034 502874
rect 92138 502846 92428 502874
rect 93242 502846 93808 502874
rect 86960 499588 87012 499594
rect 86960 499530 87012 499536
rect 87788 499588 87840 499594
rect 87788 499530 87840 499536
rect 88892 499588 88944 499594
rect 88892 499530 88944 499536
rect 89628 499588 89680 499594
rect 89628 499530 89680 499536
rect 89996 499588 90048 499594
rect 89996 499530 90048 499536
rect 86972 493338 87000 499530
rect 86960 493332 87012 493338
rect 86960 493274 87012 493280
rect 88524 489524 88576 489530
rect 88524 489466 88576 489472
rect 86868 488844 86920 488850
rect 86868 488786 86920 488792
rect 88536 486948 88564 489466
rect 89640 488986 89668 499530
rect 90928 489802 90956 502846
rect 91008 499588 91060 499594
rect 91008 499530 91060 499536
rect 90916 489796 90968 489802
rect 90916 489738 90968 489744
rect 90272 489456 90324 489462
rect 90272 489398 90324 489404
rect 89628 488980 89680 488986
rect 89628 488922 89680 488928
rect 90284 486948 90312 489398
rect 91020 488918 91048 499530
rect 92112 490680 92164 490686
rect 92112 490622 92164 490628
rect 91008 488912 91060 488918
rect 91008 488854 91060 488860
rect 92124 486948 92152 490622
rect 92400 489054 92428 502846
rect 93780 489122 93808 502846
rect 94240 499594 94268 502860
rect 94504 500064 94556 500070
rect 94504 500006 94556 500012
rect 94228 499588 94280 499594
rect 94228 499530 94280 499536
rect 94516 491298 94544 500006
rect 95344 499594 95372 502860
rect 95148 499588 95200 499594
rect 95148 499530 95200 499536
rect 95332 499588 95384 499594
rect 95332 499530 95384 499536
rect 94504 491292 94556 491298
rect 94504 491234 94556 491240
rect 95160 489870 95188 499530
rect 95700 491292 95752 491298
rect 95700 491234 95752 491240
rect 95148 489864 95200 489870
rect 95148 489806 95200 489812
rect 93860 489388 93912 489394
rect 93860 489330 93912 489336
rect 93768 489116 93820 489122
rect 93768 489058 93820 489064
rect 92388 489048 92440 489054
rect 92388 488990 92440 488996
rect 93872 486948 93900 489330
rect 95712 486948 95740 491234
rect 96448 489598 96476 502860
rect 97566 502846 97948 502874
rect 98578 502846 99328 502874
rect 96528 499588 96580 499594
rect 96528 499530 96580 499536
rect 96540 489734 96568 499530
rect 96528 489728 96580 489734
rect 96528 489670 96580 489676
rect 97920 489666 97948 502846
rect 99012 492040 99064 492046
rect 99012 491982 99064 491988
rect 97908 489660 97960 489666
rect 97908 489602 97960 489608
rect 96436 489592 96488 489598
rect 96436 489534 96488 489540
rect 97448 489320 97500 489326
rect 97448 489262 97500 489268
rect 97460 486948 97488 489262
rect 99024 486962 99052 491982
rect 99300 489394 99328 502846
rect 99668 500954 99696 502860
rect 100772 500954 100800 502860
rect 101798 502846 101996 502874
rect 102902 502846 103468 502874
rect 99656 500948 99708 500954
rect 99656 500890 99708 500896
rect 100668 500948 100720 500954
rect 100668 500890 100720 500896
rect 100760 500948 100812 500954
rect 100760 500890 100812 500896
rect 100680 489462 100708 500890
rect 100668 489456 100720 489462
rect 100668 489398 100720 489404
rect 99288 489388 99340 489394
rect 99288 489330 99340 489336
rect 101968 489190 101996 502846
rect 102048 500948 102100 500954
rect 102048 500890 102100 500896
rect 102060 489530 102088 500890
rect 102140 493400 102192 493406
rect 102140 493342 102192 493348
rect 102048 489524 102100 489530
rect 102048 489466 102100 489472
rect 101036 489184 101088 489190
rect 101036 489126 101088 489132
rect 101956 489184 102008 489190
rect 101956 489126 102008 489132
rect 99024 486934 99314 486962
rect 101048 486948 101076 489126
rect 31142 486798 31708 486826
rect 102152 486826 102180 493342
rect 103440 489326 103468 502846
rect 103992 499662 104020 502860
rect 105096 500954 105124 502860
rect 105084 500948 105136 500954
rect 105084 500890 105136 500896
rect 105188 500834 105216 502982
rect 106188 500948 106240 500954
rect 106188 500890 106240 500896
rect 104912 500806 105216 500834
rect 103980 499656 104032 499662
rect 103980 499598 104032 499604
rect 104808 499656 104860 499662
rect 104808 499598 104860 499604
rect 103428 489320 103480 489326
rect 103428 489262 103480 489268
rect 104820 489258 104848 499598
rect 104912 497457 104940 500806
rect 104898 497448 104954 497457
rect 104898 497383 104954 497392
rect 104624 489252 104676 489258
rect 104624 489194 104676 489200
rect 104808 489252 104860 489258
rect 104808 489194 104860 489200
rect 104636 486948 104664 489194
rect 106200 489161 106228 500890
rect 107212 500041 107240 502860
rect 107672 502846 108330 502874
rect 109052 502846 109342 502874
rect 107198 500032 107254 500041
rect 107198 499967 107254 499976
rect 107672 497593 107700 502846
rect 109052 497729 109080 502846
rect 110432 498001 110460 502860
rect 110616 502846 111550 502874
rect 110418 497992 110474 498001
rect 110418 497927 110474 497936
rect 110616 497865 110644 502846
rect 112640 500313 112668 502860
rect 113192 502846 113666 502874
rect 113192 500449 113220 502846
rect 114560 502648 114612 502654
rect 114560 502590 114612 502596
rect 113178 500440 113234 500449
rect 113178 500375 113234 500384
rect 112626 500304 112682 500313
rect 112444 500268 112496 500274
rect 112626 500239 112682 500248
rect 112444 500210 112496 500216
rect 110602 497856 110658 497865
rect 110602 497791 110658 497800
rect 109038 497720 109094 497729
rect 109038 497655 109094 497664
rect 107658 497584 107714 497593
rect 107658 497519 107714 497528
rect 106280 497480 106332 497486
rect 106280 497422 106332 497428
rect 106186 489152 106242 489161
rect 106186 489087 106242 489096
rect 106292 486962 106320 497422
rect 112456 490618 112484 500210
rect 114572 500177 114600 502590
rect 114756 500585 114784 502860
rect 115584 502846 115874 502874
rect 115952 502846 116886 502874
rect 117332 502846 117990 502874
rect 118712 502846 119094 502874
rect 120092 502846 120198 502874
rect 120276 502846 121210 502874
rect 121472 502846 122314 502874
rect 115584 502654 115612 502846
rect 115572 502648 115624 502654
rect 115572 502590 115624 502596
rect 115952 500721 115980 502846
rect 115938 500712 115994 500721
rect 115938 500647 115994 500656
rect 114742 500576 114798 500585
rect 114742 500511 114798 500520
rect 117332 500274 117360 502846
rect 118712 500857 118740 502846
rect 120092 500857 120120 502846
rect 118698 500848 118754 500857
rect 118698 500783 118754 500792
rect 120078 500848 120134 500857
rect 120078 500783 120134 500792
rect 120276 500342 120304 502846
rect 121472 500954 121500 502846
rect 121460 500948 121512 500954
rect 121460 500890 121512 500896
rect 123404 500410 123432 502860
rect 124416 500546 124444 502860
rect 124404 500540 124456 500546
rect 124404 500482 124456 500488
rect 125520 500478 125548 502860
rect 126624 500886 126652 502860
rect 126612 500880 126664 500886
rect 126612 500822 126664 500828
rect 127728 500614 127756 502860
rect 128740 500750 128768 502860
rect 129844 500818 129872 502860
rect 129832 500812 129884 500818
rect 129832 500754 129884 500760
rect 128728 500744 128780 500750
rect 128728 500686 128780 500692
rect 130948 500682 130976 502860
rect 130936 500676 130988 500682
rect 130936 500618 130988 500624
rect 127716 500608 127768 500614
rect 127716 500550 127768 500556
rect 125508 500472 125560 500478
rect 125508 500414 125560 500420
rect 123392 500404 123444 500410
rect 123392 500346 123444 500352
rect 120264 500336 120316 500342
rect 120264 500278 120316 500284
rect 117320 500268 117372 500274
rect 117320 500210 117372 500216
rect 131960 500206 131988 502860
rect 132512 502846 133078 502874
rect 131948 500200 132000 500206
rect 114558 500168 114614 500177
rect 131948 500142 132000 500148
rect 114558 500103 114614 500112
rect 113180 498840 113232 498846
rect 113180 498782 113232 498788
rect 109960 490612 110012 490618
rect 109960 490554 110012 490560
rect 112444 490612 112496 490618
rect 112444 490554 112496 490560
rect 108212 488572 108264 488578
rect 108212 488514 108264 488520
rect 106292 486934 106490 486962
rect 108224 486948 108252 488514
rect 109972 486948 110000 490554
rect 111800 488640 111852 488646
rect 111800 488582 111852 488588
rect 111812 486948 111840 488582
rect 113192 486962 113220 498782
rect 132512 497486 132540 502846
rect 132590 500848 132646 500857
rect 132590 500783 132646 500792
rect 132604 499633 132632 500783
rect 134168 500041 134196 502860
rect 135272 500138 135300 502860
rect 135260 500132 135312 500138
rect 135260 500074 135312 500080
rect 134154 500032 134210 500041
rect 134154 499967 134210 499976
rect 136284 499905 136312 502860
rect 137388 500070 137416 502860
rect 137376 500064 137428 500070
rect 137376 500006 137428 500012
rect 136270 499896 136326 499905
rect 136270 499831 136326 499840
rect 138492 499769 138520 502860
rect 139504 499934 139532 502860
rect 140608 500002 140636 502860
rect 140596 499996 140648 500002
rect 140596 499938 140648 499944
rect 139492 499928 139544 499934
rect 139492 499870 139544 499876
rect 141712 499866 141740 502860
rect 142066 500848 142122 500857
rect 142066 500783 142122 500792
rect 141700 499860 141752 499866
rect 141700 499802 141752 499808
rect 138478 499760 138534 499769
rect 138478 499695 138534 499704
rect 142080 499633 142108 500783
rect 142816 499798 142844 502860
rect 142804 499792 142856 499798
rect 142804 499734 142856 499740
rect 143828 499730 143856 502860
rect 144642 500848 144698 500857
rect 144642 500783 144698 500792
rect 143816 499724 143868 499730
rect 143816 499666 143868 499672
rect 144656 499633 144684 500783
rect 132590 499624 132646 499633
rect 132590 499559 132646 499568
rect 142066 499624 142122 499633
rect 142066 499559 142122 499568
rect 144642 499624 144698 499633
rect 144932 499594 144960 502860
rect 146036 500721 146064 502860
rect 147048 500857 147076 502860
rect 148152 500857 148180 502860
rect 149256 500857 149284 502860
rect 150360 500857 150388 502860
rect 151372 500857 151400 502860
rect 152476 500857 152504 502860
rect 153212 502846 153594 502874
rect 154592 502846 154698 502874
rect 154960 502846 155710 502874
rect 155972 502846 156814 502874
rect 157352 502846 157918 502874
rect 158824 502846 158930 502874
rect 159744 502846 160034 502874
rect 160112 502846 161138 502874
rect 161492 502846 162242 502874
rect 162872 502846 163254 502874
rect 147034 500848 147090 500857
rect 147034 500783 147090 500792
rect 148138 500848 148194 500857
rect 148138 500783 148194 500792
rect 149242 500848 149298 500857
rect 149242 500783 149298 500792
rect 150346 500848 150402 500857
rect 150346 500783 150402 500792
rect 151358 500848 151414 500857
rect 151358 500783 151414 500792
rect 152462 500848 152518 500857
rect 152462 500783 152518 500792
rect 151912 500744 151964 500750
rect 146022 500712 146078 500721
rect 151912 500686 151964 500692
rect 146022 500647 146078 500656
rect 144642 499559 144698 499568
rect 144920 499588 144972 499594
rect 144920 499530 144972 499536
rect 132500 497480 132552 497486
rect 132500 497422 132552 497428
rect 124220 493332 124272 493338
rect 124220 493274 124272 493280
rect 117136 491972 117188 491978
rect 117136 491914 117188 491920
rect 115388 488708 115440 488714
rect 115388 488650 115440 488656
rect 113192 486934 113574 486962
rect 115400 486948 115428 488650
rect 117148 486948 117176 491914
rect 120724 490612 120776 490618
rect 120724 490554 120776 490560
rect 118976 488776 119028 488782
rect 118976 488718 119028 488724
rect 118988 486948 119016 488718
rect 120736 486948 120764 490554
rect 122564 488844 122616 488850
rect 122564 488786 122616 488792
rect 122576 486948 122604 488786
rect 124232 486962 124260 493274
rect 135076 489864 135128 489870
rect 135076 489806 135128 489812
rect 129740 489796 129792 489802
rect 129740 489738 129792 489744
rect 126152 488980 126204 488986
rect 126152 488922 126204 488928
rect 124232 486934 124338 486962
rect 126164 486948 126192 488922
rect 127900 488912 127952 488918
rect 127900 488854 127952 488860
rect 127912 486948 127940 488854
rect 129752 486948 129780 489738
rect 133328 489116 133380 489122
rect 133328 489058 133380 489064
rect 131488 489048 131540 489054
rect 131488 488990 131540 488996
rect 131500 486948 131528 488990
rect 133340 486948 133368 489058
rect 135088 486948 135116 489806
rect 136916 489728 136968 489734
rect 136916 489670 136968 489676
rect 136928 486948 136956 489670
rect 140504 489660 140556 489666
rect 140504 489602 140556 489608
rect 138664 489592 138716 489598
rect 138664 489534 138716 489540
rect 138676 486948 138704 489534
rect 140516 486948 140544 489602
rect 145840 489524 145892 489530
rect 145840 489466 145892 489472
rect 144092 489456 144144 489462
rect 144092 489398 144144 489404
rect 142252 489388 142304 489394
rect 142252 489330 142304 489336
rect 142264 486948 142292 489330
rect 144104 486948 144132 489398
rect 145852 486948 145880 489466
rect 149428 489320 149480 489326
rect 149428 489262 149480 489268
rect 147680 489184 147732 489190
rect 147680 489126 147732 489132
rect 147692 486948 147720 489126
rect 149440 486948 149468 489262
rect 151268 489252 151320 489258
rect 151268 489194 151320 489200
rect 151280 486948 151308 489194
rect 102152 486798 102902 486826
rect 151924 486577 151952 500686
rect 152004 500540 152056 500546
rect 152004 500482 152056 500488
rect 151910 486568 151966 486577
rect 151910 486503 151966 486512
rect 24124 486464 24176 486470
rect 152016 486441 152044 500482
rect 153108 500268 153160 500274
rect 153108 500210 153160 500216
rect 153014 489152 153070 489161
rect 153014 489087 153070 489096
rect 153028 486948 153056 489087
rect 24124 486406 24176 486412
rect 152002 486432 152058 486441
rect 152002 486367 152058 486376
rect 143448 401600 143500 401606
rect 121366 401568 121422 401577
rect 143448 401542 143500 401548
rect 121366 401503 121422 401512
rect 142068 401532 142120 401538
rect 115754 401432 115810 401441
rect 115754 401367 115810 401376
rect 114466 401296 114522 401305
rect 114466 401231 114522 401240
rect 111706 401024 111762 401033
rect 111706 400959 111762 400968
rect 111614 400888 111670 400897
rect 111614 400823 111670 400832
rect 77944 396636 77996 396642
rect 77944 396578 77996 396584
rect 77956 363769 77984 396578
rect 77942 363760 77998 363769
rect 77942 363695 77998 363704
rect 21362 357640 21418 357649
rect 21362 357575 21418 357584
rect 20332 357054 20668 357082
rect 20976 357054 21312 357082
rect 20640 353326 20668 357054
rect 21284 353394 21312 357054
rect 21272 353388 21324 353394
rect 21272 353330 21324 353336
rect 20628 353320 20680 353326
rect 20628 353262 20680 353268
rect 21376 322794 21404 357575
rect 21712 357054 22048 357082
rect 22448 357054 22784 357082
rect 23184 357054 23428 357082
rect 23920 357054 24256 357082
rect 24564 357054 24808 357082
rect 25300 357054 25636 357082
rect 26036 357054 26188 357082
rect 26772 357054 27108 357082
rect 22020 353462 22048 357054
rect 22008 353456 22060 353462
rect 22008 353398 22060 353404
rect 22756 353326 22784 357054
rect 23400 353394 23428 357054
rect 24228 353462 24256 357054
rect 24780 353530 24808 357054
rect 25608 354142 25636 357054
rect 25596 354136 25648 354142
rect 25596 354078 25648 354084
rect 26160 354074 26188 357054
rect 26148 354068 26200 354074
rect 26148 354010 26200 354016
rect 27080 353598 27108 357054
rect 27494 356810 27522 357068
rect 28152 357054 28488 357082
rect 27494 356782 27568 356810
rect 27068 353592 27120 353598
rect 27068 353534 27120 353540
rect 24768 353524 24820 353530
rect 24768 353466 24820 353472
rect 23940 353456 23992 353462
rect 23940 353398 23992 353404
rect 24216 353456 24268 353462
rect 24216 353398 24268 353404
rect 27068 353456 27120 353462
rect 27068 353398 27120 353404
rect 22836 353388 22888 353394
rect 22836 353330 22888 353336
rect 23388 353388 23440 353394
rect 23388 353330 23440 353336
rect 22192 353320 22244 353326
rect 22192 353262 22244 353268
rect 22744 353320 22796 353326
rect 22744 353262 22796 353268
rect 22204 348786 22232 353262
rect 22848 348922 22876 353330
rect 23952 348922 23980 353398
rect 26240 353388 26292 353394
rect 26240 353330 26292 353336
rect 25044 353320 25096 353326
rect 25044 353262 25096 353268
rect 25056 348922 25084 353262
rect 26252 348922 26280 353330
rect 27080 348922 27108 353398
rect 27540 353326 27568 356782
rect 28172 353524 28224 353530
rect 28172 353466 28224 353472
rect 27528 353320 27580 353326
rect 27528 353262 27580 353268
rect 28184 348922 28212 353466
rect 28460 353394 28488 357054
rect 28874 356810 28902 357068
rect 29624 357054 29960 357082
rect 28874 356782 28948 356810
rect 28920 353666 28948 356782
rect 29932 354550 29960 357054
rect 30300 357054 30360 357082
rect 31096 357054 31432 357082
rect 29920 354544 29972 354550
rect 29920 354486 29972 354492
rect 29276 354136 29328 354142
rect 29276 354078 29328 354084
rect 28908 353660 28960 353666
rect 28908 353602 28960 353608
rect 28448 353388 28500 353394
rect 28448 353330 28500 353336
rect 29288 348922 29316 354078
rect 30300 353734 30328 357054
rect 30380 354068 30432 354074
rect 30380 354010 30432 354016
rect 30288 353728 30340 353734
rect 30288 353670 30340 353676
rect 30392 348922 30420 354010
rect 31404 353462 31432 357054
rect 31680 357054 31740 357082
rect 32476 357054 32812 357082
rect 33212 357054 33456 357082
rect 33948 357054 34284 357082
rect 34684 357054 35020 357082
rect 35328 357054 35664 357082
rect 36064 357054 36400 357082
rect 36800 357054 37136 357082
rect 37536 357054 37872 357082
rect 38272 357054 38424 357082
rect 39008 357054 39344 357082
rect 39652 357054 39988 357082
rect 40388 357054 40724 357082
rect 41124 357054 41276 357082
rect 41860 357054 42196 357082
rect 42596 357054 42748 357082
rect 43240 357054 43576 357082
rect 43976 357054 44128 357082
rect 44712 357054 45048 357082
rect 31680 353530 31708 357054
rect 32784 354142 32812 357054
rect 32772 354136 32824 354142
rect 32772 354078 32824 354084
rect 33428 353870 33456 357054
rect 34256 354074 34284 357054
rect 34992 354482 35020 357054
rect 34980 354476 35032 354482
rect 34980 354418 35032 354424
rect 35636 354414 35664 357054
rect 35808 354544 35860 354550
rect 35808 354486 35860 354492
rect 35624 354408 35676 354414
rect 35624 354350 35676 354356
rect 34244 354068 34296 354074
rect 34244 354010 34296 354016
rect 33416 353864 33468 353870
rect 33416 353806 33468 353812
rect 34520 353728 34572 353734
rect 34520 353670 34572 353676
rect 34428 353660 34480 353666
rect 34428 353602 34480 353608
rect 31852 353592 31904 353598
rect 31852 353534 31904 353540
rect 31668 353524 31720 353530
rect 31668 353466 31720 353472
rect 31392 353456 31444 353462
rect 31392 353398 31444 353404
rect 22848 348894 23138 348922
rect 23952 348894 24242 348922
rect 25056 348894 25346 348922
rect 26252 348894 26358 348922
rect 27080 348894 27462 348922
rect 28184 348894 28566 348922
rect 29288 348894 29670 348922
rect 30392 348894 30682 348922
rect 31864 348786 31892 353534
rect 33508 353388 33560 353394
rect 33508 353330 33560 353336
rect 32588 353320 32640 353326
rect 32588 353262 32640 353268
rect 32600 348922 32628 353262
rect 33520 348922 33548 353330
rect 34440 350554 34468 353602
rect 34532 350810 34560 353670
rect 34520 350804 34572 350810
rect 34520 350746 34572 350752
rect 35820 350554 35848 354486
rect 36372 353394 36400 357054
rect 37108 353734 37136 357054
rect 37096 353728 37148 353734
rect 37096 353670 37148 353676
rect 37188 353524 37240 353530
rect 37188 353466 37240 353472
rect 37096 353456 37148 353462
rect 37096 353398 37148 353404
rect 36360 353388 36412 353394
rect 36360 353330 36412 353336
rect 37108 350810 37136 353398
rect 37200 351898 37228 353466
rect 37844 353326 37872 357054
rect 38396 354346 38424 357054
rect 38384 354340 38436 354346
rect 38384 354282 38436 354288
rect 38200 354136 38252 354142
rect 38200 354078 38252 354084
rect 37832 353320 37884 353326
rect 37832 353262 37884 353268
rect 37188 351892 37240 351898
rect 37188 351834 37240 351840
rect 38212 351150 38240 354078
rect 39212 354068 39264 354074
rect 39212 354010 39264 354016
rect 38660 353864 38712 353870
rect 38660 353806 38712 353812
rect 38672 351218 38700 353806
rect 39028 351892 39080 351898
rect 39028 351834 39080 351840
rect 38660 351212 38712 351218
rect 38660 351154 38712 351160
rect 38200 351144 38252 351150
rect 38200 351086 38252 351092
rect 36820 350804 36872 350810
rect 36820 350746 36872 350752
rect 37096 350804 37148 350810
rect 37096 350746 37148 350752
rect 37924 350804 37976 350810
rect 37924 350746 37976 350752
rect 34440 350526 34560 350554
rect 35820 350526 35940 350554
rect 34532 348922 34560 350526
rect 35912 348922 35940 350526
rect 36832 348922 36860 350746
rect 37936 348922 37964 350746
rect 39040 348922 39068 351834
rect 39224 351354 39252 354010
rect 39316 353938 39344 357054
rect 39960 354278 39988 357054
rect 40040 354476 40092 354482
rect 40040 354418 40092 354424
rect 39948 354272 40000 354278
rect 39948 354214 40000 354220
rect 39304 353932 39356 353938
rect 39304 353874 39356 353880
rect 40052 351422 40080 354418
rect 40224 354408 40276 354414
rect 40224 354350 40276 354356
rect 40040 351416 40092 351422
rect 40040 351358 40092 351364
rect 39212 351348 39264 351354
rect 39212 351290 39264 351296
rect 40236 351286 40264 354350
rect 40696 353598 40724 357054
rect 41248 354210 41276 357054
rect 41236 354204 41288 354210
rect 41236 354146 41288 354152
rect 42168 353666 42196 357054
rect 42720 354142 42748 357054
rect 42708 354136 42760 354142
rect 42708 354078 42760 354084
rect 43548 353734 43576 357054
rect 44100 354006 44128 357054
rect 45020 354074 45048 357054
rect 45434 356810 45462 357068
rect 46184 357054 46520 357082
rect 45434 356782 45508 356810
rect 45480 354550 45508 356782
rect 45468 354544 45520 354550
rect 45468 354486 45520 354492
rect 46492 354414 46520 357054
rect 46814 356810 46842 357068
rect 47564 357054 47900 357082
rect 46814 356782 46888 356810
rect 46860 354686 46888 356782
rect 46848 354680 46900 354686
rect 46848 354622 46900 354628
rect 47872 354482 47900 357054
rect 48240 357054 48300 357082
rect 49036 357054 49372 357082
rect 49772 357054 50108 357082
rect 50416 357054 50752 357082
rect 51152 357054 51488 357082
rect 51888 357054 52224 357082
rect 52624 357054 52960 357082
rect 53360 357054 53696 357082
rect 54004 357054 54340 357082
rect 54740 357054 55076 357082
rect 55476 357054 55812 357082
rect 56212 357054 56548 357082
rect 56948 357054 57284 357082
rect 57684 357054 57836 357082
rect 58328 357054 58664 357082
rect 59064 357054 59308 357082
rect 59800 357054 60136 357082
rect 60536 357054 60688 357082
rect 61272 357054 61608 357082
rect 61916 357054 62068 357082
rect 62652 357054 62988 357082
rect 48240 354634 48268 357054
rect 48240 354618 48360 354634
rect 48240 354612 48372 354618
rect 48240 354606 48320 354612
rect 48320 354554 48372 354560
rect 47860 354476 47912 354482
rect 47860 354418 47912 354424
rect 46480 354408 46532 354414
rect 46480 354350 46532 354356
rect 49344 354346 49372 357054
rect 48596 354340 48648 354346
rect 48596 354282 48648 354288
rect 49332 354340 49384 354346
rect 49332 354282 49384 354288
rect 45008 354068 45060 354074
rect 45008 354010 45060 354016
rect 44088 354000 44140 354006
rect 44088 353942 44140 353948
rect 42248 353728 42300 353734
rect 42248 353670 42300 353676
rect 43536 353728 43588 353734
rect 43536 353670 43588 353676
rect 42156 353660 42208 353666
rect 42156 353602 42208 353608
rect 40684 353592 40736 353598
rect 40684 353534 40736 353540
rect 41604 353388 41656 353394
rect 41604 353330 41656 353336
rect 40224 351280 40276 351286
rect 40224 351222 40276 351228
rect 41616 351218 41644 353330
rect 42260 351354 42288 353670
rect 42800 353320 42852 353326
rect 42800 353262 42852 353268
rect 42812 351694 42840 353262
rect 42800 351688 42852 351694
rect 42800 351630 42852 351636
rect 47676 351688 47728 351694
rect 47676 351630 47728 351636
rect 43260 351416 43312 351422
rect 43260 351358 43312 351364
rect 42156 351348 42208 351354
rect 42156 351290 42208 351296
rect 42248 351348 42300 351354
rect 42248 351290 42300 351296
rect 41512 351212 41564 351218
rect 41512 351154 41564 351160
rect 41604 351212 41656 351218
rect 41604 351154 41656 351160
rect 40132 351144 40184 351150
rect 40132 351086 40184 351092
rect 40144 348922 40172 351086
rect 32600 348894 32890 348922
rect 33520 348894 33902 348922
rect 34532 348894 35006 348922
rect 35912 348894 36110 348922
rect 36832 348894 37214 348922
rect 37936 348894 38226 348922
rect 39040 348894 39330 348922
rect 40144 348894 40434 348922
rect 41524 348786 41552 351154
rect 42168 348922 42196 351290
rect 43272 348922 43300 351358
rect 46572 351348 46624 351354
rect 46572 351290 46624 351296
rect 44364 351280 44416 351286
rect 44364 351222 44416 351228
rect 44376 348922 44404 351222
rect 45652 351212 45704 351218
rect 45652 351154 45704 351160
rect 45664 348922 45692 351154
rect 46584 348922 46612 351290
rect 47688 348922 47716 351630
rect 48608 348922 48636 354282
rect 49700 353932 49752 353938
rect 49700 353874 49752 353880
rect 49712 348922 49740 353874
rect 50080 353530 50108 357054
rect 50724 353938 50752 357054
rect 50988 354272 51040 354278
rect 50988 354214 51040 354220
rect 50712 353932 50764 353938
rect 50712 353874 50764 353880
rect 50068 353524 50120 353530
rect 50068 353466 50120 353472
rect 51000 351778 51028 354214
rect 51460 353870 51488 357054
rect 51448 353864 51500 353870
rect 51448 353806 51500 353812
rect 51908 353592 51960 353598
rect 51908 353534 51960 353540
rect 51000 351750 51120 351778
rect 51092 348922 51120 351750
rect 51920 348922 51948 353534
rect 52196 351354 52224 357054
rect 52932 354278 52960 357054
rect 52920 354272 52972 354278
rect 52920 354214 52972 354220
rect 53012 354204 53064 354210
rect 53012 354146 53064 354152
rect 52184 351348 52236 351354
rect 52184 351290 52236 351296
rect 53024 348922 53052 354146
rect 53668 351286 53696 357054
rect 54116 353660 54168 353666
rect 54116 353602 54168 353608
rect 53656 351280 53708 351286
rect 53656 351222 53708 351228
rect 54128 348922 54156 353602
rect 54312 353326 54340 357054
rect 54300 353320 54352 353326
rect 54300 353262 54352 353268
rect 55048 351218 55076 357054
rect 55784 354210 55812 357054
rect 55772 354204 55824 354210
rect 55772 354146 55824 354152
rect 55128 354136 55180 354142
rect 55128 354078 55180 354084
rect 55140 351234 55168 354078
rect 56140 353728 56192 353734
rect 56140 353670 56192 353676
rect 55036 351212 55088 351218
rect 55140 351206 55260 351234
rect 55036 351154 55088 351160
rect 55232 348922 55260 351206
rect 56152 348922 56180 353670
rect 56520 350606 56548 357054
rect 57256 354090 57284 357054
rect 57520 354544 57572 354550
rect 57520 354486 57572 354492
rect 56784 354068 56836 354074
rect 57256 354062 57376 354090
rect 56784 354010 56836 354016
rect 56796 351898 56824 354010
rect 57244 354000 57296 354006
rect 57244 353942 57296 353948
rect 56784 351892 56836 351898
rect 56784 351834 56836 351840
rect 56508 350600 56560 350606
rect 56508 350542 56560 350548
rect 57256 348922 57284 353942
rect 57348 352782 57376 354062
rect 57336 352776 57388 352782
rect 57336 352718 57388 352724
rect 57532 351490 57560 354486
rect 57520 351484 57572 351490
rect 57520 351426 57572 351432
rect 57808 350674 57836 357054
rect 58532 354680 58584 354686
rect 58532 354622 58584 354628
rect 58072 354408 58124 354414
rect 58072 354350 58124 354356
rect 57888 353320 57940 353326
rect 57888 353262 57940 353268
rect 57900 352850 57928 353262
rect 57888 352844 57940 352850
rect 57888 352786 57940 352792
rect 58084 351830 58112 354350
rect 58348 351892 58400 351898
rect 58348 351834 58400 351840
rect 58072 351824 58124 351830
rect 58072 351766 58124 351772
rect 57796 350668 57848 350674
rect 57796 350610 57848 350616
rect 58360 348922 58388 351834
rect 58544 351626 58572 354622
rect 58636 354142 58664 357054
rect 58624 354136 58676 354142
rect 58624 354078 58676 354084
rect 58532 351620 58584 351626
rect 58532 351562 58584 351568
rect 59280 350742 59308 357054
rect 59636 354612 59688 354618
rect 59636 354554 59688 354560
rect 59360 354476 59412 354482
rect 59360 354418 59412 354424
rect 59372 351762 59400 354418
rect 59360 351756 59412 351762
rect 59360 351698 59412 351704
rect 59648 351558 59676 354554
rect 60108 352714 60136 357054
rect 60096 352708 60148 352714
rect 60096 352650 60148 352656
rect 59636 351552 59688 351558
rect 59636 351494 59688 351500
rect 59452 351484 59504 351490
rect 59452 351426 59504 351432
rect 59268 350736 59320 350742
rect 59268 350678 59320 350684
rect 59464 348922 59492 351426
rect 60660 350810 60688 357054
rect 61580 354074 61608 357054
rect 61568 354068 61620 354074
rect 61568 354010 61620 354016
rect 60740 351824 60792 351830
rect 60740 351766 60792 351772
rect 60648 350804 60700 350810
rect 60648 350746 60700 350752
rect 60752 348922 60780 351766
rect 61660 351620 61712 351626
rect 61660 351562 61712 351568
rect 61672 348922 61700 351562
rect 62040 350946 62068 357054
rect 62212 353932 62264 353938
rect 62212 353874 62264 353880
rect 62120 353524 62172 353530
rect 62120 353466 62172 353472
rect 62132 351898 62160 353466
rect 62120 351892 62172 351898
rect 62120 351834 62172 351840
rect 62224 351694 62252 353874
rect 62960 352646 62988 357054
rect 63374 356810 63402 357068
rect 64124 357054 64460 357082
rect 63374 356782 63448 356810
rect 62948 352640 63000 352646
rect 62948 352582 63000 352588
rect 62764 351756 62816 351762
rect 62764 351698 62816 351704
rect 62212 351688 62264 351694
rect 62212 351630 62264 351636
rect 62028 350940 62080 350946
rect 62028 350882 62080 350888
rect 62776 348922 62804 351698
rect 63420 350878 63448 356782
rect 64432 354006 64460 357054
rect 64800 357054 64860 357082
rect 65504 357054 65840 357082
rect 64420 354000 64472 354006
rect 64420 353942 64472 353948
rect 63500 353864 63552 353870
rect 63500 353806 63552 353812
rect 63512 351422 63540 353806
rect 63684 351552 63736 351558
rect 63684 351494 63736 351500
rect 63500 351416 63552 351422
rect 63500 351358 63552 351364
rect 63408 350872 63460 350878
rect 63408 350814 63460 350820
rect 63696 348922 63724 351494
rect 64800 351150 64828 357054
rect 64972 354340 65024 354346
rect 64972 354282 65024 354288
rect 64788 351144 64840 351150
rect 64788 351086 64840 351092
rect 64984 348922 65012 354282
rect 65812 352578 65840 357054
rect 66180 357054 66240 357082
rect 66976 357054 67312 357082
rect 67712 357054 68048 357082
rect 68448 357054 68784 357082
rect 69092 357054 69428 357082
rect 69828 357054 70164 357082
rect 70564 357054 70900 357082
rect 71300 357054 71636 357082
rect 72036 357054 72372 357082
rect 72680 357054 73016 357082
rect 73416 357054 73752 357082
rect 74152 357054 74488 357082
rect 74888 357054 75224 357082
rect 75624 357054 75868 357082
rect 65800 352572 65852 352578
rect 65800 352514 65852 352520
rect 66180 351082 66208 357054
rect 66352 351892 66404 351898
rect 66352 351834 66404 351840
rect 66168 351076 66220 351082
rect 66168 351018 66220 351024
rect 42168 348894 42550 348922
rect 43272 348894 43654 348922
rect 44376 348894 44758 348922
rect 45664 348894 45770 348922
rect 46584 348894 46874 348922
rect 47688 348894 47978 348922
rect 48608 348894 48990 348922
rect 49712 348894 50094 348922
rect 51092 348894 51198 348922
rect 51920 348894 52302 348922
rect 53024 348894 53314 348922
rect 54128 348894 54418 348922
rect 55232 348894 55522 348922
rect 56152 348894 56534 348922
rect 57256 348894 57638 348922
rect 58360 348894 58742 348922
rect 59464 348894 59846 348922
rect 60752 348894 60858 348922
rect 61672 348894 61962 348922
rect 62776 348894 63066 348922
rect 63696 348894 64078 348922
rect 64984 348894 65182 348922
rect 66364 348786 66392 351834
rect 66996 351688 67048 351694
rect 66996 351630 67048 351636
rect 67008 348922 67036 351630
rect 67284 351014 67312 357054
rect 68020 351898 68048 357054
rect 68008 351892 68060 351898
rect 68008 351834 68060 351840
rect 68756 351830 68784 357054
rect 68744 351824 68796 351830
rect 68744 351766 68796 351772
rect 69400 351626 69428 357054
rect 70136 351762 70164 357054
rect 70400 354272 70452 354278
rect 70400 354214 70452 354220
rect 70124 351756 70176 351762
rect 70124 351698 70176 351704
rect 69388 351620 69440 351626
rect 69388 351562 69440 351568
rect 68100 351416 68152 351422
rect 68100 351358 68152 351364
rect 67272 351008 67324 351014
rect 67272 350950 67324 350956
rect 68112 348922 68140 351358
rect 69204 351348 69256 351354
rect 69204 351290 69256 351296
rect 69216 348922 69244 351290
rect 70412 348922 70440 354214
rect 70872 351694 70900 357054
rect 70860 351688 70912 351694
rect 70860 351630 70912 351636
rect 71608 351490 71636 357054
rect 71596 351484 71648 351490
rect 71596 351426 71648 351432
rect 72344 351422 72372 357054
rect 72424 352844 72476 352850
rect 72424 352786 72476 352792
rect 72332 351416 72384 351422
rect 72332 351358 72384 351364
rect 71228 351280 71280 351286
rect 71228 351222 71280 351228
rect 71240 348922 71268 351222
rect 72436 348922 72464 352786
rect 72988 351354 73016 357054
rect 73724 351558 73752 357054
rect 73712 351552 73764 351558
rect 73712 351494 73764 351500
rect 72976 351348 73028 351354
rect 72976 351290 73028 351296
rect 74460 351218 74488 357054
rect 74724 354204 74776 354210
rect 74724 354146 74776 354152
rect 73436 351212 73488 351218
rect 73436 351154 73488 351160
rect 74448 351212 74500 351218
rect 74448 351154 74500 351160
rect 73448 348922 73476 351154
rect 74736 348922 74764 354146
rect 75196 351286 75224 357054
rect 75184 351280 75236 351286
rect 75184 351222 75236 351228
rect 75840 351121 75868 357054
rect 78772 354136 78824 354142
rect 78772 354078 78824 354084
rect 76748 352776 76800 352782
rect 76748 352718 76800 352724
rect 75826 351112 75882 351121
rect 75826 351047 75882 351056
rect 76012 350600 76064 350606
rect 76012 350542 76064 350548
rect 67008 348894 67390 348922
rect 68112 348894 68402 348922
rect 69216 348894 69506 348922
rect 70412 348894 70610 348922
rect 71240 348894 71622 348922
rect 72436 348894 72726 348922
rect 73448 348894 73830 348922
rect 74736 348894 74934 348922
rect 76024 348786 76052 350542
rect 76760 348922 76788 352718
rect 77852 350668 77904 350674
rect 77852 350610 77904 350616
rect 77864 348922 77892 350610
rect 78784 348922 78812 354078
rect 83188 354068 83240 354074
rect 83188 354010 83240 354016
rect 80980 352708 81032 352714
rect 80980 352650 81032 352656
rect 80060 350736 80112 350742
rect 80060 350678 80112 350684
rect 80072 348922 80100 350678
rect 80992 348922 81020 352650
rect 82084 350804 82136 350810
rect 82084 350746 82136 350752
rect 82096 348922 82124 350746
rect 83200 348922 83228 354010
rect 87420 354000 87472 354006
rect 87420 353942 87472 353948
rect 85580 352640 85632 352646
rect 85580 352582 85632 352588
rect 84384 350940 84436 350946
rect 84384 350882 84436 350888
rect 84396 348922 84424 350882
rect 85592 348922 85620 352582
rect 86316 350872 86368 350878
rect 86316 350814 86368 350820
rect 86328 348922 86356 350814
rect 87432 348922 87460 353942
rect 89720 352572 89772 352578
rect 89720 352514 89772 352520
rect 88524 351144 88576 351150
rect 88524 351086 88576 351092
rect 88536 348922 88564 351086
rect 89732 348922 89760 352514
rect 92940 351892 92992 351898
rect 92940 351834 92992 351840
rect 90732 351076 90784 351082
rect 90732 351018 90784 351024
rect 90744 348922 90772 351018
rect 91836 351008 91888 351014
rect 91836 350950 91888 350956
rect 91848 348922 91876 350950
rect 92952 348922 92980 351834
rect 94044 351824 94096 351830
rect 94044 351766 94096 351772
rect 94056 348922 94084 351766
rect 96068 351756 96120 351762
rect 96068 351698 96120 351704
rect 95240 351620 95292 351626
rect 95240 351562 95292 351568
rect 95252 348922 95280 351562
rect 96080 348922 96108 351698
rect 97172 351688 97224 351694
rect 97172 351630 97224 351636
rect 97184 348922 97212 351630
rect 101404 351552 101456 351558
rect 101404 351494 101456 351500
rect 109590 351520 109646 351529
rect 98276 351484 98328 351490
rect 98276 351426 98328 351432
rect 98288 348922 98316 351426
rect 99380 351416 99432 351422
rect 99380 351358 99432 351364
rect 99392 348922 99420 351358
rect 100852 351348 100904 351354
rect 100852 351290 100904 351296
rect 76760 348894 77050 348922
rect 77864 348894 78154 348922
rect 78784 348894 79166 348922
rect 80072 348894 80270 348922
rect 80992 348894 81374 348922
rect 82096 348894 82478 348922
rect 83200 348894 83490 348922
rect 84396 348894 84594 348922
rect 85592 348894 85698 348922
rect 86328 348894 86710 348922
rect 87432 348894 87814 348922
rect 88536 348894 88918 348922
rect 89732 348894 90022 348922
rect 90744 348894 91034 348922
rect 91848 348894 92138 348922
rect 92952 348894 93242 348922
rect 94056 348894 94254 348922
rect 95252 348894 95358 348922
rect 96080 348894 96462 348922
rect 97184 348894 97566 348922
rect 98288 348894 98578 348922
rect 99392 348894 99682 348922
rect 100864 348786 100892 351290
rect 101416 348922 101444 351494
rect 109590 351455 109646 351464
rect 107566 351384 107622 351393
rect 107566 351319 107622 351328
rect 103704 351280 103756 351286
rect 103704 351222 103756 351228
rect 102508 351212 102560 351218
rect 102508 351154 102560 351160
rect 102520 348922 102548 351154
rect 103716 348922 103744 351222
rect 104898 351112 104954 351121
rect 104898 351047 104954 351056
rect 106186 351112 106242 351121
rect 106186 351047 106242 351056
rect 104912 348922 104940 351047
rect 101416 348894 101798 348922
rect 102520 348894 102902 348922
rect 103716 348894 104006 348922
rect 104912 348894 105110 348922
rect 106200 348786 106228 351047
rect 107580 348786 107608 351319
rect 108670 351248 108726 351257
rect 108670 351183 108726 351192
rect 108684 348786 108712 351183
rect 109604 348786 109632 351455
rect 110696 351008 110748 351014
rect 110696 350950 110748 350956
rect 110708 348786 110736 350950
rect 111628 348786 111656 400823
rect 111720 351014 111748 400959
rect 112902 351656 112958 351665
rect 112902 351591 112958 351600
rect 111708 351008 111760 351014
rect 111708 350950 111760 350956
rect 112916 348786 112944 351591
rect 114480 351490 114508 401231
rect 115768 351490 115796 401367
rect 115846 401160 115902 401169
rect 115846 401095 115902 401104
rect 114008 351484 114060 351490
rect 114008 351426 114060 351432
rect 114468 351484 114520 351490
rect 114468 351426 114520 351432
rect 115112 351484 115164 351490
rect 115112 351426 115164 351432
rect 115756 351484 115808 351490
rect 115756 351426 115808 351432
rect 114020 348786 114048 351426
rect 115124 348786 115152 351426
rect 115860 349058 115888 401095
rect 121276 400988 121328 400994
rect 121276 400930 121328 400936
rect 118608 400920 118660 400926
rect 118608 400862 118660 400868
rect 118620 351490 118648 400862
rect 119342 351792 119398 351801
rect 119342 351727 119398 351736
rect 118148 351484 118200 351490
rect 118148 351426 118200 351432
rect 118608 351484 118660 351490
rect 118608 351426 118660 351432
rect 117134 350976 117190 350985
rect 117134 350911 117190 350920
rect 115768 349030 115888 349058
rect 115768 348922 115796 349030
rect 115768 348894 115874 348922
rect 117148 348786 117176 350911
rect 118160 348786 118188 351426
rect 119356 348786 119384 351727
rect 120448 350872 120500 350878
rect 120448 350814 120500 350820
rect 120460 348786 120488 350814
rect 121288 348786 121316 400930
rect 121380 350878 121408 401503
rect 142068 401474 142120 401480
rect 140688 401464 140740 401470
rect 140688 401406 140740 401412
rect 140596 401396 140648 401402
rect 140596 401338 140648 401344
rect 137928 401328 137980 401334
rect 137928 401270 137980 401276
rect 136456 401260 136508 401266
rect 136456 401202 136508 401208
rect 133788 401192 133840 401198
rect 133788 401134 133840 401140
rect 132408 401124 132460 401130
rect 132408 401066 132460 401072
rect 128268 401056 128320 401062
rect 128268 400998 128320 401004
rect 122470 351792 122526 351801
rect 122470 351727 122526 351736
rect 121368 350872 121420 350878
rect 121368 350814 121420 350820
rect 122484 348786 122512 351727
rect 125416 351280 125468 351286
rect 125416 351222 125468 351228
rect 123760 351212 123812 351218
rect 123760 351154 123812 351160
rect 123772 348786 123800 351154
rect 124678 350568 124734 350577
rect 124678 350503 124734 350512
rect 124692 348786 124720 350503
rect 125428 348922 125456 351222
rect 126886 350704 126942 350713
rect 126886 350639 126942 350648
rect 125428 348894 125534 348922
rect 126900 348786 126928 350639
rect 22126 348758 22232 348786
rect 31786 348758 31892 348786
rect 41446 348758 41552 348786
rect 66286 348758 66392 348786
rect 75946 348758 76052 348786
rect 100786 348758 100892 348786
rect 106122 348758 106228 348786
rect 107226 348758 107608 348786
rect 108330 348758 108712 348786
rect 109342 348758 109632 348786
rect 110446 348758 110736 348786
rect 111550 348758 111656 348786
rect 112654 348758 112944 348786
rect 113666 348758 114048 348786
rect 114770 348758 115152 348786
rect 116886 348758 117176 348786
rect 117990 348758 118188 348786
rect 119094 348758 119384 348786
rect 120198 348758 120488 348786
rect 121210 348758 121316 348786
rect 122314 348758 122512 348786
rect 123418 348758 123800 348786
rect 124430 348758 124720 348786
rect 126638 348758 126928 348786
rect 128280 348650 128308 400998
rect 130200 351416 130252 351422
rect 130200 351358 130252 351364
rect 129094 350840 129150 350849
rect 129094 350775 129150 350784
rect 129738 350840 129794 350849
rect 129738 350775 129794 350784
rect 129108 348786 129136 350775
rect 129752 350577 129780 350775
rect 129738 350568 129794 350577
rect 129738 350503 129794 350512
rect 130212 348786 130240 351358
rect 131028 351348 131080 351354
rect 131028 351290 131080 351296
rect 131040 348786 131068 351290
rect 132420 348786 132448 401066
rect 133800 351490 133828 401134
rect 135166 400752 135222 400761
rect 135166 400687 135222 400696
rect 133328 351484 133380 351490
rect 133328 351426 133380 351432
rect 133788 351484 133840 351490
rect 133788 351426 133840 351432
rect 133340 348786 133368 351426
rect 135180 350810 135208 400687
rect 136468 350946 136496 401202
rect 136546 400616 136602 400625
rect 136546 400551 136602 400560
rect 135536 350940 135588 350946
rect 135536 350882 135588 350888
rect 136456 350940 136508 350946
rect 136456 350882 136508 350888
rect 134432 350804 134484 350810
rect 134432 350746 134484 350752
rect 135168 350804 135220 350810
rect 135168 350746 135220 350752
rect 134444 348786 134472 350746
rect 135548 348786 135576 350882
rect 136560 348786 136588 400551
rect 137940 348922 137968 401270
rect 139306 400480 139362 400489
rect 139306 400415 139362 400424
rect 139320 351490 139348 400415
rect 138848 351484 138900 351490
rect 138848 351426 138900 351432
rect 139308 351484 139360 351490
rect 139308 351426 139360 351432
rect 137756 348894 137968 348922
rect 137756 348786 137784 348894
rect 138860 348786 138888 351426
rect 139768 350804 139820 350810
rect 139768 350746 139820 350752
rect 139780 348786 139808 350746
rect 140608 349058 140636 401338
rect 140700 350810 140728 401406
rect 140688 350804 140740 350810
rect 140688 350746 140740 350752
rect 140608 349030 140728 349058
rect 140700 348786 140728 349030
rect 142080 348786 142108 401474
rect 143460 351490 143488 401542
rect 153120 400926 153148 500210
rect 153108 400920 153160 400926
rect 153108 400862 153160 400868
rect 144828 400852 144880 400858
rect 144828 400794 144880 400800
rect 143080 351484 143132 351490
rect 143080 351426 143132 351432
rect 143448 351484 143500 351490
rect 143448 351426 143500 351432
rect 143092 348786 143120 351426
rect 144840 350674 144868 400794
rect 146116 400512 146168 400518
rect 146116 400454 146168 400460
rect 146128 351490 146156 400454
rect 146206 400344 146262 400353
rect 146206 400279 146262 400288
rect 145288 351484 145340 351490
rect 145288 351426 145340 351432
rect 146116 351484 146168 351490
rect 146116 351426 146168 351432
rect 144918 350976 144974 350985
rect 144918 350911 144974 350920
rect 144184 350668 144236 350674
rect 144184 350610 144236 350616
rect 144828 350668 144880 350674
rect 144828 350610 144880 350616
rect 144196 348786 144224 350610
rect 144932 350577 144960 350911
rect 144918 350568 144974 350577
rect 144918 350503 144974 350512
rect 145300 348786 145328 351426
rect 145562 351248 145618 351257
rect 145562 351183 145618 351192
rect 145576 350985 145604 351183
rect 145562 350976 145618 350985
rect 145562 350911 145618 350920
rect 146220 348786 146248 400279
rect 146298 351520 146354 351529
rect 146298 351455 146354 351464
rect 146942 351520 146998 351529
rect 146942 351455 146998 351464
rect 148046 351520 148102 351529
rect 148046 351455 148102 351464
rect 149426 351520 149482 351529
rect 149426 351455 149482 351464
rect 150070 351520 150126 351529
rect 150070 351455 150126 351464
rect 151174 351520 151230 351529
rect 151174 351455 151230 351464
rect 152370 351520 152426 351529
rect 152370 351455 152426 351464
rect 146312 351257 146340 351455
rect 146298 351248 146354 351257
rect 146298 351183 146354 351192
rect 146956 348922 146984 351455
rect 148060 348922 148088 351455
rect 146956 348894 147062 348922
rect 148060 348894 148166 348922
rect 149440 348786 149468 351455
rect 150084 348922 150112 351455
rect 151188 348922 151216 351455
rect 152384 348922 152412 351455
rect 153212 348922 153240 502846
rect 153476 500948 153528 500954
rect 153476 500890 153528 500896
rect 153384 500880 153436 500886
rect 153382 500848 153384 500857
rect 153436 500848 153438 500857
rect 153292 500812 153344 500818
rect 153382 500783 153438 500792
rect 153292 500754 153344 500760
rect 153304 351422 153332 500754
rect 153488 500585 153516 500890
rect 154488 500608 154540 500614
rect 153474 500576 153530 500585
rect 154488 500550 154540 500556
rect 153474 500511 153530 500520
rect 153384 500472 153436 500478
rect 153384 500414 153436 500420
rect 153292 351416 153344 351422
rect 153292 351358 153344 351364
rect 153396 351286 153424 500414
rect 153476 500404 153528 500410
rect 153476 500346 153528 500352
rect 153384 351280 153436 351286
rect 153384 351222 153436 351228
rect 153488 351218 153516 500346
rect 153844 500336 153896 500342
rect 153844 500278 153896 500284
rect 153660 499792 153712 499798
rect 153660 499734 153712 499740
rect 153568 499724 153620 499730
rect 153568 499666 153620 499672
rect 153580 400858 153608 499666
rect 153672 401606 153700 499734
rect 153752 499588 153804 499594
rect 153752 499530 153804 499536
rect 153660 401600 153712 401606
rect 153660 401542 153712 401548
rect 153568 400852 153620 400858
rect 153568 400794 153620 400800
rect 153764 400518 153792 499530
rect 153856 400994 153884 500278
rect 154396 500200 154448 500206
rect 154396 500142 154448 500148
rect 154304 500132 154356 500138
rect 154304 500074 154356 500080
rect 154120 500064 154172 500070
rect 154120 500006 154172 500012
rect 154028 499928 154080 499934
rect 154028 499870 154080 499876
rect 153936 499860 153988 499866
rect 153936 499802 153988 499808
rect 153948 401538 153976 499802
rect 153936 401532 153988 401538
rect 153936 401474 153988 401480
rect 154040 401470 154068 499870
rect 154028 401464 154080 401470
rect 154028 401406 154080 401412
rect 154132 401334 154160 500006
rect 154212 499996 154264 500002
rect 154212 499938 154264 499944
rect 154224 401402 154252 499938
rect 154212 401396 154264 401402
rect 154212 401338 154264 401344
rect 154120 401328 154172 401334
rect 154120 401270 154172 401276
rect 154316 401266 154344 500074
rect 154304 401260 154356 401266
rect 154304 401202 154356 401208
rect 154408 401130 154436 500142
rect 154396 401124 154448 401130
rect 154396 401066 154448 401072
rect 154500 401062 154528 500550
rect 154488 401056 154540 401062
rect 154488 400998 154540 401004
rect 153844 400988 153896 400994
rect 153844 400930 153896 400936
rect 153752 400512 153804 400518
rect 153752 400454 153804 400460
rect 153476 351212 153528 351218
rect 153476 351154 153528 351160
rect 154592 348922 154620 502846
rect 154764 500676 154816 500682
rect 154764 500618 154816 500624
rect 154776 351354 154804 500618
rect 154856 497480 154908 497486
rect 154856 497422 154908 497428
rect 154868 401198 154896 497422
rect 154856 401192 154908 401198
rect 154856 401134 154908 401140
rect 154764 351348 154816 351354
rect 154764 351290 154816 351296
rect 154960 348922 154988 502846
rect 155972 351490 156000 502846
rect 156052 486464 156104 486470
rect 156052 486406 156104 486412
rect 156064 465361 156092 486406
rect 156050 465352 156106 465361
rect 156050 465287 156106 465296
rect 155960 351484 156012 351490
rect 155960 351426 156012 351432
rect 156420 351484 156472 351490
rect 156420 351426 156472 351432
rect 156432 348922 156460 351426
rect 157352 348922 157380 502846
rect 158720 501220 158772 501226
rect 158720 501162 158772 501168
rect 158732 350878 158760 501162
rect 158720 350872 158772 350878
rect 158720 350814 158772 350820
rect 158824 348922 158852 502846
rect 159744 501226 159772 502846
rect 159732 501220 159784 501226
rect 159732 501162 159784 501168
rect 160112 351490 160140 502846
rect 161492 351490 161520 502846
rect 160100 351484 160152 351490
rect 160100 351426 160152 351432
rect 160836 351484 160888 351490
rect 160836 351426 160888 351432
rect 161480 351484 161532 351490
rect 161480 351426 161532 351432
rect 161940 351484 161992 351490
rect 161940 351426 161992 351432
rect 159732 350872 159784 350878
rect 159732 350814 159784 350820
rect 159744 348922 159772 350814
rect 160848 348922 160876 351426
rect 161952 348922 161980 351426
rect 162872 348922 162900 502846
rect 164240 501220 164292 501226
rect 164240 501162 164292 501168
rect 164252 350674 164280 501162
rect 164240 350668 164292 350674
rect 164240 350610 164292 350616
rect 164344 349058 164372 502860
rect 165080 502846 165462 502874
rect 165632 502846 166474 502874
rect 167012 502846 167578 502874
rect 168392 502846 168682 502874
rect 165080 501226 165108 502846
rect 165068 501220 165120 501226
rect 165068 501162 165120 501168
rect 165632 351490 165660 502846
rect 165620 351484 165672 351490
rect 165620 351426 165672 351432
rect 166172 351484 166224 351490
rect 166172 351426 166224 351432
rect 165068 350668 165120 350674
rect 165068 350610 165120 350616
rect 164252 349030 164372 349058
rect 164252 348922 164280 349030
rect 165080 348922 165108 350610
rect 166184 348922 166212 351426
rect 150084 348894 150374 348922
rect 151188 348894 151386 348922
rect 152384 348894 152490 348922
rect 153212 348894 153594 348922
rect 154592 348894 154698 348922
rect 154960 348894 155710 348922
rect 156432 348894 156814 348922
rect 157352 348894 157918 348922
rect 158824 348894 158930 348922
rect 159744 348894 160034 348922
rect 160848 348894 161138 348922
rect 161952 348894 162242 348922
rect 162872 348894 163254 348922
rect 164252 348894 164358 348922
rect 165080 348894 165462 348922
rect 166184 348894 166474 348922
rect 128754 348758 129136 348786
rect 129858 348758 130240 348786
rect 130962 348758 131068 348786
rect 131974 348758 132448 348786
rect 133078 348758 133368 348786
rect 134182 348758 134472 348786
rect 135286 348758 135576 348786
rect 136298 348758 136588 348786
rect 137402 348758 137784 348786
rect 138506 348758 138888 348786
rect 139518 348758 139808 348786
rect 140622 348758 140728 348786
rect 141726 348758 142108 348786
rect 142830 348758 143120 348786
rect 143842 348758 144224 348786
rect 144946 348758 145328 348786
rect 146050 348758 146248 348786
rect 149270 348758 149468 348786
rect 167012 348786 167040 502846
rect 168392 348922 168420 502846
rect 169772 349058 169800 502860
rect 169864 502846 170798 502874
rect 171152 502846 171902 502874
rect 172532 502846 173006 502874
rect 169864 351490 169892 502846
rect 171152 351490 171180 502846
rect 169852 351484 169904 351490
rect 169852 351426 169904 351432
rect 170404 351484 170456 351490
rect 170404 351426 170456 351432
rect 171140 351484 171192 351490
rect 171140 351426 171192 351432
rect 171600 351484 171652 351490
rect 171600 351426 171652 351432
rect 169772 349030 169892 349058
rect 168392 348894 168682 348922
rect 169864 348786 169892 349030
rect 170416 348922 170444 351426
rect 171612 348922 171640 351426
rect 172532 348922 172560 502846
rect 173900 501220 173952 501226
rect 173900 501162 173952 501168
rect 173912 351014 173940 501162
rect 173900 351008 173952 351014
rect 173900 350950 173952 350956
rect 174004 349058 174032 502860
rect 174832 502846 175122 502874
rect 175292 502846 176226 502874
rect 176672 502846 177330 502874
rect 178052 502846 178342 502874
rect 179446 502846 179552 502874
rect 174832 501226 174860 502846
rect 174820 501220 174872 501226
rect 174820 501162 174872 501168
rect 175292 351490 175320 502846
rect 176672 351490 176700 502846
rect 175280 351484 175332 351490
rect 175280 351426 175332 351432
rect 175924 351484 175976 351490
rect 175924 351426 175976 351432
rect 176660 351484 176712 351490
rect 176660 351426 176712 351432
rect 177120 351484 177172 351490
rect 177120 351426 177172 351432
rect 174820 351008 174872 351014
rect 174820 350950 174872 350956
rect 173912 349030 174032 349058
rect 173912 348922 173940 349030
rect 174832 348922 174860 350950
rect 175936 348922 175964 351426
rect 177132 348922 177160 351426
rect 178052 348922 178080 502846
rect 170416 348894 170798 348922
rect 171612 348894 171902 348922
rect 172532 348894 173006 348922
rect 173912 348894 174018 348922
rect 174832 348894 175122 348922
rect 175936 348894 176226 348922
rect 177132 348894 177330 348922
rect 178052 348894 178342 348922
rect 179524 348786 179552 502846
rect 179616 502846 180550 502874
rect 180812 502846 181562 502874
rect 182192 502846 182666 502874
rect 183572 502846 183770 502874
rect 184584 502846 184874 502874
rect 184952 502846 185886 502874
rect 186332 502846 186990 502874
rect 187712 502846 188094 502874
rect 179616 351490 179644 502846
rect 180812 351490 180840 502846
rect 179604 351484 179656 351490
rect 179604 351426 179656 351432
rect 180156 351484 180208 351490
rect 180156 351426 180208 351432
rect 180800 351484 180852 351490
rect 180800 351426 180852 351432
rect 181260 351484 181312 351490
rect 181260 351426 181312 351432
rect 180168 348922 180196 351426
rect 181272 348922 181300 351426
rect 182192 349058 182220 502846
rect 182192 349030 182404 349058
rect 182376 348922 182404 349030
rect 183572 348922 183600 502846
rect 184584 501226 184612 502846
rect 183652 501220 183704 501226
rect 183652 501162 183704 501168
rect 184572 501220 184624 501226
rect 184572 501162 184624 501168
rect 183664 499474 183692 501162
rect 183664 499446 183784 499474
rect 183756 489954 183784 499446
rect 183756 489926 183876 489954
rect 183848 480282 183876 489926
rect 183652 480276 183704 480282
rect 183652 480218 183704 480224
rect 183836 480276 183888 480282
rect 183836 480218 183888 480224
rect 183664 480162 183692 480218
rect 183664 480134 183784 480162
rect 183756 470642 183784 480134
rect 183756 470614 183876 470642
rect 183848 460970 183876 470614
rect 183652 460964 183704 460970
rect 183652 460906 183704 460912
rect 183836 460964 183888 460970
rect 183836 460906 183888 460912
rect 183664 460850 183692 460906
rect 183664 460822 183784 460850
rect 183756 451330 183784 460822
rect 183756 451302 183876 451330
rect 183848 441658 183876 451302
rect 183652 441652 183704 441658
rect 183652 441594 183704 441600
rect 183836 441652 183888 441658
rect 183836 441594 183888 441600
rect 183664 441538 183692 441594
rect 183664 441510 183784 441538
rect 183756 432018 183784 441510
rect 183756 431990 183876 432018
rect 183848 422346 183876 431990
rect 183652 422340 183704 422346
rect 183652 422282 183704 422288
rect 183836 422340 183888 422346
rect 183836 422282 183888 422288
rect 183664 422226 183692 422282
rect 183664 422198 183784 422226
rect 183756 412706 183784 422198
rect 183756 412678 183876 412706
rect 183848 403034 183876 412678
rect 183652 403028 183704 403034
rect 183652 402970 183704 402976
rect 183836 403028 183888 403034
rect 183836 402970 183888 402976
rect 183664 402914 183692 402970
rect 183664 402886 183784 402914
rect 183756 393394 183784 402886
rect 183756 393366 183876 393394
rect 183848 383722 183876 393366
rect 183652 383716 183704 383722
rect 183652 383658 183704 383664
rect 183836 383716 183888 383722
rect 183836 383658 183888 383664
rect 183664 383602 183692 383658
rect 183664 383574 183784 383602
rect 183756 374082 183784 383574
rect 183756 374054 183876 374082
rect 183848 364410 183876 374054
rect 183652 364404 183704 364410
rect 183652 364346 183704 364352
rect 183836 364404 183888 364410
rect 183836 364346 183888 364352
rect 183664 354634 183692 364346
rect 183664 354606 183876 354634
rect 183848 351082 183876 354606
rect 184952 351490 184980 502846
rect 185584 485104 185636 485110
rect 185584 485046 185636 485052
rect 185596 450945 185624 485046
rect 185582 450936 185638 450945
rect 185582 450871 185638 450880
rect 184940 351484 184992 351490
rect 184940 351426 184992 351432
rect 185492 351484 185544 351490
rect 185492 351426 185544 351432
rect 183836 351076 183888 351082
rect 183836 351018 183888 351024
rect 184572 351076 184624 351082
rect 184572 351018 184624 351024
rect 184584 348922 184612 351018
rect 185504 348922 185532 351426
rect 186332 349058 186360 502846
rect 186332 349030 186636 349058
rect 186608 348922 186636 349030
rect 187712 348922 187740 502846
rect 189092 500721 189120 502860
rect 190196 500857 190224 502860
rect 191300 500857 191328 502860
rect 190182 500848 190238 500857
rect 190182 500783 190238 500792
rect 191286 500848 191342 500857
rect 191286 500783 191342 500792
rect 189078 500712 189134 500721
rect 189078 500647 189134 500656
rect 192404 500478 192432 502860
rect 187792 500472 187844 500478
rect 187792 500414 187844 500420
rect 192392 500472 192444 500478
rect 192392 500414 192444 500420
rect 187804 358358 187832 500414
rect 193416 500274 193444 502860
rect 187884 500268 187936 500274
rect 187884 500210 187936 500216
rect 193404 500268 193456 500274
rect 193404 500210 193456 500216
rect 187792 358352 187844 358358
rect 187792 358294 187844 358300
rect 187896 358154 187924 500210
rect 194520 500177 194548 502860
rect 195244 500948 195296 500954
rect 195244 500890 195296 500896
rect 194506 500168 194562 500177
rect 194506 500103 194562 500112
rect 191840 500064 191892 500070
rect 191840 500006 191892 500012
rect 190920 494012 190972 494018
rect 190920 493954 190972 493960
rect 189724 493400 189776 493406
rect 189724 493342 189776 493348
rect 188620 493060 188672 493066
rect 188620 493002 188672 493008
rect 188632 491572 188660 493002
rect 189736 491572 189764 493342
rect 190932 491572 190960 493954
rect 191852 491586 191880 500006
rect 191932 499792 191984 499798
rect 191932 499734 191984 499740
rect 191944 493066 191972 499734
rect 193312 493672 193364 493678
rect 193312 493614 193364 493620
rect 191932 493060 191984 493066
rect 191932 493002 191984 493008
rect 191852 491558 192142 491586
rect 193324 491572 193352 493614
rect 194508 493536 194560 493542
rect 194508 493478 194560 493484
rect 194520 491572 194548 493478
rect 195256 493406 195284 500890
rect 195336 500880 195388 500886
rect 195336 500822 195388 500828
rect 195348 494018 195376 500822
rect 195624 500274 195652 502860
rect 196072 500540 196124 500546
rect 196072 500482 196124 500488
rect 195612 500268 195664 500274
rect 195612 500210 195664 500216
rect 195336 494012 195388 494018
rect 195336 493954 195388 493960
rect 196084 493678 196112 500482
rect 196636 499798 196664 502860
rect 197740 500954 197768 502860
rect 197728 500948 197780 500954
rect 197728 500890 197780 500896
rect 198844 500886 198872 502860
rect 198832 500880 198884 500886
rect 198832 500822 198884 500828
rect 197176 500744 197228 500750
rect 197176 500686 197228 500692
rect 196624 499792 196676 499798
rect 196624 499734 196676 499740
rect 196900 494012 196952 494018
rect 196900 493954 196952 493960
rect 196072 493672 196124 493678
rect 196072 493614 196124 493620
rect 195244 493400 195296 493406
rect 195244 493342 195296 493348
rect 195704 493196 195756 493202
rect 195704 493138 195756 493144
rect 195716 491572 195744 493138
rect 196912 491572 196940 493954
rect 197188 493542 197216 500686
rect 199476 500472 199528 500478
rect 199476 500414 199528 500420
rect 199488 494018 199516 500414
rect 199948 500070 199976 502860
rect 200212 500880 200264 500886
rect 200212 500822 200264 500828
rect 199936 500064 199988 500070
rect 199936 500006 199988 500012
rect 199476 494012 199528 494018
rect 199476 493954 199528 493960
rect 200224 493610 200252 500822
rect 200960 500546 200988 502860
rect 201684 500948 201736 500954
rect 201684 500890 201736 500896
rect 201592 500608 201644 500614
rect 201592 500550 201644 500556
rect 200948 500540 201000 500546
rect 200948 500482 201000 500488
rect 200488 494012 200540 494018
rect 200488 493954 200540 493960
rect 198096 493604 198148 493610
rect 198096 493546 198148 493552
rect 200212 493604 200264 493610
rect 200212 493546 200264 493552
rect 197176 493536 197228 493542
rect 197176 493478 197228 493484
rect 198108 491572 198136 493546
rect 199292 493332 199344 493338
rect 199292 493274 199344 493280
rect 199304 491572 199332 493274
rect 200500 491572 200528 493954
rect 201604 493338 201632 500550
rect 201696 494034 201724 500890
rect 202064 500750 202092 502860
rect 203168 500954 203196 502860
rect 203156 500948 203208 500954
rect 203156 500890 203208 500896
rect 202052 500744 202104 500750
rect 202052 500686 202104 500692
rect 204180 500478 204208 502860
rect 204628 500948 204680 500954
rect 204628 500890 204680 500896
rect 204168 500472 204220 500478
rect 204168 500414 204220 500420
rect 203708 499656 203760 499662
rect 203708 499598 203760 499604
rect 201696 494006 201908 494034
rect 203720 494018 203748 499598
rect 201684 493876 201736 493882
rect 201684 493818 201736 493824
rect 201592 493332 201644 493338
rect 201592 493274 201644 493280
rect 201696 491572 201724 493818
rect 201880 493202 201908 494006
rect 203708 494012 203760 494018
rect 203708 493954 203760 493960
rect 204640 493882 204668 500890
rect 205284 500886 205312 502860
rect 205272 500880 205324 500886
rect 205272 500822 205324 500828
rect 205640 500880 205692 500886
rect 205640 500822 205692 500828
rect 205272 494012 205324 494018
rect 205272 493954 205324 493960
rect 204628 493876 204680 493882
rect 204628 493818 204680 493824
rect 204076 493672 204128 493678
rect 204076 493614 204128 493620
rect 202880 493468 202932 493474
rect 202880 493410 202932 493416
rect 201868 493196 201920 493202
rect 201868 493138 201920 493144
rect 202892 491572 202920 493410
rect 204088 491572 204116 493614
rect 205284 491572 205312 493954
rect 205652 493474 205680 500822
rect 206388 500614 206416 502860
rect 206376 500608 206428 500614
rect 206376 500550 206428 500556
rect 206376 499724 206428 499730
rect 206376 499666 206428 499672
rect 206388 493678 206416 499666
rect 207492 499662 207520 502860
rect 208504 500954 208532 502860
rect 208492 500948 208544 500954
rect 208492 500890 208544 500896
rect 209608 500886 209636 502860
rect 209596 500880 209648 500886
rect 209596 500822 209648 500828
rect 209872 500472 209924 500478
rect 209872 500414 209924 500420
rect 209136 500404 209188 500410
rect 209136 500346 209188 500352
rect 207480 499656 207532 499662
rect 207480 499598 207532 499604
rect 207756 499656 207808 499662
rect 207756 499598 207808 499604
rect 207768 494018 207796 499598
rect 207756 494012 207808 494018
rect 207756 493954 207808 493960
rect 209148 493746 209176 500346
rect 206468 493740 206520 493746
rect 206468 493682 206520 493688
rect 209136 493740 209188 493746
rect 209136 493682 209188 493688
rect 206376 493672 206428 493678
rect 206376 493614 206428 493620
rect 205640 493468 205692 493474
rect 205640 493410 205692 493416
rect 206480 491572 206508 493682
rect 209884 493474 209912 500414
rect 210712 499730 210740 502860
rect 211344 500744 211396 500750
rect 211344 500686 211396 500692
rect 210700 499724 210752 499730
rect 210700 499666 210752 499672
rect 210056 493876 210108 493882
rect 210056 493818 210108 493824
rect 207664 493468 207716 493474
rect 207664 493410 207716 493416
rect 209872 493468 209924 493474
rect 209872 493410 209924 493416
rect 207676 491572 207704 493410
rect 208860 493196 208912 493202
rect 208860 493138 208912 493144
rect 208872 491572 208900 493138
rect 210068 491572 210096 493818
rect 211252 493672 211304 493678
rect 211252 493614 211304 493620
rect 211264 491572 211292 493614
rect 211356 493202 211384 500686
rect 211724 499662 211752 502860
rect 212828 500410 212856 502860
rect 213460 500880 213512 500886
rect 213460 500822 213512 500828
rect 212816 500404 212868 500410
rect 212816 500346 212868 500352
rect 211712 499656 211764 499662
rect 211712 499598 211764 499604
rect 213472 493882 213500 500822
rect 213932 500478 213960 502860
rect 214656 500948 214708 500954
rect 214656 500890 214708 500896
rect 213920 500472 213972 500478
rect 213920 500414 213972 500420
rect 213644 494012 213696 494018
rect 213644 493954 213696 493960
rect 213460 493876 213512 493882
rect 213460 493818 213512 493824
rect 212448 493740 212500 493746
rect 212448 493682 212500 493688
rect 211344 493196 211396 493202
rect 211344 493138 211396 493144
rect 212460 491572 212488 493682
rect 213656 491572 213684 493954
rect 214668 493678 214696 500890
rect 214932 500812 214984 500818
rect 214932 500754 214984 500760
rect 214944 493746 214972 500754
rect 215036 500750 215064 502860
rect 216048 500886 216076 502860
rect 217152 500954 217180 502860
rect 217140 500948 217192 500954
rect 217140 500890 217192 500896
rect 216036 500880 216088 500886
rect 216036 500822 216088 500828
rect 218256 500818 218284 502860
rect 218244 500812 218296 500818
rect 218244 500754 218296 500760
rect 215024 500744 215076 500750
rect 215024 500686 215076 500692
rect 219268 500614 219296 502860
rect 215300 500608 215352 500614
rect 215300 500550 215352 500556
rect 219256 500608 219308 500614
rect 219256 500550 219308 500556
rect 219532 500608 219584 500614
rect 219532 500550 219584 500556
rect 215312 494018 215340 500550
rect 218152 500472 218204 500478
rect 218152 500414 218204 500420
rect 216680 499656 216732 499662
rect 216680 499598 216732 499604
rect 215300 494012 215352 494018
rect 215300 493954 215352 493960
rect 216036 494012 216088 494018
rect 216036 493954 216088 493960
rect 214932 493740 214984 493746
rect 214932 493682 214984 493688
rect 214656 493672 214708 493678
rect 214656 493614 214708 493620
rect 214840 493264 214892 493270
rect 214840 493206 214892 493212
rect 214852 491572 214880 493206
rect 216048 491572 216076 493954
rect 216692 493270 216720 499598
rect 218164 494018 218192 500414
rect 218152 494012 218204 494018
rect 218152 493954 218204 493960
rect 218428 493604 218480 493610
rect 218428 493546 218480 493552
rect 217232 493536 217284 493542
rect 217232 493478 217284 493484
rect 216680 493264 216732 493270
rect 216680 493206 216732 493212
rect 217244 491572 217272 493478
rect 218440 491572 218468 493546
rect 219544 493542 219572 500550
rect 220372 499662 220400 502860
rect 221476 500478 221504 502860
rect 222580 500614 222608 502860
rect 223488 500676 223540 500682
rect 223488 500618 223540 500624
rect 222568 500608 222620 500614
rect 222568 500550 222620 500556
rect 221464 500472 221516 500478
rect 221464 500414 221516 500420
rect 220820 500132 220872 500138
rect 220820 500074 220872 500080
rect 220360 499656 220412 499662
rect 220360 499598 220412 499604
rect 219624 493876 219676 493882
rect 219624 493818 219676 493824
rect 219532 493536 219584 493542
rect 219532 493478 219584 493484
rect 219636 491572 219664 493818
rect 220832 493610 220860 500074
rect 223500 493882 223528 500618
rect 223592 500138 223620 502860
rect 224696 500682 224724 502860
rect 225800 500954 225828 502860
rect 224868 500948 224920 500954
rect 224868 500890 224920 500896
rect 225788 500948 225840 500954
rect 225788 500890 225840 500896
rect 224684 500676 224736 500682
rect 224684 500618 224736 500624
rect 224224 500472 224276 500478
rect 224224 500414 224276 500420
rect 223580 500132 223632 500138
rect 223580 500074 223632 500080
rect 223580 499928 223632 499934
rect 223580 499870 223632 499876
rect 223488 493876 223540 493882
rect 223488 493818 223540 493824
rect 222016 493672 222068 493678
rect 222016 493614 222068 493620
rect 220820 493604 220872 493610
rect 220820 493546 220872 493552
rect 220820 493468 220872 493474
rect 220820 493410 220872 493416
rect 220832 491572 220860 493410
rect 222028 491572 222056 493614
rect 223212 492924 223264 492930
rect 223212 492866 223264 492872
rect 223224 491572 223252 492866
rect 223592 492794 223620 499870
rect 224236 493678 224264 500414
rect 224224 493672 224276 493678
rect 224224 493614 224276 493620
rect 224880 493474 224908 500890
rect 226812 500478 226840 502860
rect 226800 500472 226852 500478
rect 226800 500414 226852 500420
rect 226800 493944 226852 493950
rect 226800 493886 226852 493892
rect 225604 493604 225656 493610
rect 225604 493546 225656 493552
rect 224868 493468 224920 493474
rect 224868 493410 224920 493416
rect 223580 492788 223632 492794
rect 223580 492730 223632 492736
rect 224408 492788 224460 492794
rect 224408 492730 224460 492736
rect 224420 491572 224448 492730
rect 225616 491572 225644 493546
rect 226812 491572 226840 493886
rect 227916 492930 227944 502860
rect 229020 499934 229048 502860
rect 230124 500954 230152 502860
rect 229100 500948 229152 500954
rect 229100 500890 229152 500896
rect 230112 500948 230164 500954
rect 230112 500890 230164 500896
rect 230572 500948 230624 500954
rect 230572 500890 230624 500896
rect 229008 499928 229060 499934
rect 229008 499870 229060 499876
rect 229112 499610 229140 500890
rect 229020 499582 229140 499610
rect 230388 499588 230440 499594
rect 229020 493610 229048 499582
rect 230388 499530 230440 499536
rect 230400 493950 230428 499530
rect 230388 493944 230440 493950
rect 230388 493886 230440 493892
rect 229192 493876 229244 493882
rect 229192 493818 229244 493824
rect 229008 493604 229060 493610
rect 229008 493546 229060 493552
rect 227996 493060 228048 493066
rect 227996 493002 228048 493008
rect 227904 492924 227956 492930
rect 227904 492866 227956 492872
rect 228008 491572 228036 493002
rect 229204 491572 229232 493818
rect 230388 493604 230440 493610
rect 230388 493546 230440 493552
rect 230400 491572 230428 493546
rect 230584 493066 230612 500890
rect 231136 499594 231164 502860
rect 232240 500954 232268 502860
rect 233252 502846 233358 502874
rect 232228 500948 232280 500954
rect 232228 500890 232280 500896
rect 233252 500834 233280 502846
rect 233160 500806 233280 500834
rect 233056 499792 233108 499798
rect 233056 499734 233108 499740
rect 231124 499588 231176 499594
rect 231124 499530 231176 499536
rect 231584 494012 231636 494018
rect 231584 493954 231636 493960
rect 230572 493060 230624 493066
rect 230572 493002 230624 493008
rect 231596 491572 231624 493954
rect 232780 493944 232832 493950
rect 232780 493886 232832 493892
rect 232792 491572 232820 493886
rect 233068 493610 233096 499734
rect 233160 493882 233188 500806
rect 234356 499798 234384 502860
rect 235460 500954 235488 502860
rect 236564 500954 236592 502860
rect 237484 502846 237682 502874
rect 237944 502846 238694 502874
rect 238772 502846 239798 502874
rect 240152 502846 240902 502874
rect 241532 502846 241914 502874
rect 234528 500948 234580 500954
rect 234528 500890 234580 500896
rect 235448 500948 235500 500954
rect 235448 500890 235500 500896
rect 235908 500948 235960 500954
rect 235908 500890 235960 500896
rect 236552 500948 236604 500954
rect 236552 500890 236604 500896
rect 234344 499792 234396 499798
rect 234344 499734 234396 499740
rect 234540 494018 234568 500890
rect 234528 494012 234580 494018
rect 234528 493954 234580 493960
rect 235172 494012 235224 494018
rect 235172 493954 235224 493960
rect 233148 493876 233200 493882
rect 233148 493818 233200 493824
rect 233056 493604 233108 493610
rect 233056 493546 233108 493552
rect 233976 493604 234028 493610
rect 233976 493546 234028 493552
rect 233988 491572 234016 493546
rect 235184 491572 235212 493954
rect 235920 493950 235948 500890
rect 237484 500834 237512 502846
rect 237944 501242 237972 502846
rect 237300 500806 237512 500834
rect 237576 501214 237972 501242
rect 235908 493944 235960 493950
rect 235908 493886 235960 493892
rect 236368 493808 236420 493814
rect 236368 493750 236420 493756
rect 236380 491572 236408 493750
rect 237300 493610 237328 500806
rect 237576 494018 237604 501214
rect 237564 494012 237616 494018
rect 237564 493954 237616 493960
rect 237564 493876 237616 493882
rect 237564 493818 237616 493824
rect 237288 493604 237340 493610
rect 237288 493546 237340 493552
rect 237576 491572 237604 493818
rect 238772 493814 238800 502846
rect 240152 493882 240180 502846
rect 241152 494012 241204 494018
rect 241152 493954 241204 493960
rect 240140 493876 240192 493882
rect 240140 493818 240192 493824
rect 238760 493808 238812 493814
rect 238760 493750 238812 493756
rect 239956 493536 240008 493542
rect 239956 493478 240008 493484
rect 238760 493468 238812 493474
rect 238760 493410 238812 493416
rect 238772 491572 238800 493410
rect 239968 491572 239996 493478
rect 241164 491572 241192 493954
rect 241532 493474 241560 502846
rect 243004 500018 243032 502860
rect 242820 499990 243032 500018
rect 243096 502846 244122 502874
rect 244292 502846 245226 502874
rect 245672 502846 246238 502874
rect 247236 502846 247342 502874
rect 242820 493542 242848 499990
rect 243096 494018 243124 502846
rect 243084 494012 243136 494018
rect 243084 493954 243136 493960
rect 242808 493536 242860 493542
rect 242808 493478 242860 493484
rect 241520 493468 241572 493474
rect 241520 493410 241572 493416
rect 243544 493468 243596 493474
rect 243544 493410 243596 493416
rect 242348 493264 242400 493270
rect 242348 493206 242400 493212
rect 242360 491572 242388 493206
rect 243556 491572 243584 493410
rect 244292 493270 244320 502846
rect 245672 493474 245700 502846
rect 247040 499588 247092 499594
rect 247040 499530 247092 499536
rect 245936 494012 245988 494018
rect 245936 493954 245988 493960
rect 245660 493468 245712 493474
rect 245660 493410 245712 493416
rect 244740 493332 244792 493338
rect 244740 493274 244792 493280
rect 244280 493264 244332 493270
rect 244280 493206 244332 493212
rect 244752 491572 244780 493274
rect 245948 491572 245976 493954
rect 247052 491586 247080 499530
rect 247236 493338 247264 502846
rect 248432 494018 248460 502860
rect 249444 499594 249472 502860
rect 249812 502846 250562 502874
rect 251284 502846 251666 502874
rect 249432 499588 249484 499594
rect 249432 499530 249484 499536
rect 248420 494012 248472 494018
rect 248420 493954 248472 493960
rect 249812 493814 249840 502846
rect 251180 500880 251232 500886
rect 251180 500822 251232 500828
rect 248328 493808 248380 493814
rect 248328 493750 248380 493756
rect 249800 493808 249852 493814
rect 249800 493750 249852 493756
rect 247224 493332 247276 493338
rect 247224 493274 247276 493280
rect 247052 491558 247158 491586
rect 248340 491572 248368 493750
rect 249524 493332 249576 493338
rect 249524 493274 249576 493280
rect 249536 491572 249564 493274
rect 250720 492992 250772 492998
rect 250720 492934 250772 492940
rect 250732 491572 250760 492934
rect 251192 491722 251220 500822
rect 251284 493338 251312 502846
rect 252652 499656 252704 499662
rect 252652 499598 252704 499604
rect 251272 493332 251324 493338
rect 251272 493274 251324 493280
rect 251192 491694 251496 491722
rect 251468 491586 251496 491694
rect 252664 491586 252692 499598
rect 252756 492998 252784 502860
rect 253768 500886 253796 502860
rect 253756 500880 253808 500886
rect 253756 500822 253808 500828
rect 253940 500880 253992 500886
rect 253940 500822 253992 500828
rect 252744 492992 252796 492998
rect 252744 492934 252796 492940
rect 253952 491586 253980 500822
rect 254872 499662 254900 502860
rect 255320 500948 255372 500954
rect 255320 500890 255372 500896
rect 254860 499656 254912 499662
rect 254860 499598 254912 499604
rect 255332 491586 255360 500890
rect 255976 500886 256004 502860
rect 256988 500954 257016 502860
rect 256976 500948 257028 500954
rect 256976 500890 257028 500896
rect 255964 500880 256016 500886
rect 255964 500822 256016 500828
rect 258092 499610 258120 502860
rect 256792 499588 256844 499594
rect 256792 499530 256844 499536
rect 258000 499582 258120 499610
rect 259196 499594 259224 502860
rect 259460 500948 259512 500954
rect 259460 500890 259512 500896
rect 259368 499792 259420 499798
rect 259368 499734 259420 499740
rect 259184 499588 259236 499594
rect 256804 494018 256832 499530
rect 256792 494012 256844 494018
rect 256792 493954 256844 493960
rect 257896 494012 257948 494018
rect 257896 493954 257948 493960
rect 256700 493196 256752 493202
rect 256700 493138 256752 493144
rect 251468 491558 251942 491586
rect 252664 491558 253138 491586
rect 253952 491558 254334 491586
rect 255332 491558 255530 491586
rect 256712 491572 256740 493138
rect 257908 491572 257936 493954
rect 258000 493202 258028 499582
rect 259184 499530 259236 499536
rect 257988 493196 258040 493202
rect 257988 493138 258040 493144
rect 259380 491586 259408 499734
rect 259472 494018 259500 500890
rect 260300 499798 260328 502860
rect 261312 500954 261340 502860
rect 261300 500948 261352 500954
rect 261300 500890 261352 500896
rect 262312 500948 262364 500954
rect 262312 500890 262364 500896
rect 260840 500880 260892 500886
rect 260840 500822 260892 500828
rect 260288 499792 260340 499798
rect 260288 499734 260340 499740
rect 259460 494012 259512 494018
rect 259460 493954 259512 493960
rect 260288 494012 260340 494018
rect 260288 493954 260340 493960
rect 259118 491558 259408 491586
rect 260300 491572 260328 493954
rect 260852 491450 260880 500822
rect 262324 491586 262352 500890
rect 262416 500886 262444 502860
rect 263520 500954 263548 502860
rect 263508 500948 263560 500954
rect 263508 500890 263560 500896
rect 262404 500880 262456 500886
rect 262404 500822 262456 500828
rect 264532 499798 264560 502860
rect 264992 502846 265650 502874
rect 266372 502846 266754 502874
rect 263600 499792 263652 499798
rect 263600 499734 263652 499740
rect 264520 499792 264572 499798
rect 264520 499734 264572 499740
rect 263612 491586 263640 499734
rect 264992 491586 265020 502846
rect 266372 500936 266400 502846
rect 266280 500908 266400 500936
rect 262324 491558 262706 491586
rect 263612 491558 263902 491586
rect 264992 491558 265098 491586
rect 266280 491572 266308 500908
rect 267844 499594 267872 502860
rect 268856 500954 268884 502860
rect 269960 500954 269988 502860
rect 270512 502846 271078 502874
rect 271892 502846 272090 502874
rect 267924 500948 267976 500954
rect 267924 500890 267976 500896
rect 268844 500948 268896 500954
rect 268844 500890 268896 500896
rect 269120 500948 269172 500954
rect 269120 500890 269172 500896
rect 269948 500948 270000 500954
rect 269948 500890 270000 500896
rect 266360 499588 266412 499594
rect 266360 499530 266412 499536
rect 267832 499588 267884 499594
rect 267832 499530 267884 499536
rect 266372 494018 266400 499530
rect 267936 495258 267964 500890
rect 267936 495230 268332 495258
rect 266360 494012 266412 494018
rect 266360 493954 266412 493960
rect 267464 494012 267516 494018
rect 267464 493954 267516 493960
rect 267476 491572 267504 493954
rect 268304 491586 268332 495230
rect 269132 494034 269160 500890
rect 270512 494306 270540 502846
rect 270512 494278 270724 494306
rect 269132 494006 269620 494034
rect 269592 491586 269620 494006
rect 270696 491586 270724 494278
rect 271892 491586 271920 502846
rect 273180 499662 273208 502860
rect 274298 502846 274588 502874
rect 271972 499656 272024 499662
rect 271972 499598 272024 499604
rect 273168 499656 273220 499662
rect 273168 499598 273220 499604
rect 271984 492862 272012 499598
rect 274560 493218 274588 502846
rect 274744 502846 275402 502874
rect 276032 502846 276414 502874
rect 277412 502846 277518 502874
rect 274560 493190 274680 493218
rect 271972 492856 272024 492862
rect 271972 492798 272024 492804
rect 273444 492856 273496 492862
rect 273444 492798 273496 492804
rect 268304 491558 268686 491586
rect 269592 491558 269882 491586
rect 270696 491558 271078 491586
rect 271892 491558 272274 491586
rect 273456 491572 273484 492798
rect 274652 491572 274680 493190
rect 274744 491450 274772 502846
rect 276032 491450 276060 502846
rect 277412 491586 277440 502846
rect 278608 499594 278636 502860
rect 277584 499588 277636 499594
rect 277584 499530 277636 499536
rect 278596 499588 278648 499594
rect 278596 499530 278648 499536
rect 277596 493202 277624 499530
rect 277584 493196 277636 493202
rect 277584 493138 277636 493144
rect 279424 493196 279476 493202
rect 279424 493138 279476 493144
rect 277412 491558 278254 491586
rect 279436 491572 279464 493138
rect 260852 491422 261510 491450
rect 274744 491422 275862 491450
rect 276032 491422 277058 491450
rect 279528 463570 279556 552026
rect 280526 528456 280582 528465
rect 280526 528391 280582 528400
rect 280540 518945 280568 528391
rect 280526 518936 280582 518945
rect 280526 518871 280582 518880
rect 281552 515953 281580 569162
rect 281538 515944 281594 515953
rect 281538 515879 281594 515888
rect 279608 500268 279660 500274
rect 279608 500210 279660 500216
rect 279620 471889 279648 500210
rect 280342 495544 280398 495553
rect 280342 495479 280398 495488
rect 280356 489977 280384 495479
rect 280342 489968 280398 489977
rect 280342 489903 280398 489912
rect 280158 480040 280214 480049
rect 280158 479975 280214 479984
rect 279606 471880 279662 471889
rect 279606 471815 279662 471824
rect 280172 470665 280200 479975
rect 280158 470656 280214 470665
rect 280158 470591 280214 470600
rect 279700 463684 279752 463690
rect 279700 463626 279752 463632
rect 279712 463570 279740 463626
rect 279528 463542 279740 463570
rect 280250 451208 280306 451217
rect 280250 451143 280306 451152
rect 280264 445777 280292 451143
rect 280250 445768 280306 445777
rect 280250 445703 280306 445712
rect 280342 439512 280398 439521
rect 280342 439447 280398 439456
rect 280356 434761 280384 439447
rect 280342 434752 280398 434761
rect 280342 434687 280398 434696
rect 281552 430545 281580 515879
rect 281538 430536 281594 430545
rect 281538 430471 281594 430480
rect 281632 421592 281684 421598
rect 281632 421534 281684 421540
rect 281644 421297 281672 421534
rect 281630 421288 281686 421297
rect 281630 421223 281686 421232
rect 191932 358352 191984 358358
rect 191932 358294 191984 358300
rect 187884 358148 187936 358154
rect 188048 358142 188384 358170
rect 189244 358142 189580 358170
rect 187884 358090 187936 358096
rect 188356 354754 188384 358142
rect 189552 354890 189580 358142
rect 190380 358142 190440 358170
rect 191636 358142 191788 358170
rect 189540 354884 189592 354890
rect 189540 354826 189592 354832
rect 190380 354822 190408 358142
rect 191760 355978 191788 358142
rect 191748 355972 191800 355978
rect 191748 355914 191800 355920
rect 190368 354816 190420 354822
rect 190368 354758 190420 354764
rect 188344 354748 188396 354754
rect 188344 354690 188396 354696
rect 189446 351792 189502 351801
rect 189446 351727 189502 351736
rect 191194 351792 191250 351801
rect 191194 351727 191250 351736
rect 180168 348894 180550 348922
rect 181272 348894 181562 348922
rect 182376 348894 182666 348922
rect 183572 348894 183770 348922
rect 184584 348894 184874 348922
rect 185504 348894 185886 348922
rect 186608 348894 186990 348922
rect 187712 348894 188094 348922
rect 189460 348786 189488 351727
rect 189906 351656 189962 351665
rect 189906 351591 189962 351600
rect 189920 348922 189948 351591
rect 191208 348922 191236 351727
rect 191944 349058 191972 358294
rect 245456 358278 245608 358306
rect 192924 358142 193168 358170
rect 193140 355910 193168 358142
rect 193312 358148 193364 358154
rect 194120 358142 194456 358170
rect 195316 358142 195652 358170
rect 196512 358142 196848 358170
rect 197800 358142 198136 358170
rect 198996 358142 199332 358170
rect 200192 358142 200528 358170
rect 193312 358090 193364 358096
rect 193128 355904 193180 355910
rect 193128 355846 193180 355852
rect 191944 349030 192156 349058
rect 192128 348922 192156 349030
rect 193324 348922 193352 358090
rect 194138 357504 194194 357513
rect 194138 357439 194194 357448
rect 193680 354884 193732 354890
rect 193680 354826 193732 354832
rect 193692 351490 193720 354826
rect 193864 354816 193916 354822
rect 193864 354758 193916 354764
rect 193680 351484 193732 351490
rect 193680 351426 193732 351432
rect 193876 351422 193904 354758
rect 193864 351416 193916 351422
rect 193864 351358 193916 351364
rect 194152 348922 194180 357439
rect 194428 356046 194456 358142
rect 194416 356040 194468 356046
rect 194416 355982 194468 355988
rect 195624 354754 195652 358142
rect 196820 355638 196848 358142
rect 198108 355706 198136 358142
rect 198924 356040 198976 356046
rect 198924 355982 198976 355988
rect 198648 355972 198700 355978
rect 198648 355914 198700 355920
rect 198096 355700 198148 355706
rect 198096 355642 198148 355648
rect 196808 355632 196860 355638
rect 196808 355574 196860 355580
rect 195244 354748 195296 354754
rect 195244 354690 195296 354696
rect 195612 354748 195664 354754
rect 195612 354690 195664 354696
rect 195256 348922 195284 354690
rect 196348 351484 196400 351490
rect 196348 351426 196400 351432
rect 196360 348922 196388 351426
rect 197452 351416 197504 351422
rect 197452 351358 197504 351364
rect 197464 348922 197492 351358
rect 198660 350554 198688 355914
rect 198936 351898 198964 355982
rect 199304 355774 199332 358142
rect 200500 355978 200528 358142
rect 201420 358142 201480 358170
rect 202676 358142 202828 358170
rect 203872 358142 204208 358170
rect 205068 358142 205404 358170
rect 206356 358142 206692 358170
rect 207552 358142 207888 358170
rect 208748 358142 209084 358170
rect 210036 358142 210372 358170
rect 211232 358142 211568 358170
rect 201420 356046 201448 358142
rect 201408 356040 201460 356046
rect 201408 355982 201460 355988
rect 200488 355972 200540 355978
rect 200488 355914 200540 355920
rect 199660 355904 199712 355910
rect 199660 355846 199712 355852
rect 199292 355768 199344 355774
rect 199292 355710 199344 355716
rect 198924 351892 198976 351898
rect 198924 351834 198976 351840
rect 198660 350526 198780 350554
rect 198752 348922 198780 350526
rect 199672 348922 199700 355846
rect 201500 355632 201552 355638
rect 201500 355574 201552 355580
rect 201408 354748 201460 354754
rect 201408 354690 201460 354696
rect 200580 351892 200632 351898
rect 200580 351834 200632 351840
rect 200592 348922 200620 351834
rect 201420 350554 201448 354690
rect 201512 350946 201540 355574
rect 202800 355230 202828 358142
rect 204180 355910 204208 358142
rect 204168 355904 204220 355910
rect 204168 355846 204220 355852
rect 204996 355768 205048 355774
rect 204996 355710 205048 355716
rect 203892 355700 203944 355706
rect 203892 355642 203944 355648
rect 202788 355224 202840 355230
rect 202788 355166 202840 355172
rect 201500 350940 201552 350946
rect 201500 350882 201552 350888
rect 202880 350940 202932 350946
rect 202880 350882 202932 350888
rect 201420 350526 201632 350554
rect 201604 348922 201632 350526
rect 202892 348922 202920 350882
rect 203904 348922 203932 355642
rect 205008 348922 205036 355710
rect 205376 354754 205404 358142
rect 206100 355972 206152 355978
rect 206100 355914 206152 355920
rect 205364 354748 205416 354754
rect 205364 354690 205416 354696
rect 206112 348922 206140 355914
rect 206664 354822 206692 358142
rect 206928 356040 206980 356046
rect 206928 355982 206980 355988
rect 206652 354816 206704 354822
rect 206652 354758 206704 354764
rect 206940 350554 206968 355982
rect 207860 355434 207888 358142
rect 209056 355774 209084 358142
rect 210344 356046 210372 358142
rect 210332 356040 210384 356046
rect 210332 355982 210384 355988
rect 209228 355904 209280 355910
rect 209228 355846 209280 355852
rect 209044 355768 209096 355774
rect 209044 355710 209096 355716
rect 207848 355428 207900 355434
rect 207848 355370 207900 355376
rect 208308 355224 208360 355230
rect 208308 355166 208360 355172
rect 208320 350554 208348 355166
rect 206940 350526 207152 350554
rect 208320 350526 208440 350554
rect 207124 348922 207152 350526
rect 208412 348922 208440 350526
rect 209240 348922 209268 355846
rect 211540 355842 211568 358142
rect 212368 358142 212428 358170
rect 213624 358142 213868 358170
rect 214912 358142 215248 358170
rect 216108 358142 216444 358170
rect 217304 358142 217640 358170
rect 218592 358142 218928 358170
rect 219788 358142 220124 358170
rect 220984 358142 221320 358170
rect 211528 355836 211580 355842
rect 211528 355778 211580 355784
rect 212368 355026 212396 358142
rect 213840 355910 213868 358142
rect 215220 356046 215248 358142
rect 214748 356040 214800 356046
rect 214748 355982 214800 355988
rect 215208 356040 215260 356046
rect 215208 355982 215260 355988
rect 213828 355904 213880 355910
rect 213828 355846 213880 355852
rect 214012 355768 214064 355774
rect 214012 355710 214064 355716
rect 212632 355428 212684 355434
rect 212632 355370 212684 355376
rect 212356 355020 212408 355026
rect 212356 354962 212408 354968
rect 211436 354816 211488 354822
rect 211436 354758 211488 354764
rect 210332 354748 210384 354754
rect 210332 354690 210384 354696
rect 210344 348922 210372 354690
rect 211448 348922 211476 354758
rect 212644 348922 212672 355370
rect 189920 348894 190210 348922
rect 191208 348894 191314 348922
rect 192128 348894 192418 348922
rect 193324 348894 193430 348922
rect 194152 348894 194534 348922
rect 195256 348894 195638 348922
rect 196360 348894 196650 348922
rect 197464 348894 197754 348922
rect 198752 348894 198858 348922
rect 199672 348894 199962 348922
rect 200592 348894 200974 348922
rect 201604 348894 202078 348922
rect 202892 348894 203182 348922
rect 203904 348894 204194 348922
rect 205008 348894 205298 348922
rect 206112 348894 206402 348922
rect 207124 348894 207506 348922
rect 208412 348894 208518 348922
rect 209240 348894 209622 348922
rect 210344 348894 210726 348922
rect 211448 348894 211738 348922
rect 212644 348894 212842 348922
rect 214024 348786 214052 355710
rect 214760 348922 214788 355982
rect 215668 355836 215720 355842
rect 215668 355778 215720 355784
rect 215680 348922 215708 355778
rect 216416 354754 216444 358142
rect 217612 355706 217640 358142
rect 218060 355904 218112 355910
rect 218060 355846 218112 355852
rect 217600 355700 217652 355706
rect 217600 355642 217652 355648
rect 216772 355020 216824 355026
rect 216772 354962 216824 354968
rect 216404 354748 216456 354754
rect 216404 354690 216456 354696
rect 216784 348922 216812 354962
rect 218072 348922 218100 355846
rect 218900 355570 218928 358142
rect 218980 356040 219032 356046
rect 218980 355982 219032 355988
rect 218888 355564 218940 355570
rect 218888 355506 218940 355512
rect 218992 348922 219020 355982
rect 220096 355910 220124 358142
rect 221292 356046 221320 358142
rect 222120 358142 222180 358170
rect 223408 358142 223468 358170
rect 224664 358142 224908 358170
rect 225860 358142 226196 358170
rect 227148 358142 227484 358170
rect 228344 358142 228680 358170
rect 229540 358142 229876 358170
rect 230736 358142 231072 358170
rect 232024 358142 232360 358170
rect 221280 356040 221332 356046
rect 221280 355982 221332 355988
rect 222120 355978 222148 358142
rect 223212 356040 223264 356046
rect 223212 355982 223264 355988
rect 222108 355972 222160 355978
rect 222108 355914 222160 355920
rect 220084 355904 220136 355910
rect 220084 355846 220136 355852
rect 221188 355700 221240 355706
rect 221188 355642 221240 355648
rect 220084 354748 220136 354754
rect 220084 354690 220136 354696
rect 220096 348922 220124 354690
rect 221200 348922 221228 355642
rect 222384 355564 222436 355570
rect 222384 355506 222436 355512
rect 222396 348922 222424 355506
rect 223224 350810 223252 355982
rect 223408 354822 223436 358142
rect 223672 355904 223724 355910
rect 223672 355846 223724 355852
rect 223396 354816 223448 354822
rect 223396 354758 223448 354764
rect 223212 350804 223264 350810
rect 223212 350746 223264 350752
rect 214760 348894 215050 348922
rect 215680 348894 216062 348922
rect 216784 348894 217166 348922
rect 218072 348894 218270 348922
rect 218992 348894 219282 348922
rect 220096 348894 220386 348922
rect 221200 348894 221490 348922
rect 222396 348894 222594 348922
rect 223684 348786 223712 355846
rect 224880 355570 224908 358142
rect 226168 356046 226196 358142
rect 226156 356040 226208 356046
rect 226156 355982 226208 355988
rect 226984 356040 227036 356046
rect 226984 355982 227036 355988
rect 225420 355972 225472 355978
rect 225420 355914 225472 355920
rect 224868 355564 224920 355570
rect 224868 355506 224920 355512
rect 224316 350804 224368 350810
rect 224316 350746 224368 350752
rect 224328 348922 224356 350746
rect 225432 348922 225460 355914
rect 226524 354816 226576 354822
rect 226524 354758 226576 354764
rect 226536 348922 226564 354758
rect 226996 351286 227024 355982
rect 227456 355434 227484 358142
rect 227720 355564 227772 355570
rect 227720 355506 227772 355512
rect 227444 355428 227496 355434
rect 227444 355370 227496 355376
rect 226984 351280 227036 351286
rect 226984 351222 227036 351228
rect 227732 348922 227760 355506
rect 228652 354754 228680 358142
rect 229848 355842 229876 358142
rect 231044 355910 231072 358142
rect 232332 355978 232360 358142
rect 233160 358142 233220 358170
rect 234416 358142 234568 358170
rect 235704 358142 235856 358170
rect 236900 358142 237236 358170
rect 238096 358142 238432 358170
rect 239292 358142 239628 358170
rect 240580 358142 240916 358170
rect 241776 358142 242112 358170
rect 242972 358142 243308 358170
rect 233160 356046 233188 358142
rect 234540 356046 234568 358142
rect 233148 356040 233200 356046
rect 233148 355982 233200 355988
rect 233700 356040 233752 356046
rect 233700 355982 233752 355988
rect 234528 356040 234580 356046
rect 234528 355982 234580 355988
rect 232320 355972 232372 355978
rect 232320 355914 232372 355920
rect 231032 355904 231084 355910
rect 231032 355846 231084 355852
rect 233148 355904 233200 355910
rect 233148 355846 233200 355852
rect 229836 355836 229888 355842
rect 229836 355778 229888 355784
rect 230480 355836 230532 355842
rect 230480 355778 230532 355784
rect 228824 355428 228876 355434
rect 228824 355370 228876 355376
rect 228640 354748 228692 354754
rect 228640 354690 228692 354696
rect 228732 351280 228784 351286
rect 228732 351222 228784 351228
rect 228744 348922 228772 351222
rect 228836 351218 228864 355370
rect 230388 354748 230440 354754
rect 230388 354690 230440 354696
rect 228824 351212 228876 351218
rect 228824 351154 228876 351160
rect 229836 351212 229888 351218
rect 229836 351154 229888 351160
rect 229848 348922 229876 351154
rect 230400 350554 230428 354690
rect 230492 351014 230520 355778
rect 230480 351008 230532 351014
rect 230480 350950 230532 350956
rect 231860 351008 231912 351014
rect 231860 350950 231912 350956
rect 230400 350526 230704 350554
rect 230676 348922 230704 350526
rect 231872 348922 231900 350950
rect 233160 350554 233188 355846
rect 233712 350946 233740 355982
rect 234068 355972 234120 355978
rect 234068 355914 234120 355920
rect 233700 350940 233752 350946
rect 233700 350882 233752 350888
rect 233160 350526 233280 350554
rect 233252 348922 233280 350526
rect 234080 348922 234108 355914
rect 235828 355842 235856 358142
rect 235908 356040 235960 356046
rect 235908 355982 235960 355988
rect 235816 355836 235868 355842
rect 235816 355778 235868 355784
rect 235172 350940 235224 350946
rect 235172 350882 235224 350888
rect 235184 348922 235212 350882
rect 235920 350554 235948 355982
rect 237208 355026 237236 358142
rect 237288 355836 237340 355842
rect 237288 355778 237340 355784
rect 237196 355020 237248 355026
rect 237196 354962 237248 354968
rect 237300 350554 237328 355778
rect 238300 355020 238352 355026
rect 238300 354962 238352 354968
rect 235920 350526 236224 350554
rect 237300 350526 237420 350554
rect 236196 348922 236224 350526
rect 237392 348922 237420 350526
rect 238312 348922 238340 354962
rect 238404 354822 238432 358142
rect 239600 356046 239628 358142
rect 239588 356040 239640 356046
rect 239588 355982 239640 355988
rect 240508 356040 240560 356046
rect 240508 355982 240560 355988
rect 238392 354816 238444 354822
rect 238392 354758 238444 354764
rect 239404 354816 239456 354822
rect 239404 354758 239456 354764
rect 239416 348922 239444 354758
rect 240520 348922 240548 355982
rect 240888 355842 240916 358142
rect 242084 356046 242112 358142
rect 242072 356040 242124 356046
rect 242072 355982 242124 355988
rect 242900 356040 242952 356046
rect 242900 355982 242952 355988
rect 240876 355836 240928 355842
rect 240876 355778 240928 355784
rect 241704 355836 241756 355842
rect 241704 355778 241756 355784
rect 241716 348922 241744 355778
rect 242912 348922 242940 355982
rect 243280 355366 243308 358142
rect 244108 358142 244168 358170
rect 244108 355366 244136 358142
rect 245580 355994 245608 358278
rect 246652 358142 246896 358170
rect 247848 358142 248092 358170
rect 246868 355994 246896 358142
rect 245580 355966 245884 355994
rect 246868 355966 247080 355994
rect 243268 355360 243320 355366
rect 243268 355302 243320 355308
rect 243820 355360 243872 355366
rect 243820 355302 243872 355308
rect 244096 355360 244148 355366
rect 244096 355302 244148 355308
rect 244924 355360 244976 355366
rect 244924 355302 244976 355308
rect 243832 348922 243860 355302
rect 244936 348922 244964 355302
rect 245856 348922 245884 355966
rect 247052 348922 247080 355966
rect 248064 354822 248092 358142
rect 249122 357898 249150 358156
rect 250272 358142 250332 358170
rect 251192 358142 251528 358170
rect 252572 358142 252724 358170
rect 249122 357870 249196 357898
rect 248052 354816 248104 354822
rect 248052 354758 248104 354764
rect 248604 354816 248656 354822
rect 248604 354758 248656 354764
rect 224328 348894 224710 348922
rect 225432 348894 225814 348922
rect 226536 348894 226826 348922
rect 227732 348894 227930 348922
rect 228744 348894 229034 348922
rect 229848 348894 230138 348922
rect 230676 348894 231150 348922
rect 231872 348894 232254 348922
rect 233252 348894 233358 348922
rect 234080 348894 234370 348922
rect 235184 348894 235474 348922
rect 236196 348894 236578 348922
rect 237392 348894 237682 348922
rect 238312 348894 238694 348922
rect 239416 348894 239798 348922
rect 240520 348894 240902 348922
rect 241716 348894 241914 348922
rect 242912 348894 243018 348922
rect 243832 348894 244122 348922
rect 244936 348894 245226 348922
rect 245856 348894 246238 348922
rect 247052 348894 247342 348922
rect 248616 348786 248644 354758
rect 249168 348922 249196 357870
rect 250272 348922 250300 358142
rect 249168 348894 249458 348922
rect 250272 348894 250562 348922
rect 167012 348758 167578 348786
rect 169786 348758 169892 348786
rect 179446 348758 179552 348786
rect 189106 348758 189488 348786
rect 213946 348758 214052 348786
rect 223606 348758 223712 348786
rect 248446 348758 248644 348786
rect 251192 348786 251220 358142
rect 252572 348922 252600 358142
rect 253998 357898 254026 358156
rect 254872 358142 255208 358170
rect 256068 358142 256404 358170
rect 257356 358142 257692 358170
rect 258552 358142 258888 358170
rect 259564 358142 260084 358170
rect 261036 358142 261280 358170
rect 262232 358142 262568 358170
rect 263612 358142 263764 358170
rect 264624 358142 264960 358170
rect 265912 358142 266248 358170
rect 267108 358142 267444 358170
rect 268304 358142 268640 358170
rect 269500 358142 269836 358170
rect 270512 358142 271124 358170
rect 271892 358142 272320 358170
rect 273364 358142 273516 358170
rect 274652 358142 274804 358170
rect 275664 358142 276000 358170
rect 276860 358142 277196 358170
rect 278056 358142 278392 358170
rect 279344 358142 279680 358170
rect 280540 358142 280876 358170
rect 281736 358142 282072 358170
rect 253998 357870 254072 357898
rect 254044 355994 254072 357870
rect 253860 355966 254072 355994
rect 252572 348894 252770 348922
rect 253860 348786 253888 355966
rect 254872 355162 254900 358142
rect 256068 355706 256096 358142
rect 255320 355700 255372 355706
rect 255320 355642 255372 355648
rect 256056 355700 256108 355706
rect 256056 355642 256108 355648
rect 254124 355156 254176 355162
rect 254124 355098 254176 355104
rect 254860 355156 254912 355162
rect 254860 355098 254912 355104
rect 251192 348758 251666 348786
rect 253782 348758 253888 348786
rect 254136 348786 254164 355098
rect 255332 348786 255360 355642
rect 257356 355434 257384 358142
rect 258552 356046 258580 358142
rect 258080 356040 258132 356046
rect 258080 355982 258132 355988
rect 258540 356040 258592 356046
rect 259564 355994 259592 358142
rect 258540 355982 258592 355988
rect 256700 355428 256752 355434
rect 256700 355370 256752 355376
rect 257344 355428 257396 355434
rect 257344 355370 257396 355376
rect 256712 348922 256740 355370
rect 258092 349058 258120 355982
rect 259380 355966 259592 355994
rect 258092 349030 258212 349058
rect 256712 348894 257002 348922
rect 258184 348786 258212 349030
rect 259380 348786 259408 355966
rect 261036 354754 261064 358142
rect 262232 356046 262260 358142
rect 263612 356046 263640 358142
rect 261576 356040 261628 356046
rect 261576 355982 261628 355988
rect 262220 356040 262272 356046
rect 262220 355982 262272 355988
rect 262680 356040 262732 356046
rect 262680 355982 262732 355988
rect 263600 356040 263652 356046
rect 263600 355982 263652 355988
rect 260564 354748 260616 354754
rect 260564 354690 260616 354696
rect 261024 354748 261076 354754
rect 261024 354690 261076 354696
rect 260576 348786 260604 354690
rect 261588 348786 261616 355982
rect 262692 348786 262720 355982
rect 264624 355570 264652 358142
rect 263416 355564 263468 355570
rect 263416 355506 263468 355512
rect 264612 355564 264664 355570
rect 264612 355506 264664 355512
rect 263428 348922 263456 355506
rect 265912 355298 265940 358142
rect 267108 355434 267136 358142
rect 266084 355428 266136 355434
rect 266084 355370 266136 355376
rect 267096 355428 267148 355434
rect 267096 355370 267148 355376
rect 264888 355292 264940 355298
rect 264888 355234 264940 355240
rect 265900 355292 265952 355298
rect 265900 355234 265952 355240
rect 263428 348894 263534 348922
rect 264900 348786 264928 355234
rect 266096 348786 266124 355370
rect 268200 355156 268252 355162
rect 268200 355098 268252 355104
rect 267096 354748 267148 354754
rect 267096 354690 267148 354696
rect 267108 348786 267136 354690
rect 268212 348786 268240 355098
rect 268304 354754 268332 358142
rect 269500 355162 269528 358142
rect 269488 355156 269540 355162
rect 269488 355098 269540 355104
rect 268292 354748 268344 354754
rect 268292 354690 268344 354696
rect 270512 351490 270540 358142
rect 271328 351552 271380 351558
rect 271328 351494 271380 351500
rect 269028 351484 269080 351490
rect 269028 351426 269080 351432
rect 270500 351484 270552 351490
rect 270500 351426 270552 351432
rect 269040 348786 269068 351426
rect 270224 351416 270276 351422
rect 270224 351358 270276 351364
rect 270236 348786 270264 351358
rect 271340 348786 271368 351494
rect 271892 351422 271920 358142
rect 273364 351558 273392 358142
rect 274548 351892 274600 351898
rect 274548 351834 274600 351840
rect 273352 351552 273404 351558
rect 273352 351494 273404 351500
rect 273076 351484 273128 351490
rect 273076 351426 273128 351432
rect 271880 351416 271932 351422
rect 271880 351358 271932 351364
rect 272432 350940 272484 350946
rect 272432 350882 272484 350888
rect 272444 348786 272472 350882
rect 273088 348922 273116 351426
rect 273088 348894 273194 348922
rect 274560 348786 274588 351834
rect 274652 350946 274680 358142
rect 275664 351490 275692 358142
rect 276860 351898 276888 358142
rect 276848 351892 276900 351898
rect 276848 351834 276900 351840
rect 278056 351830 278084 358142
rect 278780 354748 278832 354754
rect 278780 354690 278832 354696
rect 275744 351824 275796 351830
rect 275744 351766 275796 351772
rect 278044 351824 278096 351830
rect 278044 351766 278096 351772
rect 275652 351484 275704 351490
rect 275652 351426 275704 351432
rect 274640 350940 274692 350946
rect 274640 350882 274692 350888
rect 275756 348786 275784 351766
rect 276664 351756 276716 351762
rect 276664 351698 276716 351704
rect 276676 348786 276704 351698
rect 278792 351694 278820 354690
rect 279344 351762 279372 358142
rect 280540 354754 280568 358142
rect 280528 354748 280580 354754
rect 280528 354690 280580 354696
rect 279332 351756 279384 351762
rect 279332 351698 279384 351704
rect 277768 351688 277820 351694
rect 277768 351630 277820 351636
rect 278780 351688 278832 351694
rect 278780 351630 278832 351636
rect 277780 348786 277808 351630
rect 281736 351626 281764 358142
rect 278688 351620 278740 351626
rect 278688 351562 278740 351568
rect 281724 351620 281776 351626
rect 281724 351562 281776 351568
rect 278700 348786 278728 351562
rect 254136 348758 254886 348786
rect 255332 348758 255990 348786
rect 258106 348758 258212 348786
rect 259210 348758 259408 348786
rect 260314 348758 260604 348786
rect 261326 348758 261616 348786
rect 262430 348758 262720 348786
rect 264546 348758 264928 348786
rect 265650 348758 266124 348786
rect 266754 348758 267136 348786
rect 267858 348758 268240 348786
rect 268870 348758 269068 348786
rect 269974 348758 270264 348786
rect 271078 348758 271368 348786
rect 272090 348758 272472 348786
rect 274298 348758 274588 348786
rect 275402 348758 275784 348786
rect 276414 348758 276704 348786
rect 277518 348758 277808 348786
rect 278622 348758 278728 348786
rect 127742 348622 128308 348650
rect 280342 347576 280398 347585
rect 280342 347511 280398 347520
rect 280356 338201 280384 347511
rect 280342 338192 280398 338201
rect 280342 338127 280398 338136
rect 280342 327040 280398 327049
rect 280342 326975 280398 326984
rect 21364 322788 21416 322794
rect 21364 322730 21416 322736
rect 22112 320958 22140 322932
rect 22192 322788 22244 322794
rect 22192 322730 22244 322736
rect 22100 320952 22152 320958
rect 22100 320894 22152 320900
rect 22008 320204 22060 320210
rect 22008 320146 22060 320152
rect 20628 318776 20680 318782
rect 20628 318718 20680 318724
rect 20640 315588 20668 318718
rect 22020 315602 22048 320146
rect 22204 319462 22232 322730
rect 22192 319456 22244 319462
rect 22192 319398 22244 319404
rect 23124 318782 23152 322932
rect 23388 320476 23440 320482
rect 23388 320418 23440 320424
rect 23112 318776 23164 318782
rect 23112 318718 23164 318724
rect 23400 315602 23428 320418
rect 24228 320210 24256 322932
rect 24768 320884 24820 320890
rect 24768 320826 24820 320832
rect 24216 320204 24268 320210
rect 24216 320146 24268 320152
rect 24780 315602 24808 320826
rect 25332 320482 25360 322932
rect 26344 320890 26372 322932
rect 26332 320884 26384 320890
rect 26332 320826 26384 320832
rect 25320 320476 25372 320482
rect 25320 320418 25372 320424
rect 27448 320346 27476 322932
rect 25320 320340 25372 320346
rect 25320 320282 25372 320288
rect 27436 320340 27488 320346
rect 27436 320282 27488 320288
rect 21758 315574 22048 315602
rect 22954 315574 23428 315602
rect 24596 315574 24808 315602
rect 25332 315588 25360 320282
rect 27712 320272 27764 320278
rect 27712 320214 27764 320220
rect 26516 320204 26568 320210
rect 26516 320146 26568 320152
rect 26528 315588 26556 320146
rect 27724 315588 27752 320214
rect 28552 320210 28580 322932
rect 29656 320278 29684 322932
rect 29644 320272 29696 320278
rect 29644 320214 29696 320220
rect 30288 320272 30340 320278
rect 30288 320214 30340 320220
rect 28540 320204 28592 320210
rect 28540 320146 28592 320152
rect 28908 320204 28960 320210
rect 28908 320146 28960 320152
rect 28920 315588 28948 320146
rect 30300 315602 30328 320214
rect 30668 320210 30696 322932
rect 31772 320278 31800 322932
rect 31760 320272 31812 320278
rect 31760 320214 31812 320220
rect 32876 320210 32904 322932
rect 33692 320272 33744 320278
rect 33692 320214 33744 320220
rect 30656 320204 30708 320210
rect 30656 320146 30708 320152
rect 31668 320204 31720 320210
rect 31668 320146 31720 320152
rect 32864 320204 32916 320210
rect 32864 320146 32916 320152
rect 33048 320204 33100 320210
rect 33048 320146 33100 320152
rect 31680 315602 31708 320146
rect 30130 315574 30328 315602
rect 31326 315574 31708 315602
rect 24596 315466 24624 315574
rect 33060 315466 33088 320146
rect 33704 315588 33732 320214
rect 33888 320210 33916 322932
rect 34992 320278 35020 322932
rect 35912 322918 36110 322946
rect 35912 320906 35940 322918
rect 35820 320878 35940 320906
rect 34980 320272 35032 320278
rect 34980 320214 35032 320220
rect 33876 320204 33928 320210
rect 33876 320146 33928 320152
rect 35820 318442 35848 320878
rect 37200 320210 37228 322932
rect 38212 320210 38240 322932
rect 39316 320210 39344 322932
rect 40052 322918 40434 322946
rect 40052 320226 40080 322918
rect 41432 320226 41460 322932
rect 35900 320204 35952 320210
rect 35900 320146 35952 320152
rect 37188 320204 37240 320210
rect 37188 320146 37240 320152
rect 37280 320204 37332 320210
rect 37280 320146 37332 320152
rect 38200 320204 38252 320210
rect 38200 320146 38252 320152
rect 38568 320204 38620 320210
rect 38568 320146 38620 320152
rect 39304 320204 39356 320210
rect 39304 320146 39356 320152
rect 39960 320198 40080 320226
rect 41340 320198 41460 320226
rect 42536 320210 42564 322932
rect 42892 320884 42944 320890
rect 42892 320826 42944 320832
rect 42524 320204 42576 320210
rect 34888 318436 34940 318442
rect 34888 318378 34940 318384
rect 35808 318436 35860 318442
rect 35808 318378 35860 318384
rect 34900 315588 34928 318378
rect 35912 315602 35940 320146
rect 36544 319456 36596 319462
rect 36544 319398 36596 319404
rect 35912 315574 36110 315602
rect 24150 315438 24624 315466
rect 32522 315438 33088 315466
rect 36556 315382 36584 319398
rect 37292 315588 37320 320146
rect 38580 315602 38608 320146
rect 39960 315602 39988 320198
rect 38502 315574 38608 315602
rect 39698 315574 39988 315602
rect 41340 315466 41368 320198
rect 42524 320146 42576 320152
rect 42800 320204 42852 320210
rect 42800 320146 42852 320152
rect 41420 320136 41472 320142
rect 41420 320078 41472 320084
rect 40894 315438 41368 315466
rect 41432 315466 41460 320078
rect 42812 315602 42840 320146
rect 42904 318102 42932 320826
rect 43640 320210 43668 322932
rect 44192 322918 44758 322946
rect 45572 322918 45770 322946
rect 46492 322918 46874 322946
rect 43628 320204 43680 320210
rect 43628 320146 43680 320152
rect 42892 318096 42944 318102
rect 42892 318038 42944 318044
rect 44192 315602 44220 322918
rect 45572 315602 45600 322918
rect 46492 315602 46520 322918
rect 47964 320210 47992 322932
rect 48332 322918 48990 322946
rect 49712 322918 50094 322946
rect 51092 322918 51198 322946
rect 52302 322918 52408 322946
rect 53314 322918 53788 322946
rect 46940 320204 46992 320210
rect 46940 320146 46992 320152
rect 47952 320204 48004 320210
rect 47952 320146 48004 320152
rect 42812 315574 43286 315602
rect 44192 315574 44482 315602
rect 45572 315574 45678 315602
rect 46492 315574 46874 315602
rect 46952 315466 46980 320146
rect 48332 315466 48360 322918
rect 49712 315466 49740 322918
rect 51092 315466 51120 322918
rect 52380 320226 52408 322918
rect 53760 320226 53788 322918
rect 54404 320346 54432 322932
rect 55324 322918 55522 322946
rect 54392 320340 54444 320346
rect 54392 320282 54444 320288
rect 55220 320340 55272 320346
rect 55220 320282 55272 320288
rect 52380 320198 52500 320226
rect 53760 320198 53880 320226
rect 52472 315602 52500 320198
rect 53852 315602 53880 320198
rect 52472 315574 52854 315602
rect 53852 315574 54050 315602
rect 55232 315588 55260 320282
rect 55324 315738 55352 322918
rect 56520 320226 56548 322932
rect 57638 322918 57928 322946
rect 58742 322918 59308 322946
rect 57900 320226 57928 322918
rect 59280 320226 59308 322918
rect 56520 320198 56640 320226
rect 57900 320198 58020 320226
rect 59280 320198 59400 320226
rect 59832 320210 59860 322932
rect 60844 320210 60872 322932
rect 61948 320278 61976 322932
rect 61936 320272 61988 320278
rect 61936 320214 61988 320220
rect 63052 320210 63080 322932
rect 64064 320890 64092 322932
rect 64052 320884 64104 320890
rect 64052 320826 64104 320832
rect 64880 320884 64932 320890
rect 64880 320826 64932 320832
rect 63500 320272 63552 320278
rect 63500 320214 63552 320220
rect 55324 315710 55996 315738
rect 55968 315466 55996 315710
rect 56612 315466 56640 320198
rect 57992 315466 58020 320198
rect 59372 315466 59400 320198
rect 59820 320204 59872 320210
rect 59820 320146 59872 320152
rect 60740 320204 60792 320210
rect 60740 320146 60792 320152
rect 60832 320204 60884 320210
rect 60832 320146 60884 320152
rect 62120 320204 62172 320210
rect 62120 320146 62172 320152
rect 63040 320204 63092 320210
rect 63040 320146 63092 320152
rect 60752 315466 60780 320146
rect 62132 315602 62160 320146
rect 63512 315602 63540 320214
rect 64328 320204 64380 320210
rect 64328 320146 64380 320152
rect 64340 315602 64368 320146
rect 64892 315738 64920 320826
rect 65168 320210 65196 322932
rect 66272 320346 66300 322932
rect 66260 320340 66312 320346
rect 66260 320282 66312 320288
rect 67376 320210 67404 322932
rect 67640 320340 67692 320346
rect 67640 320282 67692 320288
rect 65156 320204 65208 320210
rect 65156 320146 65208 320152
rect 66260 320204 66312 320210
rect 66260 320146 66312 320152
rect 67364 320204 67416 320210
rect 67364 320146 67416 320152
rect 64892 315710 65564 315738
rect 62132 315574 62422 315602
rect 63512 315574 63618 315602
rect 64340 315574 64814 315602
rect 65536 315466 65564 315710
rect 66272 315466 66300 320146
rect 67652 315466 67680 320282
rect 68388 320278 68416 322932
rect 69492 320346 69520 322932
rect 69480 320340 69532 320346
rect 69480 320282 69532 320288
rect 70596 320278 70624 322932
rect 68376 320272 68428 320278
rect 68376 320214 68428 320220
rect 70400 320272 70452 320278
rect 70400 320214 70452 320220
rect 70584 320272 70636 320278
rect 70584 320214 70636 320220
rect 69020 320204 69072 320210
rect 69020 320146 69072 320152
rect 69032 315466 69060 320146
rect 70412 315602 70440 320214
rect 71608 320210 71636 322932
rect 72712 320890 72740 322932
rect 72700 320884 72752 320890
rect 72700 320826 72752 320832
rect 73816 320822 73844 322932
rect 74540 320884 74592 320890
rect 74540 320826 74592 320832
rect 73804 320816 73856 320822
rect 73804 320758 73856 320764
rect 71780 320340 71832 320346
rect 71780 320282 71832 320288
rect 71596 320204 71648 320210
rect 71596 320146 71648 320152
rect 71792 315602 71820 320282
rect 73160 320272 73212 320278
rect 73160 320214 73212 320220
rect 70412 315574 70794 315602
rect 71792 315574 71990 315602
rect 73172 315588 73200 320214
rect 73252 320204 73304 320210
rect 73252 320146 73304 320152
rect 73264 315738 73292 320146
rect 73264 315710 73844 315738
rect 73816 315466 73844 315710
rect 74552 315466 74580 320826
rect 74920 320210 74948 322932
rect 75932 320958 75960 322932
rect 75920 320952 75972 320958
rect 75920 320894 75972 320900
rect 75920 320816 75972 320822
rect 75920 320758 75972 320764
rect 74908 320204 74960 320210
rect 74908 320146 74960 320152
rect 75932 315466 75960 320758
rect 77036 320278 77064 322932
rect 78140 320414 78168 322932
rect 78680 320952 78732 320958
rect 78680 320894 78732 320900
rect 78128 320408 78180 320414
rect 78128 320350 78180 320356
rect 77024 320272 77076 320278
rect 77024 320214 77076 320220
rect 77300 320204 77352 320210
rect 77300 320146 77352 320152
rect 77312 315466 77340 320146
rect 78692 315602 78720 320894
rect 79152 320210 79180 322932
rect 80256 320346 80284 322932
rect 81256 320408 81308 320414
rect 81256 320350 81308 320356
rect 80244 320340 80296 320346
rect 80244 320282 80296 320288
rect 79968 320272 80020 320278
rect 79968 320214 80020 320220
rect 79140 320204 79192 320210
rect 79140 320146 79192 320152
rect 79980 318730 80008 320214
rect 81268 318730 81296 320350
rect 81360 320278 81388 322932
rect 82464 320890 82492 322932
rect 82452 320884 82504 320890
rect 82452 320826 82504 320832
rect 83476 320822 83504 322932
rect 83464 320816 83516 320822
rect 83464 320758 83516 320764
rect 82820 320340 82872 320346
rect 82820 320282 82872 320288
rect 81348 320272 81400 320278
rect 81348 320214 81400 320220
rect 81624 320204 81676 320210
rect 81624 320146 81676 320152
rect 79980 318702 80376 318730
rect 81268 318702 81572 318730
rect 78692 315574 79166 315602
rect 80348 315588 80376 318702
rect 81544 315588 81572 318702
rect 81636 315738 81664 320146
rect 81636 315710 82308 315738
rect 82280 315466 82308 315710
rect 82832 315466 82860 320282
rect 83096 320272 83148 320278
rect 83096 320214 83148 320220
rect 83108 317558 83136 320214
rect 84580 320210 84608 322932
rect 85120 320884 85172 320890
rect 85120 320826 85172 320832
rect 84568 320204 84620 320210
rect 84568 320146 84620 320152
rect 85132 318442 85160 320826
rect 85684 320278 85712 322932
rect 85764 320816 85816 320822
rect 85764 320758 85816 320764
rect 85672 320272 85724 320278
rect 85672 320214 85724 320220
rect 85120 318436 85172 318442
rect 85120 318378 85172 318384
rect 85776 318374 85804 320758
rect 86696 320346 86724 322932
rect 87800 320414 87828 322932
rect 88904 320482 88932 322932
rect 88892 320476 88944 320482
rect 88892 320418 88944 320424
rect 87788 320408 87840 320414
rect 87788 320350 87840 320356
rect 86684 320340 86736 320346
rect 86684 320282 86736 320288
rect 89628 320272 89680 320278
rect 89628 320214 89680 320220
rect 88064 320204 88116 320210
rect 88064 320146 88116 320152
rect 88076 318442 88104 320146
rect 89640 318730 89668 320214
rect 90008 320210 90036 322932
rect 91020 320822 91048 322932
rect 92124 321094 92152 322932
rect 92112 321088 92164 321094
rect 92112 321030 92164 321036
rect 93228 320890 93256 322932
rect 93216 320884 93268 320890
rect 93216 320826 93268 320832
rect 91008 320816 91060 320822
rect 91008 320758 91060 320764
rect 94240 320482 94268 322932
rect 95240 320816 95292 320822
rect 95240 320758 95292 320764
rect 91284 320476 91336 320482
rect 91284 320418 91336 320424
rect 94228 320476 94280 320482
rect 94228 320418 94280 320424
rect 90088 320408 90140 320414
rect 90088 320350 90140 320356
rect 89996 320204 90048 320210
rect 89996 320146 90048 320152
rect 89640 318702 89944 318730
rect 86316 318436 86368 318442
rect 86316 318378 86368 318384
rect 88064 318436 88116 318442
rect 88064 318378 88116 318384
rect 88708 318436 88760 318442
rect 88708 318378 88760 318384
rect 85764 318368 85816 318374
rect 85764 318310 85816 318316
rect 83096 317552 83148 317558
rect 83096 317494 83148 317500
rect 85120 317552 85172 317558
rect 85120 317494 85172 317500
rect 85132 315588 85160 317494
rect 86328 315588 86356 318378
rect 87512 318368 87564 318374
rect 87512 318310 87564 318316
rect 87524 315588 87552 318310
rect 88720 315588 88748 318378
rect 89916 315588 89944 318702
rect 90100 318034 90128 320350
rect 91100 320340 91152 320346
rect 91100 320282 91152 320288
rect 90088 318028 90140 318034
rect 90088 317970 90140 317976
rect 91112 315588 91140 320282
rect 91296 318782 91324 320418
rect 92664 320204 92716 320210
rect 92664 320146 92716 320152
rect 91284 318776 91336 318782
rect 91284 318718 91336 318724
rect 92296 318028 92348 318034
rect 92296 317970 92348 317976
rect 92308 315588 92336 317970
rect 92676 317490 92704 320146
rect 93492 318776 93544 318782
rect 93492 318718 93544 318724
rect 92664 317484 92716 317490
rect 92664 317426 92716 317432
rect 93504 315588 93532 318718
rect 94688 317484 94740 317490
rect 94688 317426 94740 317432
rect 94700 315588 94728 317426
rect 95252 315466 95280 320758
rect 95344 320210 95372 322932
rect 96448 320278 96476 322932
rect 96620 321088 96672 321094
rect 96620 321030 96672 321036
rect 96436 320272 96488 320278
rect 96436 320214 96488 320220
rect 95332 320204 95384 320210
rect 95332 320146 95384 320152
rect 96632 315466 96660 321030
rect 97552 320414 97580 322932
rect 98000 320884 98052 320890
rect 98000 320826 98052 320832
rect 97540 320408 97592 320414
rect 97540 320350 97592 320356
rect 98012 315602 98040 320826
rect 98564 320346 98592 322932
rect 99668 320482 99696 322932
rect 100772 321298 100800 322932
rect 100760 321292 100812 321298
rect 100760 321234 100812 321240
rect 101784 321026 101812 322932
rect 101772 321020 101824 321026
rect 101772 320962 101824 320968
rect 102888 320958 102916 322932
rect 102876 320952 102928 320958
rect 102876 320894 102928 320900
rect 99472 320476 99524 320482
rect 99472 320418 99524 320424
rect 99656 320476 99708 320482
rect 99656 320418 99708 320424
rect 98552 320340 98604 320346
rect 98552 320282 98604 320288
rect 99104 320204 99156 320210
rect 99104 320146 99156 320152
rect 99116 318782 99144 320146
rect 99104 318776 99156 318782
rect 99104 318718 99156 318724
rect 98012 315574 98302 315602
rect 99484 315588 99512 320418
rect 102140 320408 102192 320414
rect 102140 320350 102192 320356
rect 100760 320272 100812 320278
rect 100760 320214 100812 320220
rect 100668 318776 100720 318782
rect 100668 318718 100720 318724
rect 100680 315588 100708 318718
rect 100772 315466 100800 320214
rect 102152 315466 102180 320350
rect 103992 320346 104020 322932
rect 104900 320476 104952 320482
rect 104900 320418 104952 320424
rect 103520 320340 103572 320346
rect 103520 320282 103572 320288
rect 103980 320340 104032 320346
rect 103980 320282 104032 320288
rect 103532 315466 103560 320282
rect 104912 315466 104940 320418
rect 105096 320278 105124 322932
rect 106108 320890 106136 322932
rect 106280 321292 106332 321298
rect 106280 321234 106332 321240
rect 106096 320884 106148 320890
rect 106096 320826 106148 320832
rect 105084 320272 105136 320278
rect 105084 320214 105136 320220
rect 106292 315602 106320 321234
rect 106372 321020 106424 321026
rect 106372 320962 106424 320968
rect 106384 318578 106412 320962
rect 107212 320210 107240 322932
rect 108316 321162 108344 322932
rect 108304 321156 108356 321162
rect 108304 321098 108356 321104
rect 109328 321026 109356 322932
rect 109316 321020 109368 321026
rect 109316 320962 109368 320968
rect 108948 320952 109000 320958
rect 108948 320894 109000 320900
rect 107200 320204 107252 320210
rect 107200 320146 107252 320152
rect 108960 318730 108988 320894
rect 110432 320550 110460 322932
rect 111536 321094 111564 322932
rect 112654 322918 113128 322946
rect 111524 321088 111576 321094
rect 111524 321030 111576 321036
rect 110420 320544 110472 320550
rect 110420 320486 110472 320492
rect 109776 320340 109828 320346
rect 109776 320282 109828 320288
rect 108960 318702 109080 318730
rect 106372 318572 106424 318578
rect 106372 318514 106424 318520
rect 107844 318572 107896 318578
rect 107844 318514 107896 318520
rect 106292 315574 106674 315602
rect 107856 315588 107884 318514
rect 109052 315588 109080 318702
rect 109788 315602 109816 320282
rect 110420 320272 110472 320278
rect 110420 320214 110472 320220
rect 110432 316010 110460 320214
rect 112444 320204 112496 320210
rect 112444 320146 112496 320152
rect 110432 315982 111012 316010
rect 109788 315574 110262 315602
rect 110984 315466 111012 315982
rect 41432 315438 42090 315466
rect 46952 315438 48070 315466
rect 48332 315438 49266 315466
rect 49712 315438 50462 315466
rect 51092 315438 51658 315466
rect 55968 315438 56442 315466
rect 56612 315438 57638 315466
rect 57992 315438 58834 315466
rect 59372 315438 60030 315466
rect 60752 315438 61226 315466
rect 65536 315438 66010 315466
rect 66272 315438 67206 315466
rect 67652 315438 68402 315466
rect 69032 315438 69598 315466
rect 73816 315438 74382 315466
rect 74552 315438 75578 315466
rect 75932 315438 76774 315466
rect 77312 315438 77970 315466
rect 82280 315438 82754 315466
rect 82832 315438 83950 315466
rect 95252 315438 95910 315466
rect 96632 315438 97106 315466
rect 100772 315438 101890 315466
rect 102152 315438 103086 315466
rect 103532 315438 104282 315466
rect 104912 315438 105478 315466
rect 110984 315438 111458 315466
rect 36544 315376 36596 315382
rect 36544 315318 36596 315324
rect 111800 315376 111852 315382
rect 111800 315318 111852 315324
rect 14556 315308 14608 315314
rect 14556 315250 14608 315256
rect 111812 313274 111840 315318
rect 111800 313268 111852 313274
rect 111800 313210 111852 313216
rect 17132 276004 17184 276010
rect 17132 275946 17184 275952
rect 17144 274961 17172 275946
rect 17130 274952 17186 274961
rect 17130 274887 17186 274896
rect 67178 236056 67234 236065
rect 67178 235991 67234 236000
rect 67192 230450 67220 235991
rect 67180 230444 67232 230450
rect 67180 230386 67232 230392
rect 72424 230444 72476 230450
rect 72424 230386 72476 230392
rect 72436 227118 72464 230386
rect 72424 227112 72476 227118
rect 72424 227054 72476 227060
rect 79324 227112 79376 227118
rect 79324 227054 79376 227060
rect 79336 224330 79364 227054
rect 112456 224398 112484 320146
rect 113100 224602 113128 322918
rect 113652 320210 113680 322932
rect 113824 320544 113876 320550
rect 113824 320486 113876 320492
rect 113640 320204 113692 320210
rect 113640 320146 113692 320152
rect 113364 318096 113416 318102
rect 113364 318038 113416 318044
rect 113376 306406 113404 318038
rect 113180 306400 113232 306406
rect 113180 306342 113232 306348
rect 113364 306400 113416 306406
rect 113364 306342 113416 306348
rect 113192 296698 113220 306342
rect 113192 296670 113404 296698
rect 113376 295361 113404 296670
rect 113362 295352 113418 295361
rect 113362 295287 113418 295296
rect 113088 224596 113140 224602
rect 113088 224538 113140 224544
rect 113836 224466 113864 320486
rect 114756 320210 114784 322932
rect 115768 322918 115874 322946
rect 116886 322918 117268 322946
rect 117990 322918 118648 322946
rect 115204 321156 115256 321162
rect 115204 321098 115256 321104
rect 114468 320204 114520 320210
rect 114468 320146 114520 320152
rect 114744 320204 114796 320210
rect 114744 320146 114796 320152
rect 114376 313268 114428 313274
rect 114376 313210 114428 313216
rect 114388 310826 114416 313210
rect 114376 310820 114428 310826
rect 114376 310762 114428 310768
rect 114480 224942 114508 320146
rect 114468 224936 114520 224942
rect 114468 224878 114520 224884
rect 115216 224806 115244 321098
rect 115204 224800 115256 224806
rect 115204 224742 115256 224748
rect 113824 224460 113876 224466
rect 113824 224402 113876 224408
rect 112444 224392 112496 224398
rect 112444 224334 112496 224340
rect 115768 224330 115796 322918
rect 115848 320204 115900 320210
rect 115848 320146 115900 320152
rect 115860 224670 115888 320146
rect 116584 310820 116636 310826
rect 116584 310762 116636 310768
rect 115848 224664 115900 224670
rect 115848 224606 115900 224612
rect 79324 224324 79376 224330
rect 79324 224266 79376 224272
rect 100300 224324 100352 224330
rect 100300 224266 100352 224272
rect 115756 224324 115808 224330
rect 115756 224266 115808 224272
rect 55220 220856 55272 220862
rect 55220 220798 55272 220804
rect 14464 220108 14516 220114
rect 14464 220050 14516 220056
rect 55232 219708 55260 220798
rect 100312 133906 100340 224266
rect 116398 221232 116454 221241
rect 116398 221167 116454 221176
rect 116412 220862 116440 221167
rect 116400 220856 116452 220862
rect 116400 220798 116452 220804
rect 116122 220008 116178 220017
rect 116122 219943 116178 219952
rect 116136 219502 116164 219943
rect 116124 219496 116176 219502
rect 116124 219438 116176 219444
rect 104808 219428 104860 219434
rect 104808 219370 104860 219376
rect 104820 219337 104848 219370
rect 104806 219328 104862 219337
rect 104806 219263 104862 219272
rect 116398 218920 116454 218929
rect 116398 218855 116454 218864
rect 116412 218074 116440 218855
rect 116400 218068 116452 218074
rect 116400 218010 116452 218016
rect 104808 218000 104860 218006
rect 104806 217968 104808 217977
rect 104860 217968 104862 217977
rect 104806 217903 104862 217912
rect 116398 217696 116454 217705
rect 116398 217631 116454 217640
rect 116412 216646 116440 217631
rect 104808 216640 104860 216646
rect 104806 216608 104808 216617
rect 116400 216640 116452 216646
rect 104860 216608 104862 216617
rect 104806 216543 104862 216552
rect 115938 216608 115994 216617
rect 116400 216582 116452 216588
rect 115938 216543 115994 216552
rect 115952 215966 115980 216543
rect 104808 215960 104860 215966
rect 104808 215902 104860 215908
rect 115940 215960 115992 215966
rect 115940 215902 115992 215908
rect 104820 215665 104848 215902
rect 104806 215656 104862 215665
rect 104806 215591 104862 215600
rect 116398 215384 116454 215393
rect 116398 215319 116400 215328
rect 116452 215319 116454 215328
rect 116400 215290 116452 215296
rect 104808 215280 104860 215286
rect 104808 215222 104860 215228
rect 104820 214713 104848 215222
rect 104806 214704 104862 214713
rect 104806 214639 104862 214648
rect 116398 214160 116454 214169
rect 116398 214095 116454 214104
rect 116412 213994 116440 214095
rect 116400 213988 116452 213994
rect 116400 213930 116452 213936
rect 104808 213920 104860 213926
rect 104808 213862 104860 213868
rect 104820 213489 104848 213862
rect 104806 213480 104862 213489
rect 104806 213415 104862 213424
rect 115938 213072 115994 213081
rect 115938 213007 115994 213016
rect 115952 212566 115980 213007
rect 115940 212560 115992 212566
rect 115940 212502 115992 212508
rect 104440 212492 104492 212498
rect 104440 212434 104492 212440
rect 104452 212129 104480 212434
rect 104438 212120 104494 212129
rect 104438 212055 104494 212064
rect 116306 211848 116362 211857
rect 116306 211783 116362 211792
rect 116320 211206 116348 211783
rect 116308 211200 116360 211206
rect 116308 211142 116360 211148
rect 104808 211132 104860 211138
rect 104808 211074 104860 211080
rect 104820 210905 104848 211074
rect 104806 210896 104862 210905
rect 104806 210831 104862 210840
rect 116306 210760 116362 210769
rect 116306 210695 116362 210704
rect 116320 209846 116348 210695
rect 116308 209840 116360 209846
rect 116308 209782 116360 209788
rect 104808 209772 104860 209778
rect 104808 209714 104860 209720
rect 104820 209545 104848 209714
rect 104806 209536 104862 209545
rect 104806 209471 104862 209480
rect 116030 209536 116086 209545
rect 116030 209471 116086 209480
rect 116044 208418 116072 209471
rect 116032 208412 116084 208418
rect 116032 208354 116084 208360
rect 104808 208344 104860 208350
rect 104808 208286 104860 208292
rect 116398 208312 116454 208321
rect 104820 208185 104848 208286
rect 116398 208247 116454 208256
rect 104806 208176 104862 208185
rect 104806 208111 104862 208120
rect 116306 207224 116362 207233
rect 116306 207159 116362 207168
rect 113824 207120 113876 207126
rect 113824 207062 113876 207068
rect 104716 206984 104768 206990
rect 104716 206926 104768 206932
rect 104806 206952 104862 206961
rect 104728 206281 104756 206926
rect 113836 206922 113864 207062
rect 116320 207058 116348 207159
rect 116412 207126 116440 208247
rect 116400 207120 116452 207126
rect 116400 207062 116452 207068
rect 116308 207052 116360 207058
rect 116308 206994 116360 207000
rect 104806 206887 104808 206896
rect 104860 206887 104862 206896
rect 113824 206916 113876 206922
rect 104808 206858 104860 206864
rect 113824 206858 113876 206864
rect 104714 206272 104770 206281
rect 104714 206207 104770 206216
rect 115938 206000 115994 206009
rect 115938 205935 115994 205944
rect 115952 205698 115980 205935
rect 115940 205692 115992 205698
rect 115940 205634 115992 205640
rect 104808 205624 104860 205630
rect 104808 205566 104860 205572
rect 104820 205057 104848 205566
rect 104806 205048 104862 205057
rect 104806 204983 104862 204992
rect 116398 204912 116454 204921
rect 116398 204847 116454 204856
rect 116412 204338 116440 204847
rect 116400 204332 116452 204338
rect 116400 204274 116452 204280
rect 104808 204264 104860 204270
rect 104808 204206 104860 204212
rect 104820 203697 104848 204206
rect 104806 203688 104862 203697
rect 104806 203623 104862 203632
rect 116306 203688 116362 203697
rect 116306 203623 116362 203632
rect 116320 202910 116348 203623
rect 116308 202904 116360 202910
rect 116308 202846 116360 202852
rect 104808 202836 104860 202842
rect 104808 202778 104860 202784
rect 104820 202473 104848 202778
rect 104806 202464 104862 202473
rect 104806 202399 104862 202408
rect 116122 202464 116178 202473
rect 116122 202399 116178 202408
rect 116136 201550 116164 202399
rect 116124 201544 116176 201550
rect 116124 201486 116176 201492
rect 104808 201476 104860 201482
rect 104808 201418 104860 201424
rect 104820 201113 104848 201418
rect 116122 201376 116178 201385
rect 116122 201311 116178 201320
rect 104806 201104 104862 201113
rect 104806 201039 104862 201048
rect 116136 200258 116164 201311
rect 116124 200252 116176 200258
rect 116124 200194 116176 200200
rect 113272 200184 113324 200190
rect 115940 200184 115992 200190
rect 113272 200126 113324 200132
rect 115938 200152 115940 200161
rect 115992 200152 115994 200161
rect 104808 200116 104860 200122
rect 104808 200058 104860 200064
rect 104820 199889 104848 200058
rect 104806 199880 104862 199889
rect 104806 199815 104862 199824
rect 113284 198694 113312 200126
rect 115938 200087 115994 200096
rect 115938 199064 115994 199073
rect 115938 198999 115994 199008
rect 115952 198762 115980 198999
rect 114468 198756 114520 198762
rect 114468 198698 114520 198704
rect 115940 198756 115992 198762
rect 115940 198698 115992 198704
rect 104808 198688 104860 198694
rect 104808 198630 104860 198636
rect 113272 198688 113324 198694
rect 113272 198630 113324 198636
rect 104820 198529 104848 198630
rect 104806 198520 104862 198529
rect 104806 198455 104862 198464
rect 104716 197328 104768 197334
rect 104716 197270 104768 197276
rect 104806 197296 104862 197305
rect 104728 196625 104756 197270
rect 114480 197266 114508 198698
rect 116122 197840 116178 197849
rect 116122 197775 116178 197784
rect 116136 197402 116164 197775
rect 116124 197396 116176 197402
rect 116124 197338 116176 197344
rect 104806 197231 104808 197240
rect 104860 197231 104862 197240
rect 114468 197260 114520 197266
rect 104808 197202 104860 197208
rect 114468 197202 114520 197208
rect 116398 196752 116454 196761
rect 116398 196687 116454 196696
rect 104714 196616 104770 196625
rect 104714 196551 104770 196560
rect 116412 196042 116440 196687
rect 116400 196036 116452 196042
rect 116400 195978 116452 195984
rect 104808 195968 104860 195974
rect 104808 195910 104860 195916
rect 104820 195401 104848 195910
rect 115938 195528 115994 195537
rect 115938 195463 115994 195472
rect 104806 195392 104862 195401
rect 104806 195327 104862 195336
rect 115952 194614 115980 195463
rect 115940 194608 115992 194614
rect 115940 194550 115992 194556
rect 104808 194540 104860 194546
rect 104808 194482 104860 194488
rect 104820 194041 104848 194482
rect 116122 194304 116178 194313
rect 116122 194239 116178 194248
rect 104806 194032 104862 194041
rect 104806 193967 104862 193976
rect 116136 193254 116164 194239
rect 116124 193248 116176 193254
rect 116124 193190 116176 193196
rect 116398 193216 116454 193225
rect 104440 193180 104492 193186
rect 116398 193151 116454 193160
rect 104440 193122 104492 193128
rect 104452 192817 104480 193122
rect 104438 192808 104494 192817
rect 104438 192743 104494 192752
rect 116412 192030 116440 193151
rect 113916 192024 113968 192030
rect 116400 192024 116452 192030
rect 113916 191966 113968 191972
rect 116030 191992 116086 192001
rect 113180 191956 113232 191962
rect 113180 191898 113232 191904
rect 104440 191820 104492 191826
rect 104440 191762 104492 191768
rect 104452 191457 104480 191762
rect 104438 191448 104494 191457
rect 104438 191383 104494 191392
rect 113192 190466 113220 191898
rect 113928 191826 113956 191966
rect 116400 191966 116452 191972
rect 116030 191927 116032 191936
rect 116084 191927 116086 191936
rect 116032 191898 116084 191904
rect 113916 191820 113968 191826
rect 113916 191762 113968 191768
rect 116490 190904 116546 190913
rect 116490 190839 116546 190848
rect 116504 190670 116532 190839
rect 113272 190664 113324 190670
rect 113272 190606 113324 190612
rect 116492 190664 116544 190670
rect 116492 190606 116544 190612
rect 104716 190460 104768 190466
rect 104716 190402 104768 190408
rect 113180 190460 113232 190466
rect 113180 190402 113232 190408
rect 104728 190233 104756 190402
rect 104714 190224 104770 190233
rect 104714 190159 104770 190168
rect 113284 189038 113312 190606
rect 116398 189680 116454 189689
rect 116398 189615 116454 189624
rect 116412 189106 116440 189615
rect 114468 189100 114520 189106
rect 114468 189042 114520 189048
rect 116400 189100 116452 189106
rect 116400 189042 116452 189048
rect 104808 189032 104860 189038
rect 104808 188974 104860 188980
rect 113272 189032 113324 189038
rect 113272 188974 113324 188980
rect 104820 188873 104848 188974
rect 104806 188864 104862 188873
rect 104806 188799 104862 188808
rect 114100 187740 114152 187746
rect 114100 187682 114152 187688
rect 104808 187672 104860 187678
rect 104808 187614 104860 187620
rect 104820 187513 104848 187614
rect 104806 187504 104862 187513
rect 104806 187439 104862 187448
rect 104716 186312 104768 186318
rect 104716 186254 104768 186260
rect 104806 186280 104862 186289
rect 104728 185609 104756 186254
rect 114112 186250 114140 187682
rect 114480 187678 114508 189042
rect 116398 188456 116454 188465
rect 116398 188391 116454 188400
rect 116412 187746 116440 188391
rect 116400 187740 116452 187746
rect 116400 187682 116452 187688
rect 114468 187672 114520 187678
rect 114468 187614 114520 187620
rect 115938 187368 115994 187377
rect 115938 187303 115994 187312
rect 115952 186386 115980 187303
rect 115940 186380 115992 186386
rect 115940 186322 115992 186328
rect 104806 186215 104808 186224
rect 104860 186215 104862 186224
rect 114100 186244 114152 186250
rect 104808 186186 104860 186192
rect 114100 186186 114152 186192
rect 116030 186144 116086 186153
rect 116030 186079 116086 186088
rect 104714 185600 104770 185609
rect 104714 185535 104770 185544
rect 114468 185020 114520 185026
rect 114468 184962 114520 184968
rect 104808 184884 104860 184890
rect 104808 184826 104860 184832
rect 104820 184385 104848 184826
rect 104806 184376 104862 184385
rect 104806 184311 104862 184320
rect 114376 183592 114428 183598
rect 114376 183534 114428 183540
rect 104808 183524 104860 183530
rect 104808 183466 104860 183472
rect 104820 183025 104848 183466
rect 104806 183016 104862 183025
rect 104806 182951 104862 182960
rect 113180 182232 113232 182238
rect 113180 182174 113232 182180
rect 104808 182164 104860 182170
rect 104808 182106 104860 182112
rect 104820 181801 104848 182106
rect 104806 181792 104862 181801
rect 104806 181727 104862 181736
rect 113192 180810 113220 182174
rect 114388 182170 114416 183534
rect 114480 183530 114508 184962
rect 116044 184958 116072 186079
rect 116398 185056 116454 185065
rect 116398 184991 116400 185000
rect 116452 184991 116454 185000
rect 116400 184962 116452 184968
rect 116032 184952 116084 184958
rect 116032 184894 116084 184900
rect 116398 183832 116454 183841
rect 116398 183767 116454 183776
rect 116412 183598 116440 183767
rect 116400 183592 116452 183598
rect 116400 183534 116452 183540
rect 114468 183524 114520 183530
rect 114468 183466 114520 183472
rect 115938 182608 115994 182617
rect 115938 182543 115994 182552
rect 115952 182238 115980 182543
rect 115940 182232 115992 182238
rect 115940 182174 115992 182180
rect 114376 182164 114428 182170
rect 114376 182106 114428 182112
rect 115938 181520 115994 181529
rect 115938 181455 115994 181464
rect 115952 181150 115980 181455
rect 113272 181144 113324 181150
rect 113272 181086 113324 181092
rect 115940 181144 115992 181150
rect 115940 181086 115992 181092
rect 104808 180804 104860 180810
rect 104808 180746 104860 180752
rect 113180 180804 113232 180810
rect 113180 180746 113232 180752
rect 104820 180441 104848 180746
rect 104806 180432 104862 180441
rect 104806 180367 104862 180376
rect 113284 179382 113312 181086
rect 116398 180296 116454 180305
rect 116398 180231 116454 180240
rect 116412 179450 116440 180231
rect 113916 179444 113968 179450
rect 113916 179386 113968 179392
rect 116400 179444 116452 179450
rect 116400 179386 116452 179392
rect 104808 179376 104860 179382
rect 104808 179318 104860 179324
rect 113272 179376 113324 179382
rect 113272 179318 113324 179324
rect 104820 179081 104848 179318
rect 104806 179072 104862 179081
rect 104806 179007 104862 179016
rect 113928 178022 113956 179386
rect 115938 179208 115994 179217
rect 115938 179143 115994 179152
rect 115952 178090 115980 179143
rect 114192 178084 114244 178090
rect 114192 178026 114244 178032
rect 115940 178084 115992 178090
rect 115940 178026 115992 178032
rect 104164 178016 104216 178022
rect 104164 177958 104216 177964
rect 113916 178016 113968 178022
rect 113916 177958 113968 177964
rect 104176 177857 104204 177958
rect 104162 177848 104218 177857
rect 104162 177783 104218 177792
rect 114100 176792 114152 176798
rect 114100 176734 114152 176740
rect 104164 176656 104216 176662
rect 104164 176598 104216 176604
rect 104176 176497 104204 176598
rect 104162 176488 104218 176497
rect 104162 176423 104218 176432
rect 104806 175264 104862 175273
rect 114112 175234 114140 176734
rect 114204 176662 114232 178026
rect 115938 177984 115994 177993
rect 115938 177919 115994 177928
rect 115952 176798 115980 177919
rect 116398 176896 116454 176905
rect 116398 176831 116454 176840
rect 115940 176792 115992 176798
rect 115940 176734 115992 176740
rect 116412 176730 116440 176831
rect 114468 176724 114520 176730
rect 114468 176666 114520 176672
rect 116400 176724 116452 176730
rect 116400 176666 116452 176672
rect 114192 176656 114244 176662
rect 114192 176598 114244 176604
rect 114284 175296 114336 175302
rect 114284 175238 114336 175244
rect 104806 175199 104808 175208
rect 104860 175199 104862 175208
rect 114100 175228 114152 175234
rect 104808 175170 104860 175176
rect 114100 175170 114152 175176
rect 104532 175160 104584 175166
rect 104532 175102 104584 175108
rect 104544 174593 104572 175102
rect 104530 174584 104586 174593
rect 104530 174519 104586 174528
rect 114296 173874 114324 175238
rect 114480 175166 114508 176666
rect 116398 175672 116454 175681
rect 116398 175607 116454 175616
rect 116412 175302 116440 175607
rect 116400 175296 116452 175302
rect 116400 175238 116452 175244
rect 114468 175160 114520 175166
rect 114468 175102 114520 175108
rect 115938 174448 115994 174457
rect 115938 174383 115994 174392
rect 115952 173942 115980 174383
rect 114376 173936 114428 173942
rect 114376 173878 114428 173884
rect 115940 173936 115992 173942
rect 115940 173878 115992 173884
rect 104808 173868 104860 173874
rect 104808 173810 104860 173816
rect 114284 173868 114336 173874
rect 114284 173810 114336 173816
rect 104820 173369 104848 173810
rect 104806 173360 104862 173369
rect 104806 173295 104862 173304
rect 113180 172576 113232 172582
rect 113180 172518 113232 172524
rect 104440 172508 104492 172514
rect 104440 172450 104492 172456
rect 104452 172145 104480 172450
rect 104438 172136 104494 172145
rect 104438 172071 104494 172080
rect 113192 171086 113220 172518
rect 114388 172514 114416 173878
rect 116398 173360 116454 173369
rect 116398 173295 116454 173304
rect 116412 172582 116440 173295
rect 116400 172576 116452 172582
rect 116400 172518 116452 172524
rect 114376 172508 114428 172514
rect 114376 172450 114428 172456
rect 116122 172136 116178 172145
rect 116122 172071 116178 172080
rect 116136 171630 116164 172071
rect 113272 171624 113324 171630
rect 113272 171566 113324 171572
rect 116124 171624 116176 171630
rect 116124 171566 116176 171572
rect 104808 171080 104860 171086
rect 104808 171022 104860 171028
rect 113180 171080 113232 171086
rect 113180 171022 113232 171028
rect 104820 170785 104848 171022
rect 104806 170776 104862 170785
rect 104806 170711 104862 170720
rect 104256 169788 104308 169794
rect 104256 169730 104308 169736
rect 104164 168360 104216 168366
rect 104164 168302 104216 168308
rect 104176 168201 104204 168302
rect 104162 168192 104218 168201
rect 104162 168127 104218 168136
rect 104268 166977 104296 169730
rect 113284 169726 113312 171566
rect 116306 171048 116362 171057
rect 116306 170983 116362 170992
rect 116320 169862 116348 170983
rect 113916 169856 113968 169862
rect 113916 169798 113968 169804
rect 116308 169856 116360 169862
rect 116308 169798 116360 169804
rect 116398 169824 116454 169833
rect 104808 169720 104860 169726
rect 104808 169662 104860 169668
rect 113272 169720 113324 169726
rect 113272 169662 113324 169668
rect 104820 169425 104848 169662
rect 104806 169416 104862 169425
rect 104806 169351 104862 169360
rect 104808 168428 104860 168434
rect 104808 168370 104860 168376
rect 104254 166968 104310 166977
rect 104254 166903 104310 166912
rect 104820 165617 104848 168370
rect 113928 168366 113956 169798
rect 116398 169759 116400 169768
rect 116452 169759 116454 169768
rect 116400 169730 116452 169736
rect 116398 168600 116454 168609
rect 116398 168535 116454 168544
rect 116412 168434 116440 168535
rect 116400 168428 116452 168434
rect 116400 168370 116452 168376
rect 113916 168360 113968 168366
rect 113916 168302 113968 168308
rect 115938 167512 115994 167521
rect 115938 167447 115994 167456
rect 115952 167074 115980 167447
rect 114468 167068 114520 167074
rect 114468 167010 114520 167016
rect 115940 167068 115992 167074
rect 115940 167010 115992 167016
rect 113824 165640 113876 165646
rect 104806 165608 104862 165617
rect 104624 165572 104676 165578
rect 113824 165582 113876 165588
rect 104806 165543 104862 165552
rect 104624 165514 104676 165520
rect 104636 164937 104664 165514
rect 104622 164928 104678 164937
rect 104622 164863 104678 164872
rect 113836 164218 113864 165582
rect 114480 165578 114508 167010
rect 115938 166288 115994 166297
rect 115938 166223 115994 166232
rect 115952 165646 115980 166223
rect 115940 165640 115992 165646
rect 115940 165582 115992 165588
rect 114468 165572 114520 165578
rect 114468 165514 114520 165520
rect 116122 165200 116178 165209
rect 116122 165135 116178 165144
rect 116136 164286 116164 165135
rect 114468 164280 114520 164286
rect 114468 164222 114520 164228
rect 116124 164280 116176 164286
rect 116124 164222 116176 164228
rect 104808 164212 104860 164218
rect 104808 164154 104860 164160
rect 113824 164212 113876 164218
rect 113824 164154 113876 164160
rect 104820 163713 104848 164154
rect 104806 163704 104862 163713
rect 104806 163639 104862 163648
rect 113180 162920 113232 162926
rect 113180 162862 113232 162868
rect 104808 162852 104860 162858
rect 104808 162794 104860 162800
rect 104820 162353 104848 162794
rect 104806 162344 104862 162353
rect 104806 162279 104862 162288
rect 103704 161492 103756 161498
rect 103704 161434 103756 161440
rect 103716 158681 103744 161434
rect 113192 161430 113220 162862
rect 114480 162858 114508 164222
rect 116398 163976 116454 163985
rect 116398 163911 116454 163920
rect 116412 162926 116440 163911
rect 116400 162920 116452 162926
rect 116400 162862 116452 162868
rect 114468 162852 114520 162858
rect 114468 162794 114520 162800
rect 116214 162752 116270 162761
rect 116214 162687 116270 162696
rect 116228 162042 116256 162687
rect 113272 162036 113324 162042
rect 113272 161978 113324 161984
rect 116216 162036 116268 162042
rect 116216 161978 116268 161984
rect 104808 161424 104860 161430
rect 104808 161366 104860 161372
rect 113180 161424 113232 161430
rect 113180 161366 113232 161372
rect 104820 160993 104848 161366
rect 104806 160984 104862 160993
rect 104806 160919 104862 160928
rect 104256 160132 104308 160138
rect 104256 160074 104308 160080
rect 103702 158672 103758 158681
rect 103702 158607 103758 158616
rect 104268 157321 104296 160074
rect 113284 160070 113312 161978
rect 116398 161664 116454 161673
rect 116398 161599 116454 161608
rect 116412 161498 116440 161599
rect 116400 161492 116452 161498
rect 116400 161434 116452 161440
rect 116398 160440 116454 160449
rect 116398 160375 116454 160384
rect 116412 160138 116440 160375
rect 116400 160132 116452 160138
rect 116400 160074 116452 160080
rect 104808 160064 104860 160070
rect 104808 160006 104860 160012
rect 113272 160064 113324 160070
rect 113272 160006 113324 160012
rect 104820 159769 104848 160006
rect 104806 159760 104862 159769
rect 104806 159695 104862 159704
rect 116398 159352 116454 159361
rect 116398 159287 116454 159296
rect 116412 158778 116440 159287
rect 104808 158772 104860 158778
rect 104808 158714 104860 158720
rect 116400 158772 116452 158778
rect 116400 158714 116452 158720
rect 104348 157412 104400 157418
rect 104348 157354 104400 157360
rect 104254 157312 104310 157321
rect 104254 157247 104310 157256
rect 104256 154624 104308 154630
rect 104256 154566 104308 154572
rect 103796 153264 103848 153270
rect 103796 153206 103848 153212
rect 103704 151836 103756 151842
rect 103704 151778 103756 151784
rect 103716 149025 103744 151778
rect 103808 150385 103836 153206
rect 104268 151609 104296 154566
rect 104360 154465 104388 157354
rect 104820 155961 104848 158714
rect 116398 158128 116454 158137
rect 116398 158063 116454 158072
rect 116412 157418 116440 158063
rect 116400 157412 116452 157418
rect 116400 157354 116452 157360
rect 116030 157040 116086 157049
rect 116030 156975 116086 156984
rect 116044 155990 116072 156975
rect 114284 155984 114336 155990
rect 104806 155952 104862 155961
rect 114284 155926 114336 155932
rect 116032 155984 116084 155990
rect 116032 155926 116084 155932
rect 104806 155887 104862 155896
rect 113456 154692 113508 154698
rect 113456 154634 113508 154640
rect 104624 154556 104676 154562
rect 104624 154498 104676 154504
rect 104346 154456 104402 154465
rect 104346 154391 104402 154400
rect 104636 153921 104664 154498
rect 104622 153912 104678 153921
rect 104622 153847 104678 153856
rect 113468 153202 113496 154634
rect 114296 154562 114324 155926
rect 116030 155816 116086 155825
rect 116030 155751 116086 155760
rect 116044 154698 116072 155751
rect 116032 154692 116084 154698
rect 116032 154634 116084 154640
rect 116400 154624 116452 154630
rect 116398 154592 116400 154601
rect 116452 154592 116454 154601
rect 114284 154556 114336 154562
rect 116398 154527 116454 154536
rect 114284 154498 114336 154504
rect 115938 153504 115994 153513
rect 115938 153439 115994 153448
rect 115952 153270 115980 153439
rect 115940 153264 115992 153270
rect 115940 153206 115992 153212
rect 104808 153196 104860 153202
rect 104808 153138 104860 153144
rect 113456 153196 113508 153202
rect 113456 153138 113508 153144
rect 104820 152697 104848 153138
rect 104806 152688 104862 152697
rect 104806 152623 104862 152632
rect 116398 152280 116454 152289
rect 116398 152215 116454 152224
rect 116412 151842 116440 152215
rect 116400 151836 116452 151842
rect 116400 151778 116452 151784
rect 104254 151600 104310 151609
rect 104254 151535 104310 151544
rect 116398 151192 116454 151201
rect 116398 151127 116454 151136
rect 116412 150482 116440 151127
rect 104348 150476 104400 150482
rect 104348 150418 104400 150424
rect 116400 150476 116452 150482
rect 116400 150418 116452 150424
rect 103794 150376 103850 150385
rect 103794 150311 103850 150320
rect 103702 149016 103758 149025
rect 103702 148951 103758 148960
rect 104360 147665 104388 150418
rect 116398 149968 116454 149977
rect 116398 149903 116454 149912
rect 116412 149122 116440 149903
rect 104808 149116 104860 149122
rect 104808 149058 104860 149064
rect 116400 149116 116452 149122
rect 116400 149058 116452 149064
rect 104716 147688 104768 147694
rect 104346 147656 104402 147665
rect 104716 147630 104768 147636
rect 104346 147591 104402 147600
rect 104532 146328 104584 146334
rect 104532 146270 104584 146276
rect 104164 144968 104216 144974
rect 104164 144910 104216 144916
rect 103520 143608 103572 143614
rect 103520 143550 103572 143556
rect 103532 140593 103560 143550
rect 103704 142180 103756 142186
rect 103704 142122 103756 142128
rect 103518 140584 103574 140593
rect 103518 140519 103574 140528
rect 103716 139369 103744 142122
rect 104176 141817 104204 144910
rect 104544 143041 104572 146270
rect 104624 144900 104676 144906
rect 104624 144842 104676 144848
rect 104636 144265 104664 144842
rect 104728 144809 104756 147630
rect 104820 146305 104848 149058
rect 116398 148744 116454 148753
rect 116398 148679 116454 148688
rect 116412 147694 116440 148679
rect 116400 147688 116452 147694
rect 115938 147656 115994 147665
rect 116400 147630 116452 147636
rect 115938 147591 115994 147600
rect 115952 146402 115980 147591
rect 116398 146432 116454 146441
rect 113640 146396 113692 146402
rect 113640 146338 113692 146344
rect 115940 146396 115992 146402
rect 116398 146367 116454 146376
rect 115940 146338 115992 146344
rect 104806 146296 104862 146305
rect 104806 146231 104862 146240
rect 113652 144906 113680 146338
rect 116412 146334 116440 146367
rect 116400 146328 116452 146334
rect 116400 146270 116452 146276
rect 116030 145344 116086 145353
rect 116030 145279 116086 145288
rect 116044 144974 116072 145279
rect 116032 144968 116084 144974
rect 116032 144910 116084 144916
rect 113640 144900 113692 144906
rect 113640 144842 113692 144848
rect 104714 144800 104770 144809
rect 104714 144735 104770 144744
rect 104622 144256 104678 144265
rect 104622 144191 104678 144200
rect 116398 144120 116454 144129
rect 116398 144055 116454 144064
rect 116412 143614 116440 144055
rect 116400 143608 116452 143614
rect 116400 143550 116452 143556
rect 104530 143032 104586 143041
rect 104530 142967 104586 142976
rect 116398 142896 116454 142905
rect 116398 142831 116454 142840
rect 116412 142186 116440 142831
rect 116400 142180 116452 142186
rect 116400 142122 116452 142128
rect 104162 141808 104218 141817
rect 104162 141743 104218 141752
rect 116398 141808 116454 141817
rect 116398 141743 116454 141752
rect 116412 140826 116440 141743
rect 104348 140820 104400 140826
rect 104348 140762 104400 140768
rect 116400 140820 116452 140826
rect 116400 140762 116452 140768
rect 103702 139360 103758 139369
rect 103702 139295 103758 139304
rect 104360 138009 104388 140762
rect 116398 140584 116454 140593
rect 116398 140519 116454 140528
rect 113548 139528 113600 139534
rect 116308 139528 116360 139534
rect 113548 139470 113600 139476
rect 116306 139496 116308 139505
rect 116360 139496 116362 139505
rect 104808 139460 104860 139466
rect 104808 139402 104860 139408
rect 104346 138000 104402 138009
rect 104346 137935 104402 137944
rect 104716 136672 104768 136678
rect 104820 136649 104848 139402
rect 104716 136614 104768 136620
rect 104806 136640 104862 136649
rect 104348 135312 104400 135318
rect 104348 135254 104400 135260
rect 100484 133952 100536 133958
rect 100312 133900 100484 133906
rect 100312 133894 100536 133900
rect 103612 133952 103664 133958
rect 103612 133894 103664 133900
rect 100312 133878 100524 133894
rect 100392 131164 100444 131170
rect 100392 131106 100444 131112
rect 10416 129260 10468 129266
rect 10416 129202 10468 129208
rect 10324 126948 10376 126954
rect 10324 126890 10376 126896
rect 32232 125089 32260 127228
rect 78232 125526 78260 127228
rect 100404 125526 100432 131106
rect 103624 127634 103652 133894
rect 104360 132025 104388 135254
rect 104728 133249 104756 136614
rect 104806 136575 104862 136584
rect 113560 135250 113588 139470
rect 116412 139466 116440 140519
rect 116306 139431 116362 139440
rect 116400 139460 116452 139466
rect 116400 139402 116452 139408
rect 115846 138272 115902 138281
rect 115846 138207 115902 138216
rect 104808 135244 104860 135250
rect 104808 135186 104860 135192
rect 113548 135244 113600 135250
rect 113548 135186 113600 135192
rect 104820 135153 104848 135186
rect 104806 135144 104862 135153
rect 104806 135079 104862 135088
rect 109868 133952 109920 133958
rect 109868 133894 109920 133900
rect 104808 133884 104860 133890
rect 104808 133826 104860 133832
rect 104820 133793 104848 133826
rect 104806 133784 104862 133793
rect 104806 133719 104862 133728
rect 104714 133240 104770 133249
rect 104714 133175 104770 133184
rect 104346 132016 104402 132025
rect 104346 131951 104402 131960
rect 109880 130762 109908 133894
rect 115860 133890 115888 138207
rect 116398 137184 116454 137193
rect 116398 137119 116454 137128
rect 116412 136678 116440 137119
rect 116400 136672 116452 136678
rect 116400 136614 116452 136620
rect 115938 135960 115994 135969
rect 115938 135895 115994 135904
rect 115952 135318 115980 135895
rect 115940 135312 115992 135318
rect 115940 135254 115992 135260
rect 116398 134736 116454 134745
rect 116398 134671 116454 134680
rect 116412 133958 116440 134671
rect 116400 133952 116452 133958
rect 116400 133894 116452 133900
rect 115848 133884 115900 133890
rect 115848 133826 115900 133832
rect 114560 132932 114612 132938
rect 114560 132874 114612 132880
rect 113916 131232 113968 131238
rect 113916 131174 113968 131180
rect 103980 130756 104032 130762
rect 103980 130698 104032 130704
rect 109868 130756 109920 130762
rect 109868 130698 109920 130704
rect 103992 130665 104020 130698
rect 103978 130656 104034 130665
rect 103978 130591 104034 130600
rect 104808 129736 104860 129742
rect 104808 129678 104860 129684
rect 104820 129305 104848 129678
rect 104806 129296 104862 129305
rect 104806 129231 104862 129240
rect 113928 128246 113956 131174
rect 114572 129742 114600 132874
rect 116398 132424 116454 132433
rect 116398 132359 116454 132368
rect 115938 131336 115994 131345
rect 115938 131271 115994 131280
rect 115952 131170 115980 131271
rect 116412 131238 116440 132359
rect 116400 131232 116452 131238
rect 116400 131174 116452 131180
rect 115940 131164 115992 131170
rect 115940 131106 115992 131112
rect 114560 129736 114612 129742
rect 114560 129678 114612 129684
rect 116400 129328 116452 129334
rect 116400 129270 116452 129276
rect 116412 128897 116440 129270
rect 116398 128888 116454 128897
rect 116398 128823 116454 128832
rect 116400 128308 116452 128314
rect 116400 128250 116452 128256
rect 104808 128240 104860 128246
rect 104808 128182 104860 128188
rect 113916 128240 113968 128246
rect 113916 128182 113968 128188
rect 104820 128081 104848 128182
rect 104806 128072 104862 128081
rect 104806 128007 104862 128016
rect 116412 127809 116440 128250
rect 116398 127800 116454 127809
rect 116398 127735 116454 127744
rect 103612 127628 103664 127634
rect 103612 127570 103664 127576
rect 116308 127628 116360 127634
rect 116308 127570 116360 127576
rect 78220 125520 78272 125526
rect 78220 125462 78272 125468
rect 100392 125520 100444 125526
rect 100392 125462 100444 125468
rect 32218 125080 32274 125089
rect 32218 125015 32274 125024
rect 116320 124273 116348 127570
rect 116400 126948 116452 126954
rect 116400 126890 116452 126896
rect 116412 126585 116440 126890
rect 116398 126576 116454 126585
rect 116398 126511 116454 126520
rect 116400 125588 116452 125594
rect 116400 125530 116452 125536
rect 116412 125497 116440 125530
rect 116398 125488 116454 125497
rect 116398 125423 116454 125432
rect 116306 124264 116362 124273
rect 116306 124199 116362 124208
rect 116596 123049 116624 310762
rect 117240 224534 117268 322918
rect 117964 321088 118016 321094
rect 117964 321030 118016 321036
rect 117228 224528 117280 224534
rect 117228 224470 117280 224476
rect 117976 223922 118004 321030
rect 118620 224194 118648 322918
rect 119080 320210 119108 322932
rect 119344 321020 119396 321026
rect 119344 320962 119396 320968
rect 119068 320204 119120 320210
rect 119068 320146 119120 320152
rect 119356 224874 119384 320962
rect 120184 320210 120212 322932
rect 121210 322918 121316 322946
rect 122314 322918 122788 322946
rect 123418 322918 124168 322946
rect 119988 320204 120040 320210
rect 119988 320146 120040 320152
rect 120172 320204 120224 320210
rect 120172 320146 120224 320152
rect 119344 224868 119396 224874
rect 119344 224810 119396 224816
rect 118608 224188 118660 224194
rect 118608 224130 118660 224136
rect 120000 224058 120028 320146
rect 121288 224262 121316 322918
rect 121552 320884 121604 320890
rect 121552 320826 121604 320832
rect 121368 320204 121420 320210
rect 121368 320146 121420 320152
rect 120080 224256 120132 224262
rect 120080 224198 120132 224204
rect 121276 224256 121328 224262
rect 121276 224198 121328 224204
rect 119988 224052 120040 224058
rect 119988 223994 120040 224000
rect 117964 223916 118016 223922
rect 117964 223858 118016 223864
rect 120092 221748 120120 224198
rect 121380 223990 121408 320146
rect 121368 223984 121420 223990
rect 121368 223926 121420 223932
rect 121092 223644 121144 223650
rect 121092 223586 121144 223592
rect 121104 221748 121132 223586
rect 121564 221626 121592 320826
rect 122760 224738 122788 322918
rect 122748 224732 122800 224738
rect 122748 224674 122800 224680
rect 123208 224392 123260 224398
rect 123208 224334 123260 224340
rect 123220 221748 123248 224334
rect 124140 223854 124168 322918
rect 124416 320210 124444 322932
rect 124404 320204 124456 320210
rect 124404 320146 124456 320152
rect 125416 320204 125468 320210
rect 125416 320146 125468 320152
rect 125428 226658 125456 320146
rect 125244 226630 125456 226658
rect 124312 224800 124364 224806
rect 124312 224742 124364 224748
rect 124128 223848 124180 223854
rect 124128 223790 124180 223796
rect 124324 221748 124352 224742
rect 125244 224126 125272 226630
rect 125520 225010 125548 322932
rect 126638 322918 126928 322946
rect 127742 322918 128308 322946
rect 125508 225004 125560 225010
rect 125508 224946 125560 224952
rect 125416 224868 125468 224874
rect 125416 224810 125468 224816
rect 125232 224120 125284 224126
rect 125232 224062 125284 224068
rect 125428 221748 125456 224810
rect 126428 224460 126480 224466
rect 126428 224402 126480 224408
rect 126440 221748 126468 224402
rect 126900 224398 126928 322918
rect 128280 224874 128308 322918
rect 128740 320210 128768 322932
rect 129844 320210 129872 322932
rect 130962 322918 131068 322946
rect 131974 322918 132448 322946
rect 128728 320204 128780 320210
rect 128728 320146 128780 320152
rect 129648 320204 129700 320210
rect 129648 320146 129700 320152
rect 129832 320204 129884 320210
rect 129832 320146 129884 320152
rect 130936 320204 130988 320210
rect 130936 320146 130988 320152
rect 128268 224868 128320 224874
rect 128268 224810 128320 224816
rect 129372 224596 129424 224602
rect 129372 224538 129424 224544
rect 128636 224460 128688 224466
rect 128636 224402 128688 224408
rect 126888 224392 126940 224398
rect 126888 224334 126940 224340
rect 127532 223916 127584 223922
rect 127532 223858 127584 223864
rect 127544 221748 127572 223858
rect 128648 221748 128676 224402
rect 129384 221762 129412 224538
rect 129660 223718 129688 320146
rect 130948 224942 130976 320146
rect 130936 224936 130988 224942
rect 130936 224878 130988 224884
rect 131040 224670 131068 322918
rect 130752 224664 130804 224670
rect 130752 224606 130804 224612
rect 131028 224664 131080 224670
rect 131028 224606 131080 224612
rect 129648 223712 129700 223718
rect 129648 223654 129700 223660
rect 129384 221734 129674 221762
rect 130764 221748 130792 224606
rect 132420 224602 132448 322918
rect 133064 320210 133092 322932
rect 134168 320210 134196 322932
rect 135272 320210 135300 322932
rect 136298 322918 136496 322946
rect 137402 322918 137968 322946
rect 133052 320204 133104 320210
rect 133052 320146 133104 320152
rect 133788 320204 133840 320210
rect 133788 320146 133840 320152
rect 134156 320204 134208 320210
rect 134156 320146 134208 320152
rect 135168 320204 135220 320210
rect 135168 320146 135220 320152
rect 135260 320204 135312 320210
rect 135260 320146 135312 320152
rect 132868 224800 132920 224806
rect 132868 224742 132920 224748
rect 132408 224596 132460 224602
rect 132408 224538 132460 224544
rect 131764 224324 131816 224330
rect 131764 224266 131816 224272
rect 131776 221748 131804 224266
rect 132880 221748 132908 224742
rect 133800 223786 133828 320146
rect 133972 224528 134024 224534
rect 133972 224470 134024 224476
rect 133788 223780 133840 223786
rect 133788 223722 133840 223728
rect 133984 221748 134012 224470
rect 134984 224052 135036 224058
rect 134984 223994 135036 224000
rect 134996 221748 135024 223994
rect 135180 223854 135208 320146
rect 136468 224330 136496 322918
rect 136548 320204 136600 320210
rect 136548 320146 136600 320152
rect 136456 224324 136508 224330
rect 136456 224266 136508 224272
rect 136560 224058 136588 320146
rect 137940 224534 137968 322918
rect 138492 320210 138520 322932
rect 139504 320210 139532 322932
rect 138480 320204 138532 320210
rect 138480 320146 138532 320152
rect 139308 320204 139360 320210
rect 139308 320146 139360 320152
rect 139492 320204 139544 320210
rect 139492 320146 139544 320152
rect 138204 224732 138256 224738
rect 138204 224674 138256 224680
rect 137928 224528 137980 224534
rect 137928 224470 137980 224476
rect 137192 224256 137244 224262
rect 137192 224198 137244 224204
rect 136548 224052 136600 224058
rect 136548 223994 136600 224000
rect 136088 223984 136140 223990
rect 136088 223926 136140 223932
rect 135168 223848 135220 223854
rect 135168 223790 135220 223796
rect 136100 221748 136128 223926
rect 137204 221748 137232 224198
rect 138216 221748 138244 224674
rect 139320 224210 139348 320146
rect 140608 224262 140636 322932
rect 141726 322918 142108 322946
rect 142830 322918 143488 322946
rect 140688 320204 140740 320210
rect 140688 320146 140740 320152
rect 140596 224256 140648 224262
rect 139320 224182 139440 224210
rect 140596 224198 140648 224204
rect 139308 224120 139360 224126
rect 139308 224062 139360 224068
rect 139320 221748 139348 224062
rect 139412 223922 139440 224182
rect 140320 224188 140372 224194
rect 140320 224130 140372 224136
rect 139400 223916 139452 223922
rect 139400 223858 139452 223864
rect 140332 221748 140360 224130
rect 140700 224126 140728 320146
rect 142080 224398 142108 322918
rect 142528 224460 142580 224466
rect 142528 224402 142580 224408
rect 141424 224392 141476 224398
rect 141424 224334 141476 224340
rect 142068 224392 142120 224398
rect 142068 224334 142120 224340
rect 140688 224120 140740 224126
rect 140688 224062 140740 224068
rect 141436 221748 141464 224334
rect 142540 221748 142568 224402
rect 143460 223990 143488 322918
rect 143828 320210 143856 322932
rect 144932 320210 144960 322932
rect 146050 322918 146248 322946
rect 147062 322918 147628 322946
rect 143816 320204 143868 320210
rect 143816 320146 143868 320152
rect 144828 320204 144880 320210
rect 144828 320146 144880 320152
rect 144920 320204 144972 320210
rect 144920 320146 144972 320152
rect 146116 320204 146168 320210
rect 146116 320146 146168 320152
rect 143540 224868 143592 224874
rect 143540 224810 143592 224816
rect 143448 223984 143500 223990
rect 143448 223926 143500 223932
rect 143552 221748 143580 224810
rect 144840 224194 144868 320146
rect 146024 254176 146076 254182
rect 146022 254144 146024 254153
rect 146076 254144 146078 254153
rect 146022 254079 146078 254088
rect 145748 224936 145800 224942
rect 145748 224878 145800 224884
rect 144828 224188 144880 224194
rect 144828 224130 144880 224136
rect 144644 223712 144696 223718
rect 144644 223654 144696 223660
rect 144656 221748 144684 223654
rect 145760 221748 145788 224878
rect 146128 224806 146156 320146
rect 146116 224800 146168 224806
rect 146116 224742 146168 224748
rect 146220 224466 146248 322918
rect 147600 224670 147628 322918
rect 148152 320210 148180 322932
rect 149256 320210 149284 322932
rect 148140 320204 148192 320210
rect 148140 320146 148192 320152
rect 148968 320204 149020 320210
rect 148968 320146 149020 320152
rect 149244 320204 149296 320210
rect 149244 320146 149296 320152
rect 150256 320204 150308 320210
rect 150256 320146 150308 320152
rect 146760 224664 146812 224670
rect 146760 224606 146812 224612
rect 147588 224664 147640 224670
rect 147588 224606 147640 224612
rect 146208 224460 146260 224466
rect 146208 224402 146260 224408
rect 146772 221748 146800 224606
rect 147864 224596 147916 224602
rect 147864 224538 147916 224544
rect 147876 221748 147904 224538
rect 148980 223786 149008 320146
rect 149520 254176 149572 254182
rect 149518 254144 149520 254153
rect 149572 254144 149574 254153
rect 149518 254079 149574 254088
rect 150268 224874 150296 320146
rect 150256 224868 150308 224874
rect 150256 224810 150308 224816
rect 150360 224602 150388 322932
rect 151386 322918 151768 322946
rect 152490 322918 153148 322946
rect 151740 224738 151768 322918
rect 151728 224732 151780 224738
rect 151728 224674 151780 224680
rect 150348 224596 150400 224602
rect 150348 224538 150400 224544
rect 152096 224324 152148 224330
rect 152096 224266 152148 224272
rect 151084 224052 151136 224058
rect 151084 223994 151136 224000
rect 149980 223848 150032 223854
rect 149980 223790 150032 223796
rect 148876 223780 148928 223786
rect 148876 223722 148928 223728
rect 148968 223780 149020 223786
rect 148968 223722 149020 223728
rect 148888 221748 148916 223722
rect 149992 221748 150020 223790
rect 151096 221748 151124 223994
rect 152108 221748 152136 224266
rect 153120 224058 153148 322918
rect 153580 320210 153608 322932
rect 154684 320210 154712 322932
rect 155710 322918 155908 322946
rect 156814 322918 157288 322946
rect 153568 320204 153620 320210
rect 153568 320146 153620 320152
rect 154488 320204 154540 320210
rect 154488 320146 154540 320152
rect 154672 320204 154724 320210
rect 154672 320146 154724 320152
rect 155776 320204 155828 320210
rect 155776 320146 155828 320152
rect 153200 224528 153252 224534
rect 153200 224470 153252 224476
rect 153108 224052 153160 224058
rect 153108 223994 153160 224000
rect 153212 221748 153240 224470
rect 154304 223916 154356 223922
rect 154304 223858 154356 223864
rect 154316 221748 154344 223858
rect 154500 223854 154528 320146
rect 155788 224942 155816 320146
rect 155776 224936 155828 224942
rect 155776 224878 155828 224884
rect 155880 224534 155908 322918
rect 155868 224528 155920 224534
rect 155868 224470 155920 224476
rect 156420 224256 156472 224262
rect 156420 224198 156472 224204
rect 155316 224120 155368 224126
rect 155316 224062 155368 224068
rect 154488 223848 154540 223854
rect 154488 223790 154540 223796
rect 155328 221748 155356 224062
rect 156432 221748 156460 224198
rect 157260 223718 157288 322918
rect 157904 320210 157932 322932
rect 158916 320210 158944 322932
rect 157892 320204 157944 320210
rect 157892 320146 157944 320152
rect 158628 320204 158680 320210
rect 158628 320146 158680 320152
rect 158904 320204 158956 320210
rect 158904 320146 158956 320152
rect 159916 320204 159968 320210
rect 159916 320146 159968 320152
rect 157432 224392 157484 224398
rect 157432 224334 157484 224340
rect 157248 223712 157300 223718
rect 157248 223654 157300 223660
rect 157444 221748 157472 224334
rect 158640 223990 158668 320146
rect 159928 224194 159956 320146
rect 160020 224262 160048 322932
rect 161138 322918 161428 322946
rect 162242 322918 162808 322946
rect 161400 224806 161428 322918
rect 160652 224800 160704 224806
rect 160652 224742 160704 224748
rect 161388 224800 161440 224806
rect 161388 224742 161440 224748
rect 160008 224256 160060 224262
rect 160008 224198 160060 224204
rect 159640 224188 159692 224194
rect 159640 224130 159692 224136
rect 159916 224188 159968 224194
rect 159916 224130 159968 224136
rect 158536 223984 158588 223990
rect 158536 223926 158588 223932
rect 158628 223984 158680 223990
rect 158628 223926 158680 223932
rect 158548 221748 158576 223926
rect 159652 221748 159680 224130
rect 160664 221748 160692 224742
rect 161756 224460 161808 224466
rect 161756 224402 161808 224408
rect 161768 221748 161796 224402
rect 162780 223922 162808 322918
rect 163240 320278 163268 322932
rect 163228 320272 163280 320278
rect 163228 320214 163280 320220
rect 164344 320210 164372 322932
rect 165462 322918 165568 322946
rect 166474 322918 166948 322946
rect 167578 322918 168328 322946
rect 164332 320204 164384 320210
rect 164332 320146 164384 320152
rect 165436 320204 165488 320210
rect 165436 320146 165488 320152
rect 164976 224868 165028 224874
rect 164976 224810 165028 224816
rect 162860 224664 162912 224670
rect 162860 224606 162912 224612
rect 162768 223916 162820 223922
rect 162768 223858 162820 223864
rect 162872 221748 162900 224606
rect 163872 223780 163924 223786
rect 163872 223722 163924 223728
rect 163884 221748 163912 223722
rect 164988 221748 165016 224810
rect 165448 224670 165476 320146
rect 165436 224664 165488 224670
rect 165436 224606 165488 224612
rect 165540 224330 165568 322918
rect 166080 224596 166132 224602
rect 166080 224538 166132 224544
rect 165528 224324 165580 224330
rect 165528 224266 165580 224272
rect 166092 221748 166120 224538
rect 166920 224126 166948 322918
rect 167644 320272 167696 320278
rect 167644 320214 167696 320220
rect 167656 224874 167684 320214
rect 167644 224868 167696 224874
rect 167644 224810 167696 224816
rect 167092 224732 167144 224738
rect 167092 224674 167144 224680
rect 166908 224120 166960 224126
rect 166908 224062 166960 224068
rect 167104 221748 167132 224674
rect 168196 224052 168248 224058
rect 168196 223994 168248 224000
rect 168208 221748 168236 223994
rect 168300 223786 168328 322918
rect 168668 320210 168696 322932
rect 169772 320210 169800 322932
rect 170798 322918 171088 322946
rect 171902 322918 172468 322946
rect 168656 320204 168708 320210
rect 168656 320146 168708 320152
rect 169668 320204 169720 320210
rect 169668 320146 169720 320152
rect 169760 320204 169812 320210
rect 169760 320146 169812 320152
rect 170956 320204 171008 320210
rect 170956 320146 171008 320152
rect 169680 224058 169708 320146
rect 170312 224936 170364 224942
rect 170312 224878 170364 224884
rect 169668 224052 169720 224058
rect 169668 223994 169720 224000
rect 169208 223848 169260 223854
rect 169208 223790 169260 223796
rect 168288 223780 168340 223786
rect 168288 223722 168340 223728
rect 169220 221748 169248 223790
rect 170324 221748 170352 224878
rect 170968 224738 170996 320146
rect 170956 224732 171008 224738
rect 170956 224674 171008 224680
rect 171060 224398 171088 322918
rect 171416 224528 171468 224534
rect 171416 224470 171468 224476
rect 171048 224392 171100 224398
rect 171048 224334 171100 224340
rect 171428 221748 171456 224470
rect 172440 223802 172468 322918
rect 172992 320210 173020 322932
rect 174004 320210 174032 322932
rect 175122 322918 175228 322946
rect 176226 322918 176608 322946
rect 177330 322918 177988 322946
rect 172980 320204 173032 320210
rect 172980 320146 173032 320152
rect 173808 320204 173860 320210
rect 173808 320146 173860 320152
rect 173992 320204 174044 320210
rect 173992 320146 174044 320152
rect 175096 320204 175148 320210
rect 175096 320146 175148 320152
rect 173820 223990 173848 320146
rect 175108 224602 175136 320146
rect 175096 224596 175148 224602
rect 175096 224538 175148 224544
rect 175200 224466 175228 322918
rect 175188 224460 175240 224466
rect 175188 224402 175240 224408
rect 175648 224256 175700 224262
rect 175648 224198 175700 224204
rect 174636 224188 174688 224194
rect 174636 224130 174688 224136
rect 173532 223984 173584 223990
rect 173532 223926 173584 223932
rect 173808 223984 173860 223990
rect 173808 223926 173860 223932
rect 172440 223774 172560 223802
rect 172532 223718 172560 223774
rect 172428 223712 172480 223718
rect 172428 223654 172480 223660
rect 172520 223712 172572 223718
rect 172520 223654 172572 223660
rect 172440 221748 172468 223654
rect 173544 221748 173572 223926
rect 174648 221748 174676 224130
rect 175660 221748 175688 224198
rect 176580 223854 176608 322918
rect 176752 224800 176804 224806
rect 176752 224742 176804 224748
rect 176568 223848 176620 223854
rect 176568 223790 176620 223796
rect 176764 221748 176792 224742
rect 177960 224194 177988 322918
rect 178328 320210 178356 322932
rect 179432 320210 179460 322932
rect 180550 322918 180656 322946
rect 181562 322918 182128 322946
rect 178316 320204 178368 320210
rect 178316 320146 178368 320152
rect 179328 320204 179380 320210
rect 179328 320146 179380 320152
rect 179420 320204 179472 320210
rect 179420 320146 179472 320152
rect 179340 224942 179368 320146
rect 179328 224936 179380 224942
rect 179328 224878 179380 224884
rect 178868 224868 178920 224874
rect 178868 224810 178920 224816
rect 177948 224188 178000 224194
rect 177948 224130 178000 224136
rect 177764 223916 177816 223922
rect 177764 223858 177816 223864
rect 177776 221748 177804 223858
rect 178880 221748 178908 224810
rect 179972 224664 180024 224670
rect 179972 224606 180024 224612
rect 179984 221748 180012 224606
rect 180628 224262 180656 322918
rect 180708 320204 180760 320210
rect 180708 320146 180760 320152
rect 180720 224874 180748 320146
rect 180708 224868 180760 224874
rect 180708 224810 180760 224816
rect 180984 224324 181036 224330
rect 180984 224266 181036 224272
rect 180616 224256 180668 224262
rect 180616 224198 180668 224204
rect 180996 221748 181024 224266
rect 182100 224210 182128 322918
rect 182652 320210 182680 322932
rect 183756 320210 183784 322932
rect 182640 320204 182692 320210
rect 182640 320146 182692 320152
rect 183468 320204 183520 320210
rect 183468 320146 183520 320152
rect 183744 320204 183796 320210
rect 183744 320146 183796 320152
rect 184756 320204 184808 320210
rect 184756 320146 184808 320152
rect 183480 224806 183508 320146
rect 183468 224800 183520 224806
rect 183468 224742 183520 224748
rect 184768 224534 184796 320146
rect 184756 224528 184808 224534
rect 184756 224470 184808 224476
rect 184860 224330 184888 322932
rect 185886 322918 186268 322946
rect 186990 322918 187648 322946
rect 188094 322918 188476 322946
rect 185584 315308 185636 315314
rect 185584 315250 185636 315256
rect 185596 274961 185624 315250
rect 185582 274952 185638 274961
rect 185582 274887 185638 274896
rect 185308 224732 185360 224738
rect 185308 224674 185360 224680
rect 184848 224324 184900 224330
rect 184848 224266 184900 224272
rect 182100 224182 182220 224210
rect 182192 224126 182220 224182
rect 182088 224120 182140 224126
rect 182088 224062 182140 224068
rect 182180 224120 182232 224126
rect 182180 224062 182232 224068
rect 182100 221748 182128 224062
rect 184204 224052 184256 224058
rect 184204 223994 184256 224000
rect 183192 223780 183244 223786
rect 183192 223722 183244 223728
rect 183204 221748 183232 223722
rect 184216 221748 184244 223994
rect 185320 221748 185348 224674
rect 186240 224670 186268 322918
rect 187620 224738 187648 322918
rect 187608 224732 187660 224738
rect 187608 224674 187660 224680
rect 186228 224664 186280 224670
rect 186228 224606 186280 224612
rect 188448 224398 188476 322918
rect 189092 320521 189120 322932
rect 189078 320512 189134 320521
rect 189078 320447 189134 320456
rect 190196 320249 190224 322932
rect 191300 320249 191328 322932
rect 192404 320385 192432 322932
rect 192390 320376 192446 320385
rect 192390 320311 192446 320320
rect 190182 320240 190238 320249
rect 190182 320175 190238 320184
rect 191286 320240 191342 320249
rect 191286 320175 191342 320184
rect 191840 320204 191892 320210
rect 191840 320146 191892 320152
rect 191196 318776 191248 318782
rect 191196 318718 191248 318724
rect 190000 318096 190052 318102
rect 190000 318038 190052 318044
rect 188896 317552 188948 317558
rect 188896 317494 188948 317500
rect 188908 315602 188936 317494
rect 190012 315602 190040 318038
rect 191208 315602 191236 318718
rect 191852 317558 191880 320146
rect 193416 319433 193444 322932
rect 194520 320249 194548 322932
rect 195624 320822 195652 322932
rect 195612 320816 195664 320822
rect 195612 320758 195664 320764
rect 194506 320240 194562 320249
rect 196636 320210 196664 322932
rect 197372 322918 197754 322946
rect 197372 320362 197400 322918
rect 197188 320334 197400 320362
rect 198740 320340 198792 320346
rect 194506 320175 194562 320184
rect 196624 320204 196676 320210
rect 196624 320146 196676 320152
rect 193402 319424 193458 319433
rect 193402 319359 193458 319368
rect 192392 318572 192444 318578
rect 192392 318514 192444 318520
rect 191840 317552 191892 317558
rect 191840 317494 191892 317500
rect 192404 315602 192432 318514
rect 193588 318504 193640 318510
rect 193588 318446 193640 318452
rect 193600 315602 193628 318446
rect 194508 318436 194560 318442
rect 194508 318378 194560 318384
rect 194520 315602 194548 318378
rect 195796 318300 195848 318306
rect 195796 318242 195848 318248
rect 195808 315602 195836 318242
rect 197188 318102 197216 320334
rect 198740 320282 198792 320288
rect 197544 320272 197596 320278
rect 197544 320214 197596 320220
rect 197268 320204 197320 320210
rect 197268 320146 197320 320152
rect 197280 318782 197308 320146
rect 197268 318776 197320 318782
rect 197268 318718 197320 318724
rect 197556 318578 197584 320214
rect 197544 318572 197596 318578
rect 197544 318514 197596 318520
rect 198752 318510 198780 320282
rect 198844 320210 198872 322932
rect 199948 320278 199976 322932
rect 200120 320408 200172 320414
rect 200120 320350 200172 320356
rect 199936 320272 199988 320278
rect 199936 320214 199988 320220
rect 198832 320204 198884 320210
rect 198832 320146 198884 320152
rect 199016 320204 199068 320210
rect 199016 320146 199068 320152
rect 198740 318504 198792 318510
rect 198740 318446 198792 318452
rect 199028 318442 199056 320146
rect 199016 318436 199068 318442
rect 199016 318378 199068 318384
rect 200132 318306 200160 320350
rect 200960 320346 200988 322932
rect 200948 320340 201000 320346
rect 200948 320282 201000 320288
rect 201500 320272 201552 320278
rect 201500 320214 201552 320220
rect 200764 318776 200816 318782
rect 200764 318718 200816 318724
rect 200120 318300 200172 318306
rect 200120 318242 200172 318248
rect 198372 318232 198424 318238
rect 198372 318174 198424 318180
rect 197176 318096 197228 318102
rect 197176 318038 197228 318044
rect 197176 317960 197228 317966
rect 197176 317902 197228 317908
rect 197188 315602 197216 317902
rect 198384 315602 198412 318174
rect 199568 317756 199620 317762
rect 199568 317698 199620 317704
rect 199580 315602 199608 317698
rect 200776 315602 200804 318718
rect 201512 317966 201540 320214
rect 202064 320210 202092 322932
rect 203168 320414 203196 322932
rect 203156 320408 203208 320414
rect 203156 320350 203208 320356
rect 204180 320278 204208 322932
rect 204260 320612 204312 320618
rect 204260 320554 204312 320560
rect 204168 320272 204220 320278
rect 204168 320214 204220 320220
rect 202052 320204 202104 320210
rect 202052 320146 202104 320152
rect 202880 320204 202932 320210
rect 202880 320146 202932 320152
rect 201960 318708 202012 318714
rect 201960 318650 202012 318656
rect 201500 317960 201552 317966
rect 201500 317902 201552 317908
rect 201972 315602 202000 318650
rect 202892 318238 202920 320146
rect 204168 318300 204220 318306
rect 204168 318242 204220 318248
rect 202880 318232 202932 318238
rect 202880 318174 202932 318180
rect 202788 318164 202840 318170
rect 202788 318106 202840 318112
rect 188600 315574 188936 315602
rect 189704 315574 190040 315602
rect 190900 315574 191236 315602
rect 192096 315574 192432 315602
rect 193292 315574 193628 315602
rect 194488 315574 194548 315602
rect 195684 315574 195836 315602
rect 196880 315574 197216 315602
rect 198076 315574 198412 315602
rect 199272 315574 199608 315602
rect 200468 315574 200804 315602
rect 201664 315574 202000 315602
rect 202800 315602 202828 318106
rect 204180 315602 204208 318242
rect 204272 317762 204300 320554
rect 205284 320210 205312 322932
rect 206388 320618 206416 322932
rect 207032 322918 207506 322946
rect 208412 322918 208518 322946
rect 206376 320612 206428 320618
rect 206376 320554 206428 320560
rect 205272 320204 205324 320210
rect 207032 320192 207060 322918
rect 208412 320770 208440 322918
rect 208320 320742 208440 320770
rect 205272 320146 205324 320152
rect 206940 320164 207060 320192
rect 207112 320204 207164 320210
rect 206940 318782 206968 320164
rect 207112 320146 207164 320152
rect 206928 318776 206980 318782
rect 206928 318718 206980 318724
rect 207124 318170 207152 320146
rect 208320 318714 208348 320742
rect 208400 320612 208452 320618
rect 208400 320554 208452 320560
rect 208308 318708 208360 318714
rect 208308 318650 208360 318656
rect 208412 318306 208440 320554
rect 209608 320210 209636 322932
rect 210712 320618 210740 322932
rect 211172 322918 211738 322946
rect 212552 322918 212842 322946
rect 210700 320612 210752 320618
rect 210700 320554 210752 320560
rect 211172 320226 211200 322918
rect 212552 320226 212580 322918
rect 213932 320498 213960 322932
rect 209596 320204 209648 320210
rect 209596 320146 209648 320152
rect 211080 320198 211200 320226
rect 212460 320198 212580 320226
rect 213840 320470 213960 320498
rect 209136 318436 209188 318442
rect 209136 318378 209188 318384
rect 208400 318300 208452 318306
rect 208400 318242 208452 318248
rect 207112 318164 207164 318170
rect 207112 318106 207164 318112
rect 207940 318164 207992 318170
rect 207940 318106 207992 318112
rect 204260 317756 204312 317762
rect 204260 317698 204312 317704
rect 206744 317620 206796 317626
rect 206744 317562 206796 317568
rect 205364 317552 205416 317558
rect 205364 317494 205416 317500
rect 205376 315602 205404 317494
rect 206756 315602 206784 317562
rect 207952 315602 207980 318106
rect 209148 315602 209176 318378
rect 210332 317756 210384 317762
rect 210332 317698 210384 317704
rect 210344 315602 210372 317698
rect 211080 317558 211108 320198
rect 211528 318776 211580 318782
rect 211528 318718 211580 318724
rect 211068 317552 211120 317558
rect 211068 317494 211120 317500
rect 211540 315602 211568 318718
rect 212460 317626 212488 320198
rect 213840 318170 213868 320470
rect 215036 318442 215064 322932
rect 215024 318436 215076 318442
rect 215024 318378 215076 318384
rect 213828 318164 213880 318170
rect 213828 318106 213880 318112
rect 213828 317960 213880 317966
rect 213828 317902 213880 317908
rect 212448 317620 212500 317626
rect 212448 317562 212500 317568
rect 212448 317484 212500 317490
rect 212448 317426 212500 317432
rect 212460 315602 212488 317426
rect 213840 315602 213868 317902
rect 216048 317762 216076 322932
rect 217152 318782 217180 322932
rect 218072 322918 218270 322946
rect 218072 320226 218100 322918
rect 217980 320198 218100 320226
rect 217140 318776 217192 318782
rect 217140 318718 217192 318724
rect 217508 318300 217560 318306
rect 217508 318242 217560 318248
rect 216036 317756 216088 317762
rect 216036 317698 216088 317704
rect 216312 317620 216364 317626
rect 216312 317562 216364 317568
rect 215116 317484 215168 317490
rect 215116 317426 215168 317432
rect 215128 315602 215156 317426
rect 216324 315602 216352 317562
rect 217520 315602 217548 318242
rect 217980 317558 218008 320198
rect 218704 318232 218756 318238
rect 218704 318174 218756 318180
rect 217968 317552 218020 317558
rect 217968 317494 218020 317500
rect 218716 315602 218744 318174
rect 219268 317966 219296 322932
rect 219900 320204 219952 320210
rect 219900 320146 219952 320152
rect 219256 317960 219308 317966
rect 219256 317902 219308 317908
rect 219912 315602 219940 320146
rect 220372 317490 220400 322932
rect 220636 318708 220688 318714
rect 220636 318650 220688 318656
rect 220360 317484 220412 317490
rect 220360 317426 220412 317432
rect 202800 315574 202860 315602
rect 204056 315574 204208 315602
rect 205252 315574 205404 315602
rect 206448 315574 206784 315602
rect 207644 315574 207980 315602
rect 208840 315574 209176 315602
rect 210036 315574 210372 315602
rect 211232 315574 211568 315602
rect 212428 315574 212488 315602
rect 213624 315574 213868 315602
rect 214820 315574 215156 315602
rect 216016 315574 216352 315602
rect 217212 315574 217548 315602
rect 218408 315574 218744 315602
rect 219604 315574 219940 315602
rect 220648 315602 220676 318650
rect 221476 317626 221504 322932
rect 222580 318306 222608 322932
rect 223488 318776 223540 318782
rect 223488 318718 223540 318724
rect 222568 318300 222620 318306
rect 222568 318242 222620 318248
rect 222016 317960 222068 317966
rect 222016 317902 222068 317908
rect 221464 317620 221516 317626
rect 221464 317562 221516 317568
rect 222028 315602 222056 317902
rect 223500 315602 223528 318718
rect 223592 318238 223620 322932
rect 224696 320210 224724 322932
rect 224684 320204 224736 320210
rect 224684 320146 224736 320152
rect 224868 320204 224920 320210
rect 224868 320146 224920 320152
rect 223580 318232 223632 318238
rect 223580 318174 223632 318180
rect 220648 315574 220800 315602
rect 221996 315574 222056 315602
rect 223192 315574 223528 315602
rect 224880 315466 224908 320146
rect 225800 318714 225828 322932
rect 226248 320680 226300 320686
rect 226248 320622 226300 320628
rect 225788 318708 225840 318714
rect 225788 318650 225840 318656
rect 226260 315602 226288 320622
rect 226812 317966 226840 322932
rect 227076 320816 227128 320822
rect 227076 320758 227128 320764
rect 226800 317960 226852 317966
rect 226800 317902 226852 317908
rect 227088 315602 227116 320758
rect 227916 318782 227944 322932
rect 228272 321020 228324 321026
rect 228272 320962 228324 320968
rect 227904 318776 227956 318782
rect 227904 318718 227956 318724
rect 228284 315602 228312 320962
rect 229020 320210 229048 322932
rect 230124 320686 230152 322932
rect 231136 320822 231164 322932
rect 231768 321224 231820 321230
rect 231768 321166 231820 321172
rect 231124 320816 231176 320822
rect 231124 320758 231176 320764
rect 230112 320680 230164 320686
rect 230112 320622 230164 320628
rect 229468 320340 229520 320346
rect 229468 320282 229520 320288
rect 229008 320204 229060 320210
rect 229008 320146 229060 320152
rect 229480 315602 229508 320282
rect 230296 320204 230348 320210
rect 230296 320146 230348 320152
rect 226076 315574 226288 315602
rect 226780 315574 227116 315602
rect 227976 315574 228312 315602
rect 229172 315574 229508 315602
rect 230308 315602 230336 320146
rect 231780 315602 231808 321166
rect 232240 321026 232268 322932
rect 232228 321020 232280 321026
rect 232228 320962 232280 320968
rect 233344 320346 233372 322932
rect 233332 320340 233384 320346
rect 233332 320282 233384 320288
rect 233148 320272 233200 320278
rect 233148 320214 233200 320220
rect 233160 315602 233188 320214
rect 234356 320210 234384 322932
rect 235460 321230 235488 322932
rect 235448 321224 235500 321230
rect 235448 321166 235500 321172
rect 235448 320476 235500 320482
rect 235448 320418 235500 320424
rect 234344 320204 234396 320210
rect 234344 320146 234396 320152
rect 234528 320204 234580 320210
rect 234528 320146 234580 320152
rect 230308 315574 230368 315602
rect 231564 315574 231808 315602
rect 232760 315574 233188 315602
rect 226076 315466 226104 315574
rect 234540 315466 234568 320146
rect 235460 315602 235488 320418
rect 236564 320278 236592 322932
rect 236644 320408 236696 320414
rect 236644 320350 236696 320356
rect 236552 320272 236604 320278
rect 236552 320214 236604 320220
rect 236656 315602 236684 320350
rect 237668 320210 237696 322932
rect 238680 320482 238708 322932
rect 238668 320476 238720 320482
rect 238668 320418 238720 320424
rect 239784 320414 239812 322932
rect 239772 320408 239824 320414
rect 239772 320350 239824 320356
rect 238668 320340 238720 320346
rect 238668 320282 238720 320288
rect 237840 320272 237892 320278
rect 237840 320214 237892 320220
rect 237656 320204 237708 320210
rect 237656 320146 237708 320152
rect 237852 315602 237880 320214
rect 235152 315574 235488 315602
rect 236348 315574 236684 315602
rect 237544 315574 237880 315602
rect 238680 315602 238708 320282
rect 240888 320278 240916 322932
rect 241900 320346 241928 322932
rect 241888 320340 241940 320346
rect 241888 320282 241940 320288
rect 242624 320340 242676 320346
rect 242624 320282 242676 320288
rect 240876 320272 240928 320278
rect 240876 320214 240928 320220
rect 241428 320272 241480 320278
rect 241428 320214 241480 320220
rect 240048 320204 240100 320210
rect 240048 320146 240100 320152
rect 240060 315602 240088 320146
rect 241440 315602 241468 320214
rect 242636 315602 242664 320282
rect 243004 320210 243032 322932
rect 244108 320278 244136 322932
rect 245212 320346 245240 322932
rect 246120 320476 246172 320482
rect 246120 320418 246172 320424
rect 245200 320340 245252 320346
rect 245200 320282 245252 320288
rect 244096 320272 244148 320278
rect 244096 320214 244148 320220
rect 245016 320272 245068 320278
rect 245016 320214 245068 320220
rect 242992 320204 243044 320210
rect 242992 320146 243044 320152
rect 243820 320204 243872 320210
rect 243820 320146 243872 320152
rect 243832 315602 243860 320146
rect 245028 315602 245056 320214
rect 246132 318186 246160 320418
rect 246224 320210 246252 322932
rect 247328 320278 247356 322932
rect 248236 320816 248288 320822
rect 248236 320758 248288 320764
rect 247316 320272 247368 320278
rect 247316 320214 247368 320220
rect 247408 320272 247460 320278
rect 247408 320214 247460 320220
rect 246212 320204 246264 320210
rect 246212 320146 246264 320152
rect 246132 318158 246252 318186
rect 246224 315602 246252 318158
rect 247420 315602 247448 320214
rect 238680 315574 238740 315602
rect 239936 315574 240088 315602
rect 241132 315574 241468 315602
rect 242328 315574 242664 315602
rect 243524 315574 243860 315602
rect 244720 315574 245056 315602
rect 245916 315574 246252 315602
rect 247112 315574 247448 315602
rect 248248 315602 248276 320758
rect 248432 320482 248460 322932
rect 248420 320476 248472 320482
rect 248420 320418 248472 320424
rect 249444 320278 249472 322932
rect 250548 320822 250576 322932
rect 250536 320816 250588 320822
rect 250536 320758 250588 320764
rect 249432 320272 249484 320278
rect 249432 320214 249484 320220
rect 251088 320272 251140 320278
rect 251088 320214 251140 320220
rect 249708 320204 249760 320210
rect 249708 320146 249760 320152
rect 249720 315602 249748 320146
rect 251100 315602 251128 320214
rect 251652 320210 251680 322932
rect 252756 320278 252784 322932
rect 253388 320340 253440 320346
rect 253388 320282 253440 320288
rect 252744 320272 252796 320278
rect 252744 320214 252796 320220
rect 251640 320204 251692 320210
rect 251640 320146 251692 320152
rect 252468 320204 252520 320210
rect 252468 320146 252520 320152
rect 248248 315574 248308 315602
rect 249504 315574 249748 315602
rect 250700 315574 251128 315602
rect 252480 315466 252508 320146
rect 253400 315602 253428 320282
rect 253768 320210 253796 322932
rect 254872 320346 254900 322932
rect 254860 320340 254912 320346
rect 254860 320282 254912 320288
rect 255976 320278 256004 322932
rect 256608 320816 256660 320822
rect 256608 320758 256660 320764
rect 254584 320272 254636 320278
rect 254584 320214 254636 320220
rect 255964 320272 256016 320278
rect 255964 320214 256016 320220
rect 253756 320204 253808 320210
rect 253756 320146 253808 320152
rect 254596 315602 254624 320214
rect 255780 320204 255832 320210
rect 255780 320146 255832 320152
rect 255792 315602 255820 320146
rect 253092 315574 253428 315602
rect 254288 315574 254624 315602
rect 255484 315574 255820 315602
rect 256620 315602 256648 320758
rect 256988 320210 257016 322932
rect 258092 320822 258120 322932
rect 258080 320816 258132 320822
rect 258080 320758 258132 320764
rect 259196 320278 259224 322932
rect 257988 320272 258040 320278
rect 257988 320214 258040 320220
rect 259184 320272 259236 320278
rect 259184 320214 259236 320220
rect 256976 320204 257028 320210
rect 256976 320146 257028 320152
rect 258000 315602 258028 320214
rect 260300 320210 260328 322932
rect 260852 322918 261326 322946
rect 262232 322918 262430 322946
rect 259368 320204 259420 320210
rect 259368 320146 259420 320152
rect 260288 320204 260340 320210
rect 260852 320192 260880 322918
rect 262232 320192 262260 322918
rect 263520 320210 263548 322932
rect 264532 320210 264560 322932
rect 264992 322918 265650 322946
rect 266372 322918 266754 322946
rect 267752 322918 267858 322946
rect 260288 320146 260340 320152
rect 260760 320164 260880 320192
rect 262140 320164 262260 320192
rect 263508 320204 263560 320210
rect 259380 315602 259408 320146
rect 256620 315574 256680 315602
rect 257876 315574 258028 315602
rect 259072 315574 259408 315602
rect 260760 315466 260788 320164
rect 262140 315466 262168 320164
rect 263508 320146 263560 320152
rect 263600 320204 263652 320210
rect 263600 320146 263652 320152
rect 264520 320204 264572 320210
rect 264520 320146 264572 320152
rect 262220 320068 262272 320074
rect 262220 320010 262272 320016
rect 262232 315602 262260 320010
rect 263612 315602 263640 320146
rect 264992 315602 265020 322918
rect 266372 320192 266400 322918
rect 267752 320906 267780 322918
rect 266280 320164 266400 320192
rect 267660 320878 267780 320906
rect 266280 315602 266308 320164
rect 267660 315602 267688 320878
rect 268856 320210 268884 322932
rect 269960 320210 269988 322932
rect 270512 322918 271078 322946
rect 271892 322918 272090 322946
rect 267740 320204 267792 320210
rect 267740 320146 267792 320152
rect 268844 320204 268896 320210
rect 268844 320146 268896 320152
rect 269120 320204 269172 320210
rect 269120 320146 269172 320152
rect 269948 320204 270000 320210
rect 269948 320146 270000 320152
rect 262232 315574 262660 315602
rect 263612 315574 263856 315602
rect 264992 315574 265052 315602
rect 266248 315574 266308 315602
rect 267444 315574 267688 315602
rect 224388 315438 224908 315466
rect 225584 315438 226104 315466
rect 233956 315438 234568 315466
rect 251896 315438 252508 315466
rect 260268 315438 260788 315466
rect 261464 315438 262168 315466
rect 267752 315466 267780 320146
rect 269132 315466 269160 320146
rect 270512 315466 270540 322918
rect 271892 315602 271920 322918
rect 273180 320226 273208 322932
rect 273180 320198 273300 320226
rect 273272 315602 273300 320198
rect 274284 315602 274312 322932
rect 275388 315602 275416 322932
rect 276032 322918 276414 322946
rect 277412 322918 277518 322946
rect 278622 322918 278728 322946
rect 276032 320210 276060 322918
rect 277412 320210 277440 322918
rect 278700 320210 278728 322918
rect 279516 320884 279568 320890
rect 279516 320826 279568 320832
rect 276020 320204 276072 320210
rect 276020 320146 276072 320152
rect 276664 320204 276716 320210
rect 276664 320146 276716 320152
rect 277400 320204 277452 320210
rect 277400 320146 277452 320152
rect 277860 320204 277912 320210
rect 277860 320146 277912 320152
rect 278688 320204 278740 320210
rect 278688 320146 278740 320152
rect 279056 320204 279108 320210
rect 279056 320146 279108 320152
rect 276676 315602 276704 320146
rect 277872 315602 277900 320146
rect 279068 315602 279096 320146
rect 271892 315574 272228 315602
rect 273272 315574 273424 315602
rect 274284 315574 274620 315602
rect 275388 315574 275816 315602
rect 276676 315574 277012 315602
rect 277872 315574 278208 315602
rect 279068 315574 279404 315602
rect 267752 315438 268640 315466
rect 269132 315438 269836 315466
rect 270512 315438 271032 315466
rect 279528 295905 279556 320826
rect 280356 317665 280384 326975
rect 282196 322153 282224 700470
rect 282460 700460 282512 700466
rect 282460 700402 282512 700408
rect 282368 700392 282420 700398
rect 282368 700334 282420 700340
rect 282276 700324 282328 700330
rect 282276 700266 282328 700272
rect 282288 586129 282316 700266
rect 282380 614106 282408 700334
rect 282368 614100 282420 614106
rect 282368 614042 282420 614048
rect 282274 586120 282330 586129
rect 282274 586055 282330 586064
rect 282276 569900 282328 569906
rect 282276 569842 282328 569848
rect 282288 569226 282316 569842
rect 282276 569220 282328 569226
rect 282276 569162 282328 569168
rect 282274 430536 282330 430545
rect 282274 430471 282330 430480
rect 282288 421598 282316 430471
rect 282276 421592 282328 421598
rect 282276 421534 282328 421540
rect 282276 377052 282328 377058
rect 282276 376994 282328 377000
rect 282288 360194 282316 376994
rect 282472 369889 282500 700402
rect 283944 698290 283972 703446
rect 332520 700602 332548 703520
rect 348804 700641 348832 703520
rect 348790 700632 348846 700641
rect 305644 700596 305696 700602
rect 305644 700538 305696 700544
rect 332508 700596 332560 700602
rect 348790 700567 348846 700576
rect 332508 700538 332560 700544
rect 301504 700528 301556 700534
rect 301504 700470 301556 700476
rect 283288 698284 283340 698290
rect 283288 698226 283340 698232
rect 283932 698284 283984 698290
rect 283932 698226 283984 698232
rect 283300 694142 283328 698226
rect 283104 694136 283156 694142
rect 283104 694078 283156 694084
rect 283288 694136 283340 694142
rect 283288 694078 283340 694084
rect 283116 692782 283144 694078
rect 283104 692776 283156 692782
rect 283104 692718 283156 692724
rect 283288 692776 283340 692782
rect 283288 692718 283340 692724
rect 283300 683233 283328 692718
rect 282918 683224 282974 683233
rect 282918 683159 282974 683168
rect 283286 683224 283342 683233
rect 283286 683159 283342 683168
rect 282932 683126 282960 683159
rect 282920 683120 282972 683126
rect 282920 683062 282972 683068
rect 287704 667956 287756 667962
rect 287704 667898 287756 667904
rect 283380 666596 283432 666602
rect 283380 666538 283432 666544
rect 283392 659682 283420 666538
rect 283208 659654 283420 659682
rect 283208 647290 283236 659654
rect 283104 647284 283156 647290
rect 283104 647226 283156 647232
rect 283196 647284 283248 647290
rect 283196 647226 283248 647232
rect 283116 640422 283144 647226
rect 283104 640416 283156 640422
rect 283104 640358 283156 640364
rect 283196 640416 283248 640422
rect 283196 640358 283248 640364
rect 283208 630698 283236 640358
rect 283012 630692 283064 630698
rect 283012 630634 283064 630640
rect 283196 630692 283248 630698
rect 283196 630634 283248 630640
rect 283024 630578 283052 630634
rect 283024 630550 283144 630578
rect 283116 621058 283144 630550
rect 283116 621030 283236 621058
rect 283208 611386 283236 621030
rect 283012 611380 283064 611386
rect 283012 611322 283064 611328
rect 283196 611380 283248 611386
rect 283196 611322 283248 611328
rect 283024 611266 283052 611322
rect 283024 611238 283144 611266
rect 283116 601746 283144 611238
rect 284298 608832 284354 608841
rect 284298 608767 284354 608776
rect 283116 601718 283236 601746
rect 283208 598942 283236 601718
rect 283196 598936 283248 598942
rect 283196 598878 283248 598884
rect 283012 589348 283064 589354
rect 283012 589290 283064 589296
rect 283024 579698 283052 589290
rect 283012 579692 283064 579698
rect 283012 579634 283064 579640
rect 283104 579692 283156 579698
rect 283104 579634 283156 579640
rect 283116 578241 283144 579634
rect 283102 578232 283158 578241
rect 283102 578167 283158 578176
rect 283286 578232 283342 578241
rect 283286 578167 283342 578176
rect 283300 560318 283328 578167
rect 284312 569906 284340 608767
rect 284300 569900 284352 569906
rect 284300 569842 284352 569848
rect 286324 569220 286376 569226
rect 286324 569162 286376 569168
rect 283196 560312 283248 560318
rect 283196 560254 283248 560260
rect 283288 560312 283340 560318
rect 283288 560254 283340 560260
rect 283208 553330 283236 560254
rect 283116 553302 283236 553330
rect 283116 550633 283144 553302
rect 282918 550624 282974 550633
rect 282918 550559 282974 550568
rect 283102 550624 283158 550633
rect 283102 550559 283158 550568
rect 282932 541006 282960 550559
rect 282920 541000 282972 541006
rect 282920 540942 282972 540948
rect 283196 541000 283248 541006
rect 283196 540942 283248 540948
rect 282826 527368 282882 527377
rect 282826 527303 282882 527312
rect 282840 527218 282868 527303
rect 283010 527232 283066 527241
rect 282840 527190 283010 527218
rect 283010 527167 283066 527176
rect 283208 518945 283236 540942
rect 282918 518936 282974 518945
rect 282918 518871 282974 518880
rect 283194 518936 283250 518945
rect 283194 518871 283250 518880
rect 282932 514758 282960 518871
rect 282920 514752 282972 514758
rect 282920 514694 282972 514700
rect 283104 514752 283156 514758
rect 283104 514694 283156 514700
rect 283116 509250 283144 514694
rect 283104 509244 283156 509250
rect 283104 509186 283156 509192
rect 283012 499588 283064 499594
rect 283012 499530 283064 499536
rect 283024 495446 283052 499530
rect 283012 495440 283064 495446
rect 283012 495382 283064 495388
rect 283196 495440 283248 495446
rect 283196 495382 283248 495388
rect 283208 492658 283236 495382
rect 282920 492652 282972 492658
rect 282920 492594 282972 492600
rect 283196 492652 283248 492658
rect 283196 492594 283248 492600
rect 282932 483041 282960 492594
rect 282918 483032 282974 483041
rect 282918 482967 282974 482976
rect 283102 483032 283158 483041
rect 283102 482967 283158 482976
rect 283116 473226 283144 482967
rect 283116 473198 283328 473226
rect 283300 471986 283328 473198
rect 283104 471980 283156 471986
rect 283104 471922 283156 471928
rect 283288 471980 283340 471986
rect 283288 471922 283340 471928
rect 283116 462330 283144 471922
rect 283104 462324 283156 462330
rect 283104 462266 283156 462272
rect 283196 452668 283248 452674
rect 283196 452610 283248 452616
rect 283208 447166 283236 452610
rect 283012 447160 283064 447166
rect 283012 447102 283064 447108
rect 283196 447160 283248 447166
rect 283196 447102 283248 447108
rect 283024 437578 283052 447102
rect 283012 437572 283064 437578
rect 283012 437514 283064 437520
rect 282920 434852 282972 434858
rect 282920 434794 282972 434800
rect 282932 433294 282960 434794
rect 282920 433288 282972 433294
rect 282920 433230 282972 433236
rect 283012 423700 283064 423706
rect 283012 423642 283064 423648
rect 283024 418146 283052 423642
rect 283024 418118 283144 418146
rect 283116 415410 283144 418118
rect 283104 415404 283156 415410
rect 283104 415346 283156 415352
rect 283196 405748 283248 405754
rect 283196 405690 283248 405696
rect 283208 402354 283236 405690
rect 283196 402348 283248 402354
rect 283196 402290 283248 402296
rect 284298 392728 284354 392737
rect 284298 392663 284354 392672
rect 284312 377058 284340 392663
rect 284300 377052 284352 377058
rect 284300 376994 284352 377000
rect 282458 369880 282514 369889
rect 282458 369815 282514 369824
rect 282276 360188 282328 360194
rect 282276 360130 282328 360136
rect 282552 360188 282604 360194
rect 282552 360130 282604 360136
rect 282564 360097 282592 360130
rect 282550 360088 282606 360097
rect 282550 360023 282606 360032
rect 282564 357406 282592 360023
rect 282552 357400 282604 357406
rect 282552 357342 282604 357348
rect 282368 347812 282420 347818
rect 282368 347754 282420 347760
rect 282380 340898 282408 347754
rect 282288 340870 282408 340898
rect 282288 336025 282316 340870
rect 282274 336016 282330 336025
rect 282274 335951 282330 335960
rect 282182 322144 282238 322153
rect 282182 322079 282238 322088
rect 282288 321994 282316 335951
rect 282104 321966 282316 321994
rect 280342 317656 280398 317665
rect 280342 317591 280398 317600
rect 280342 317384 280398 317393
rect 280342 317319 280398 317328
rect 280356 309641 280384 317319
rect 280342 309632 280398 309641
rect 280342 309567 280398 309576
rect 282104 309126 282132 321966
rect 282092 309120 282144 309126
rect 282092 309062 282144 309068
rect 282552 299532 282604 299538
rect 282552 299474 282604 299480
rect 279514 295896 279570 295905
rect 279514 295831 279570 295840
rect 280710 295080 280766 295089
rect 280710 295015 280766 295024
rect 280724 277681 280752 295015
rect 282564 292602 282592 299474
rect 282368 292596 282420 292602
rect 282368 292538 282420 292544
rect 282552 292596 282604 292602
rect 282552 292538 282604 292544
rect 282380 278798 282408 292538
rect 282276 278792 282328 278798
rect 282276 278734 282328 278740
rect 282368 278792 282420 278798
rect 282368 278734 282420 278740
rect 280710 277672 280766 277681
rect 280710 277607 280766 277616
rect 282288 273306 282316 278734
rect 282288 273278 282408 273306
rect 282380 263634 282408 273278
rect 282184 263628 282236 263634
rect 282184 263570 282236 263576
rect 282368 263628 282420 263634
rect 282368 263570 282420 263576
rect 282196 255105 282224 263570
rect 282182 255096 282238 255105
rect 282182 255031 282238 255040
rect 280526 251152 280582 251161
rect 280526 251087 280582 251096
rect 280540 241641 280568 251087
rect 280526 241632 280582 241641
rect 280526 241567 280582 241576
rect 209778 235240 209834 235249
rect 209778 235175 209834 235184
rect 250442 235240 250498 235249
rect 250442 235175 250498 235184
rect 205822 233880 205878 233889
rect 205822 233815 205878 233824
rect 205730 229800 205786 229809
rect 205730 229735 205786 229744
rect 204534 228304 204590 228313
rect 204534 228239 204590 228248
rect 193864 224936 193916 224942
rect 193864 224878 193916 224884
rect 189540 224596 189592 224602
rect 189540 224538 189592 224544
rect 186320 224392 186372 224398
rect 186320 224334 186372 224340
rect 188436 224392 188488 224398
rect 188436 224334 188488 224340
rect 186332 221748 186360 224334
rect 188528 223984 188580 223990
rect 188528 223926 188580 223932
rect 187424 223712 187476 223718
rect 187424 223654 187476 223660
rect 187436 221748 187464 223654
rect 188540 221748 188568 223926
rect 189552 221748 189580 224538
rect 190644 224460 190696 224466
rect 190644 224402 190696 224408
rect 190656 221748 190684 224402
rect 192760 224188 192812 224194
rect 192760 224130 192812 224136
rect 191748 223848 191800 223854
rect 191748 223790 191800 223796
rect 191760 221748 191788 223790
rect 192772 221748 192800 224130
rect 193876 221748 193904 224878
rect 194876 224868 194928 224874
rect 194876 224810 194928 224816
rect 194888 221748 194916 224810
rect 198096 224800 198148 224806
rect 198096 224742 198148 224748
rect 195980 224256 196032 224262
rect 195980 224198 196032 224204
rect 195992 221748 196020 224198
rect 197084 224120 197136 224126
rect 197084 224062 197136 224068
rect 197096 221748 197124 224062
rect 198108 221748 198136 224742
rect 202420 224732 202472 224738
rect 202420 224674 202472 224680
rect 201316 224664 201368 224670
rect 201316 224606 201368 224612
rect 199200 224528 199252 224534
rect 199200 224470 199252 224476
rect 199212 221748 199240 224470
rect 200304 224324 200356 224330
rect 200304 224266 200356 224272
rect 200316 221748 200344 224266
rect 201328 221748 201356 224606
rect 202432 221748 202460 224674
rect 203432 224392 203484 224398
rect 203432 224334 203484 224340
rect 203444 221748 203472 224334
rect 204548 221748 204576 228239
rect 205744 221762 205772 229735
rect 205666 221734 205772 221762
rect 205836 221626 205864 233815
rect 207018 232520 207074 232529
rect 207018 232455 207074 232464
rect 207032 221626 207060 232455
rect 208858 223680 208914 223689
rect 208858 223615 208914 223624
rect 208872 221748 208900 223615
rect 209792 221762 209820 235175
rect 214564 233912 214616 233918
rect 214564 233854 214616 233860
rect 214576 231826 214604 233854
rect 214484 231798 214604 231826
rect 214484 225010 214512 231798
rect 214748 229764 214800 229770
rect 214748 229706 214800 229712
rect 214656 225684 214708 225690
rect 214656 225626 214708 225632
rect 214472 225004 214524 225010
rect 214472 224946 214524 224952
rect 210976 224256 211028 224262
rect 210976 224198 211028 224204
rect 209792 221734 209898 221762
rect 210988 221748 211016 224198
rect 214472 222216 214524 222222
rect 214472 222158 214524 222164
rect 214484 222086 214512 222158
rect 214472 222080 214524 222086
rect 214472 222022 214524 222028
rect 121564 221598 122222 221626
rect 205836 221598 206678 221626
rect 207032 221598 207782 221626
rect 213918 221368 213974 221377
rect 213918 221303 213974 221312
rect 213932 220862 213960 221303
rect 213920 220856 213972 220862
rect 213920 220798 213972 220804
rect 214010 220552 214066 220561
rect 214010 220487 214066 220496
rect 214024 220182 214052 220487
rect 214012 220176 214064 220182
rect 214012 220118 214064 220124
rect 116676 220108 116728 220114
rect 116676 220050 116728 220056
rect 213920 220108 213972 220114
rect 213920 220050 213972 220056
rect 116688 130121 116716 220050
rect 213932 219745 213960 220050
rect 213918 219736 213974 219745
rect 213918 219671 213974 219680
rect 213918 218920 213974 218929
rect 213918 218855 213974 218864
rect 213932 218822 213960 218855
rect 213920 218816 213972 218822
rect 213920 218758 213972 218764
rect 214012 218748 214064 218754
rect 214012 218690 214064 218696
rect 214024 218249 214052 218690
rect 214010 218240 214066 218249
rect 214010 218175 214066 218184
rect 213918 217424 213974 217433
rect 213918 217359 213974 217368
rect 213932 217326 213960 217359
rect 213920 217320 213972 217326
rect 213920 217262 213972 217268
rect 213920 216640 213972 216646
rect 213918 216608 213920 216617
rect 213972 216608 213974 216617
rect 213918 216543 213974 216552
rect 213920 215960 213972 215966
rect 213920 215902 213972 215908
rect 213932 215801 213960 215902
rect 213918 215792 213974 215801
rect 213918 215727 213974 215736
rect 213920 215280 213972 215286
rect 213920 215222 213972 215228
rect 213932 215121 213960 215222
rect 214012 215212 214064 215218
rect 214012 215154 214064 215160
rect 213918 215112 213974 215121
rect 213918 215047 213974 215056
rect 214024 214305 214052 215154
rect 214010 214296 214066 214305
rect 214010 214231 214066 214240
rect 213920 213920 213972 213926
rect 213920 213862 213972 213868
rect 213932 213489 213960 213862
rect 214012 213852 214064 213858
rect 214012 213794 214064 213800
rect 213918 213480 213974 213489
rect 213918 213415 213974 213424
rect 214024 212673 214052 213794
rect 214010 212664 214066 212673
rect 214010 212599 214066 212608
rect 214564 212560 214616 212566
rect 214484 212508 214564 212514
rect 214484 212502 214616 212508
rect 213920 212492 213972 212498
rect 213920 212434 213972 212440
rect 214484 212486 214604 212502
rect 213932 211993 213960 212434
rect 214012 212424 214064 212430
rect 214012 212366 214064 212372
rect 213918 211984 213974 211993
rect 213918 211919 213974 211928
rect 214024 211177 214052 212366
rect 214010 211168 214066 211177
rect 213920 211132 213972 211138
rect 214010 211103 214066 211112
rect 213920 211074 213972 211080
rect 213932 210361 213960 211074
rect 213918 210352 213974 210361
rect 213918 210287 213974 210296
rect 214012 209772 214064 209778
rect 214012 209714 214064 209720
rect 213920 209704 213972 209710
rect 213920 209646 213972 209652
rect 213932 209545 213960 209646
rect 213918 209536 213974 209545
rect 213918 209471 213974 209480
rect 214024 208865 214052 209714
rect 214010 208856 214066 208865
rect 214010 208791 214066 208800
rect 214012 208344 214064 208350
rect 214012 208286 214064 208292
rect 213920 208276 213972 208282
rect 213920 208218 213972 208224
rect 213932 208049 213960 208218
rect 213918 208040 213974 208049
rect 213918 207975 213974 207984
rect 214024 207233 214052 208286
rect 214010 207224 214066 207233
rect 214010 207159 214066 207168
rect 213920 206984 213972 206990
rect 213920 206926 213972 206932
rect 213932 206417 213960 206926
rect 214012 206916 214064 206922
rect 214012 206858 214064 206864
rect 213918 206408 213974 206417
rect 213918 206343 213974 206352
rect 214024 205737 214052 206858
rect 214010 205728 214066 205737
rect 214484 205698 214512 212486
rect 214010 205663 214066 205672
rect 214472 205692 214524 205698
rect 214472 205634 214524 205640
rect 213920 205624 213972 205630
rect 213920 205566 213972 205572
rect 213932 204921 213960 205566
rect 213918 204912 213974 204921
rect 213918 204847 213974 204856
rect 214012 204264 214064 204270
rect 214012 204206 214064 204212
rect 213920 204196 213972 204202
rect 213920 204138 213972 204144
rect 213932 204105 213960 204138
rect 213918 204096 213974 204105
rect 213918 204031 213974 204040
rect 214024 203289 214052 204206
rect 214010 203280 214066 203289
rect 214010 203215 214066 203224
rect 214472 202904 214524 202910
rect 214472 202846 214524 202852
rect 213920 202836 213972 202842
rect 213920 202778 213972 202784
rect 213932 202473 213960 202778
rect 214012 202768 214064 202774
rect 214012 202710 214064 202716
rect 213918 202464 213974 202473
rect 213918 202399 213974 202408
rect 214024 201793 214052 202710
rect 214010 201784 214066 201793
rect 214010 201719 214066 201728
rect 213920 201476 213972 201482
rect 213920 201418 213972 201424
rect 213932 200977 213960 201418
rect 214012 201408 214064 201414
rect 214012 201350 214064 201356
rect 213918 200968 213974 200977
rect 213918 200903 213974 200912
rect 214024 200161 214052 201350
rect 214484 200598 214512 202846
rect 214472 200592 214524 200598
rect 214472 200534 214524 200540
rect 214010 200152 214066 200161
rect 213920 200116 213972 200122
rect 214010 200087 214066 200096
rect 213920 200058 213972 200064
rect 213932 199345 213960 200058
rect 213918 199336 213974 199345
rect 213918 199271 213974 199280
rect 214012 198688 214064 198694
rect 213918 198656 213974 198665
rect 214012 198630 214064 198636
rect 213918 198591 213920 198600
rect 213972 198591 213974 198600
rect 213920 198562 213972 198568
rect 214024 197849 214052 198630
rect 214010 197840 214066 197849
rect 214010 197775 214066 197784
rect 214012 197328 214064 197334
rect 214012 197270 214064 197276
rect 213920 197260 213972 197266
rect 213920 197202 213972 197208
rect 213932 197033 213960 197202
rect 213918 197024 213974 197033
rect 213918 196959 213974 196968
rect 214024 196217 214052 197270
rect 214010 196208 214066 196217
rect 214010 196143 214066 196152
rect 213920 195968 213972 195974
rect 213920 195910 213972 195916
rect 213932 195537 213960 195910
rect 214012 195900 214064 195906
rect 214012 195842 214064 195848
rect 213918 195528 213974 195537
rect 213918 195463 213974 195472
rect 214024 194721 214052 195842
rect 214010 194712 214066 194721
rect 214010 194647 214066 194656
rect 214196 194608 214248 194614
rect 214196 194550 214248 194556
rect 213920 194540 213972 194546
rect 213920 194482 213972 194488
rect 213932 193905 213960 194482
rect 213918 193896 213974 193905
rect 213918 193831 213974 193840
rect 213920 193180 213972 193186
rect 213920 193122 213972 193128
rect 213932 193089 213960 193122
rect 214012 193112 214064 193118
rect 213918 193080 213974 193089
rect 214012 193054 214064 193060
rect 213918 193015 213974 193024
rect 214024 192409 214052 193054
rect 214010 192400 214066 192409
rect 214010 192335 214066 192344
rect 214104 191888 214156 191894
rect 214104 191830 214156 191836
rect 214012 191820 214064 191826
rect 214012 191762 214064 191768
rect 213920 191752 213972 191758
rect 213920 191694 213972 191700
rect 213932 191593 213960 191694
rect 213918 191584 213974 191593
rect 213918 191519 213974 191528
rect 214024 190777 214052 191762
rect 214010 190768 214066 190777
rect 214010 190703 214066 190712
rect 214012 190460 214064 190466
rect 214012 190402 214064 190408
rect 213920 190392 213972 190398
rect 213920 190334 213972 190340
rect 213932 189961 213960 190334
rect 213918 189952 213974 189961
rect 213918 189887 213974 189896
rect 214024 189281 214052 190402
rect 214010 189272 214066 189281
rect 214010 189207 214066 189216
rect 213920 189032 213972 189038
rect 213920 188974 213972 188980
rect 213932 188465 213960 188974
rect 213918 188456 213974 188465
rect 213918 188391 213974 188400
rect 213918 186824 213974 186833
rect 213918 186759 213974 186768
rect 213932 186590 213960 186759
rect 213920 186584 213972 186590
rect 213920 186526 213972 186532
rect 213918 185328 213974 185337
rect 213918 185263 213974 185272
rect 213932 185094 213960 185263
rect 213920 185088 213972 185094
rect 213920 185030 213972 185036
rect 214012 184952 214064 184958
rect 214012 184894 214064 184900
rect 213920 183592 213972 183598
rect 213920 183534 213972 183540
rect 213932 180690 213960 183534
rect 214024 180826 214052 184894
rect 214116 184521 214144 191830
rect 214208 187649 214236 194550
rect 214472 193248 214524 193254
rect 214472 193190 214524 193196
rect 214288 190596 214340 190602
rect 214288 190538 214340 190544
rect 214194 187640 214250 187649
rect 214194 187575 214250 187584
rect 214196 186380 214248 186386
rect 214196 186322 214248 186328
rect 214102 184512 214158 184521
rect 214102 184447 214158 184456
rect 214208 181506 214236 186322
rect 214300 181937 214328 190538
rect 214380 189100 214432 189106
rect 214380 189042 214432 189048
rect 214286 181928 214342 181937
rect 214286 181863 214342 181872
rect 214208 181478 214328 181506
rect 214024 180798 214236 180826
rect 213932 180662 214144 180690
rect 213920 180600 213972 180606
rect 213918 180568 213920 180577
rect 213972 180568 213974 180577
rect 213918 180503 213974 180512
rect 214012 179376 214064 179382
rect 214012 179318 214064 179324
rect 213920 179104 213972 179110
rect 213918 179072 213920 179081
rect 213972 179072 213974 179081
rect 213918 179007 213974 179016
rect 214024 178265 214052 179318
rect 214010 178256 214066 178265
rect 214010 178191 214066 178200
rect 213920 178016 213972 178022
rect 213920 177958 213972 177964
rect 213932 177449 213960 177958
rect 213918 177440 213974 177449
rect 213918 177375 213974 177384
rect 214116 177290 214144 180662
rect 213932 177262 214144 177290
rect 213932 174434 213960 177262
rect 214012 176656 214064 176662
rect 214012 176598 214064 176604
rect 214024 175953 214052 176598
rect 214010 175944 214066 175953
rect 214010 175879 214066 175888
rect 214208 175137 214236 180798
rect 214300 176633 214328 181478
rect 214392 179761 214420 189042
rect 214484 186017 214512 193190
rect 214470 186008 214526 186017
rect 214470 185943 214526 185952
rect 214472 182368 214524 182374
rect 214472 182310 214524 182316
rect 214378 179752 214434 179761
rect 214378 179687 214434 179696
rect 214484 178140 214512 182310
rect 214392 178112 214512 178140
rect 214286 176624 214342 176633
rect 214286 176559 214342 176568
rect 214194 175128 214250 175137
rect 214194 175063 214250 175072
rect 213932 174406 214052 174434
rect 213918 174312 213974 174321
rect 213918 174247 213974 174256
rect 213932 174214 213960 174247
rect 213920 174208 213972 174214
rect 213920 174150 213972 174156
rect 213920 173868 213972 173874
rect 213920 173810 213972 173816
rect 213932 172825 213960 173810
rect 214024 173505 214052 174406
rect 214194 173904 214250 173913
rect 214194 173839 214250 173848
rect 214010 173496 214066 173505
rect 214010 173431 214066 173440
rect 213918 172816 213974 172825
rect 213918 172751 213974 172760
rect 213920 172508 213972 172514
rect 213920 172450 213972 172456
rect 213932 171193 213960 172450
rect 213918 171184 213974 171193
rect 213918 171119 213974 171128
rect 213918 169552 213974 169561
rect 213918 169487 213974 169496
rect 213932 169114 213960 169487
rect 213920 169108 213972 169114
rect 213920 169050 213972 169056
rect 213920 168360 213972 168366
rect 213920 168302 213972 168308
rect 213932 168065 213960 168302
rect 213918 168056 213974 168065
rect 213918 167991 213974 168000
rect 213920 167000 213972 167006
rect 213920 166942 213972 166948
rect 213932 166433 213960 166942
rect 214208 166938 214236 173839
rect 214392 172009 214420 178112
rect 214472 173936 214524 173942
rect 214470 173904 214472 173913
rect 214524 173904 214526 173913
rect 214470 173839 214526 173848
rect 214378 172000 214434 172009
rect 214378 171935 214434 171944
rect 214196 166932 214248 166938
rect 214196 166874 214248 166880
rect 214472 166932 214524 166938
rect 214472 166874 214524 166880
rect 214012 166592 214064 166598
rect 214012 166534 214064 166540
rect 213918 166424 213974 166433
rect 213918 166359 213974 166368
rect 214024 165753 214052 166534
rect 214010 165744 214066 165753
rect 214010 165679 214066 165688
rect 213920 165572 213972 165578
rect 213920 165514 213972 165520
rect 213932 164937 213960 165514
rect 213918 164928 213974 164937
rect 213918 164863 213974 164872
rect 214484 164234 214512 166874
rect 214484 164206 214604 164234
rect 213920 164144 213972 164150
rect 213918 164112 213920 164121
rect 213972 164112 213974 164121
rect 213918 164047 213974 164056
rect 213920 163600 213972 163606
rect 213920 163542 213972 163548
rect 213932 163305 213960 163542
rect 213918 163296 213974 163305
rect 213918 163231 213974 163240
rect 213920 162852 213972 162858
rect 213920 162794 213972 162800
rect 213932 162625 213960 162794
rect 213918 162616 213974 162625
rect 213918 162551 213974 162560
rect 213920 162308 213972 162314
rect 213920 162250 213972 162256
rect 213932 161809 213960 162250
rect 213918 161800 213974 161809
rect 213918 161735 213974 161744
rect 213920 161424 213972 161430
rect 213920 161366 213972 161372
rect 213932 160993 213960 161366
rect 213918 160984 213974 160993
rect 213918 160919 213974 160928
rect 213920 160880 213972 160886
rect 213920 160822 213972 160828
rect 213932 160177 213960 160822
rect 213918 160168 213974 160177
rect 213918 160103 213974 160112
rect 213918 157040 213974 157049
rect 213918 156975 213974 156984
rect 213932 155990 213960 156975
rect 214102 156360 214158 156369
rect 214102 156295 214158 156304
rect 213920 155984 213972 155990
rect 213920 155926 213972 155932
rect 213918 155544 213974 155553
rect 213918 155479 213974 155488
rect 213932 154630 213960 155479
rect 213920 154624 213972 154630
rect 213920 154566 213972 154572
rect 214010 153912 214066 153921
rect 214010 153847 214066 153856
rect 213920 153332 213972 153338
rect 213920 153274 213972 153280
rect 213932 153241 213960 153274
rect 214024 153270 214052 153847
rect 214012 153264 214064 153270
rect 213918 153232 213974 153241
rect 214012 153206 214064 153212
rect 213918 153167 213974 153176
rect 213918 152416 213974 152425
rect 213918 152351 213974 152360
rect 213932 151910 213960 152351
rect 213920 151904 213972 151910
rect 213920 151846 213972 151852
rect 213918 151600 213974 151609
rect 213918 151535 213974 151544
rect 213932 150890 213960 151535
rect 213920 150884 213972 150890
rect 213920 150826 213972 150832
rect 213918 150784 213974 150793
rect 213918 150719 213974 150728
rect 213932 150482 213960 150719
rect 213920 150476 213972 150482
rect 213920 150418 213972 150424
rect 213918 149968 213974 149977
rect 213918 149903 213974 149912
rect 213932 149394 213960 149903
rect 213920 149388 213972 149394
rect 213920 149330 213972 149336
rect 213918 149288 213974 149297
rect 213918 149223 213974 149232
rect 213932 149122 213960 149223
rect 213920 149116 213972 149122
rect 213920 149058 213972 149064
rect 214116 149054 214144 156295
rect 214104 149048 214156 149054
rect 214104 148990 214156 148996
rect 213918 148472 213974 148481
rect 213918 148407 213974 148416
rect 213932 148034 213960 148407
rect 214576 148374 214604 164206
rect 214564 148368 214616 148374
rect 214564 148310 214616 148316
rect 213920 148028 213972 148034
rect 213920 147970 213972 147976
rect 214010 147656 214066 147665
rect 214010 147591 214066 147600
rect 213918 146840 213974 146849
rect 213918 146775 213974 146784
rect 213932 146402 213960 146775
rect 213920 146396 213972 146402
rect 213920 146338 213972 146344
rect 214024 146334 214052 147591
rect 214012 146328 214064 146334
rect 214012 146270 214064 146276
rect 214010 146160 214066 146169
rect 214010 146095 214066 146104
rect 213918 145344 213974 145353
rect 213918 145279 213974 145288
rect 213932 145042 213960 145279
rect 213920 145036 213972 145042
rect 213920 144978 213972 144984
rect 214024 144974 214052 146095
rect 214012 144968 214064 144974
rect 214012 144910 214064 144916
rect 214010 144528 214066 144537
rect 214010 144463 214066 144472
rect 213918 143712 213974 143721
rect 213918 143647 213920 143656
rect 213972 143647 213974 143656
rect 213920 143618 213972 143624
rect 214024 143614 214052 144463
rect 214012 143608 214064 143614
rect 214012 143550 214064 143556
rect 214562 143576 214618 143585
rect 214562 143511 214618 143520
rect 214576 143478 214604 143511
rect 214380 143472 214432 143478
rect 214380 143414 214432 143420
rect 214564 143472 214616 143478
rect 214564 143414 214616 143420
rect 214010 143032 214066 143041
rect 214010 142967 214066 142976
rect 213920 142248 213972 142254
rect 213918 142216 213920 142225
rect 213972 142216 213974 142225
rect 214024 142186 214052 142967
rect 213918 142151 213974 142160
rect 214012 142180 214064 142186
rect 214012 142122 214064 142128
rect 213918 141400 213974 141409
rect 213918 141335 213974 141344
rect 213932 140826 213960 141335
rect 213920 140820 213972 140826
rect 213920 140762 213972 140768
rect 214010 140584 214066 140593
rect 214010 140519 214066 140528
rect 213918 139904 213974 139913
rect 213918 139839 213974 139848
rect 213932 139534 213960 139839
rect 213920 139528 213972 139534
rect 213920 139470 213972 139476
rect 214024 139466 214052 140519
rect 214012 139460 214064 139466
rect 214012 139402 214064 139408
rect 214010 139088 214066 139097
rect 214010 139023 214066 139032
rect 213918 138272 213974 138281
rect 213918 138207 213974 138216
rect 213932 138038 213960 138207
rect 214024 138106 214052 139023
rect 214012 138100 214064 138106
rect 214012 138042 214064 138048
rect 213920 138032 213972 138038
rect 213920 137974 213972 137980
rect 214010 137456 214066 137465
rect 214010 137391 214066 137400
rect 213918 136776 213974 136785
rect 213918 136711 213920 136720
rect 213972 136711 213974 136720
rect 213920 136682 213972 136688
rect 214024 136678 214052 137391
rect 214012 136672 214064 136678
rect 214012 136614 214064 136620
rect 213918 135960 213974 135969
rect 213918 135895 213974 135904
rect 213932 135318 213960 135895
rect 213920 135312 213972 135318
rect 213920 135254 213972 135260
rect 214010 135144 214066 135153
rect 214392 135130 214420 143414
rect 214392 135102 214512 135130
rect 214010 135079 214066 135088
rect 213918 134328 213974 134337
rect 213918 134263 213974 134272
rect 213932 133958 213960 134263
rect 214024 134026 214052 135079
rect 214012 134020 214064 134026
rect 214012 133962 214064 133968
rect 213920 133952 213972 133958
rect 213920 133894 213972 133900
rect 117134 133648 117190 133657
rect 117134 133583 117190 133592
rect 117148 132938 117176 133583
rect 214010 133512 214066 133521
rect 214010 133447 214066 133456
rect 117136 132932 117188 132938
rect 117136 132874 117188 132880
rect 213918 132832 213974 132841
rect 213918 132767 213974 132776
rect 213932 132598 213960 132767
rect 213920 132592 213972 132598
rect 213920 132534 213972 132540
rect 214024 132530 214052 133447
rect 214012 132524 214064 132530
rect 214012 132466 214064 132472
rect 214010 132016 214066 132025
rect 214010 131951 214066 131960
rect 213920 131232 213972 131238
rect 213918 131200 213920 131209
rect 213972 131200 213974 131209
rect 214024 131170 214052 131951
rect 213918 131135 213974 131144
rect 214012 131164 214064 131170
rect 214012 131106 214064 131112
rect 213918 130384 213974 130393
rect 213918 130319 213974 130328
rect 116674 130112 116730 130121
rect 116674 130047 116730 130056
rect 213932 129810 213960 130319
rect 213920 129804 213972 129810
rect 213920 129746 213972 129752
rect 213918 129704 213974 129713
rect 213918 129639 213974 129648
rect 213932 129062 213960 129639
rect 213920 129056 213972 129062
rect 213920 128998 213972 129004
rect 213918 128888 213974 128897
rect 213918 128823 213974 128832
rect 213932 128382 213960 128823
rect 213920 128376 213972 128382
rect 213920 128318 213972 128324
rect 213918 128072 213974 128081
rect 213918 128007 213974 128016
rect 213932 127634 213960 128007
rect 213920 127628 213972 127634
rect 213920 127570 213972 127576
rect 213918 127256 213974 127265
rect 213918 127191 213974 127200
rect 213932 127022 213960 127191
rect 213920 127016 213972 127022
rect 213920 126958 213972 126964
rect 213918 126576 213974 126585
rect 213918 126511 213974 126520
rect 213932 126274 213960 126511
rect 213920 126268 213972 126274
rect 213920 126210 213972 126216
rect 213918 125760 213974 125769
rect 213918 125695 213974 125704
rect 213932 125662 213960 125695
rect 213920 125656 213972 125662
rect 213920 125598 213972 125604
rect 214484 125594 214512 135102
rect 214380 125588 214432 125594
rect 214380 125530 214432 125536
rect 214472 125588 214524 125594
rect 214472 125530 214524 125536
rect 213918 124944 213974 124953
rect 213918 124879 213920 124888
rect 213972 124879 213974 124888
rect 213920 124850 213972 124856
rect 213920 124160 213972 124166
rect 213918 124128 213920 124137
rect 213972 124128 213974 124137
rect 213918 124063 213974 124072
rect 213920 123480 213972 123486
rect 213918 123448 213920 123457
rect 213972 123448 213974 123457
rect 213918 123383 213974 123392
rect 116582 123040 116638 123049
rect 116582 122975 116638 122984
rect 213920 122800 213972 122806
rect 213920 122742 213972 122748
rect 213932 122641 213960 122742
rect 213918 122632 213974 122641
rect 213918 122567 213974 122576
rect 213920 122120 213972 122126
rect 213920 122062 213972 122068
rect 116398 121952 116454 121961
rect 116398 121887 116454 121896
rect 116412 121514 116440 121887
rect 213932 121825 213960 122062
rect 213918 121816 213974 121825
rect 213918 121751 213974 121760
rect 50988 121508 51040 121514
rect 50988 121450 51040 121456
rect 116400 121508 116452 121514
rect 116400 121450 116452 121456
rect 51000 99362 51028 121450
rect 213920 121440 213972 121446
rect 213920 121382 213972 121388
rect 213932 121009 213960 121382
rect 213918 121000 213974 121009
rect 213918 120935 213974 120944
rect 213920 120760 213972 120766
rect 116398 120728 116454 120737
rect 213920 120702 213972 120708
rect 116398 120663 116454 120672
rect 116412 120154 116440 120663
rect 213932 120329 213960 120702
rect 213918 120320 213974 120329
rect 213918 120255 213974 120264
rect 94504 120148 94556 120154
rect 94504 120090 94556 120096
rect 116400 120148 116452 120154
rect 116400 120090 116452 120096
rect 94412 111852 94464 111858
rect 94412 111794 94464 111800
rect 94320 104916 94372 104922
rect 94320 104858 94372 104864
rect 94228 102196 94280 102202
rect 94228 102138 94280 102144
rect 50646 99334 51028 99362
rect 94136 98048 94188 98054
rect 94136 97990 94188 97996
rect 94148 81977 94176 97990
rect 94240 85513 94268 102138
rect 94332 87281 94360 104858
rect 94424 92721 94452 111794
rect 94516 98977 94544 120090
rect 213920 120080 213972 120086
rect 213920 120022 213972 120028
rect 116398 119640 116454 119649
rect 116398 119575 116454 119584
rect 116412 118726 116440 119575
rect 213932 119513 213960 120022
rect 213918 119504 213974 119513
rect 213918 119439 213974 119448
rect 94688 118720 94740 118726
rect 94688 118662 94740 118668
rect 116400 118720 116452 118726
rect 116400 118662 116452 118668
rect 213918 118688 213974 118697
rect 94596 117360 94648 117366
rect 94596 117302 94648 117308
rect 94502 98968 94558 98977
rect 94502 98903 94558 98912
rect 94608 97209 94636 117302
rect 94700 98025 94728 118662
rect 213918 118623 213920 118632
rect 213972 118623 213974 118632
rect 214392 118640 214420 125530
rect 214392 118612 214512 118640
rect 213920 118594 213972 118600
rect 214012 118584 214064 118590
rect 214012 118526 214064 118532
rect 116398 118416 116454 118425
rect 116398 118351 116454 118360
rect 116412 117366 116440 118351
rect 214024 117881 214052 118526
rect 214010 117872 214066 117881
rect 214010 117807 214066 117816
rect 116400 117360 116452 117366
rect 116400 117302 116452 117308
rect 214012 117292 214064 117298
rect 214012 117234 214064 117240
rect 213920 117224 213972 117230
rect 116398 117192 116454 117201
rect 213920 117166 213972 117172
rect 116398 117127 116454 117136
rect 116122 116104 116178 116113
rect 94964 116068 95016 116074
rect 116122 116039 116124 116048
rect 94964 116010 95016 116016
rect 116176 116039 116178 116048
rect 116124 116010 116176 116016
rect 94780 116000 94832 116006
rect 94780 115942 94832 115948
rect 94686 98016 94742 98025
rect 94686 97951 94742 97960
rect 94594 97200 94650 97209
rect 94594 97135 94650 97144
rect 94792 96257 94820 115942
rect 94872 114572 94924 114578
rect 94872 114514 94924 114520
rect 94778 96248 94834 96257
rect 94778 96183 94834 96192
rect 94688 95260 94740 95266
rect 94688 95202 94740 95208
rect 94504 93900 94556 93906
rect 94504 93842 94556 93848
rect 94410 92712 94466 92721
rect 94410 92647 94466 92656
rect 94318 87272 94374 87281
rect 94318 87207 94374 87216
rect 94412 86624 94464 86630
rect 94412 86566 94464 86572
rect 94424 86465 94452 86566
rect 94410 86456 94466 86465
rect 94410 86391 94466 86400
rect 94226 85504 94282 85513
rect 94226 85439 94282 85448
rect 94228 83428 94280 83434
rect 94228 83370 94280 83376
rect 94240 82929 94268 83370
rect 94226 82920 94282 82929
rect 94226 82855 94282 82864
rect 94134 81968 94190 81977
rect 94134 81903 94190 81912
rect 94412 81320 94464 81326
rect 94412 81262 94464 81268
rect 94424 81025 94452 81262
rect 94410 81016 94466 81025
rect 94410 80951 94466 80960
rect 94412 80028 94464 80034
rect 94412 79970 94464 79976
rect 94424 79257 94452 79970
rect 94410 79248 94466 79257
rect 94410 79183 94466 79192
rect 94516 78441 94544 93842
rect 94596 91860 94648 91866
rect 94596 91802 94648 91808
rect 94608 91769 94636 91802
rect 94594 91760 94650 91769
rect 94594 91695 94650 91704
rect 94596 91112 94648 91118
rect 94596 91054 94648 91060
rect 94502 78432 94558 78441
rect 94502 78367 94558 78376
rect 94228 78260 94280 78266
rect 94228 78202 94280 78208
rect 94240 77489 94268 78202
rect 94226 77480 94282 77489
rect 94226 77415 94282 77424
rect 94608 76537 94636 91054
rect 94700 80209 94728 95202
rect 94884 94489 94912 114514
rect 94976 95441 95004 116010
rect 116412 116006 116440 117127
rect 213932 117065 213960 117166
rect 213918 117056 213974 117065
rect 213918 116991 213974 117000
rect 214024 116385 214052 117234
rect 214010 116376 214066 116385
rect 214010 116311 214066 116320
rect 116400 116000 116452 116006
rect 116400 115942 116452 115948
rect 214012 115932 214064 115938
rect 214012 115874 214064 115880
rect 213920 115864 213972 115870
rect 213920 115806 213972 115812
rect 213932 115569 213960 115806
rect 213918 115560 213974 115569
rect 213918 115495 213974 115504
rect 116398 114880 116454 114889
rect 116398 114815 116454 114824
rect 116412 114578 116440 114815
rect 214024 114753 214052 115874
rect 214010 114744 214066 114753
rect 214010 114679 214066 114688
rect 116400 114572 116452 114578
rect 116400 114514 116452 114520
rect 214012 114504 214064 114510
rect 214012 114446 214064 114452
rect 213920 114436 213972 114442
rect 213920 114378 213972 114384
rect 213932 113937 213960 114378
rect 213918 113928 213974 113937
rect 213918 113863 213974 113872
rect 116398 113792 116454 113801
rect 116398 113727 116454 113736
rect 116412 113218 116440 113727
rect 214024 113257 214052 114446
rect 214010 113248 214066 113257
rect 97264 113212 97316 113218
rect 97264 113154 97316 113160
rect 116400 113212 116452 113218
rect 214010 113183 214066 113192
rect 116400 113154 116452 113160
rect 95884 110492 95936 110498
rect 95884 110434 95936 110440
rect 95148 109064 95200 109070
rect 95148 109006 95200 109012
rect 95056 107704 95108 107710
rect 95056 107646 95108 107652
rect 94962 95432 95018 95441
rect 94962 95367 95018 95376
rect 94870 94480 94926 94489
rect 94870 94415 94926 94424
rect 95068 93786 95096 107646
rect 94976 93758 95096 93786
rect 94780 91044 94832 91050
rect 94780 90986 94832 90992
rect 94792 90001 94820 90986
rect 94778 89992 94834 90001
rect 94778 89927 94834 89936
rect 94976 89185 95004 93758
rect 95160 93650 95188 109006
rect 95068 93622 95188 93650
rect 95068 90953 95096 93622
rect 95148 93560 95200 93566
rect 95146 93528 95148 93537
rect 95200 93528 95202 93537
rect 95146 93463 95202 93472
rect 95896 91866 95924 110434
rect 97276 93566 97304 113154
rect 213920 113144 213972 113150
rect 213920 113086 213972 113092
rect 116398 112568 116454 112577
rect 116398 112503 116454 112512
rect 116412 111858 116440 112503
rect 213932 112441 213960 113086
rect 213918 112432 213974 112441
rect 213918 112367 213974 112376
rect 116400 111852 116452 111858
rect 116400 111794 116452 111800
rect 214012 111784 214064 111790
rect 214012 111726 214064 111732
rect 213920 111716 213972 111722
rect 213920 111658 213972 111664
rect 213932 111625 213960 111658
rect 213918 111616 213974 111625
rect 213918 111551 213974 111560
rect 116398 111480 116454 111489
rect 116398 111415 116454 111424
rect 116412 110498 116440 111415
rect 214024 110809 214052 111726
rect 214010 110800 214066 110809
rect 214010 110735 214066 110744
rect 116400 110492 116452 110498
rect 116400 110434 116452 110440
rect 214012 110424 214064 110430
rect 214012 110366 214064 110372
rect 213920 110356 213972 110362
rect 213920 110298 213972 110304
rect 116398 110256 116454 110265
rect 116398 110191 116454 110200
rect 116412 109070 116440 110191
rect 213932 110129 213960 110298
rect 213918 110120 213974 110129
rect 213918 110055 213974 110064
rect 214024 109313 214052 110366
rect 214010 109304 214066 109313
rect 214010 109239 214066 109248
rect 116400 109064 116452 109070
rect 116306 109032 116362 109041
rect 214484 109041 214512 118612
rect 116400 109006 116452 109012
rect 214470 109032 214526 109041
rect 116306 108967 116362 108976
rect 214012 108996 214064 109002
rect 116320 107778 116348 108967
rect 214470 108967 214526 108976
rect 214012 108938 214064 108944
rect 213920 108928 213972 108934
rect 213920 108870 213972 108876
rect 213932 108497 213960 108870
rect 213918 108488 213974 108497
rect 213918 108423 213974 108432
rect 116398 107944 116454 107953
rect 116398 107879 116454 107888
rect 102784 107772 102836 107778
rect 102784 107714 102836 107720
rect 116308 107772 116360 107778
rect 116308 107714 116360 107720
rect 98644 106344 98696 106350
rect 98644 106286 98696 106292
rect 97356 99408 97408 99414
rect 97356 99350 97408 99356
rect 97264 93560 97316 93566
rect 97264 93502 97316 93508
rect 95976 92540 96028 92546
rect 95976 92482 96028 92488
rect 95884 91860 95936 91866
rect 95884 91802 95936 91808
rect 95054 90944 95110 90953
rect 95054 90879 95110 90888
rect 94962 89176 95018 89185
rect 94962 89111 95018 89120
rect 94964 88392 95016 88398
rect 94964 88334 95016 88340
rect 94780 85604 94832 85610
rect 94780 85546 94832 85552
rect 94686 80200 94742 80209
rect 94686 80135 94742 80144
rect 94688 77308 94740 77314
rect 94688 77250 94740 77256
rect 94594 76528 94650 76537
rect 94594 76463 94650 76472
rect 94596 75744 94648 75750
rect 94594 75712 94596 75721
rect 94648 75712 94650 75721
rect 94594 75647 94650 75656
rect 94504 74588 94556 74594
rect 94504 74530 94556 74536
rect 94412 72956 94464 72962
rect 94412 72898 94464 72904
rect 94424 72185 94452 72898
rect 94410 72176 94466 72185
rect 94410 72111 94466 72120
rect 94412 69080 94464 69086
rect 94412 69022 94464 69028
rect 93860 68536 93912 68542
rect 93858 68504 93860 68513
rect 93912 68504 93914 68513
rect 93858 68439 93914 68448
rect 94320 64932 94372 64938
rect 94320 64874 94372 64880
rect 94228 63708 94280 63714
rect 94228 63650 94280 63656
rect 93952 62076 94004 62082
rect 93952 62018 94004 62024
rect 93964 61441 93992 62018
rect 93950 61432 94006 61441
rect 93950 61367 94006 61376
rect 94240 57769 94268 63650
rect 94226 57760 94282 57769
rect 94226 57695 94282 57704
rect 94332 56953 94360 64874
rect 94424 59537 94452 69022
rect 94516 64025 94544 74530
rect 94596 74316 94648 74322
rect 94596 74258 94648 74264
rect 94608 73953 94636 74258
rect 94594 73944 94650 73953
rect 94594 73879 94650 73888
rect 94596 70440 94648 70446
rect 94596 70382 94648 70388
rect 94502 64016 94558 64025
rect 94502 63951 94558 63960
rect 94504 62144 94556 62150
rect 94504 62086 94556 62092
rect 94410 59528 94466 59537
rect 94410 59463 94466 59472
rect 94412 57996 94464 58002
rect 94412 57938 94464 57944
rect 94318 56944 94374 56953
rect 94318 56879 94374 56888
rect 93860 56636 93912 56642
rect 93860 56578 93912 56584
rect 93872 50697 93900 56578
rect 94044 55344 94096 55350
rect 94044 55286 94096 55292
rect 93952 55276 94004 55282
rect 93952 55218 94004 55224
rect 93858 50688 93914 50697
rect 93858 50623 93914 50632
rect 93964 49745 93992 55218
rect 93950 49736 94006 49745
rect 93950 49671 94006 49680
rect 94056 48929 94084 55286
rect 94424 51513 94452 57938
rect 94516 54233 94544 62086
rect 94608 60489 94636 70382
rect 94700 65929 94728 77250
rect 94792 73001 94820 85546
rect 94872 84244 94924 84250
rect 94872 84186 94924 84192
rect 94778 72992 94834 73001
rect 94778 72927 94834 72936
rect 94884 71233 94912 84186
rect 94976 74769 95004 88334
rect 95148 88256 95200 88262
rect 95146 88224 95148 88233
rect 95200 88224 95202 88233
rect 95146 88159 95202 88168
rect 95148 85536 95200 85542
rect 95148 85478 95200 85484
rect 95160 84697 95188 85478
rect 95146 84688 95202 84697
rect 95146 84623 95202 84632
rect 95148 84176 95200 84182
rect 95148 84118 95200 84124
rect 95160 83745 95188 84118
rect 95146 83736 95202 83745
rect 95146 83671 95202 83680
rect 95884 82884 95936 82890
rect 95884 82826 95936 82832
rect 95056 81456 95108 81462
rect 95056 81398 95108 81404
rect 94962 74760 95018 74769
rect 94962 74695 95018 74704
rect 94964 71800 95016 71806
rect 94964 71742 95016 71748
rect 94870 71224 94926 71233
rect 94870 71159 94926 71168
rect 94872 70304 94924 70310
rect 94870 70272 94872 70281
rect 94924 70272 94926 70281
rect 94870 70207 94926 70216
rect 94872 67652 94924 67658
rect 94872 67594 94924 67600
rect 94780 66292 94832 66298
rect 94780 66234 94832 66240
rect 94686 65920 94742 65929
rect 94686 65855 94742 65864
rect 94688 65340 94740 65346
rect 94688 65282 94740 65288
rect 94700 64977 94728 65282
rect 94686 64968 94742 64977
rect 94686 64903 94742 64912
rect 94792 63714 94820 66234
rect 94780 63708 94832 63714
rect 94780 63650 94832 63656
rect 94884 63594 94912 67594
rect 94792 63566 94912 63594
rect 94688 62212 94740 62218
rect 94688 62154 94740 62160
rect 94594 60480 94650 60489
rect 94594 60415 94650 60424
rect 94700 55185 94728 62154
rect 94792 58721 94820 63566
rect 94872 63504 94924 63510
rect 94872 63446 94924 63452
rect 94884 63209 94912 63446
rect 94870 63200 94926 63209
rect 94870 63135 94926 63144
rect 94976 62257 95004 71742
rect 95068 69465 95096 81398
rect 95148 78736 95200 78742
rect 95148 78678 95200 78684
rect 95054 69456 95110 69465
rect 95054 69391 95110 69400
rect 95160 67697 95188 78678
rect 95896 70310 95924 82826
rect 95988 78266 96016 92482
rect 97264 87032 97316 87038
rect 97264 86974 97316 86980
rect 95976 78260 96028 78266
rect 95976 78202 96028 78208
rect 97276 74322 97304 86974
rect 97368 83434 97396 99350
rect 98656 88262 98684 106286
rect 101404 103556 101456 103562
rect 101404 103498 101456 103504
rect 100024 96688 100076 96694
rect 100024 96630 100076 96636
rect 98736 90364 98788 90370
rect 98736 90306 98788 90312
rect 98644 88256 98696 88262
rect 98644 88198 98696 88204
rect 97356 83428 97408 83434
rect 97356 83370 97408 83376
rect 98644 80096 98696 80102
rect 98644 80038 98696 80044
rect 97356 75948 97408 75954
rect 97356 75890 97408 75896
rect 97264 74316 97316 74322
rect 97264 74258 97316 74264
rect 95976 73228 96028 73234
rect 95976 73170 96028 73176
rect 95884 70304 95936 70310
rect 95884 70246 95936 70252
rect 95146 67688 95202 67697
rect 95146 67623 95202 67632
rect 95148 66904 95200 66910
rect 95148 66846 95200 66852
rect 95160 66745 95188 66846
rect 95146 66736 95202 66745
rect 95146 66671 95202 66680
rect 95148 63572 95200 63578
rect 95148 63514 95200 63520
rect 94962 62248 95018 62257
rect 94962 62183 95018 62192
rect 94964 60784 95016 60790
rect 94964 60726 95016 60732
rect 94778 58712 94834 58721
rect 94778 58647 94834 58656
rect 94686 55176 94742 55185
rect 94686 55111 94742 55120
rect 94502 54224 94558 54233
rect 94502 54159 94558 54168
rect 94780 53848 94832 53854
rect 94780 53790 94832 53796
rect 94410 51504 94466 51513
rect 94410 51439 94466 51448
rect 94228 51128 94280 51134
rect 94228 51070 94280 51076
rect 94042 48920 94098 48929
rect 94042 48855 94098 48864
rect 94136 46980 94188 46986
rect 94136 46922 94188 46928
rect 93952 45620 94004 45626
rect 93952 45562 94004 45568
rect 93964 41721 93992 45562
rect 94148 42537 94176 46922
rect 94240 46209 94268 51070
rect 94504 48408 94556 48414
rect 94504 48350 94556 48356
rect 94412 48340 94464 48346
rect 94412 48282 94464 48288
rect 94226 46200 94282 46209
rect 94226 46135 94282 46144
rect 94424 44441 94452 48282
rect 94410 44432 94466 44441
rect 94410 44367 94466 44376
rect 94516 43489 94544 48350
rect 94792 47977 94820 53790
rect 94976 53281 95004 60726
rect 95056 59424 95108 59430
rect 95056 59366 95108 59372
rect 94962 53272 95018 53281
rect 94962 53207 95018 53216
rect 95068 52465 95096 59366
rect 95160 56001 95188 63514
rect 95988 63510 96016 73170
rect 97368 65346 97396 75890
rect 98656 68542 98684 80038
rect 98748 80034 98776 90306
rect 100036 81326 100064 96630
rect 101416 86630 101444 103498
rect 102796 91050 102824 107714
rect 116412 107710 116440 107879
rect 116400 107704 116452 107710
rect 214024 107681 214052 108938
rect 116400 107646 116452 107652
rect 214010 107672 214066 107681
rect 213920 107636 213972 107642
rect 214010 107607 214066 107616
rect 213920 107578 213972 107584
rect 213932 107001 213960 107578
rect 213918 106992 213974 107001
rect 213918 106927 213974 106936
rect 116398 106720 116454 106729
rect 116398 106655 116454 106664
rect 116412 106350 116440 106655
rect 116400 106344 116452 106350
rect 116400 106286 116452 106292
rect 213920 106276 213972 106282
rect 213920 106218 213972 106224
rect 213932 106185 213960 106218
rect 214012 106208 214064 106214
rect 213918 106176 213974 106185
rect 214012 106150 214064 106156
rect 213918 106111 213974 106120
rect 116398 105632 116454 105641
rect 116398 105567 116454 105576
rect 116412 104922 116440 105567
rect 214024 105369 214052 106150
rect 214010 105360 214066 105369
rect 214010 105295 214066 105304
rect 116400 104916 116452 104922
rect 116400 104858 116452 104864
rect 214012 104848 214064 104854
rect 214012 104790 214064 104796
rect 213920 104780 213972 104786
rect 213920 104722 213972 104728
rect 213932 104553 213960 104722
rect 213918 104544 213974 104553
rect 213918 104479 213974 104488
rect 116398 104408 116454 104417
rect 116398 104343 116454 104352
rect 116412 103562 116440 104343
rect 214024 103873 214052 104790
rect 214668 104122 214696 225626
rect 214760 158681 214788 229706
rect 250456 229158 250484 235175
rect 245568 229152 245620 229158
rect 245568 229094 245620 229100
rect 250444 229152 250496 229158
rect 250444 229094 250496 229100
rect 214932 228404 214984 228410
rect 214932 228346 214984 228352
rect 214840 200592 214892 200598
rect 214840 200534 214892 200540
rect 214852 179586 214880 200534
rect 214840 179580 214892 179586
rect 214840 179522 214892 179528
rect 214840 179444 214892 179450
rect 214840 179386 214892 179392
rect 214852 167249 214880 179386
rect 214838 167240 214894 167249
rect 214838 167175 214894 167184
rect 214746 158672 214802 158681
rect 214746 158607 214802 158616
rect 214944 157865 214972 228346
rect 229744 223644 229796 223650
rect 229744 223586 229796 223592
rect 229008 222896 229060 222902
rect 229008 222838 229060 222844
rect 229020 221377 229048 222838
rect 229006 221368 229062 221377
rect 229006 221303 229062 221312
rect 226340 220856 226392 220862
rect 226338 220824 226340 220833
rect 226392 220824 226394 220833
rect 226338 220759 226394 220768
rect 226340 220176 226392 220182
rect 226338 220144 226340 220153
rect 226392 220144 226394 220153
rect 226338 220079 226394 220088
rect 226432 220108 226484 220114
rect 226432 220050 226484 220056
rect 226444 219609 226472 220050
rect 226430 219600 226486 219609
rect 226430 219535 226486 219544
rect 226338 219056 226394 219065
rect 226338 218991 226394 219000
rect 226352 218822 226380 218991
rect 226340 218816 226392 218822
rect 226340 218758 226392 218764
rect 226432 218748 226484 218754
rect 226432 218690 226484 218696
rect 226444 218385 226472 218690
rect 226430 218376 226486 218385
rect 226430 218311 226486 218320
rect 226338 217832 226394 217841
rect 226338 217767 226394 217776
rect 226352 217326 226380 217767
rect 226340 217320 226392 217326
rect 226340 217262 226392 217268
rect 226430 217288 226486 217297
rect 226430 217223 226486 217232
rect 226444 216646 226472 217223
rect 226432 216640 226484 216646
rect 226338 216608 226394 216617
rect 226432 216582 226484 216588
rect 226338 216543 226394 216552
rect 226352 215966 226380 216543
rect 226430 216064 226486 216073
rect 226430 215999 226486 216008
rect 226340 215960 226392 215966
rect 226340 215902 226392 215908
rect 226338 215520 226394 215529
rect 226338 215455 226394 215464
rect 226352 215218 226380 215455
rect 226444 215286 226472 215999
rect 226432 215280 226484 215286
rect 226432 215222 226484 215228
rect 226340 215212 226392 215218
rect 226340 215154 226392 215160
rect 226430 214840 226486 214849
rect 226430 214775 226486 214784
rect 226338 214296 226394 214305
rect 226338 214231 226394 214240
rect 226352 213858 226380 214231
rect 226444 213926 226472 214775
rect 226432 213920 226484 213926
rect 226432 213862 226484 213868
rect 226340 213852 226392 213858
rect 226340 213794 226392 213800
rect 226430 213616 226486 213625
rect 226430 213551 226486 213560
rect 226338 213072 226394 213081
rect 226338 213007 226394 213016
rect 226352 212430 226380 213007
rect 226444 212498 226472 213551
rect 226522 212528 226578 212537
rect 226432 212492 226484 212498
rect 226522 212463 226578 212472
rect 226432 212434 226484 212440
rect 226340 212424 226392 212430
rect 226340 212366 226392 212372
rect 226062 211848 226118 211857
rect 226062 211783 226118 211792
rect 225970 210760 226026 210769
rect 225970 210695 226026 210704
rect 225984 208282 226012 210695
rect 226076 209710 226104 211783
rect 226246 211304 226302 211313
rect 226246 211239 226302 211248
rect 226154 210080 226210 210089
rect 226154 210015 226210 210024
rect 226064 209704 226116 209710
rect 226064 209646 226116 209652
rect 226062 209536 226118 209545
rect 226062 209471 226118 209480
rect 225972 208276 226024 208282
rect 225972 208218 226024 208224
rect 225786 207768 225842 207777
rect 225786 207703 225842 207712
rect 225602 205320 225658 205329
rect 225602 205255 225658 205264
rect 225616 201482 225644 205255
rect 225694 204776 225750 204785
rect 225694 204711 225750 204720
rect 225604 201476 225656 201482
rect 225604 201418 225656 201424
rect 225708 201414 225736 204711
rect 225800 204202 225828 207703
rect 225970 207224 226026 207233
rect 225970 207159 226026 207168
rect 225878 206544 225934 206553
rect 225878 206479 225934 206488
rect 225788 204196 225840 204202
rect 225788 204138 225840 204144
rect 225892 202842 225920 206479
rect 225984 204270 226012 207159
rect 226076 206990 226104 209471
rect 226168 208350 226196 210015
rect 226260 209778 226288 211239
rect 226536 211138 226564 212463
rect 226524 211132 226576 211138
rect 226524 211074 226576 211080
rect 226248 209772 226300 209778
rect 226248 209714 226300 209720
rect 226246 208992 226302 209001
rect 226246 208927 226302 208936
rect 226156 208344 226208 208350
rect 226156 208286 226208 208292
rect 226154 208040 226210 208049
rect 226154 207975 226210 207984
rect 226064 206984 226116 206990
rect 226064 206926 226116 206932
rect 226168 205630 226196 207975
rect 226260 206922 226288 208927
rect 226248 206916 226300 206922
rect 226248 206858 226300 206864
rect 226246 206000 226302 206009
rect 226246 205935 226302 205944
rect 226156 205624 226208 205630
rect 226156 205566 226208 205572
rect 226260 204354 226288 205935
rect 226168 204326 226288 204354
rect 225972 204264 226024 204270
rect 225972 204206 226024 204212
rect 226062 203552 226118 203561
rect 226062 203487 226118 203496
rect 225970 203008 226026 203017
rect 225970 202943 226026 202952
rect 225880 202836 225932 202842
rect 225880 202778 225932 202784
rect 225786 202464 225842 202473
rect 225786 202399 225842 202408
rect 225696 201408 225748 201414
rect 225696 201350 225748 201356
rect 225694 200016 225750 200025
rect 225694 199951 225750 199960
rect 224132 198824 224184 198830
rect 224132 198766 224184 198772
rect 223948 198756 224000 198762
rect 223948 198698 224000 198704
rect 221464 194676 221516 194682
rect 221464 194618 221516 194624
rect 220084 193316 220136 193322
rect 220084 193258 220136 193264
rect 215300 191956 215352 191962
rect 215300 191898 215352 191904
rect 215024 190528 215076 190534
rect 215024 190470 215076 190476
rect 215036 182889 215064 190470
rect 215312 184362 215340 191898
rect 218704 189168 218756 189174
rect 218704 189110 218756 189116
rect 215944 187740 215996 187746
rect 215944 187682 215996 187688
rect 215220 184334 215340 184362
rect 215220 183705 215248 184334
rect 215300 184204 215352 184210
rect 215300 184146 215352 184152
rect 215206 183696 215262 183705
rect 215206 183631 215262 183640
rect 215022 182880 215078 182889
rect 215022 182815 215078 182824
rect 215024 182300 215076 182306
rect 215024 182242 215076 182248
rect 215036 170377 215064 182242
rect 215206 182200 215262 182209
rect 215312 182186 215340 184146
rect 215262 182158 215340 182186
rect 215206 182135 215262 182144
rect 215116 180872 215168 180878
rect 215116 180814 215168 180820
rect 215022 170368 215078 170377
rect 215022 170303 215078 170312
rect 215128 168881 215156 180814
rect 215956 179110 215984 187682
rect 218716 180606 218744 189110
rect 220096 185094 220124 193258
rect 221476 186590 221504 194618
rect 223960 193118 223988 198698
rect 224040 197396 224092 197402
rect 224040 197338 224092 197344
rect 223948 193112 224000 193118
rect 223948 193054 224000 193060
rect 224052 191826 224080 197338
rect 224144 193186 224172 198766
rect 224500 197464 224552 197470
rect 224500 197406 224552 197412
rect 224316 196104 224368 196110
rect 224316 196046 224368 196052
rect 224224 194744 224276 194750
rect 224224 194686 224276 194692
rect 224132 193180 224184 193186
rect 224132 193122 224184 193128
rect 224040 191820 224092 191826
rect 224040 191762 224092 191768
rect 224236 189038 224264 194686
rect 224328 190398 224356 196046
rect 224408 196036 224460 196042
rect 224408 195978 224460 195984
rect 224420 190466 224448 195978
rect 224512 191758 224540 197406
rect 225708 194546 225736 199951
rect 225800 197266 225828 202399
rect 225878 200696 225934 200705
rect 225878 200631 225934 200640
rect 225788 197260 225840 197266
rect 225788 197202 225840 197208
rect 225892 195906 225920 200631
rect 225984 198694 226012 202943
rect 225972 198688 226024 198694
rect 225972 198630 226024 198636
rect 226076 198626 226104 203487
rect 226168 202774 226196 204326
rect 226246 204232 226302 204241
rect 226246 204167 226302 204176
rect 226156 202768 226208 202774
rect 226156 202710 226208 202716
rect 226154 201784 226210 201793
rect 226154 201719 226210 201728
rect 226064 198620 226116 198626
rect 226064 198562 226116 198568
rect 226168 197334 226196 201719
rect 226260 200122 226288 204167
rect 226338 201240 226394 201249
rect 226338 201175 226394 201184
rect 226248 200116 226300 200122
rect 226248 200058 226300 200064
rect 226352 200002 226380 201175
rect 226260 199974 226380 200002
rect 226156 197328 226208 197334
rect 226156 197270 226208 197276
rect 226260 195974 226288 199974
rect 226430 199472 226486 199481
rect 226430 199407 226486 199416
rect 226338 198928 226394 198937
rect 226338 198863 226394 198872
rect 226352 198762 226380 198863
rect 226444 198830 226472 199407
rect 226432 198824 226484 198830
rect 226432 198766 226484 198772
rect 226340 198756 226392 198762
rect 226340 198698 226392 198704
rect 226430 198248 226486 198257
rect 226430 198183 226486 198192
rect 226338 197704 226394 197713
rect 226338 197639 226394 197648
rect 226352 197402 226380 197639
rect 226444 197470 226472 198183
rect 226432 197464 226484 197470
rect 226432 197406 226484 197412
rect 226340 197396 226392 197402
rect 226340 197338 226392 197344
rect 226338 197024 226394 197033
rect 226338 196959 226394 196968
rect 226352 196110 226380 196959
rect 226706 196480 226762 196489
rect 226706 196415 226762 196424
rect 226340 196104 226392 196110
rect 226340 196046 226392 196052
rect 226720 196042 226748 196415
rect 226708 196036 226760 196042
rect 226708 195978 226760 195984
rect 226248 195968 226300 195974
rect 226248 195910 226300 195916
rect 226522 195936 226578 195945
rect 225880 195900 225932 195906
rect 226522 195871 226578 195880
rect 225880 195842 225932 195848
rect 226338 195256 226394 195265
rect 226338 195191 226394 195200
rect 226352 194614 226380 195191
rect 226536 194750 226564 195871
rect 226524 194744 226576 194750
rect 226430 194712 226486 194721
rect 226524 194686 226576 194692
rect 226430 194647 226432 194656
rect 226484 194647 226486 194656
rect 226432 194618 226484 194624
rect 226340 194608 226392 194614
rect 226340 194550 226392 194556
rect 225696 194540 225748 194546
rect 225696 194482 225748 194488
rect 226338 194168 226394 194177
rect 226338 194103 226394 194112
rect 226352 193254 226380 194103
rect 226430 193488 226486 193497
rect 226430 193423 226486 193432
rect 226444 193322 226472 193423
rect 226432 193316 226484 193322
rect 226432 193258 226484 193264
rect 226340 193248 226392 193254
rect 226340 193190 226392 193196
rect 226430 192944 226486 192953
rect 226430 192879 226486 192888
rect 226338 192400 226394 192409
rect 226338 192335 226394 192344
rect 226352 191962 226380 192335
rect 226340 191956 226392 191962
rect 226340 191898 226392 191904
rect 226444 191894 226472 192879
rect 226432 191888 226484 191894
rect 226432 191830 226484 191836
rect 224500 191752 224552 191758
rect 224500 191694 224552 191700
rect 226430 191720 226486 191729
rect 226430 191655 226486 191664
rect 226340 190596 226392 190602
rect 226340 190538 226392 190544
rect 226352 190505 226380 190538
rect 226444 190534 226472 191655
rect 226522 191176 226578 191185
rect 226522 191111 226578 191120
rect 226432 190528 226484 190534
rect 226338 190496 226394 190505
rect 224408 190460 224460 190466
rect 226432 190470 226484 190476
rect 226338 190431 226394 190440
rect 224408 190402 224460 190408
rect 224316 190392 224368 190398
rect 224316 190334 224368 190340
rect 226430 189952 226486 189961
rect 226430 189887 226486 189896
rect 226338 189408 226394 189417
rect 226338 189343 226394 189352
rect 226352 189106 226380 189343
rect 226444 189174 226472 189887
rect 226432 189168 226484 189174
rect 226432 189110 226484 189116
rect 226340 189100 226392 189106
rect 226340 189042 226392 189048
rect 224224 189032 224276 189038
rect 224224 188974 224276 188980
rect 226338 188728 226394 188737
rect 226338 188663 226394 188672
rect 222936 187808 222988 187814
rect 222936 187750 222988 187756
rect 221464 186584 221516 186590
rect 221464 186526 221516 186532
rect 220084 185088 220136 185094
rect 220084 185030 220136 185036
rect 220176 185020 220228 185026
rect 220176 184962 220228 184968
rect 218704 180600 218756 180606
rect 218704 180542 218756 180548
rect 215944 179104 215996 179110
rect 215944 179046 215996 179052
rect 218704 176724 218756 176730
rect 218704 176666 218756 176672
rect 218060 170400 218112 170406
rect 218060 170342 218112 170348
rect 215114 168872 215170 168881
rect 215114 168807 215170 168816
rect 218072 162314 218100 170342
rect 218716 164150 218744 176666
rect 220188 174214 220216 184962
rect 221464 181280 221516 181286
rect 221464 181222 221516 181228
rect 220176 174208 220228 174214
rect 220176 174150 220228 174156
rect 220084 174072 220136 174078
rect 220084 174014 220136 174020
rect 218796 171828 218848 171834
rect 218796 171770 218848 171776
rect 218704 164144 218756 164150
rect 218704 164086 218756 164092
rect 218060 162308 218112 162314
rect 218060 162250 218112 162256
rect 218808 160886 218836 171770
rect 220096 163606 220124 174014
rect 221476 169114 221504 181222
rect 222844 179512 222896 179518
rect 222844 179454 222896 179460
rect 221556 178152 221608 178158
rect 221556 178094 221608 178100
rect 221464 169108 221516 169114
rect 221464 169050 221516 169056
rect 221568 166598 221596 178094
rect 222856 168366 222884 179454
rect 222948 179382 222976 187750
rect 226352 187746 226380 188663
rect 226430 188184 226486 188193
rect 226430 188119 226486 188128
rect 226444 187814 226472 188119
rect 226432 187808 226484 187814
rect 226432 187750 226484 187756
rect 226340 187740 226392 187746
rect 226340 187682 226392 187688
rect 226338 186960 226394 186969
rect 226338 186895 226394 186904
rect 224408 186448 224460 186454
rect 224408 186390 224460 186396
rect 222936 179376 222988 179382
rect 222936 179318 222988 179324
rect 224316 178084 224368 178090
rect 224316 178026 224368 178032
rect 224224 175296 224276 175302
rect 224224 175238 224276 175244
rect 223580 174140 223632 174146
rect 223580 174082 223632 174088
rect 223592 171834 223620 174082
rect 223580 171828 223632 171834
rect 223580 171770 223632 171776
rect 222844 168360 222896 168366
rect 222844 168302 222896 168308
rect 221556 166592 221608 166598
rect 221556 166534 221608 166540
rect 220084 163600 220136 163606
rect 220084 163542 220136 163548
rect 224236 162858 224264 175238
rect 224328 167006 224356 178026
rect 224420 176662 224448 186390
rect 226352 186386 226380 186895
rect 226432 186448 226484 186454
rect 226430 186416 226432 186425
rect 226484 186416 226486 186425
rect 226340 186380 226392 186386
rect 226430 186351 226486 186360
rect 226340 186322 226392 186328
rect 226338 185872 226394 185881
rect 226338 185807 226394 185816
rect 226352 184958 226380 185807
rect 226430 185192 226486 185201
rect 226430 185127 226486 185136
rect 226444 185026 226472 185127
rect 226432 185020 226484 185026
rect 226432 184962 226484 184968
rect 226340 184952 226392 184958
rect 226340 184894 226392 184900
rect 226338 184648 226394 184657
rect 226338 184583 226394 184592
rect 226352 183598 226380 184583
rect 226536 184210 226564 191111
rect 227074 187640 227130 187649
rect 227074 187575 227130 187584
rect 226524 184204 226576 184210
rect 226524 184146 226576 184152
rect 226982 184104 227038 184113
rect 226982 184039 227038 184048
rect 226340 183592 226392 183598
rect 226340 183534 226392 183540
rect 226430 183424 226486 183433
rect 226430 183359 226486 183368
rect 225694 182880 225750 182889
rect 225694 182815 225750 182824
rect 225602 178120 225658 178129
rect 225602 178055 225658 178064
rect 224408 176656 224460 176662
rect 224408 176598 224460 176604
rect 224316 167000 224368 167006
rect 224316 166942 224368 166948
rect 225616 165578 225644 178055
rect 225708 172514 225736 182815
rect 226444 182374 226472 183359
rect 226432 182368 226484 182374
rect 226432 182310 226484 182316
rect 226340 182300 226392 182306
rect 226340 182242 226392 182248
rect 226352 182209 226380 182242
rect 226338 182200 226394 182209
rect 226338 182135 226394 182144
rect 226338 181656 226394 181665
rect 226338 181591 226394 181600
rect 226352 181286 226380 181591
rect 226340 181280 226392 181286
rect 226340 181222 226392 181228
rect 226338 181112 226394 181121
rect 226338 181047 226394 181056
rect 226352 180878 226380 181047
rect 226340 180872 226392 180878
rect 226340 180814 226392 180820
rect 226430 180432 226486 180441
rect 226430 180367 226486 180376
rect 226338 179888 226394 179897
rect 226338 179823 226394 179832
rect 226352 179450 226380 179823
rect 226444 179518 226472 180367
rect 226432 179512 226484 179518
rect 226432 179454 226484 179460
rect 226340 179444 226392 179450
rect 226340 179386 226392 179392
rect 226338 179344 226394 179353
rect 226338 179279 226394 179288
rect 226352 178090 226380 179279
rect 226430 178664 226486 178673
rect 226430 178599 226486 178608
rect 226444 178158 226472 178599
rect 226432 178152 226484 178158
rect 226432 178094 226484 178100
rect 226340 178084 226392 178090
rect 226340 178026 226392 178032
rect 226338 177576 226394 177585
rect 226338 177511 226394 177520
rect 226352 176730 226380 177511
rect 226430 176896 226486 176905
rect 226430 176831 226486 176840
rect 226340 176724 226392 176730
rect 226340 176666 226392 176672
rect 226444 174078 226472 176831
rect 226890 176352 226946 176361
rect 226890 176287 226946 176296
rect 226904 175302 226932 176287
rect 226892 175296 226944 175302
rect 226892 175238 226944 175244
rect 226432 174072 226484 174078
rect 226432 174014 226484 174020
rect 226996 173874 227024 184039
rect 227088 178022 227116 187575
rect 227720 180872 227772 180878
rect 227720 180814 227772 180820
rect 227076 178016 227128 178022
rect 227076 177958 227128 177964
rect 227442 175808 227498 175817
rect 227442 175743 227498 175752
rect 226984 173868 227036 173874
rect 226984 173810 227036 173816
rect 225696 172508 225748 172514
rect 225696 172450 225748 172456
rect 227456 170406 227484 175743
rect 227732 174146 227760 180814
rect 227720 174140 227772 174146
rect 227720 174082 227772 174088
rect 227444 170400 227496 170406
rect 227444 170342 227496 170348
rect 225604 165572 225656 165578
rect 225604 165514 225656 165520
rect 224224 162852 224276 162858
rect 224224 162794 224276 162800
rect 229756 161430 229784 223586
rect 245580 222970 245608 229094
rect 286336 224262 286364 569162
rect 287716 474706 287744 667898
rect 298192 531072 298244 531078
rect 298192 531014 298244 531020
rect 298100 531004 298152 531010
rect 298100 530946 298152 530952
rect 298112 530890 298140 530946
rect 298204 530890 298232 531014
rect 298112 530862 298232 530890
rect 296626 527504 296682 527513
rect 296626 527439 296682 527448
rect 298098 527504 298154 527513
rect 298098 527439 298100 527448
rect 296640 527270 296668 527439
rect 298152 527439 298154 527448
rect 298100 527410 298152 527416
rect 288532 527264 288584 527270
rect 288530 527232 288532 527241
rect 296628 527264 296680 527270
rect 288584 527232 288586 527241
rect 296628 527206 296680 527212
rect 288530 527167 288586 527176
rect 289728 500268 289780 500274
rect 289728 500210 289780 500216
rect 287704 474700 287756 474706
rect 287704 474642 287756 474648
rect 289636 425740 289688 425746
rect 289636 425682 289688 425688
rect 288898 317112 288954 317121
rect 288898 317047 288954 317056
rect 288912 316742 288940 317047
rect 288900 316736 288952 316742
rect 288900 316678 288952 316684
rect 289648 308961 289676 425682
rect 289740 325281 289768 500210
rect 299388 496120 299440 496126
rect 299388 496062 299440 496068
rect 299400 495514 299428 496062
rect 298100 495508 298152 495514
rect 298100 495450 298152 495456
rect 299388 495508 299440 495514
rect 299388 495450 299440 495456
rect 292580 421592 292632 421598
rect 292580 421534 292632 421540
rect 292592 329338 292620 421534
rect 298112 329338 298140 495450
rect 292592 329310 292988 329338
rect 298112 329310 298508 329338
rect 292960 329066 292988 329310
rect 298480 329066 298508 329310
rect 292960 329038 293526 329066
rect 298480 329038 298954 329066
rect 289726 325272 289782 325281
rect 289726 325207 289782 325216
rect 289634 308952 289690 308961
rect 289634 308887 289690 308896
rect 300860 305652 300912 305658
rect 300860 305594 300912 305600
rect 300872 305561 300900 305594
rect 300858 305552 300914 305561
rect 300858 305487 300914 305496
rect 292592 302841 292620 304844
rect 296180 303618 296208 304844
rect 299492 304830 299782 304858
rect 296168 303612 296220 303618
rect 296168 303554 296220 303560
rect 292578 302832 292634 302841
rect 292578 302767 292634 302776
rect 299492 225622 299520 304830
rect 301516 228410 301544 700470
rect 304264 556232 304316 556238
rect 304264 556174 304316 556180
rect 302976 527468 303028 527474
rect 302976 527410 303028 527416
rect 302988 527241 303016 527410
rect 302974 527232 303030 527241
rect 302974 527167 303030 527176
rect 304276 328273 304304 556174
rect 304356 415472 304408 415478
rect 304356 415414 304408 415420
rect 304262 328264 304318 328273
rect 304262 328199 304318 328208
rect 303620 327072 303672 327078
rect 303620 327014 303672 327020
rect 303632 326369 303660 327014
rect 303618 326360 303674 326369
rect 303618 326295 303674 326304
rect 303620 325644 303672 325650
rect 303620 325586 303672 325592
rect 303632 324465 303660 325586
rect 303618 324456 303674 324465
rect 303618 324391 303674 324400
rect 304368 322561 304396 415414
rect 304448 368552 304500 368558
rect 304448 368494 304500 368500
rect 304354 322552 304410 322561
rect 304354 322487 304410 322496
rect 303620 321632 303672 321638
rect 303620 321574 303672 321580
rect 303632 318753 303660 321574
rect 304460 320657 304488 368494
rect 304446 320648 304502 320657
rect 304446 320583 304502 320592
rect 303618 318744 303674 318753
rect 303618 318679 303674 318688
rect 304354 316976 304410 316985
rect 304354 316911 304410 316920
rect 304262 315072 304318 315081
rect 304262 315007 304318 315016
rect 303618 313168 303674 313177
rect 303618 313103 303674 313112
rect 303632 311914 303660 313103
rect 303620 311908 303672 311914
rect 303620 311850 303672 311856
rect 303618 311264 303674 311273
rect 303618 311199 303674 311208
rect 303632 310554 303660 311199
rect 303620 310548 303672 310554
rect 303620 310490 303672 310496
rect 303618 309360 303674 309369
rect 303618 309295 303674 309304
rect 303632 309194 303660 309295
rect 303620 309188 303672 309194
rect 303620 309130 303672 309136
rect 303618 307456 303674 307465
rect 303618 307391 303674 307400
rect 303632 306406 303660 307391
rect 303620 306400 303672 306406
rect 303620 306342 303672 306348
rect 304276 229090 304304 315007
rect 304368 276010 304396 316911
rect 304356 276004 304408 276010
rect 304356 275946 304408 275952
rect 305656 229770 305684 700538
rect 397472 700534 397500 703520
rect 397460 700528 397512 700534
rect 397460 700470 397512 700476
rect 413664 700466 413692 703520
rect 313924 700460 313976 700466
rect 313924 700402 313976 700408
rect 413652 700460 413704 700466
rect 413652 700402 413704 700408
rect 312544 700392 312596 700398
rect 312544 700334 312596 700340
rect 305644 229764 305696 229770
rect 305644 229706 305696 229712
rect 304264 229084 304316 229090
rect 304264 229026 304316 229032
rect 301504 228404 301556 228410
rect 301504 228346 301556 228352
rect 312556 225690 312584 700334
rect 313280 614100 313332 614106
rect 313280 614042 313332 614048
rect 313292 613465 313320 614042
rect 313278 613456 313334 613465
rect 313278 613391 313334 613400
rect 313280 463684 313332 463690
rect 313280 463626 313332 463632
rect 313292 462777 313320 463626
rect 313278 462768 313334 462777
rect 313278 462703 313334 462712
rect 312544 225684 312596 225690
rect 312544 225626 312596 225632
rect 299480 225616 299532 225622
rect 299480 225558 299532 225564
rect 286324 224256 286376 224262
rect 286324 224198 286376 224204
rect 283380 223644 283432 223650
rect 283380 223586 283432 223592
rect 231124 222964 231176 222970
rect 231124 222906 231176 222912
rect 245568 222964 245620 222970
rect 245568 222906 245620 222912
rect 230848 180872 230900 180878
rect 231136 180826 231164 222906
rect 283392 221612 283420 223586
rect 313936 222902 313964 700402
rect 462332 700398 462360 703520
rect 478524 700505 478552 703520
rect 478510 700496 478566 700505
rect 478510 700431 478566 700440
rect 462320 700392 462372 700398
rect 462320 700334 462372 700340
rect 527192 700330 527220 703520
rect 543476 700369 543504 703520
rect 543462 700360 543518 700369
rect 315304 700324 315356 700330
rect 315304 700266 315356 700272
rect 527180 700324 527232 700330
rect 543462 700295 543518 700304
rect 527180 700266 527232 700272
rect 314658 515808 314714 515817
rect 314658 515743 314714 515752
rect 314672 439657 314700 515743
rect 314658 439648 314714 439657
rect 314658 439583 314714 439592
rect 314672 426426 314700 439583
rect 314660 426420 314712 426426
rect 314660 426362 314712 426368
rect 314672 425746 314700 426362
rect 314660 425740 314712 425746
rect 314660 425682 314712 425688
rect 315316 233918 315344 700266
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 576124 696992 576176 696998
rect 576124 696934 576176 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 453304 681760 453356 681766
rect 453304 681702 453356 681708
rect 453316 616826 453344 681702
rect 506018 663912 506074 663921
rect 506018 663847 506074 663856
rect 506032 662388 506060 663847
rect 552018 641744 552074 641753
rect 552018 641679 552074 641688
rect 551650 639568 551706 639577
rect 551650 639503 551706 639512
rect 456062 635216 456118 635225
rect 456062 635151 456118 635160
rect 453304 616820 453356 616826
rect 453304 616762 453356 616768
rect 455418 591696 455474 591705
rect 455418 591631 455474 591640
rect 316894 570030 317368 570058
rect 317340 552702 317368 570030
rect 318536 570030 318642 570058
rect 318536 569974 318564 570030
rect 318524 569968 318576 569974
rect 318524 569910 318576 569916
rect 318708 569968 318760 569974
rect 318708 569910 318760 569916
rect 317328 552696 317380 552702
rect 317328 552638 317380 552644
rect 318720 533798 318748 569910
rect 320376 567254 320404 570044
rect 322230 570030 322888 570058
rect 323978 570030 324176 570058
rect 320364 567248 320416 567254
rect 320364 567190 320416 567196
rect 321468 567248 321520 567254
rect 321468 567190 321520 567196
rect 318708 533792 318760 533798
rect 318708 533734 318760 533740
rect 321284 533588 321336 533594
rect 321284 533530 321336 533536
rect 320732 533520 320784 533526
rect 320732 533462 320784 533468
rect 319628 533452 319680 533458
rect 319628 533394 319680 533400
rect 318524 533384 318576 533390
rect 318524 533326 318576 533332
rect 318536 528850 318564 533326
rect 319640 528850 319668 533394
rect 320744 528850 320772 533462
rect 318228 528822 318564 528850
rect 319332 528822 319668 528850
rect 320436 528822 320772 528850
rect 321296 528714 321324 533530
rect 321480 532438 321508 567190
rect 322860 541686 322888 570030
rect 322848 541680 322900 541686
rect 322848 541622 322900 541628
rect 323952 533724 324004 533730
rect 323952 533666 324004 533672
rect 322848 533656 322900 533662
rect 322848 533598 322900 533604
rect 321468 532432 321520 532438
rect 321468 532374 321520 532380
rect 322860 528850 322888 533598
rect 323964 528850 323992 533666
rect 324148 532574 324176 570030
rect 325804 568342 325832 570044
rect 327552 568546 327580 570044
rect 327540 568540 327592 568546
rect 327540 568482 327592 568488
rect 328276 568540 328328 568546
rect 328276 568482 328328 568488
rect 325792 568336 325844 568342
rect 325792 568278 325844 568284
rect 326894 567896 326950 567905
rect 326894 567831 326950 567840
rect 324136 532568 324188 532574
rect 324136 532510 324188 532516
rect 325054 532128 325110 532137
rect 325054 532063 325110 532072
rect 325068 528850 325096 532063
rect 326908 531146 326936 567831
rect 328288 533866 328316 568482
rect 329392 568478 329420 570044
rect 331048 570030 331154 570058
rect 329380 568472 329432 568478
rect 329380 568414 329432 568420
rect 328368 567860 328420 567866
rect 328368 567802 328420 567808
rect 328276 533860 328328 533866
rect 328276 533802 328328 533808
rect 326988 532024 327040 532030
rect 326988 531966 327040 531972
rect 326068 531140 326120 531146
rect 326068 531082 326120 531088
rect 326896 531140 326948 531146
rect 326896 531082 326948 531088
rect 326080 528850 326108 531082
rect 327000 528850 327028 531966
rect 328380 528850 328408 567802
rect 331048 533934 331076 570030
rect 332416 567996 332468 568002
rect 332416 567938 332468 567944
rect 331128 567928 331180 567934
rect 331128 567870 331180 567876
rect 331036 533928 331088 533934
rect 331036 533870 331088 533876
rect 329288 532092 329340 532098
rect 329288 532034 329340 532040
rect 329300 528850 329328 532034
rect 331140 531146 331168 567870
rect 331496 532160 331548 532166
rect 331496 532102 331548 532108
rect 330392 531140 330444 531146
rect 330392 531082 330444 531088
rect 331128 531140 331180 531146
rect 331128 531082 331180 531088
rect 330404 528850 330432 531082
rect 331508 528850 331536 532102
rect 332428 528850 332456 567938
rect 332980 567730 333008 570044
rect 334742 570030 335216 570058
rect 332968 567724 333020 567730
rect 332968 567666 333020 567672
rect 335188 534002 335216 570030
rect 336476 570030 336582 570058
rect 335268 568064 335320 568070
rect 335268 568006 335320 568012
rect 335176 533996 335228 534002
rect 335176 533938 335228 533944
rect 333612 532228 333664 532234
rect 333612 532170 333664 532176
rect 333624 528850 333652 532170
rect 335280 531146 335308 568006
rect 336476 567662 336504 570030
rect 338316 568546 338344 570044
rect 338304 568540 338356 568546
rect 338304 568482 338356 568488
rect 339316 568540 339368 568546
rect 339316 568482 339368 568488
rect 336556 568132 336608 568138
rect 336556 568074 336608 568080
rect 336464 567656 336516 567662
rect 336464 567598 336516 567604
rect 335820 532296 335872 532302
rect 335820 532238 335872 532244
rect 334716 531140 334768 531146
rect 334716 531082 334768 531088
rect 335268 531140 335320 531146
rect 335268 531082 335320 531088
rect 334728 528850 334756 531082
rect 335832 528850 335860 532238
rect 336568 528850 336596 568074
rect 339328 534070 339356 568482
rect 339408 568200 339460 568206
rect 339408 568142 339460 568148
rect 339316 534064 339368 534070
rect 339316 534006 339368 534012
rect 337936 532364 337988 532370
rect 337936 532306 337988 532312
rect 337948 528850 337976 532306
rect 339420 528986 339448 568142
rect 340156 567458 340184 570044
rect 341918 570030 342116 570058
rect 341984 568268 342036 568274
rect 341984 568210 342036 568216
rect 340144 567452 340196 567458
rect 340144 567394 340196 567400
rect 340144 532500 340196 532506
rect 340144 532442 340196 532448
rect 339500 531616 339552 531622
rect 339500 531558 339552 531564
rect 339512 531214 339540 531558
rect 339500 531208 339552 531214
rect 339500 531150 339552 531156
rect 339144 528958 339448 528986
rect 339144 528850 339172 528958
rect 340156 528850 340184 532442
rect 341996 531146 342024 568210
rect 342088 533322 342116 570030
rect 343548 568404 343600 568410
rect 343548 568346 343600 568352
rect 342076 533316 342128 533322
rect 342076 533258 342128 533264
rect 342168 532636 342220 532642
rect 342168 532578 342220 532584
rect 341156 531140 341208 531146
rect 341156 531082 341208 531088
rect 341984 531140 342036 531146
rect 341984 531082 342036 531088
rect 341168 528850 341196 531082
rect 342180 528850 342208 532578
rect 322552 528822 322888 528850
rect 323656 528822 323992 528850
rect 324760 528822 325096 528850
rect 325772 528822 326108 528850
rect 326876 528822 327028 528850
rect 327980 528822 328408 528850
rect 328992 528822 329328 528850
rect 330096 528822 330432 528850
rect 331200 528822 331536 528850
rect 332304 528822 332456 528850
rect 333316 528822 333652 528850
rect 334420 528822 334756 528850
rect 335524 528822 335860 528850
rect 336536 528822 336596 528850
rect 337640 528822 337976 528850
rect 338744 528822 339172 528850
rect 339848 528822 340184 528850
rect 340860 528822 341196 528850
rect 341964 528822 342208 528850
rect 343560 528714 343588 568346
rect 343744 567390 343772 570044
rect 345506 570030 346256 570058
rect 346124 568540 346176 568546
rect 346124 568482 346176 568488
rect 343732 567384 343784 567390
rect 343732 567326 343784 567332
rect 344376 532704 344428 532710
rect 344376 532646 344428 532652
rect 344388 528850 344416 532646
rect 344928 531548 344980 531554
rect 344928 531490 344980 531496
rect 344940 531010 344968 531490
rect 346136 531146 346164 568482
rect 346228 533254 346256 570030
rect 347332 567322 347360 570044
rect 347688 567792 347740 567798
rect 347688 567734 347740 567740
rect 347320 567316 347372 567322
rect 347320 567258 347372 567264
rect 346216 533248 346268 533254
rect 346216 533190 346268 533196
rect 346308 531956 346360 531962
rect 346308 531898 346360 531904
rect 345480 531140 345532 531146
rect 345480 531082 345532 531088
rect 346124 531140 346176 531146
rect 346124 531082 346176 531088
rect 344928 531004 344980 531010
rect 344928 530946 344980 530952
rect 345492 528850 345520 531082
rect 346320 528850 346348 531898
rect 347700 528850 347728 567734
rect 349080 533186 349108 570044
rect 350448 567588 350500 567594
rect 350448 567530 350500 567536
rect 349068 533180 349120 533186
rect 349068 533122 349120 533128
rect 348700 531888 348752 531894
rect 348700 531830 348752 531836
rect 347780 531480 347832 531486
rect 347780 531422 347832 531428
rect 347792 531214 347820 531422
rect 347780 531208 347832 531214
rect 347780 531150 347832 531156
rect 348712 528850 348740 531830
rect 350460 531146 350488 567530
rect 350920 567254 350948 570044
rect 352682 570030 353248 570058
rect 351736 567520 351788 567526
rect 351736 567462 351788 567468
rect 350908 567248 350960 567254
rect 350908 567190 350960 567196
rect 350908 531820 350960 531826
rect 350908 531762 350960 531768
rect 349804 531140 349856 531146
rect 349804 531082 349856 531088
rect 350448 531140 350500 531146
rect 350448 531082 350500 531088
rect 349816 528850 349844 531082
rect 350920 528850 350948 531762
rect 351748 528850 351776 567462
rect 353220 535226 353248 570030
rect 354416 570030 354522 570058
rect 354416 569974 354444 570030
rect 354404 569968 354456 569974
rect 354404 569910 354456 569916
rect 354588 569968 354640 569974
rect 354588 569910 354640 569916
rect 354496 543040 354548 543046
rect 354496 542982 354548 542988
rect 353208 535220 353260 535226
rect 353208 535162 353260 535168
rect 353024 531752 353076 531758
rect 353024 531694 353076 531700
rect 353036 528850 353064 531694
rect 353208 531412 353260 531418
rect 353208 531354 353260 531360
rect 353220 531282 353248 531354
rect 353208 531276 353260 531282
rect 353208 531218 353260 531224
rect 354508 531146 354536 542982
rect 354600 533118 354628 569910
rect 356256 567254 356284 570044
rect 356244 567248 356296 567254
rect 356244 567190 356296 567196
rect 357348 567248 357400 567254
rect 357348 567190 357400 567196
rect 355876 563712 355928 563718
rect 355876 563654 355928 563660
rect 354588 533112 354640 533118
rect 354588 533054 354640 533060
rect 355232 531684 355284 531690
rect 355232 531626 355284 531632
rect 354036 531140 354088 531146
rect 354036 531082 354088 531088
rect 354496 531140 354548 531146
rect 354496 531082 354548 531088
rect 354048 528850 354076 531082
rect 355244 528850 355272 531626
rect 355888 529122 355916 563654
rect 357360 562986 357388 567190
rect 358096 565214 358124 570044
rect 359844 567254 359872 570044
rect 361592 570030 361698 570058
rect 362972 570030 363446 570058
rect 364352 570030 365194 570058
rect 365732 570030 367034 570058
rect 368492 570030 368782 570058
rect 369872 570030 370622 570058
rect 371344 570030 372370 570058
rect 374012 570030 374210 570058
rect 375392 570030 375958 570058
rect 376772 570030 377798 570058
rect 358820 567248 358872 567254
rect 358820 567190 358872 567196
rect 359832 567248 359884 567254
rect 359832 567190 359884 567196
rect 358084 565208 358136 565214
rect 358084 565150 358136 565156
rect 357268 562958 357388 562986
rect 357268 553466 357296 562958
rect 358832 558210 358860 567190
rect 361592 566506 361620 570030
rect 361580 566500 361632 566506
rect 361580 566442 361632 566448
rect 362972 562358 363000 570030
rect 364352 563106 364380 570030
rect 364340 563100 364392 563106
rect 364340 563042 364392 563048
rect 365732 562358 365760 570030
rect 368388 565888 368440 565894
rect 368388 565830 368440 565836
rect 362960 562352 363012 562358
rect 362960 562294 363012 562300
rect 364248 562352 364300 562358
rect 364248 562294 364300 562300
rect 365720 562352 365772 562358
rect 365720 562294 365772 562300
rect 367008 562352 367060 562358
rect 367008 562294 367060 562300
rect 362868 560992 362920 560998
rect 362868 560934 362920 560940
rect 358820 558204 358872 558210
rect 358820 558146 358872 558152
rect 360108 558204 360160 558210
rect 360108 558146 360160 558152
rect 357176 553438 357296 553466
rect 357176 536178 357204 553438
rect 358728 540252 358780 540258
rect 358728 540194 358780 540200
rect 357164 536172 357216 536178
rect 357164 536114 357216 536120
rect 357348 531616 357400 531622
rect 357348 531558 357400 531564
rect 355888 529094 355962 529122
rect 344080 528822 344416 528850
rect 345184 528822 345520 528850
rect 346288 528822 346348 528850
rect 347392 528822 347728 528850
rect 348404 528822 348740 528850
rect 349508 528822 349844 528850
rect 350612 528822 350948 528850
rect 351624 528822 351776 528850
rect 352728 528822 353064 528850
rect 353832 528822 354076 528850
rect 354936 528822 355272 528850
rect 355934 528836 355962 529094
rect 357360 528850 357388 531558
rect 357052 528822 357388 528850
rect 358740 528714 358768 540194
rect 360120 537538 360148 558146
rect 360108 537532 360160 537538
rect 360108 537474 360160 537480
rect 360568 536104 360620 536110
rect 360568 536046 360620 536052
rect 359464 531548 359516 531554
rect 359464 531490 359516 531496
rect 359476 528850 359504 531490
rect 360580 528850 360608 536046
rect 361488 531480 361540 531486
rect 361488 531422 361540 531428
rect 361500 528850 361528 531422
rect 362880 528850 362908 560934
rect 364260 554062 364288 562294
rect 365628 562284 365680 562290
rect 365628 562226 365680 562232
rect 364248 554056 364300 554062
rect 364248 553998 364300 554004
rect 363788 531412 363840 531418
rect 363788 531354 363840 531360
rect 363800 528850 363828 531354
rect 365640 528986 365668 562226
rect 366916 546508 366968 546514
rect 366916 546450 366968 546456
rect 366824 538892 366876 538898
rect 366824 538834 366876 538840
rect 366836 528986 366864 538834
rect 359168 528822 359504 528850
rect 360272 528822 360608 528850
rect 361376 528822 361528 528850
rect 362480 528822 362908 528850
rect 363492 528822 363828 528850
rect 365088 528958 365668 528986
rect 366284 528958 366864 528986
rect 365088 528714 365116 528958
rect 366284 528850 366312 528958
rect 366928 528850 366956 546450
rect 367020 535294 367048 562294
rect 367008 535288 367060 535294
rect 367008 535230 367060 535236
rect 365700 528822 366312 528850
rect 366712 528822 366956 528850
rect 368400 528714 368428 565830
rect 368492 528850 368520 570030
rect 369872 565894 369900 570030
rect 369860 565888 369912 565894
rect 369860 565830 369912 565836
rect 369860 563100 369912 563106
rect 369860 563042 369912 563048
rect 369872 535378 369900 563042
rect 371240 554056 371292 554062
rect 371240 553998 371292 554004
rect 369872 535350 370544 535378
rect 369860 535288 369912 535294
rect 369860 535230 369912 535236
rect 369872 528850 369900 535230
rect 370516 528850 370544 535350
rect 371252 528986 371280 553998
rect 371344 546514 371372 570030
rect 372620 566500 372672 566506
rect 372620 566442 372672 566448
rect 371332 546508 371384 546514
rect 371332 546450 371384 546456
rect 371252 528958 371556 528986
rect 371528 528850 371556 528958
rect 368492 528822 368920 528850
rect 369872 528822 370024 528850
rect 370516 528822 371036 528850
rect 371528 528822 372140 528850
rect 321296 528686 321448 528714
rect 343068 528686 343588 528714
rect 358156 528686 358768 528714
rect 364596 528686 365116 528714
rect 367816 528686 368428 528714
rect 372632 528714 372660 566442
rect 374012 538898 374040 570030
rect 375392 562358 375420 570030
rect 375564 565140 375616 565146
rect 375564 565082 375616 565088
rect 375380 562352 375432 562358
rect 375380 562294 375432 562300
rect 374000 538892 374052 538898
rect 374000 538834 374052 538840
rect 374092 537532 374144 537538
rect 374092 537474 374144 537480
rect 374104 528850 374132 537474
rect 375576 528850 375604 565082
rect 376116 536172 376168 536178
rect 376116 536114 376168 536120
rect 374104 528822 374256 528850
rect 375360 528822 375604 528850
rect 376128 528850 376156 536114
rect 376772 531418 376800 570030
rect 379532 567610 379560 570044
rect 380912 570030 381386 570058
rect 382292 570030 383134 570058
rect 383764 570030 384974 570058
rect 386432 570030 386722 570058
rect 387904 570030 388562 570058
rect 389284 570030 390310 570058
rect 391952 570030 392150 570058
rect 393332 570030 393898 570058
rect 394804 570030 395738 570058
rect 379532 567582 379652 567610
rect 379520 567248 379572 567254
rect 379520 567190 379572 567196
rect 378232 535220 378284 535226
rect 378232 535162 378284 535168
rect 377220 533112 377272 533118
rect 377220 533054 377272 533060
rect 376760 531412 376812 531418
rect 376760 531354 376812 531360
rect 377232 528850 377260 533054
rect 378244 528850 378272 535162
rect 379532 528850 379560 567190
rect 379624 560998 379652 567582
rect 379612 560992 379664 560998
rect 379612 560934 379664 560940
rect 380440 533180 380492 533186
rect 380440 533122 380492 533128
rect 380452 528850 380480 533122
rect 380912 531486 380940 570030
rect 380992 567316 381044 567322
rect 380992 567258 381044 567264
rect 380900 531480 380952 531486
rect 380900 531422 380952 531428
rect 376128 528822 376464 528850
rect 377232 528822 377568 528850
rect 378244 528822 378580 528850
rect 379532 528822 379684 528850
rect 380452 528822 380788 528850
rect 381004 528714 381032 567258
rect 382292 536110 382320 570030
rect 383660 567384 383712 567390
rect 383660 567326 383712 567332
rect 382280 536104 382332 536110
rect 382280 536046 382332 536052
rect 382556 533248 382608 533254
rect 382556 533190 382608 533196
rect 382568 528850 382596 533190
rect 383672 528850 383700 567326
rect 383764 531554 383792 570030
rect 385040 567452 385092 567458
rect 385040 567394 385092 567400
rect 385052 533474 385080 567394
rect 386432 540258 386460 570030
rect 387800 567656 387852 567662
rect 387800 567598 387852 567604
rect 386420 540252 386472 540258
rect 386420 540194 386472 540200
rect 386880 534064 386932 534070
rect 386880 534006 386932 534012
rect 385052 533446 385632 533474
rect 385132 533316 385184 533322
rect 385132 533258 385184 533264
rect 383752 531548 383804 531554
rect 383752 531490 383804 531496
rect 385144 528850 385172 533258
rect 382568 528822 382904 528850
rect 383672 528822 384008 528850
rect 385112 528822 385172 528850
rect 385604 528714 385632 533446
rect 386892 528850 386920 534006
rect 387812 528850 387840 567598
rect 387904 531622 387932 570030
rect 389180 567724 389232 567730
rect 389180 567666 389232 567672
rect 389192 534154 389220 567666
rect 389284 563718 389312 570030
rect 389272 563712 389324 563718
rect 389272 563654 389324 563660
rect 389192 534126 389956 534154
rect 389180 533996 389232 534002
rect 389180 533938 389232 533944
rect 387892 531616 387944 531622
rect 387892 531558 387944 531564
rect 389192 528850 389220 533938
rect 389928 528986 389956 534126
rect 391204 533928 391256 533934
rect 391204 533870 391256 533876
rect 389928 528958 390140 528986
rect 390112 528850 390140 528958
rect 391216 528850 391244 533870
rect 391952 531690 391980 570030
rect 392032 568472 392084 568478
rect 392032 568414 392084 568420
rect 391940 531684 391992 531690
rect 391940 531626 391992 531632
rect 392044 528986 392072 568414
rect 393332 543046 393360 570030
rect 393320 543040 393372 543046
rect 393320 542982 393372 542988
rect 393320 533860 393372 533866
rect 393320 533802 393372 533808
rect 392044 528958 392348 528986
rect 392320 528850 392348 528958
rect 393332 528850 393360 533802
rect 394804 531758 394832 570030
rect 394884 568336 394936 568342
rect 394884 568278 394936 568284
rect 394792 531752 394844 531758
rect 394792 531694 394844 531700
rect 394896 528850 394924 568278
rect 397472 567526 397500 570044
rect 398852 570030 399326 570058
rect 397460 567520 397512 567526
rect 397460 567462 397512 567468
rect 396080 541680 396132 541686
rect 396080 541622 396132 541628
rect 395528 532568 395580 532574
rect 395528 532510 395580 532516
rect 386892 528822 387228 528850
rect 387812 528822 388332 528850
rect 389192 528822 389344 528850
rect 390112 528822 390448 528850
rect 391216 528822 391552 528850
rect 392320 528822 392656 528850
rect 393332 528822 393668 528850
rect 394772 528822 394924 528850
rect 395540 528850 395568 532510
rect 396092 528986 396120 541622
rect 397644 532432 397696 532438
rect 397644 532374 397696 532380
rect 396092 528958 396580 528986
rect 396552 528850 396580 528958
rect 397656 528850 397684 532374
rect 398852 531826 398880 570030
rect 401060 567594 401088 570044
rect 401612 570030 402914 570058
rect 401048 567588 401100 567594
rect 401048 567530 401100 567536
rect 400312 552696 400364 552702
rect 400312 552638 400364 552644
rect 398932 533792 398984 533798
rect 398932 533734 398984 533740
rect 398840 531820 398892 531826
rect 398840 531762 398892 531768
rect 398944 528850 398972 533734
rect 400324 528850 400352 552638
rect 401508 532432 401560 532438
rect 401508 532374 401560 532380
rect 401520 528850 401548 532374
rect 401612 531894 401640 570030
rect 404648 567798 404676 570044
rect 405752 570030 406502 570058
rect 404636 567792 404688 567798
rect 404636 567734 404688 567740
rect 403072 533044 403124 533050
rect 403072 532986 403124 532992
rect 401600 531888 401652 531894
rect 401600 531830 401652 531836
rect 395540 528822 395876 528850
rect 396552 528822 396888 528850
rect 397656 528822 397992 528850
rect 398944 528822 399096 528850
rect 400200 528822 400352 528850
rect 401212 528822 401548 528850
rect 403084 528850 403112 532986
rect 404452 532976 404504 532982
rect 404452 532918 404504 532924
rect 404464 528850 404492 532918
rect 405752 531962 405780 570030
rect 408236 568546 408264 570044
rect 409892 570030 409998 570058
rect 408224 568540 408276 568546
rect 408224 568482 408276 568488
rect 407396 532908 407448 532914
rect 407396 532850 407448 532856
rect 405740 531956 405792 531962
rect 405740 531898 405792 531904
rect 405188 529848 405240 529854
rect 405188 529790 405240 529796
rect 403084 528822 403420 528850
rect 404432 528822 404492 528850
rect 405200 528850 405228 529790
rect 407408 528850 407436 532850
rect 409892 532710 409920 570030
rect 411824 568410 411852 570044
rect 412652 570030 413586 570058
rect 411812 568404 411864 568410
rect 411812 568346 411864 568352
rect 409880 532704 409932 532710
rect 409880 532646 409932 532652
rect 412652 532642 412680 570030
rect 415412 568274 415440 570044
rect 416792 570030 417174 570058
rect 415400 568268 415452 568274
rect 415400 568210 415452 568216
rect 412732 532840 412784 532846
rect 412732 532782 412784 532788
rect 412640 532636 412692 532642
rect 412640 532578 412692 532584
rect 408590 531992 408646 532001
rect 408590 531927 408646 531936
rect 408604 528850 408632 531927
rect 409880 530936 409932 530942
rect 409880 530878 409932 530884
rect 409892 528850 409920 530878
rect 411628 530868 411680 530874
rect 411628 530810 411680 530816
rect 405200 528822 405536 528850
rect 407408 528822 407744 528850
rect 408604 528822 408756 528850
rect 409860 528822 409920 528850
rect 411640 528850 411668 530810
rect 412744 528850 412772 532782
rect 416792 532506 416820 570030
rect 419000 568206 419028 570044
rect 419552 570030 420762 570058
rect 418988 568200 419040 568206
rect 418988 568142 419040 568148
rect 416780 532500 416832 532506
rect 416780 532442 416832 532448
rect 419552 532370 419580 570030
rect 422588 568138 422616 570044
rect 423692 570030 424350 570058
rect 422576 568132 422628 568138
rect 422576 568074 422628 568080
rect 421378 533216 421434 533225
rect 421378 533151 421434 533160
rect 419632 532772 419684 532778
rect 419632 532714 419684 532720
rect 419540 532364 419592 532370
rect 419540 532306 419592 532312
rect 414020 530800 414072 530806
rect 414020 530742 414072 530748
rect 414032 528850 414060 530742
rect 415952 530732 416004 530738
rect 415952 530674 416004 530680
rect 415964 528850 415992 530674
rect 418252 530664 418304 530670
rect 418252 530606 418304 530612
rect 417056 529780 417108 529786
rect 417056 529722 417108 529728
rect 417068 528850 417096 529722
rect 418264 528850 418292 530606
rect 419644 528850 419672 532714
rect 420276 530596 420328 530602
rect 420276 530538 420328 530544
rect 411640 528822 411976 528850
rect 412744 528822 413080 528850
rect 414032 528822 414184 528850
rect 415964 528822 416300 528850
rect 417068 528822 417404 528850
rect 418264 528822 418508 528850
rect 419520 528822 419672 528850
rect 420288 528850 420316 530538
rect 421392 528850 421420 533151
rect 423692 532302 423720 570030
rect 426176 568070 426204 570044
rect 427832 570030 427938 570058
rect 426164 568064 426216 568070
rect 426164 568006 426216 568012
rect 425702 533080 425758 533089
rect 425702 533015 425758 533024
rect 423680 532296 423732 532302
rect 423680 532238 423732 532244
rect 422484 530528 422536 530534
rect 422484 530470 422536 530476
rect 422496 528850 422524 530470
rect 424600 530460 424652 530466
rect 424600 530402 424652 530408
rect 424612 528850 424640 530402
rect 425716 528850 425744 533015
rect 427832 532234 427860 570030
rect 429764 568002 429792 570044
rect 430592 570030 431526 570058
rect 429752 567996 429804 568002
rect 429752 567938 429804 567944
rect 430026 532944 430082 532953
rect 430026 532879 430082 532888
rect 427820 532228 427872 532234
rect 427820 532170 427872 532176
rect 429292 531072 429344 531078
rect 429292 531014 429344 531020
rect 426716 530392 426768 530398
rect 426716 530334 426768 530340
rect 426728 528850 426756 530334
rect 429304 528850 429332 531014
rect 420288 528822 420624 528850
rect 421392 528822 421728 528850
rect 422496 528822 422832 528850
rect 424612 528822 424948 528850
rect 425716 528822 426052 528850
rect 426728 528822 427064 528850
rect 429272 528822 429332 528850
rect 430040 528850 430068 532879
rect 430592 532166 430620 570030
rect 433352 567934 433380 570044
rect 434732 570030 435114 570058
rect 433340 567928 433392 567934
rect 433340 567870 433392 567876
rect 430580 532160 430632 532166
rect 430580 532102 430632 532108
rect 434732 532098 434760 570030
rect 436940 567866 436968 570044
rect 437492 570030 438702 570058
rect 436928 567860 436980 567866
rect 436928 567802 436980 567808
rect 436008 535152 436060 535158
rect 436008 535094 436060 535100
rect 434720 532092 434772 532098
rect 434720 532034 434772 532040
rect 434258 531856 434314 531865
rect 434258 531791 434314 531800
rect 433340 531004 433392 531010
rect 433340 530946 433392 530952
rect 431040 529916 431092 529922
rect 431040 529858 431092 529864
rect 431052 528850 431080 529858
rect 433352 528850 433380 530946
rect 434272 528850 434300 531791
rect 435364 531140 435416 531146
rect 435364 531082 435416 531088
rect 435376 528850 435404 531082
rect 436020 530602 436048 535094
rect 437492 532030 437520 570030
rect 440528 567905 440556 570044
rect 441632 570030 442290 570058
rect 443012 570030 444130 570058
rect 445772 570030 445878 570058
rect 447152 570030 447718 570058
rect 448532 570030 449466 570058
rect 440514 567896 440570 567905
rect 440514 567831 440570 567840
rect 441632 532137 441660 570030
rect 442908 535016 442960 535022
rect 442908 534958 442960 534964
rect 441802 532808 441858 532817
rect 441802 532743 441858 532752
rect 441618 532128 441674 532137
rect 441618 532063 441674 532072
rect 437480 532024 437532 532030
rect 437480 531966 437532 531972
rect 440790 531720 440846 531729
rect 440790 531655 440846 531664
rect 439688 531276 439740 531282
rect 439688 531218 439740 531224
rect 437664 531208 437716 531214
rect 437664 531150 437716 531156
rect 436008 530596 436060 530602
rect 436008 530538 436060 530544
rect 436468 529712 436520 529718
rect 436468 529654 436520 529660
rect 436480 528850 436508 529654
rect 437676 528850 437704 531150
rect 438952 529644 439004 529650
rect 438952 529586 439004 529592
rect 438964 528850 438992 529586
rect 430040 528822 430376 528850
rect 431052 528822 431388 528850
rect 433352 528822 433596 528850
rect 434272 528822 434608 528850
rect 435376 528822 435712 528850
rect 436480 528822 436816 528850
rect 437676 528822 437920 528850
rect 438932 528822 438992 528850
rect 439700 528850 439728 531218
rect 440804 528850 440832 531655
rect 441816 528850 441844 532743
rect 442920 531282 442948 534958
rect 443012 533730 443040 570030
rect 443000 533724 443052 533730
rect 443000 533666 443052 533672
rect 445772 533662 445800 570030
rect 446128 535084 446180 535090
rect 446128 535026 446180 535032
rect 445760 533656 445812 533662
rect 445760 533598 445812 533604
rect 442998 531584 443054 531593
rect 442998 531519 443054 531528
rect 442908 531276 442960 531282
rect 442908 531218 442960 531224
rect 443012 528850 443040 531519
rect 444380 530596 444432 530602
rect 444380 530538 444432 530544
rect 444392 528850 444420 530538
rect 445116 529576 445168 529582
rect 445116 529518 445168 529524
rect 439700 528822 440036 528850
rect 440804 528822 441140 528850
rect 441816 528822 442152 528850
rect 443012 528822 443256 528850
rect 444360 528822 444420 528850
rect 445128 528850 445156 529518
rect 446140 528850 446168 535026
rect 447152 533594 447180 570030
rect 447140 533588 447192 533594
rect 447140 533530 447192 533536
rect 448532 533526 448560 570030
rect 450452 534948 450504 534954
rect 450452 534890 450504 534896
rect 448520 533520 448572 533526
rect 448520 533462 448572 533468
rect 448520 531276 448572 531282
rect 448520 531218 448572 531224
rect 447324 529508 447376 529514
rect 447324 529450 447376 529456
rect 447336 528850 447364 529450
rect 448532 528850 448560 531218
rect 449440 529440 449492 529446
rect 449440 529382 449492 529388
rect 449452 528850 449480 529382
rect 450464 528850 450492 534890
rect 451292 533458 451320 570044
rect 452672 570030 453054 570058
rect 452568 534880 452620 534886
rect 452568 534822 452620 534828
rect 451280 533452 451332 533458
rect 451280 533394 451332 533400
rect 452580 529938 452608 534822
rect 452672 533390 452700 570030
rect 452660 533384 452712 533390
rect 452660 533326 452712 533332
rect 455432 532438 455460 591631
rect 456076 568546 456104 635151
rect 551374 632224 551430 632233
rect 551112 632182 551374 632210
rect 456800 616820 456852 616826
rect 456800 616762 456852 616768
rect 456812 616321 456840 616762
rect 456798 616312 456854 616321
rect 456798 616247 456854 616256
rect 483032 568546 483060 570044
rect 529032 568546 529060 570044
rect 550822 569800 550878 569809
rect 550822 569735 550878 569744
rect 551006 569800 551062 569809
rect 551006 569735 551062 569744
rect 550836 569537 550864 569735
rect 550822 569528 550878 569537
rect 550822 569463 550878 569472
rect 456064 568540 456116 568546
rect 456064 568482 456116 568488
rect 483020 568540 483072 568546
rect 483020 568482 483072 568488
rect 529020 568540 529072 568546
rect 529020 568482 529072 568488
rect 529848 568540 529900 568546
rect 529848 568482 529900 568488
rect 455420 532432 455472 532438
rect 455420 532374 455472 532380
rect 454774 531448 454830 531457
rect 454774 531383 454830 531392
rect 452580 529910 452700 529938
rect 451556 529372 451608 529378
rect 451556 529314 451608 529320
rect 451568 528850 451596 529314
rect 452672 528850 452700 529910
rect 454040 529168 454092 529174
rect 454040 529110 454092 529116
rect 454052 528850 454080 529110
rect 445128 528822 445464 528850
rect 446140 528822 446476 528850
rect 447336 528822 447580 528850
rect 448532 528822 448684 528850
rect 449452 528822 449788 528850
rect 450464 528822 450800 528850
rect 451568 528822 451904 528850
rect 452672 528822 453008 528850
rect 454020 528822 454080 528850
rect 454788 528850 454816 531383
rect 454788 528822 455124 528850
rect 372632 528686 373244 528714
rect 381004 528686 381800 528714
rect 385604 528686 386124 528714
rect 456076 528562 456104 568482
rect 493966 560960 494022 560969
rect 493966 560895 494022 560904
rect 483848 534812 483900 534818
rect 483848 534754 483900 534760
rect 456984 534744 457036 534750
rect 456984 534686 457036 534692
rect 456202 529100 456254 529106
rect 456202 529042 456254 529048
rect 456214 528836 456242 529042
rect 456996 528850 457024 534686
rect 459100 534676 459152 534682
rect 459100 534618 459152 534624
rect 458318 529032 458370 529038
rect 458318 528974 458370 528980
rect 456996 528822 457332 528850
rect 458330 528836 458358 528974
rect 459112 528850 459140 534618
rect 461216 534608 461268 534614
rect 461216 534550 461268 534556
rect 460204 528964 460256 528970
rect 460204 528906 460256 528912
rect 460216 528850 460244 528906
rect 461228 528850 461256 534550
rect 464528 534540 464580 534546
rect 464528 534482 464580 534488
rect 463792 530324 463844 530330
rect 463792 530266 463844 530272
rect 462320 528896 462372 528902
rect 459112 528822 459448 528850
rect 460216 528822 460552 528850
rect 461228 528822 461564 528850
rect 463804 528850 463832 530266
rect 462372 528844 462668 528850
rect 462320 528838 462668 528844
rect 462332 528822 462668 528838
rect 463772 528822 463832 528850
rect 464540 528850 464568 534482
rect 466644 534472 466696 534478
rect 466644 534414 466696 534420
rect 465540 530256 465592 530262
rect 465540 530198 465592 530204
rect 465552 528850 465580 530198
rect 466656 528850 466684 534414
rect 468760 534404 468812 534410
rect 468760 534346 468812 534352
rect 467840 530188 467892 530194
rect 467840 530130 467892 530136
rect 467852 528850 467880 530130
rect 468772 528850 468800 534346
rect 470968 534336 471020 534342
rect 470968 534278 471020 534284
rect 469864 530120 469916 530126
rect 469864 530062 469916 530068
rect 469876 528850 469904 530062
rect 470980 528850 471008 534278
rect 473452 534268 473504 534274
rect 473452 534210 473504 534216
rect 471704 530256 471756 530262
rect 471704 530198 471756 530204
rect 464540 528822 464876 528850
rect 465552 528822 465888 528850
rect 466656 528822 466992 528850
rect 467852 528822 468096 528850
rect 468772 528822 469108 528850
rect 469876 528822 470212 528850
rect 470980 528822 471316 528850
rect 315948 528556 316000 528562
rect 315948 528498 316000 528504
rect 456064 528556 456116 528562
rect 456064 528498 456116 528504
rect 315960 515817 315988 528498
rect 401968 528488 402020 528494
rect 402020 528436 402316 528442
rect 401968 528430 402316 528436
rect 401980 528414 402316 528430
rect 406304 528426 406640 528442
rect 406292 528420 406640 528426
rect 406344 528414 406640 528420
rect 406292 528362 406344 528368
rect 410616 528352 410668 528358
rect 471716 528329 471744 530198
rect 472072 530052 472124 530058
rect 472072 529994 472124 530000
rect 472084 528850 472112 529994
rect 473464 528850 473492 534210
rect 475292 534200 475344 534206
rect 475292 534142 475344 534148
rect 474188 529984 474240 529990
rect 474188 529926 474240 529932
rect 472084 528822 472420 528850
rect 473432 528822 473492 528850
rect 474200 528850 474228 529926
rect 475304 528850 475332 534142
rect 481732 530256 481784 530262
rect 477498 530224 477554 530233
rect 481732 530198 481784 530204
rect 477498 530159 477554 530168
rect 478880 530188 478932 530194
rect 477512 528850 477540 530159
rect 478880 530130 478932 530136
rect 478892 528850 478920 530130
rect 480626 530088 480682 530097
rect 480626 530023 480682 530032
rect 474200 528822 474536 528850
rect 475304 528822 475640 528850
rect 476316 528834 476652 528850
rect 476304 528828 476652 528834
rect 476356 528822 476652 528828
rect 477512 528822 477756 528850
rect 478860 528822 478920 528850
rect 480640 528850 480668 530023
rect 481548 529984 481600 529990
rect 481548 529926 481600 529932
rect 481560 529310 481588 529926
rect 481548 529304 481600 529310
rect 481548 529246 481600 529252
rect 481744 528850 481772 530198
rect 482928 530052 482980 530058
rect 482928 529994 482980 530000
rect 482940 529242 482968 529994
rect 482928 529236 482980 529242
rect 482928 529178 482980 529184
rect 483860 528850 483888 534754
rect 493782 534712 493838 534721
rect 493782 534647 493838 534656
rect 487160 534132 487212 534138
rect 487160 534074 487212 534080
rect 484952 529984 485004 529990
rect 484952 529926 485004 529932
rect 484964 528850 484992 529926
rect 487172 528850 487200 534074
rect 492034 531176 492090 531185
rect 492034 531111 492090 531120
rect 488540 530052 488592 530058
rect 488540 529994 488592 530000
rect 488552 528850 488580 529994
rect 490378 529952 490434 529961
rect 490378 529887 490434 529896
rect 480640 528822 480976 528850
rect 481744 528822 482080 528850
rect 483860 528822 484196 528850
rect 484964 528822 485300 528850
rect 487172 528822 487508 528850
rect 488520 528822 488580 528850
rect 490392 528850 490420 529887
rect 492048 528850 492076 531111
rect 493140 530188 493192 530194
rect 493140 530130 493192 530136
rect 493152 528850 493180 530130
rect 490392 528822 490728 528850
rect 491740 528822 492076 528850
rect 492844 528822 493180 528850
rect 476304 528770 476356 528776
rect 479616 528760 479668 528766
rect 493796 528714 493824 534647
rect 493980 530194 494008 560895
rect 499486 545728 499542 545737
rect 499486 545663 499542 545672
rect 498566 532400 498622 532409
rect 498566 532335 498622 532344
rect 495346 532264 495402 532273
rect 495346 532199 495402 532208
rect 493968 530188 494020 530194
rect 493968 530130 494020 530136
rect 495360 528850 495388 532199
rect 497462 532128 497518 532137
rect 497462 532063 497518 532072
rect 496358 531992 496414 532001
rect 496358 531927 496414 531936
rect 496372 528850 496400 531927
rect 497476 528850 497504 532063
rect 498580 528850 498608 532335
rect 499500 528850 499528 545663
rect 508226 533624 508282 533633
rect 508226 533559 508282 533568
rect 514668 533588 514720 533594
rect 506110 533488 506166 533497
rect 506110 533423 506166 533432
rect 501786 533352 501842 533361
rect 501786 533287 501842 533296
rect 500682 530768 500738 530777
rect 500682 530703 500738 530712
rect 500696 528850 500724 530703
rect 501800 528850 501828 533287
rect 505006 532672 505062 532681
rect 505006 532607 505062 532616
rect 503626 532536 503682 532545
rect 503626 532471 503682 532480
rect 502890 530632 502946 530641
rect 502890 530567 502946 530576
rect 502904 528850 502932 530567
rect 503640 528850 503668 532471
rect 505020 528850 505048 532607
rect 506124 528850 506152 533423
rect 507122 531040 507178 531049
rect 507122 530975 507178 530984
rect 507136 528850 507164 530975
rect 508240 528850 508268 533559
rect 514668 533530 514720 533536
rect 512552 533520 512604 533526
rect 512552 533462 512604 533468
rect 510436 533452 510488 533458
rect 510436 533394 510488 533400
rect 509054 530904 509110 530913
rect 509054 530839 509110 530848
rect 509068 528850 509096 530839
rect 510448 528850 510476 533394
rect 511448 530596 511500 530602
rect 511448 530538 511500 530544
rect 511460 528850 511488 530538
rect 512564 528850 512592 533462
rect 513656 530664 513708 530670
rect 513656 530606 513708 530612
rect 513668 528850 513696 530606
rect 514680 528850 514708 533530
rect 529860 533390 529888 568482
rect 551020 563281 551048 569735
rect 551006 563272 551062 563281
rect 551006 563207 551062 563216
rect 551006 560280 551062 560289
rect 551006 560215 551062 560224
rect 551020 555529 551048 560215
rect 551006 555520 551062 555529
rect 551006 555455 551062 555464
rect 543648 547256 543700 547262
rect 543648 547198 543700 547204
rect 540888 547188 540940 547194
rect 540888 547130 540940 547136
rect 530860 533656 530912 533662
rect 530860 533598 530912 533604
rect 529848 533384 529900 533390
rect 529848 533326 529900 533332
rect 527640 532364 527692 532370
rect 527640 532306 527692 532312
rect 525524 532228 525576 532234
rect 525524 532170 525576 532176
rect 523316 532160 523368 532166
rect 523316 532102 523368 532108
rect 521200 532092 521252 532098
rect 521200 532034 521252 532040
rect 518716 532024 518768 532030
rect 518716 531966 518768 531972
rect 516874 531856 516930 531865
rect 516874 531791 516930 531800
rect 515770 531176 515826 531185
rect 515770 531111 515826 531120
rect 515784 528850 515812 531111
rect 516888 528850 516916 531791
rect 517980 530732 518032 530738
rect 517980 530674 518032 530680
rect 517992 528850 518020 530674
rect 518728 528850 518756 531966
rect 520096 530800 520148 530806
rect 520096 530742 520148 530748
rect 520108 528850 520136 530742
rect 521212 528850 521240 532034
rect 522212 530936 522264 530942
rect 522212 530878 522264 530884
rect 522224 528850 522252 530878
rect 523328 528850 523356 532102
rect 524328 530868 524380 530874
rect 524328 530810 524380 530816
rect 524340 528850 524368 530810
rect 525536 528850 525564 532170
rect 526536 531004 526588 531010
rect 526536 530946 526588 530952
rect 526548 528850 526576 530946
rect 527652 528850 527680 532306
rect 529756 532296 529808 532302
rect 529756 532238 529808 532244
rect 528468 531072 528520 531078
rect 528468 531014 528520 531020
rect 528480 528850 528508 531014
rect 529768 528850 529796 532238
rect 530872 528850 530900 533598
rect 536288 532568 536340 532574
rect 536288 532510 536340 532516
rect 531964 532432 532016 532438
rect 531964 532374 532016 532380
rect 531976 528850 532004 532374
rect 535184 531276 535236 531282
rect 535184 531218 535236 531224
rect 533988 531208 534040 531214
rect 533988 531150 534040 531156
rect 533068 531140 533120 531146
rect 533068 531082 533120 531088
rect 533080 528850 533108 531082
rect 534000 528850 534028 531150
rect 535196 528850 535224 531218
rect 536300 528850 536328 532510
rect 538128 532500 538180 532506
rect 538128 532442 538180 532448
rect 537300 530460 537352 530466
rect 537300 530402 537352 530408
rect 537312 528850 537340 530402
rect 538140 528850 538168 532442
rect 539508 530256 539560 530262
rect 539508 530198 539560 530204
rect 539520 528850 539548 530198
rect 540900 528986 540928 547130
rect 543660 530534 543688 547198
rect 545028 547120 545080 547126
rect 545028 547062 545080 547068
rect 542728 530528 542780 530534
rect 542728 530470 542780 530476
rect 543648 530528 543700 530534
rect 543648 530470 543700 530476
rect 541624 530392 541676 530398
rect 541624 530334 541676 530340
rect 540624 528958 540928 528986
rect 540624 528850 540652 528958
rect 541636 528850 541664 530334
rect 542740 528850 542768 530470
rect 543648 530324 543700 530330
rect 543648 530266 543700 530272
rect 543660 528850 543688 530266
rect 545040 528986 545068 547062
rect 547052 532636 547104 532642
rect 547052 532578 547104 532584
rect 545946 531312 546002 531321
rect 545946 531247 546002 531256
rect 544856 528958 545068 528986
rect 544856 528850 544884 528958
rect 545960 528850 545988 531247
rect 547064 528850 547092 532578
rect 549168 532160 549220 532166
rect 549168 532102 549220 532108
rect 548156 530936 548208 530942
rect 548156 530878 548208 530884
rect 548168 528850 548196 530878
rect 549180 528850 549208 532102
rect 551112 532030 551140 632182
rect 551374 632159 551430 632168
rect 551558 628416 551614 628425
rect 551558 628351 551614 628360
rect 551374 628008 551430 628017
rect 551374 627943 551430 627952
rect 551388 627366 551416 627943
rect 551376 627360 551428 627366
rect 551376 627302 551428 627308
rect 551466 622432 551522 622441
rect 551466 622367 551522 622376
rect 551374 621344 551430 621353
rect 551296 621302 551374 621330
rect 551192 618724 551244 618730
rect 551192 618666 551244 618672
rect 551204 606558 551232 618666
rect 551192 606552 551244 606558
rect 551192 606494 551244 606500
rect 551296 606490 551324 621302
rect 551374 621279 551430 621288
rect 551374 618624 551430 618633
rect 551374 618559 551430 618568
rect 551388 617545 551416 618559
rect 551374 617536 551430 617545
rect 551374 617471 551430 617480
rect 551480 615754 551508 622367
rect 551572 618730 551600 628351
rect 551664 628017 551692 639503
rect 551650 628008 551706 628017
rect 551650 627943 551706 627952
rect 551652 627360 551704 627366
rect 551652 627302 551704 627308
rect 551560 618724 551612 618730
rect 551560 618666 551612 618672
rect 551558 618488 551614 618497
rect 551558 618423 551614 618432
rect 551388 615726 551508 615754
rect 551388 611318 551416 615726
rect 551572 615210 551600 618423
rect 551664 616457 551692 627302
rect 551650 616448 551706 616457
rect 551650 616383 551706 616392
rect 551480 615182 551600 615210
rect 551376 611312 551428 611318
rect 551376 611254 551428 611260
rect 551284 606484 551336 606490
rect 551284 606426 551336 606432
rect 551284 606348 551336 606354
rect 551284 606290 551336 606296
rect 551192 598052 551244 598058
rect 551192 597994 551244 598000
rect 551204 582418 551232 597994
rect 551296 597038 551324 606290
rect 551374 601624 551430 601633
rect 551374 601559 551430 601568
rect 551388 601458 551416 601559
rect 551376 601452 551428 601458
rect 551376 601394 551428 601400
rect 551374 599992 551430 600001
rect 551374 599927 551430 599936
rect 551284 597032 551336 597038
rect 551284 596974 551336 596980
rect 551284 596896 551336 596902
rect 551284 596838 551336 596844
rect 551296 587246 551324 596838
rect 551388 596630 551416 599927
rect 551376 596624 551428 596630
rect 551376 596566 551428 596572
rect 551376 596488 551428 596494
rect 551376 596430 551428 596436
rect 551388 595241 551416 596430
rect 551374 595232 551430 595241
rect 551374 595167 551430 595176
rect 551376 595128 551428 595134
rect 551374 595096 551376 595105
rect 551428 595096 551430 595105
rect 551374 595031 551430 595040
rect 551374 592376 551430 592385
rect 551374 592311 551376 592320
rect 551428 592311 551430 592320
rect 551376 592282 551428 592288
rect 551374 592240 551430 592249
rect 551374 592175 551376 592184
rect 551428 592175 551430 592184
rect 551376 592146 551428 592152
rect 551376 592068 551428 592074
rect 551376 592010 551428 592016
rect 551284 587240 551336 587246
rect 551284 587182 551336 587188
rect 551388 587058 551416 592010
rect 551296 587030 551416 587058
rect 551192 582412 551244 582418
rect 551192 582354 551244 582360
rect 551296 576994 551324 587030
rect 551376 586968 551428 586974
rect 551374 586936 551376 586945
rect 551428 586936 551430 586945
rect 551374 586871 551430 586880
rect 551376 586288 551428 586294
rect 551374 586256 551376 586265
rect 551428 586256 551430 586265
rect 551374 586191 551430 586200
rect 551374 582040 551430 582049
rect 551374 581975 551430 581984
rect 551388 577561 551416 581975
rect 551374 577552 551430 577561
rect 551374 577487 551430 577496
rect 551296 576966 551416 576994
rect 551192 576904 551244 576910
rect 551192 576846 551244 576852
rect 551284 576904 551336 576910
rect 551284 576846 551336 576852
rect 551100 532024 551152 532030
rect 551100 531966 551152 531972
rect 551204 531010 551232 576846
rect 551296 531078 551324 576846
rect 551388 532370 551416 576966
rect 551480 533662 551508 615182
rect 551650 613864 551706 613873
rect 551650 613799 551706 613808
rect 551558 612776 551614 612785
rect 551558 612711 551614 612720
rect 551468 533656 551520 533662
rect 551468 533598 551520 533604
rect 551572 532574 551600 612711
rect 551664 612241 551692 613799
rect 551742 613728 551798 613737
rect 551742 613663 551798 613672
rect 551650 612232 551706 612241
rect 551650 612167 551706 612176
rect 551650 611688 551706 611697
rect 551650 611623 551706 611632
rect 551560 532568 551612 532574
rect 551560 532510 551612 532516
rect 551376 532364 551428 532370
rect 551376 532306 551428 532312
rect 551376 531276 551428 531282
rect 551376 531218 551428 531224
rect 551284 531072 551336 531078
rect 551284 531014 551336 531020
rect 551192 531004 551244 531010
rect 551192 530946 551244 530952
rect 550272 530732 550324 530738
rect 550272 530674 550324 530680
rect 550284 528850 550312 530674
rect 551388 528850 551416 531218
rect 551664 530466 551692 611623
rect 551756 601225 551784 613663
rect 551836 611312 551888 611318
rect 551836 611254 551888 611260
rect 551848 606694 551876 611254
rect 551836 606688 551888 606694
rect 551836 606630 551888 606636
rect 551836 606552 551888 606558
rect 551836 606494 551888 606500
rect 551742 601216 551798 601225
rect 551742 601151 551798 601160
rect 551742 600400 551798 600409
rect 551742 600335 551798 600344
rect 551756 532642 551784 600335
rect 551848 598058 551876 606494
rect 551928 606484 551980 606490
rect 551928 606426 551980 606432
rect 551836 598052 551888 598058
rect 551836 597994 551888 598000
rect 551834 597952 551890 597961
rect 551834 597887 551890 597896
rect 551744 532636 551796 532642
rect 551744 532578 551796 532584
rect 551848 532166 551876 597887
rect 551940 596902 551968 606426
rect 551928 596896 551980 596902
rect 551928 596838 551980 596844
rect 551928 596760 551980 596766
rect 551928 596702 551980 596708
rect 551940 592074 551968 596702
rect 551928 592068 551980 592074
rect 551928 592010 551980 592016
rect 551928 587240 551980 587246
rect 551928 587182 551980 587188
rect 551940 576910 551968 587182
rect 551928 576904 551980 576910
rect 551928 576846 551980 576852
rect 551928 572620 551980 572626
rect 551928 572562 551980 572568
rect 551836 532160 551888 532166
rect 551836 532102 551888 532108
rect 551940 531282 551968 572562
rect 552032 533458 552060 641679
rect 553398 641064 553454 641073
rect 553398 640999 553454 641008
rect 552202 639976 552258 639985
rect 552202 639911 552258 639920
rect 552110 638752 552166 638761
rect 552110 638687 552166 638696
rect 552020 533452 552072 533458
rect 552020 533394 552072 533400
rect 551928 531276 551980 531282
rect 551928 531218 551980 531224
rect 552124 530670 552152 638687
rect 552216 533526 552244 639911
rect 552294 637528 552350 637537
rect 552294 637463 552350 637472
rect 552308 533594 552336 637463
rect 552386 631408 552442 631417
rect 552386 631343 552442 631352
rect 552296 533588 552348 533594
rect 552296 533530 552348 533536
rect 552204 533520 552256 533526
rect 552204 533462 552256 533468
rect 552400 531434 552428 631343
rect 552478 624064 552534 624073
rect 552478 623999 552534 624008
rect 552308 531406 552428 531434
rect 552308 530806 552336 531406
rect 552388 531276 552440 531282
rect 552388 531218 552440 531224
rect 552296 530800 552348 530806
rect 552296 530742 552348 530748
rect 552112 530664 552164 530670
rect 552112 530606 552164 530612
rect 551652 530460 551704 530466
rect 551652 530402 551704 530408
rect 552400 528850 552428 531218
rect 552492 531146 552520 623999
rect 552570 614408 552626 614417
rect 552570 614343 552626 614352
rect 552584 531214 552612 614343
rect 553030 608288 553086 608297
rect 553030 608223 553086 608232
rect 552662 604616 552718 604625
rect 552662 604551 552718 604560
rect 552572 531208 552624 531214
rect 552572 531150 552624 531156
rect 552480 531140 552532 531146
rect 552480 531082 552532 531088
rect 552676 530330 552704 604551
rect 552754 599720 552810 599729
rect 552754 599655 552810 599664
rect 552768 530942 552796 599655
rect 552846 597272 552902 597281
rect 552846 597207 552902 597216
rect 552756 530936 552808 530942
rect 552756 530878 552808 530884
rect 552860 530738 552888 597207
rect 552938 594824 552994 594833
rect 552938 594759 552994 594768
rect 552952 531282 552980 594759
rect 553044 547194 553072 608223
rect 553122 605840 553178 605849
rect 553122 605775 553178 605784
rect 553136 547262 553164 605775
rect 553214 603392 553270 603401
rect 553214 603327 553270 603336
rect 553124 547256 553176 547262
rect 553124 547198 553176 547204
rect 553032 547188 553084 547194
rect 553032 547130 553084 547136
rect 553228 547126 553256 603327
rect 553306 596048 553362 596057
rect 553306 595983 553362 595992
rect 553320 576910 553348 595983
rect 553308 576904 553360 576910
rect 553308 576846 553360 576852
rect 553306 576056 553362 576065
rect 553306 575991 553362 576000
rect 553320 575550 553348 575991
rect 553308 575544 553360 575550
rect 553308 575486 553360 575492
rect 553306 574832 553362 574841
rect 553306 574767 553362 574776
rect 553320 574258 553348 574767
rect 553308 574252 553360 574258
rect 553308 574194 553360 574200
rect 553306 574152 553362 574161
rect 553306 574087 553308 574096
rect 553360 574087 553362 574096
rect 553308 574058 553360 574064
rect 553306 572928 553362 572937
rect 553306 572863 553362 572872
rect 553320 572762 553348 572863
rect 553308 572756 553360 572762
rect 553308 572698 553360 572704
rect 553306 571704 553362 571713
rect 553306 571639 553308 571648
rect 553360 571639 553362 571648
rect 553308 571610 553360 571616
rect 553306 570072 553362 570081
rect 553306 570007 553362 570016
rect 553320 569974 553348 570007
rect 553308 569968 553360 569974
rect 553308 569910 553360 569916
rect 553216 547120 553268 547126
rect 553216 547062 553268 547068
rect 552940 531276 552992 531282
rect 552940 531218 552992 531224
rect 552848 530732 552900 530738
rect 552848 530674 552900 530680
rect 553308 530460 553360 530466
rect 553308 530402 553360 530408
rect 552664 530324 552716 530330
rect 552664 530266 552716 530272
rect 553320 528850 553348 530402
rect 553412 530398 553440 640999
rect 553490 633856 553546 633865
rect 553490 633791 553546 633800
rect 553504 530602 553532 633791
rect 553582 630184 553638 630193
rect 553582 630119 553638 630128
rect 553596 532098 553624 630119
rect 553766 627736 553822 627745
rect 553766 627671 553822 627680
rect 553674 626512 553730 626521
rect 553674 626447 553730 626456
rect 553584 532092 553636 532098
rect 553584 532034 553636 532040
rect 553492 530596 553544 530602
rect 553492 530538 553544 530544
rect 553688 530534 553716 626447
rect 553780 532234 553808 627671
rect 553858 625288 553914 625297
rect 553858 625223 553914 625232
rect 553872 532302 553900 625223
rect 553950 620392 554006 620401
rect 553950 620327 554006 620336
rect 553964 532438 553992 620327
rect 554134 617944 554190 617953
rect 554134 617879 554190 617888
rect 554042 615632 554098 615641
rect 554042 615567 554098 615576
rect 553952 532432 554004 532438
rect 553952 532374 554004 532380
rect 553860 532296 553912 532302
rect 553860 532238 553912 532244
rect 553768 532228 553820 532234
rect 553768 532170 553820 532176
rect 554056 530874 554084 615567
rect 554148 532506 554176 617879
rect 554226 616856 554282 616865
rect 554226 616791 554282 616800
rect 554136 532500 554188 532506
rect 554136 532442 554188 532448
rect 554044 530868 554096 530874
rect 554044 530810 554096 530816
rect 553676 530528 553728 530534
rect 553676 530470 553728 530476
rect 553400 530392 553452 530398
rect 553400 530334 553452 530340
rect 554240 530262 554268 616791
rect 554318 610736 554374 610745
rect 554318 610671 554374 610680
rect 554332 532710 554360 610671
rect 554410 609512 554466 609521
rect 554410 609447 554466 609456
rect 554320 532704 554372 532710
rect 554320 532646 554372 532652
rect 554228 530256 554280 530262
rect 554228 530198 554280 530204
rect 554424 530194 554452 609447
rect 554502 607064 554558 607073
rect 554502 606999 554558 607008
rect 554412 530188 554464 530194
rect 554412 530130 554464 530136
rect 554516 530126 554544 606999
rect 554594 593736 554650 593745
rect 554594 593671 554650 593680
rect 554608 590170 554636 593671
rect 554686 592512 554742 592521
rect 554686 592447 554742 592456
rect 554596 590164 554648 590170
rect 554596 590106 554648 590112
rect 554594 590064 554650 590073
rect 554594 589999 554650 590008
rect 554608 589354 554636 589999
rect 554596 589348 554648 589354
rect 554596 589290 554648 589296
rect 554594 588840 554650 588849
rect 554594 588775 554596 588784
rect 554648 588775 554650 588784
rect 554596 588746 554648 588752
rect 554594 587616 554650 587625
rect 554594 587551 554650 587560
rect 554608 587110 554636 587551
rect 554596 587104 554648 587110
rect 554596 587046 554648 587052
rect 554596 586968 554648 586974
rect 554596 586910 554648 586916
rect 554608 530466 554636 586910
rect 554596 530460 554648 530466
rect 554596 530402 554648 530408
rect 554504 530120 554556 530126
rect 554504 530062 554556 530068
rect 554700 528850 554728 592447
rect 554778 591288 554834 591297
rect 554778 591223 554834 591232
rect 495052 528822 495388 528850
rect 496064 528822 496400 528850
rect 497168 528822 497504 528850
rect 498272 528822 498608 528850
rect 499284 528822 499528 528850
rect 500388 528822 500724 528850
rect 501492 528822 501828 528850
rect 502596 528822 502932 528850
rect 503608 528822 503668 528850
rect 504712 528822 505048 528850
rect 505816 528822 506152 528850
rect 506828 528822 507164 528850
rect 507932 528822 508268 528850
rect 509036 528822 509096 528850
rect 510140 528822 510476 528850
rect 511152 528822 511488 528850
rect 512256 528822 512592 528850
rect 513360 528822 513696 528850
rect 514372 528822 514708 528850
rect 515476 528822 515812 528850
rect 516580 528822 516916 528850
rect 517684 528822 518020 528850
rect 518696 528822 518756 528850
rect 519800 528822 520136 528850
rect 520904 528822 521240 528850
rect 521916 528822 522252 528850
rect 523020 528822 523356 528850
rect 524124 528822 524368 528850
rect 525228 528822 525564 528850
rect 526240 528822 526576 528850
rect 527344 528822 527680 528850
rect 528448 528822 528508 528850
rect 529460 528822 529796 528850
rect 530564 528822 530900 528850
rect 531668 528822 532004 528850
rect 532772 528822 533108 528850
rect 533784 528822 534028 528850
rect 534888 528822 535224 528850
rect 535992 528822 536328 528850
rect 537004 528822 537340 528850
rect 538108 528822 538168 528850
rect 539212 528822 539548 528850
rect 540316 528822 540652 528850
rect 541328 528822 541664 528850
rect 542432 528822 542768 528850
rect 543536 528822 543688 528850
rect 544548 528822 544884 528850
rect 545652 528822 545988 528850
rect 546756 528822 547092 528850
rect 547860 528822 548196 528850
rect 548872 528822 549208 528850
rect 549976 528822 550312 528850
rect 551080 528822 551416 528850
rect 552092 528822 552428 528850
rect 553196 528822 553348 528850
rect 554300 528822 554728 528850
rect 554792 528714 554820 591223
rect 556160 589348 556212 589354
rect 556160 589290 556212 589296
rect 554870 586392 554926 586401
rect 554870 586327 554872 586336
rect 554924 586327 554926 586336
rect 554872 586298 554924 586304
rect 554872 585200 554924 585206
rect 554870 585168 554872 585177
rect 554924 585168 554926 585177
rect 554870 585103 554926 585112
rect 554870 583808 554926 583817
rect 554870 583743 554872 583752
rect 554924 583743 554926 583752
rect 554872 583714 554924 583720
rect 555422 582720 555478 582729
rect 555422 582655 555478 582664
rect 554870 581088 554926 581097
rect 554870 581023 554872 581032
rect 554924 581023 554926 581032
rect 554872 580994 554924 581000
rect 554870 579728 554926 579737
rect 554870 579663 554872 579672
rect 554924 579663 554926 579672
rect 554872 579634 554924 579640
rect 554870 578504 554926 578513
rect 554870 578439 554926 578448
rect 554884 578270 554912 578439
rect 554872 578264 554924 578270
rect 554872 578206 554924 578212
rect 554870 577280 554926 577289
rect 554870 577215 554926 577224
rect 554884 576910 554912 577215
rect 554872 576904 554924 576910
rect 554872 576846 554924 576852
rect 555436 530670 555464 582655
rect 555424 530664 555476 530670
rect 555424 530606 555476 530612
rect 556172 528850 556200 589290
rect 557632 588804 557684 588810
rect 557632 588746 557684 588752
rect 556804 587104 556856 587110
rect 556804 587046 556856 587052
rect 556816 530058 556844 587046
rect 556804 530052 556856 530058
rect 556804 529994 556856 530000
rect 557644 528850 557672 588746
rect 558184 586356 558236 586362
rect 558184 586298 558236 586304
rect 558196 530330 558224 586298
rect 560300 585200 560352 585206
rect 560300 585142 560352 585148
rect 558276 571668 558328 571674
rect 558276 571610 558328 571616
rect 558288 530602 558316 571610
rect 558276 530596 558328 530602
rect 558276 530538 558328 530544
rect 558184 530324 558236 530330
rect 558184 530266 558236 530272
rect 559288 530324 559340 530330
rect 559288 530266 559340 530272
rect 558276 530052 558328 530058
rect 558276 529994 558328 530000
rect 556172 528822 556416 528850
rect 557520 528822 557672 528850
rect 558288 528850 558316 529994
rect 559300 528850 559328 530266
rect 560312 528850 560340 585142
rect 561772 583772 561824 583778
rect 561772 583714 561824 583720
rect 560944 575544 560996 575550
rect 560944 575486 560996 575492
rect 560956 529990 560984 575486
rect 560944 529984 560996 529990
rect 560944 529926 560996 529932
rect 561784 529122 561812 583714
rect 563060 581052 563112 581058
rect 563060 580994 563112 581000
rect 562600 530664 562652 530670
rect 562600 530606 562652 530612
rect 561784 529094 561858 529122
rect 558288 528822 558624 528850
rect 559300 528822 559636 528850
rect 560312 528822 560740 528850
rect 561830 528836 561858 529094
rect 562612 528850 562640 530606
rect 563072 529666 563100 580994
rect 564440 579692 564492 579698
rect 564440 579634 564492 579640
rect 563072 529638 563652 529666
rect 563624 528850 563652 529638
rect 564452 528986 564480 579634
rect 565820 578264 565872 578270
rect 565820 578206 565872 578212
rect 564452 528958 564756 528986
rect 564728 528850 564756 528958
rect 565832 528850 565860 578206
rect 567292 576904 567344 576910
rect 567292 576846 567344 576852
rect 567304 528850 567332 576846
rect 568580 574252 568632 574258
rect 568580 574194 568632 574200
rect 567936 529984 567988 529990
rect 567936 529926 567988 529932
rect 562612 528822 562948 528850
rect 563624 528822 563960 528850
rect 564728 528822 565064 528850
rect 565832 528822 566168 528850
rect 567180 528822 567332 528850
rect 567948 528850 567976 529926
rect 567948 528822 568284 528850
rect 568592 528714 568620 574194
rect 569960 574116 570012 574122
rect 569960 574058 570012 574064
rect 569972 528714 570000 574058
rect 571432 572756 571484 572762
rect 571432 572698 571484 572704
rect 571444 529122 571472 572698
rect 572720 569968 572772 569974
rect 572720 569910 572772 569916
rect 572260 530596 572312 530602
rect 572260 530538 572312 530544
rect 571444 529094 571518 529122
rect 571490 528836 571518 529094
rect 572272 528850 572300 530538
rect 572732 528986 572760 569910
rect 574376 533384 574428 533390
rect 574376 533326 574428 533332
rect 572732 528958 573220 528986
rect 572272 528822 572608 528850
rect 573192 528714 573220 528958
rect 574388 528850 574416 533326
rect 574388 528822 574724 528850
rect 479668 528708 479964 528714
rect 479616 528702 479964 528708
rect 479628 528686 479964 528702
rect 483032 528698 483184 528714
rect 483020 528692 483184 528698
rect 483072 528686 483184 528692
rect 493796 528686 493948 528714
rect 554792 528686 555404 528714
rect 568592 528686 569388 528714
rect 569972 528686 570492 528714
rect 573192 528686 573712 528714
rect 483020 528634 483072 528640
rect 486056 528624 486108 528630
rect 489274 528592 489330 528601
rect 486108 528572 486404 528578
rect 486056 528566 486404 528572
rect 486068 528550 486404 528566
rect 489330 528550 489624 528578
rect 489274 528527 489330 528536
rect 471702 528320 471758 528329
rect 410668 528300 410964 528306
rect 410616 528294 410964 528300
rect 410628 528278 410964 528294
rect 414952 528290 415288 528306
rect 414940 528284 415288 528290
rect 414992 528278 415288 528284
rect 471702 528255 471758 528264
rect 414940 528226 414992 528232
rect 423680 528216 423732 528222
rect 427820 528216 427872 528222
rect 423732 528164 423844 528170
rect 423680 528158 423844 528164
rect 432144 528216 432196 528222
rect 427872 528164 428168 528170
rect 427820 528158 428168 528164
rect 432196 528164 432492 528170
rect 432144 528158 432492 528164
rect 423692 528142 423844 528158
rect 427832 528142 428168 528158
rect 432156 528142 432492 528158
rect 317418 527232 317474 527241
rect 317418 527167 317474 527176
rect 317432 526969 317460 527167
rect 317418 526960 317474 526969
rect 317418 526895 317474 526904
rect 315946 515808 316002 515817
rect 315946 515743 316002 515752
rect 416596 503056 416648 503062
rect 324332 502982 324760 503010
rect 416148 503004 416596 503010
rect 416148 502998 416648 503004
rect 418160 503056 418212 503062
rect 418804 503056 418856 503062
rect 418212 503004 418804 503010
rect 418160 502998 418856 503004
rect 420276 503056 420328 503062
rect 420328 503004 420868 503010
rect 420276 502998 420868 503004
rect 413284 502988 413336 502994
rect 317892 502846 318228 502874
rect 318812 502846 319332 502874
rect 320192 502846 320436 502874
rect 321112 502846 321448 502874
rect 321572 502846 322552 502874
rect 323320 502846 323656 502874
rect 317892 499594 317920 502846
rect 318812 499610 318840 502846
rect 320192 499610 320220 502846
rect 317328 499588 317380 499594
rect 317328 499530 317380 499536
rect 317880 499588 317932 499594
rect 317880 499530 317932 499536
rect 318720 499582 318840 499610
rect 320100 499582 320220 499610
rect 317340 476610 317368 499530
rect 318720 477018 318748 499582
rect 320100 477018 320128 499582
rect 321112 495514 321140 502846
rect 320456 495508 320508 495514
rect 320456 495450 320508 495456
rect 321100 495508 321152 495514
rect 321100 495450 321152 495456
rect 320468 495394 320496 495450
rect 320284 495366 320496 495394
rect 320284 492658 320312 495366
rect 320272 492652 320324 492658
rect 320272 492594 320324 492600
rect 320732 492652 320784 492658
rect 320732 492594 320784 492600
rect 320744 483041 320772 492594
rect 320546 483032 320602 483041
rect 320546 482967 320602 482976
rect 320730 483032 320786 483041
rect 320730 482967 320786 482976
rect 317880 477012 317932 477018
rect 317880 476954 317932 476960
rect 318708 477012 318760 477018
rect 318708 476954 318760 476960
rect 319076 477012 319128 477018
rect 319076 476954 319128 476960
rect 320088 477012 320140 477018
rect 320088 476954 320140 476960
rect 316684 476604 316736 476610
rect 316684 476546 316736 476552
rect 317328 476604 317380 476610
rect 317328 476546 317380 476552
rect 316696 474164 316724 476546
rect 317892 474164 317920 476954
rect 319088 474164 319116 476954
rect 320560 474178 320588 482967
rect 320390 474150 320588 474178
rect 321572 474164 321600 502846
rect 323320 500410 323348 502846
rect 324332 500834 324360 502982
rect 413284 502930 413336 502936
rect 416148 502982 416636 502998
rect 418172 502982 418844 502998
rect 420288 502982 420868 502998
rect 325758 502602 325786 502860
rect 324240 500806 324360 500834
rect 325712 502574 325786 502602
rect 325896 502846 326876 502874
rect 327092 502846 327980 502874
rect 328472 502846 328992 502874
rect 329852 502846 330096 502874
rect 331200 502846 331352 502874
rect 322848 500404 322900 500410
rect 322848 500346 322900 500352
rect 323308 500404 323360 500410
rect 323308 500346 323360 500352
rect 322860 474178 322888 500346
rect 324240 474178 324268 500806
rect 325712 476218 325740 502574
rect 325620 476190 325740 476218
rect 325620 474178 325648 476190
rect 322782 474150 322888 474178
rect 323978 474150 324268 474178
rect 325266 474150 325648 474178
rect 325896 474042 325924 502846
rect 327092 474042 327120 502846
rect 328472 474042 328500 502846
rect 329852 474178 329880 502846
rect 329852 474150 330142 474178
rect 331324 474164 331352 502846
rect 331416 502846 332304 502874
rect 332612 502846 333316 502874
rect 333992 502846 334420 502874
rect 335372 502846 335524 502874
rect 336536 502846 336688 502874
rect 337640 502846 338068 502874
rect 338744 502846 339448 502874
rect 339848 502846 340184 502874
rect 340860 502846 341196 502874
rect 341964 502846 342208 502874
rect 343068 502846 343220 502874
rect 344080 502846 344416 502874
rect 345184 502846 345520 502874
rect 346288 502846 346348 502874
rect 347392 502846 347728 502874
rect 348404 502846 349108 502874
rect 349508 502846 349844 502874
rect 350612 502846 350948 502874
rect 351624 502846 351776 502874
rect 352728 502846 353248 502874
rect 353832 502846 354168 502874
rect 354936 502846 355272 502874
rect 331416 476474 331444 502846
rect 332612 476882 332640 502846
rect 332600 476876 332652 476882
rect 332600 476818 332652 476824
rect 333796 476876 333848 476882
rect 333796 476818 333848 476824
rect 331404 476468 331456 476474
rect 331404 476410 331456 476416
rect 332508 476468 332560 476474
rect 332508 476410 332560 476416
rect 332520 474164 332548 476410
rect 333808 474164 333836 476818
rect 333992 476610 334020 502846
rect 335372 476882 335400 502846
rect 336660 476882 336688 502846
rect 335360 476876 335412 476882
rect 335360 476818 335412 476824
rect 336188 476876 336240 476882
rect 336188 476818 336240 476824
rect 336648 476876 336700 476882
rect 336648 476818 336700 476824
rect 337476 476876 337528 476882
rect 337476 476818 337528 476824
rect 333980 476604 334032 476610
rect 333980 476546 334032 476552
rect 334992 476604 335044 476610
rect 334992 476546 335044 476552
rect 335004 474164 335032 476546
rect 336200 474164 336228 476818
rect 337488 474164 337516 476818
rect 338040 476218 338068 502846
rect 339420 476218 339448 502846
rect 340156 500954 340184 502846
rect 341168 500954 341196 502846
rect 340144 500948 340196 500954
rect 340144 500890 340196 500896
rect 340788 500948 340840 500954
rect 340788 500890 340840 500896
rect 341156 500948 341208 500954
rect 341156 500890 341208 500896
rect 342076 500948 342128 500954
rect 342076 500890 342128 500896
rect 340800 476218 340828 500890
rect 342088 476218 342116 500890
rect 342180 476882 342208 502846
rect 343192 500954 343220 502846
rect 343180 500948 343232 500954
rect 343180 500890 343232 500896
rect 343732 500948 343784 500954
rect 343732 500890 343784 500896
rect 343744 476898 343772 500890
rect 344388 499866 344416 502846
rect 345492 500954 345520 502846
rect 345480 500948 345532 500954
rect 345480 500890 345532 500896
rect 346216 500948 346268 500954
rect 346216 500890 346268 500896
rect 344376 499860 344428 499866
rect 344376 499802 344428 499808
rect 344928 499860 344980 499866
rect 344928 499802 344980 499808
rect 344940 477494 344968 499802
rect 344928 477488 344980 477494
rect 344928 477430 344980 477436
rect 346032 477488 346084 477494
rect 346032 477430 346084 477436
rect 342168 476876 342220 476882
rect 342168 476818 342220 476824
rect 343548 476876 343600 476882
rect 343744 476870 344324 476898
rect 343548 476818 343600 476824
rect 338040 476190 338344 476218
rect 339420 476190 339540 476218
rect 340800 476190 340920 476218
rect 342088 476190 342300 476218
rect 338316 474178 338344 476190
rect 339512 474178 339540 476190
rect 340892 474178 340920 476190
rect 342272 474178 342300 476190
rect 338316 474150 338698 474178
rect 339512 474150 339894 474178
rect 340892 474150 341090 474178
rect 342272 474150 342378 474178
rect 343560 474164 343588 476818
rect 344296 474042 344324 476870
rect 346044 474164 346072 477430
rect 346228 476882 346256 500890
rect 346216 476876 346268 476882
rect 346216 476818 346268 476824
rect 346320 476338 346348 502846
rect 347228 476876 347280 476882
rect 347228 476818 347280 476824
rect 346308 476332 346360 476338
rect 346308 476274 346360 476280
rect 347240 474164 347268 476818
rect 347700 476406 347728 502846
rect 349080 476610 349108 502846
rect 349816 500410 349844 502846
rect 350920 500682 350948 502846
rect 350908 500676 350960 500682
rect 350908 500618 350960 500624
rect 349804 500404 349856 500410
rect 349804 500346 349856 500352
rect 350448 500404 350500 500410
rect 350448 500346 350500 500352
rect 350460 476882 350488 500346
rect 350448 476876 350500 476882
rect 350448 476818 350500 476824
rect 351748 476814 351776 502846
rect 351828 500676 351880 500682
rect 351828 500618 351880 500624
rect 351840 476950 351868 500618
rect 353220 477494 353248 502846
rect 354140 500954 354168 502846
rect 354128 500948 354180 500954
rect 354128 500890 354180 500896
rect 354588 500948 354640 500954
rect 354588 500890 354640 500896
rect 353208 477488 353260 477494
rect 353208 477430 353260 477436
rect 354600 477426 354628 500890
rect 355244 500818 355272 502846
rect 355934 502602 355962 502860
rect 357052 502846 357388 502874
rect 358156 502846 358768 502874
rect 359168 502846 359504 502874
rect 360272 502846 360608 502874
rect 361376 502846 361436 502874
rect 362480 502846 362908 502874
rect 363492 502846 363828 502874
rect 364596 502846 364932 502874
rect 365700 502846 366036 502874
rect 366712 502846 366956 502874
rect 367816 502846 368428 502874
rect 368920 502846 369256 502874
rect 370024 502846 370360 502874
rect 371036 502846 371096 502874
rect 372140 502846 372568 502874
rect 373244 502846 373948 502874
rect 374256 502846 374592 502874
rect 375360 502846 375696 502874
rect 376464 502846 376708 502874
rect 377568 502846 378088 502874
rect 378580 502846 378916 502874
rect 379684 502846 380020 502874
rect 355888 502574 355962 502602
rect 355232 500812 355284 500818
rect 355232 500754 355284 500760
rect 355784 477488 355836 477494
rect 355784 477430 355836 477436
rect 354588 477420 354640 477426
rect 354588 477362 354640 477368
rect 351828 476944 351880 476950
rect 351828 476886 351880 476892
rect 353300 476944 353352 476950
rect 353300 476886 353352 476892
rect 352104 476876 352156 476882
rect 352104 476818 352156 476824
rect 351736 476808 351788 476814
rect 351736 476750 351788 476756
rect 349068 476604 349120 476610
rect 349068 476546 349120 476552
rect 350908 476604 350960 476610
rect 350908 476546 350960 476552
rect 347688 476400 347740 476406
rect 347688 476342 347740 476348
rect 349620 476400 349672 476406
rect 349620 476342 349672 476348
rect 348424 476332 348476 476338
rect 348424 476274 348476 476280
rect 348436 474164 348464 476274
rect 349632 474164 349660 476342
rect 350920 474164 350948 476546
rect 352116 474164 352144 476818
rect 353312 474164 353340 476886
rect 354588 476808 354640 476814
rect 354588 476750 354640 476756
rect 354600 474164 354628 476750
rect 355796 474164 355824 477430
rect 355888 476950 355916 502574
rect 355968 500812 356020 500818
rect 355968 500754 356020 500760
rect 355876 476944 355928 476950
rect 355876 476886 355928 476892
rect 355980 476882 356008 500754
rect 356980 477420 357032 477426
rect 356980 477362 357032 477368
rect 355968 476876 356020 476882
rect 355968 476818 356020 476824
rect 356992 474164 357020 477362
rect 357360 476610 357388 502846
rect 358740 476882 358768 502846
rect 359476 500954 359504 502846
rect 359464 500948 359516 500954
rect 359464 500890 359516 500896
rect 360108 500948 360160 500954
rect 360108 500890 360160 500896
rect 359464 476944 359516 476950
rect 359464 476886 359516 476892
rect 358176 476876 358228 476882
rect 358176 476818 358228 476824
rect 358728 476876 358780 476882
rect 358728 476818 358780 476824
rect 357348 476604 357400 476610
rect 357348 476546 357400 476552
rect 358188 474164 358216 476818
rect 359476 474164 359504 476886
rect 360120 476542 360148 500890
rect 360580 500002 360608 502846
rect 360568 499996 360620 500002
rect 360568 499938 360620 499944
rect 361408 476950 361436 502846
rect 361488 499996 361540 500002
rect 361488 499938 361540 499944
rect 361396 476944 361448 476950
rect 361396 476886 361448 476892
rect 361500 476746 361528 499938
rect 362880 477222 362908 502846
rect 363800 500546 363828 502846
rect 364904 500954 364932 502846
rect 366008 500954 366036 502846
rect 364892 500948 364944 500954
rect 364892 500890 364944 500896
rect 365628 500948 365680 500954
rect 365628 500890 365680 500896
rect 365996 500948 366048 500954
rect 365996 500890 366048 500896
rect 363788 500540 363840 500546
rect 363788 500482 363840 500488
rect 364248 500540 364300 500546
rect 364248 500482 364300 500488
rect 362868 477216 362920 477222
rect 362868 477158 362920 477164
rect 364260 477018 364288 500482
rect 364248 477012 364300 477018
rect 364248 476954 364300 476960
rect 365536 476944 365588 476950
rect 365536 476886 365588 476892
rect 361856 476876 361908 476882
rect 361856 476818 361908 476824
rect 361488 476740 361540 476746
rect 361488 476682 361540 476688
rect 360660 476604 360712 476610
rect 360660 476546 360712 476552
rect 360108 476536 360160 476542
rect 360108 476478 360160 476484
rect 360672 474164 360700 476546
rect 361868 474164 361896 476818
rect 364340 476740 364392 476746
rect 364340 476682 364392 476688
rect 363052 476536 363104 476542
rect 363052 476478 363104 476484
rect 363064 474164 363092 476478
rect 364352 474164 364380 476682
rect 365548 474164 365576 476886
rect 365640 476882 365668 500890
rect 366732 477216 366784 477222
rect 366732 477158 366784 477164
rect 365628 476876 365680 476882
rect 365628 476818 365680 476824
rect 366744 474164 366772 477158
rect 366928 476610 366956 502846
rect 367008 500948 367060 500954
rect 367008 500890 367060 500896
rect 367020 476678 367048 500890
rect 368020 477012 368072 477018
rect 368020 476954 368072 476960
rect 367008 476672 367060 476678
rect 367008 476614 367060 476620
rect 366916 476604 366968 476610
rect 366916 476546 366968 476552
rect 368032 474164 368060 476954
rect 368400 476746 368428 502846
rect 369228 500138 369256 502846
rect 370332 500954 370360 502846
rect 370320 500948 370372 500954
rect 370320 500890 370372 500896
rect 369216 500132 369268 500138
rect 369216 500074 369268 500080
rect 369768 500132 369820 500138
rect 369768 500074 369820 500080
rect 369780 477494 369808 500074
rect 369768 477488 369820 477494
rect 369768 477430 369820 477436
rect 369216 476876 369268 476882
rect 369216 476818 369268 476824
rect 368388 476740 368440 476746
rect 368388 476682 368440 476688
rect 369228 474164 369256 476818
rect 371068 476814 371096 502846
rect 371148 500948 371200 500954
rect 371148 500890 371200 500896
rect 371160 477018 371188 500890
rect 371148 477012 371200 477018
rect 371148 476954 371200 476960
rect 372540 476950 372568 502846
rect 372528 476944 372580 476950
rect 372528 476886 372580 476892
rect 373920 476882 373948 502846
rect 374564 500002 374592 502846
rect 375668 500954 375696 502846
rect 375656 500948 375708 500954
rect 375656 500890 375708 500896
rect 376576 500948 376628 500954
rect 376576 500890 376628 500896
rect 374552 499996 374604 500002
rect 374552 499938 374604 499944
rect 375288 499996 375340 500002
rect 375288 499938 375340 499944
rect 374092 477488 374144 477494
rect 374092 477430 374144 477436
rect 373908 476876 373960 476882
rect 373908 476818 373960 476824
rect 371056 476808 371108 476814
rect 371056 476750 371108 476756
rect 372896 476740 372948 476746
rect 372896 476682 372948 476688
rect 370412 476672 370464 476678
rect 370412 476614 370464 476620
rect 370424 474164 370452 476614
rect 371608 476604 371660 476610
rect 371608 476546 371660 476552
rect 371620 474164 371648 476546
rect 372908 474164 372936 476682
rect 374104 474164 374132 477430
rect 375300 477154 375328 499938
rect 375288 477148 375340 477154
rect 375288 477090 375340 477096
rect 376588 477018 376616 500890
rect 375288 477012 375340 477018
rect 375288 476954 375340 476960
rect 376576 477012 376628 477018
rect 376576 476954 376628 476960
rect 375300 474164 375328 476954
rect 376576 476808 376628 476814
rect 376576 476750 376628 476756
rect 376588 474164 376616 476750
rect 376680 476270 376708 502846
rect 378060 477426 378088 502846
rect 378888 500002 378916 502846
rect 379992 500138 380020 502846
rect 380774 502602 380802 502860
rect 381800 502846 382228 502874
rect 382904 502846 383608 502874
rect 384008 502846 384344 502874
rect 385112 502846 385448 502874
rect 386124 502846 386276 502874
rect 387228 502846 387748 502874
rect 388332 502846 388668 502874
rect 389344 502846 389680 502874
rect 380728 502574 380802 502602
rect 379980 500132 380032 500138
rect 379980 500074 380032 500080
rect 378876 499996 378928 500002
rect 378876 499938 378928 499944
rect 379428 499996 379480 500002
rect 379428 499938 379480 499944
rect 378048 477420 378100 477426
rect 378048 477362 378100 477368
rect 377772 476944 377824 476950
rect 377772 476886 377824 476892
rect 376668 476264 376720 476270
rect 376668 476206 376720 476212
rect 377784 474164 377812 476886
rect 378968 476876 379020 476882
rect 378968 476818 379020 476824
rect 378980 474164 379008 476818
rect 379440 476338 379468 499938
rect 380164 477148 380216 477154
rect 380164 477090 380216 477096
rect 379428 476332 379480 476338
rect 379428 476274 379480 476280
rect 380176 474164 380204 477090
rect 380728 476882 380756 502574
rect 380808 500132 380860 500138
rect 380808 500074 380860 500080
rect 380820 476950 380848 500074
rect 382200 477018 382228 502846
rect 383580 477222 383608 502846
rect 384316 500954 384344 502846
rect 385420 500954 385448 502846
rect 384304 500948 384356 500954
rect 384304 500890 384356 500896
rect 384948 500948 385000 500954
rect 384948 500890 385000 500896
rect 385408 500948 385460 500954
rect 385408 500890 385460 500896
rect 383844 477420 383896 477426
rect 383844 477362 383896 477368
rect 383568 477216 383620 477222
rect 383568 477158 383620 477164
rect 381452 477012 381504 477018
rect 381452 476954 381504 476960
rect 382188 477012 382240 477018
rect 382188 476954 382240 476960
rect 380808 476944 380860 476950
rect 380808 476886 380860 476892
rect 380716 476876 380768 476882
rect 380716 476818 380768 476824
rect 381464 474164 381492 476954
rect 382648 476264 382700 476270
rect 382648 476206 382700 476212
rect 382660 474164 382688 476206
rect 383856 474164 383884 477362
rect 384960 476270 384988 500890
rect 386248 476814 386276 502846
rect 386328 500948 386380 500954
rect 386328 500890 386380 500896
rect 386340 477086 386368 500890
rect 386328 477080 386380 477086
rect 386328 477022 386380 477028
rect 386328 476944 386380 476950
rect 386328 476886 386380 476892
rect 386236 476808 386288 476814
rect 386236 476750 386288 476756
rect 385132 476332 385184 476338
rect 385132 476274 385184 476280
rect 384948 476264 385000 476270
rect 384948 476206 385000 476212
rect 385144 474164 385172 476274
rect 386340 474164 386368 476886
rect 387524 476876 387576 476882
rect 387524 476818 387576 476824
rect 387536 474164 387564 476818
rect 387720 476474 387748 502846
rect 388640 499934 388668 502846
rect 389652 500002 389680 502846
rect 390434 502602 390462 502860
rect 391552 502846 391888 502874
rect 392656 502846 393268 502874
rect 393668 502846 394004 502874
rect 394772 502846 395108 502874
rect 395876 502846 395936 502874
rect 396888 502846 397408 502874
rect 397992 502846 398328 502874
rect 399096 502846 399432 502874
rect 400200 502846 400536 502874
rect 401212 502846 401548 502874
rect 403420 502846 403756 502874
rect 404432 502846 404768 502874
rect 409860 502846 409920 502874
rect 390388 502574 390462 502602
rect 389640 499996 389692 500002
rect 389640 499938 389692 499944
rect 388628 499928 388680 499934
rect 388628 499870 388680 499876
rect 389088 499928 389140 499934
rect 389088 499870 389140 499876
rect 389100 477018 389128 499870
rect 390008 477216 390060 477222
rect 390008 477158 390060 477164
rect 388720 477012 388772 477018
rect 388720 476954 388772 476960
rect 389088 477012 389140 477018
rect 389088 476954 389140 476960
rect 387708 476468 387760 476474
rect 387708 476410 387760 476416
rect 388732 474164 388760 476954
rect 390020 474164 390048 477158
rect 390388 476882 390416 502574
rect 390468 499996 390520 500002
rect 390468 499938 390520 499944
rect 390480 477358 390508 499938
rect 390468 477352 390520 477358
rect 390468 477294 390520 477300
rect 391860 477222 391888 502846
rect 391848 477216 391900 477222
rect 391848 477158 391900 477164
rect 393240 477086 393268 502846
rect 393976 500002 394004 502846
rect 395080 500954 395108 502846
rect 395068 500948 395120 500954
rect 395068 500890 395120 500896
rect 393964 499996 394016 500002
rect 393964 499938 394016 499944
rect 394608 499996 394660 500002
rect 394608 499938 394660 499944
rect 392400 477080 392452 477086
rect 392400 477022 392452 477028
rect 393228 477080 393280 477086
rect 393228 477022 393280 477028
rect 390376 476876 390428 476882
rect 390376 476818 390428 476824
rect 391204 476264 391256 476270
rect 391204 476206 391256 476212
rect 391216 474164 391244 476206
rect 392412 474164 392440 477022
rect 393688 476808 393740 476814
rect 393688 476750 393740 476756
rect 393700 474164 393728 476750
rect 394620 476746 394648 499938
rect 395908 476814 395936 502846
rect 395988 500948 396040 500954
rect 395988 500890 396040 500896
rect 396000 477290 396028 500890
rect 397276 477352 397328 477358
rect 397276 477294 397328 477300
rect 395988 477284 396040 477290
rect 395988 477226 396040 477232
rect 396080 477012 396132 477018
rect 396080 476954 396132 476960
rect 395896 476808 395948 476814
rect 395896 476750 395948 476756
rect 394608 476740 394660 476746
rect 394608 476682 394660 476688
rect 394884 476468 394936 476474
rect 394884 476410 394936 476416
rect 394896 474164 394924 476410
rect 396092 474164 396120 476954
rect 397288 474164 397316 477294
rect 397380 477018 397408 502846
rect 398300 500410 398328 502846
rect 398288 500404 398340 500410
rect 398288 500346 398340 500352
rect 398748 500404 398800 500410
rect 398748 500346 398800 500352
rect 397368 477012 397420 477018
rect 397368 476954 397420 476960
rect 398760 476950 398788 500346
rect 399404 500002 399432 502846
rect 400508 500954 400536 502846
rect 400496 500948 400548 500954
rect 400496 500890 400548 500896
rect 401416 500948 401468 500954
rect 401416 500890 401468 500896
rect 399392 499996 399444 500002
rect 399392 499938 399444 499944
rect 400128 499996 400180 500002
rect 400128 499938 400180 499944
rect 400140 477222 400168 499938
rect 399760 477216 399812 477222
rect 399760 477158 399812 477164
rect 400128 477216 400180 477222
rect 400128 477158 400180 477164
rect 398748 476944 398800 476950
rect 398748 476886 398800 476892
rect 398564 476876 398616 476882
rect 398564 476818 398616 476824
rect 398576 474164 398604 476818
rect 399772 474164 399800 477158
rect 401428 477086 401456 500890
rect 400956 477080 401008 477086
rect 400956 477022 401008 477028
rect 401416 477080 401468 477086
rect 401416 477022 401468 477028
rect 400968 474164 400996 477022
rect 401520 476882 401548 502846
rect 403728 500886 403756 502846
rect 404740 500954 404768 502846
rect 404728 500948 404780 500954
rect 404728 500890 404780 500896
rect 409892 500886 409920 502846
rect 411640 502846 411976 502874
rect 411640 500954 411668 502846
rect 411628 500948 411680 500954
rect 411628 500890 411680 500896
rect 403716 500880 403768 500886
rect 403716 500822 403768 500828
rect 409880 500880 409932 500886
rect 409880 500822 409932 500828
rect 403440 477284 403492 477290
rect 403440 477226 403492 477232
rect 401508 476876 401560 476882
rect 401508 476818 401560 476824
rect 402244 476740 402296 476746
rect 402244 476682 402296 476688
rect 402256 474164 402284 476682
rect 403452 474164 403480 477226
rect 408316 477216 408368 477222
rect 408316 477158 408368 477164
rect 405832 477012 405884 477018
rect 405832 476954 405884 476960
rect 404636 476808 404688 476814
rect 404636 476750 404688 476756
rect 404648 474164 404676 476750
rect 405844 474164 405872 476954
rect 407120 476944 407172 476950
rect 407120 476886 407172 476892
rect 407132 474164 407160 476886
rect 408328 474164 408356 477158
rect 409512 477080 409564 477086
rect 409512 477022 409564 477028
rect 409524 474164 409552 477022
rect 410708 476876 410760 476882
rect 410708 476818 410760 476824
rect 410720 474164 410748 476818
rect 325896 474014 326462 474042
rect 327092 474014 327658 474042
rect 328472 474014 328946 474042
rect 344296 474014 344770 474042
rect 338118 428768 338174 428777
rect 338118 428703 338174 428712
rect 336004 311908 336056 311914
rect 336004 311850 336056 311856
rect 315304 233912 315356 233918
rect 315304 233854 315356 233860
rect 313924 222896 313976 222902
rect 313924 222838 313976 222844
rect 336016 182170 336044 311850
rect 338132 198665 338160 428703
rect 338394 428632 338450 428641
rect 338394 428567 338450 428576
rect 338118 198656 338174 198665
rect 338118 198591 338174 198600
rect 336004 182164 336056 182170
rect 336004 182106 336056 182112
rect 230900 180820 231164 180826
rect 230848 180814 231164 180820
rect 230860 180798 231164 180814
rect 283392 173913 283420 175508
rect 283378 173904 283434 173913
rect 283378 173839 283434 173848
rect 283392 173233 283420 173839
rect 232226 173224 232282 173233
rect 232226 173159 232282 173168
rect 283378 173224 283434 173233
rect 283378 173159 283434 173168
rect 232240 167006 232268 173159
rect 232228 167000 232280 167006
rect 232228 166942 232280 166948
rect 232596 167000 232648 167006
rect 232596 166942 232648 166948
rect 232608 164218 232636 166942
rect 232320 164212 232372 164218
rect 232320 164154 232372 164160
rect 232596 164212 232648 164218
rect 232596 164154 232648 164160
rect 229744 161424 229796 161430
rect 229744 161366 229796 161372
rect 218796 160880 218848 160886
rect 218796 160822 218848 160828
rect 214930 157856 214986 157865
rect 214930 157791 214986 157800
rect 224684 155984 224736 155990
rect 224684 155926 224736 155932
rect 214930 154728 214986 154737
rect 214930 154663 214986 154672
rect 214748 148368 214800 148374
rect 214748 148310 214800 148316
rect 214760 143585 214788 148310
rect 214944 147626 214972 154663
rect 224592 153332 224644 153338
rect 224592 153274 224644 153280
rect 224500 151904 224552 151910
rect 224500 151846 224552 151852
rect 215944 151836 215996 151842
rect 215944 151778 215996 151784
rect 214932 147620 214984 147626
rect 214932 147562 214984 147568
rect 214746 143576 214802 143585
rect 214746 143511 214802 143520
rect 214746 109032 214802 109041
rect 214746 108967 214802 108976
rect 214576 104094 214696 104122
rect 214010 103864 214066 103873
rect 214010 103799 214066 103808
rect 116400 103556 116452 103562
rect 116400 103498 116452 103504
rect 214012 103488 214064 103494
rect 214012 103430 214064 103436
rect 213920 103420 213972 103426
rect 213920 103362 213972 103368
rect 116306 103184 116362 103193
rect 116306 103119 116362 103128
rect 116320 102202 116348 103119
rect 213932 103057 213960 103362
rect 213918 103048 213974 103057
rect 213918 102983 213974 102992
rect 214024 102241 214052 103430
rect 214010 102232 214066 102241
rect 116308 102196 116360 102202
rect 214010 102167 214066 102176
rect 116308 102138 116360 102144
rect 213920 102128 213972 102134
rect 116306 102096 116362 102105
rect 213920 102070 213972 102076
rect 116306 102031 116362 102040
rect 105544 100836 105596 100842
rect 105544 100778 105596 100784
rect 104164 100768 104216 100774
rect 104164 100710 104216 100716
rect 102784 91044 102836 91050
rect 102784 90986 102836 90992
rect 102876 89752 102928 89758
rect 102876 89694 102928 89700
rect 101404 86624 101456 86630
rect 101404 86566 101456 86572
rect 101496 85672 101548 85678
rect 101496 85614 101548 85620
rect 100024 81320 100076 81326
rect 100024 81262 100076 81268
rect 98736 80028 98788 80034
rect 98736 79970 98788 79976
rect 100024 78804 100076 78810
rect 100024 78746 100076 78752
rect 98644 68536 98696 68542
rect 98644 68478 98696 68484
rect 100036 66910 100064 78746
rect 101508 72962 101536 85614
rect 102888 75750 102916 89694
rect 104176 85542 104204 100710
rect 104164 85536 104216 85542
rect 104164 85478 104216 85484
rect 105556 84182 105584 100778
rect 116320 100774 116348 102031
rect 213932 101425 213960 102070
rect 213918 101416 213974 101425
rect 213918 101351 213974 101360
rect 116398 100872 116454 100881
rect 116398 100807 116400 100816
rect 116452 100807 116454 100816
rect 116400 100778 116452 100784
rect 116308 100768 116360 100774
rect 116308 100710 116360 100716
rect 213920 100700 213972 100706
rect 213920 100642 213972 100648
rect 213932 100609 213960 100642
rect 214012 100632 214064 100638
rect 213918 100600 213974 100609
rect 214012 100574 214064 100580
rect 213918 100535 213974 100544
rect 214024 99929 214052 100574
rect 214010 99920 214066 99929
rect 214010 99855 214066 99864
rect 116398 99784 116454 99793
rect 116398 99719 116454 99728
rect 116412 99414 116440 99719
rect 116400 99408 116452 99414
rect 116400 99350 116452 99356
rect 116398 98560 116454 98569
rect 116398 98495 116454 98504
rect 116412 98054 116440 98495
rect 116400 98048 116452 98054
rect 116400 97990 116452 97996
rect 214104 97980 214156 97986
rect 214104 97922 214156 97928
rect 213920 97640 213972 97646
rect 213920 97582 213972 97588
rect 116398 97336 116454 97345
rect 116398 97271 116454 97280
rect 116412 96694 116440 97271
rect 213932 96801 213960 97582
rect 214116 97481 214144 97922
rect 214102 97472 214158 97481
rect 214102 97407 214158 97416
rect 213918 96792 213974 96801
rect 213918 96727 213974 96736
rect 116400 96688 116452 96694
rect 116400 96630 116452 96636
rect 116306 96248 116362 96257
rect 116306 96183 116362 96192
rect 116320 95266 116348 96183
rect 214576 95985 214604 104094
rect 214656 99340 214708 99346
rect 214656 99282 214708 99288
rect 214668 98297 214696 99282
rect 214654 98288 214710 98297
rect 214654 98223 214710 98232
rect 214562 95976 214618 95985
rect 214562 95911 214618 95920
rect 116308 95260 116360 95266
rect 116308 95202 116360 95208
rect 214760 95169 214788 108967
rect 215116 99272 215168 99278
rect 215116 99214 215168 99220
rect 215128 99113 215156 99214
rect 215114 99104 215170 99113
rect 215114 99039 215170 99048
rect 215956 97646 215984 151778
rect 216680 150884 216732 150890
rect 216680 150826 216732 150832
rect 216692 146266 216720 150826
rect 224224 150476 224276 150482
rect 224224 150418 224276 150424
rect 216772 149388 216824 149394
rect 216772 149330 216824 149336
rect 216680 146260 216732 146266
rect 216680 146202 216732 146208
rect 216784 144906 216812 149330
rect 224132 149116 224184 149122
rect 224132 149058 224184 149064
rect 216864 148028 216916 148034
rect 216864 147970 216916 147976
rect 216772 144900 216824 144906
rect 216772 144842 216824 144848
rect 216772 143676 216824 143682
rect 216772 143618 216824 143624
rect 216680 142248 216732 142254
rect 216680 142190 216732 142196
rect 216692 137970 216720 142190
rect 216784 139398 216812 143618
rect 216876 143546 216904 147970
rect 217600 146396 217652 146402
rect 217600 146338 217652 146344
rect 217324 145036 217376 145042
rect 217324 144978 217376 144984
rect 216864 143540 216916 143546
rect 216864 143482 216916 143488
rect 217336 140758 217364 144978
rect 217612 142118 217640 146338
rect 224144 143478 224172 149058
rect 224236 144838 224264 150418
rect 224512 146198 224540 151846
rect 224604 147490 224632 153274
rect 224696 150414 224724 155926
rect 224776 154624 224828 154630
rect 232332 154601 232360 164154
rect 224776 154566 224828 154572
rect 232318 154592 232374 154601
rect 224684 150408 224736 150414
rect 224684 150350 224736 150356
rect 224788 148986 224816 154566
rect 232318 154527 232374 154536
rect 232502 154592 232558 154601
rect 232502 154527 232558 154536
rect 224868 153264 224920 153270
rect 224868 153206 224920 153212
rect 224776 148980 224828 148986
rect 224776 148922 224828 148928
rect 224880 147558 224908 153206
rect 227444 150408 227496 150414
rect 227444 150350 227496 150356
rect 227456 149433 227484 150350
rect 232516 149734 232544 154527
rect 286140 151836 286192 151842
rect 286140 151778 286192 151784
rect 232136 149728 232188 149734
rect 232136 149670 232188 149676
rect 232504 149728 232556 149734
rect 232504 149670 232556 149676
rect 227442 149424 227498 149433
rect 227442 149359 227498 149368
rect 227444 149048 227496 149054
rect 227444 148990 227496 148996
rect 227456 148889 227484 148990
rect 227536 148980 227588 148986
rect 227536 148922 227588 148928
rect 227442 148880 227498 148889
rect 227442 148815 227498 148824
rect 227548 148209 227576 148922
rect 227534 148200 227590 148209
rect 227534 148135 227590 148144
rect 227442 147656 227498 147665
rect 227442 147591 227444 147600
rect 227496 147591 227498 147600
rect 227444 147562 227496 147568
rect 224868 147552 224920 147558
rect 224868 147494 224920 147500
rect 226984 147552 227036 147558
rect 226984 147494 227036 147500
rect 224592 147484 224644 147490
rect 224592 147426 224644 147432
rect 226996 146985 227024 147494
rect 227536 147484 227588 147490
rect 227536 147426 227588 147432
rect 226982 146976 227038 146985
rect 226982 146911 227038 146920
rect 227548 146441 227576 147426
rect 227534 146432 227590 146441
rect 227534 146367 227590 146376
rect 227628 146328 227680 146334
rect 227628 146270 227680 146276
rect 226708 146260 226760 146266
rect 226708 146202 226760 146208
rect 224500 146192 224552 146198
rect 224500 146134 224552 146140
rect 226720 145217 226748 146202
rect 227444 146192 227496 146198
rect 227444 146134 227496 146140
rect 227456 145897 227484 146134
rect 227442 145888 227498 145897
rect 227442 145823 227498 145832
rect 226706 145208 226762 145217
rect 226706 145143 226762 145152
rect 227260 144968 227312 144974
rect 227260 144910 227312 144916
rect 226524 144900 226576 144906
rect 226524 144842 226576 144848
rect 224224 144832 224276 144838
rect 224224 144774 224276 144780
rect 226536 143993 226564 144842
rect 226522 143984 226578 143993
rect 226522 143919 226578 143928
rect 226892 143540 226944 143546
rect 226892 143482 226944 143488
rect 224132 143472 224184 143478
rect 224132 143414 224184 143420
rect 226904 142905 226932 143482
rect 226890 142896 226946 142905
rect 226890 142831 226946 142840
rect 217600 142112 217652 142118
rect 217600 142054 217652 142060
rect 226708 142112 226760 142118
rect 226708 142054 226760 142060
rect 226720 141681 226748 142054
rect 226706 141672 226762 141681
rect 226706 141607 226762 141616
rect 227272 141001 227300 144910
rect 227444 144832 227496 144838
rect 227444 144774 227496 144780
rect 227456 144673 227484 144774
rect 227442 144664 227498 144673
rect 227442 144599 227498 144608
rect 227536 143608 227588 143614
rect 227536 143550 227588 143556
rect 227444 143472 227496 143478
rect 227442 143440 227444 143449
rect 227496 143440 227498 143449
rect 227442 143375 227498 143384
rect 227352 142180 227404 142186
rect 227352 142122 227404 142128
rect 227258 140992 227314 141001
rect 227258 140927 227314 140936
rect 226708 140820 226760 140826
rect 226708 140762 226760 140768
rect 217324 140752 217376 140758
rect 217324 140694 217376 140700
rect 226616 139528 226668 139534
rect 226616 139470 226668 139476
rect 226524 139460 226576 139466
rect 226524 139402 226576 139408
rect 216772 139392 216824 139398
rect 216772 139334 216824 139340
rect 226432 138100 226484 138106
rect 226432 138042 226484 138048
rect 216680 137964 216732 137970
rect 216680 137906 216732 137912
rect 226444 135697 226472 138042
rect 226536 136785 226564 139402
rect 226522 136776 226578 136785
rect 226522 136711 226578 136720
rect 226628 136241 226656 139470
rect 226720 137465 226748 140762
rect 227076 140752 227128 140758
rect 227076 140694 227128 140700
rect 227088 140457 227116 140694
rect 227074 140448 227130 140457
rect 227074 140383 227130 140392
rect 227364 138689 227392 142122
rect 227548 139777 227576 143550
rect 227640 142225 227668 146270
rect 227626 142216 227682 142225
rect 227626 142151 227682 142160
rect 227534 139768 227590 139777
rect 227534 139703 227590 139712
rect 227444 139392 227496 139398
rect 227444 139334 227496 139340
rect 227456 139233 227484 139334
rect 227442 139224 227498 139233
rect 227442 139159 227498 139168
rect 227350 138680 227406 138689
rect 227350 138615 227406 138624
rect 226800 138032 226852 138038
rect 226800 137974 226852 137980
rect 227442 138000 227498 138009
rect 226706 137456 226762 137465
rect 226706 137391 226762 137400
rect 226614 136232 226670 136241
rect 226614 136167 226670 136176
rect 226430 135688 226486 135697
rect 226430 135623 226486 135632
rect 226812 135017 226840 137974
rect 227442 137935 227444 137944
rect 227496 137935 227498 137944
rect 227444 137906 227496 137912
rect 227076 136740 227128 136746
rect 227076 136682 227128 136688
rect 226798 135008 226854 135017
rect 226798 134943 226854 134952
rect 227088 133793 227116 136682
rect 227444 136672 227496 136678
rect 227444 136614 227496 136620
rect 227456 134473 227484 136614
rect 227628 135312 227680 135318
rect 227628 135254 227680 135260
rect 227442 134464 227498 134473
rect 227442 134399 227498 134408
rect 227536 134020 227588 134026
rect 227536 133962 227588 133968
rect 227352 133952 227404 133958
rect 227352 133894 227404 133900
rect 227074 133784 227130 133793
rect 227074 133719 227130 133728
rect 226708 132592 226760 132598
rect 226708 132534 226760 132540
rect 226524 131232 226576 131238
rect 226524 131174 226576 131180
rect 226536 129577 226564 131174
rect 226720 130801 226748 132534
rect 227364 132025 227392 133894
rect 227548 132569 227576 133962
rect 227640 133249 227668 135254
rect 227626 133240 227682 133249
rect 227626 133175 227682 133184
rect 227534 132560 227590 132569
rect 227444 132524 227496 132530
rect 227534 132495 227590 132504
rect 227444 132466 227496 132472
rect 227350 132016 227406 132025
rect 227350 131951 227406 131960
rect 227456 131481 227484 132466
rect 227442 131472 227498 131481
rect 227442 131407 227498 131416
rect 227076 131164 227128 131170
rect 227076 131106 227128 131112
rect 226706 130792 226762 130801
rect 226706 130727 226762 130736
rect 227088 130257 227116 131106
rect 227074 130248 227130 130257
rect 227074 130183 227130 130192
rect 227536 129804 227588 129810
rect 227536 129746 227588 129752
rect 226522 129568 226578 129577
rect 226522 129503 226578 129512
rect 227444 129056 227496 129062
rect 227548 129033 227576 129746
rect 227444 128998 227496 129004
rect 227534 129024 227590 129033
rect 227456 128489 227484 128998
rect 227534 128959 227590 128968
rect 232148 128602 232176 149670
rect 286152 149668 286180 151778
rect 232056 128574 232176 128602
rect 227442 128480 227498 128489
rect 227442 128415 227498 128424
rect 226340 128376 226392 128382
rect 226340 128318 226392 128324
rect 226352 127809 226380 128318
rect 226338 127800 226394 127809
rect 226338 127735 226394 127744
rect 227444 127628 227496 127634
rect 227444 127570 227496 127576
rect 227456 127265 227484 127570
rect 227442 127256 227498 127265
rect 227442 127191 227498 127200
rect 227444 127016 227496 127022
rect 227444 126958 227496 126964
rect 227456 126585 227484 126958
rect 227442 126576 227498 126585
rect 227442 126511 227498 126520
rect 227444 126268 227496 126274
rect 227444 126210 227496 126216
rect 227456 126041 227484 126210
rect 227442 126032 227498 126041
rect 227442 125967 227498 125976
rect 227444 125656 227496 125662
rect 227444 125598 227496 125604
rect 227456 125361 227484 125598
rect 227442 125352 227498 125361
rect 227442 125287 227498 125296
rect 227260 124908 227312 124914
rect 227260 124850 227312 124856
rect 227272 124817 227300 124850
rect 227258 124808 227314 124817
rect 227258 124743 227314 124752
rect 227258 124264 227314 124273
rect 227258 124199 227314 124208
rect 227272 124166 227300 124199
rect 227260 124160 227312 124166
rect 227260 124102 227312 124108
rect 227258 123584 227314 123593
rect 227258 123519 227314 123528
rect 227272 123486 227300 123519
rect 227260 123480 227312 123486
rect 227260 123422 227312 123428
rect 227442 123040 227498 123049
rect 227442 122975 227498 122984
rect 227456 122806 227484 122975
rect 227444 122800 227496 122806
rect 227444 122742 227496 122748
rect 227442 122360 227498 122369
rect 227442 122295 227498 122304
rect 227456 122126 227484 122295
rect 227444 122120 227496 122126
rect 227444 122062 227496 122068
rect 227442 121816 227498 121825
rect 227442 121751 227498 121760
rect 227456 121446 227484 121751
rect 227444 121440 227496 121446
rect 227444 121382 227496 121388
rect 227442 121272 227498 121281
rect 227442 121207 227498 121216
rect 227456 120766 227484 121207
rect 227444 120760 227496 120766
rect 227444 120702 227496 120708
rect 227442 120592 227498 120601
rect 227442 120527 227498 120536
rect 227456 120086 227484 120527
rect 227444 120080 227496 120086
rect 226430 120048 226486 120057
rect 227444 120022 227496 120028
rect 226430 119983 226486 119992
rect 226338 119368 226394 119377
rect 226338 119303 226394 119312
rect 226246 118824 226302 118833
rect 226246 118759 226302 118768
rect 226154 117600 226210 117609
rect 226154 117535 226210 117544
rect 226168 115870 226196 117535
rect 226260 117230 226288 118759
rect 226352 118590 226380 119303
rect 226444 118658 226472 119983
rect 226432 118652 226484 118658
rect 226432 118594 226484 118600
rect 226340 118584 226392 118590
rect 226340 118526 226392 118532
rect 227442 118144 227498 118153
rect 227442 118079 227498 118088
rect 227456 117298 227484 118079
rect 227444 117292 227496 117298
rect 227444 117234 227496 117240
rect 226248 117224 226300 117230
rect 226248 117166 226300 117172
rect 227442 117056 227498 117065
rect 227442 116991 227498 117000
rect 226246 116376 226302 116385
rect 226246 116311 226302 116320
rect 226156 115864 226208 115870
rect 226156 115806 226208 115812
rect 226154 115152 226210 115161
rect 226154 115087 226210 115096
rect 226062 114608 226118 114617
rect 226062 114543 226118 114552
rect 225970 113384 226026 113393
rect 225970 113319 226026 113328
rect 225878 112160 225934 112169
rect 225878 112095 225934 112104
rect 225786 110392 225842 110401
rect 225786 110327 225842 110336
rect 225602 109168 225658 109177
rect 225602 109103 225658 109112
rect 224776 104916 224828 104922
rect 224776 104858 224828 104864
rect 224788 99278 224816 104858
rect 225616 104786 225644 109103
rect 225694 107944 225750 107953
rect 225694 107879 225750 107888
rect 225604 104780 225656 104786
rect 225604 104722 225656 104728
rect 224868 103692 224920 103698
rect 224868 103634 224920 103640
rect 224776 99272 224828 99278
rect 224776 99214 224828 99220
rect 224880 97986 224908 103634
rect 225708 103426 225736 107879
rect 225800 106282 225828 110327
rect 225892 108934 225920 112095
rect 225984 110362 226012 113319
rect 226076 111722 226104 114543
rect 226168 113150 226196 115087
rect 226260 114442 226288 116311
rect 227456 115938 227484 116991
rect 227444 115932 227496 115938
rect 227444 115874 227496 115880
rect 227074 115832 227130 115841
rect 232056 115818 232084 128574
rect 232056 115790 232176 115818
rect 227074 115767 227130 115776
rect 227088 114510 227116 115767
rect 227076 114504 227128 114510
rect 227076 114446 227128 114452
rect 226248 114436 226300 114442
rect 226248 114378 226300 114384
rect 226246 114064 226302 114073
rect 226246 113999 226302 114008
rect 226156 113144 226208 113150
rect 226156 113086 226208 113092
rect 226154 112840 226210 112849
rect 226154 112775 226210 112784
rect 226064 111716 226116 111722
rect 226064 111658 226116 111664
rect 226062 110936 226118 110945
rect 226062 110871 226118 110880
rect 225972 110356 226024 110362
rect 225972 110298 226024 110304
rect 225880 108928 225932 108934
rect 225880 108870 225932 108876
rect 226076 107642 226104 110871
rect 226168 110430 226196 112775
rect 226260 111790 226288 113999
rect 226248 111784 226300 111790
rect 226248 111726 226300 111732
rect 226246 111616 226302 111625
rect 226246 111551 226302 111560
rect 226156 110424 226208 110430
rect 226156 110366 226208 110372
rect 226260 109002 226288 111551
rect 226338 109848 226394 109857
rect 226338 109783 226394 109792
rect 226248 108996 226300 109002
rect 226248 108938 226300 108944
rect 226352 108882 226380 109783
rect 226260 108854 226380 108882
rect 226154 108624 226210 108633
rect 226154 108559 226210 108568
rect 226064 107636 226116 107642
rect 226064 107578 226116 107584
rect 225970 107400 226026 107409
rect 225970 107335 226026 107344
rect 225878 106856 225934 106865
rect 225878 106791 225934 106800
rect 225788 106276 225840 106282
rect 225788 106218 225840 106224
rect 225696 103420 225748 103426
rect 225696 103362 225748 103368
rect 225892 102134 225920 106791
rect 225984 103494 226012 107335
rect 226062 105632 226118 105641
rect 226062 105567 226118 105576
rect 225972 103488 226024 103494
rect 225972 103430 226024 103436
rect 225880 102128 225932 102134
rect 225880 102070 225932 102076
rect 226076 100638 226104 105567
rect 226168 104854 226196 108559
rect 226260 106214 226288 108854
rect 226248 106208 226300 106214
rect 226248 106150 226300 106156
rect 226246 105768 226302 105777
rect 226246 105703 226302 105712
rect 226156 104848 226208 104854
rect 226156 104790 226208 104796
rect 226260 104530 226288 105703
rect 227442 104952 227498 104961
rect 227442 104887 227444 104896
rect 227496 104887 227498 104896
rect 227444 104858 227496 104864
rect 226168 104502 226288 104530
rect 226168 100706 226196 104502
rect 226246 104408 226302 104417
rect 226246 104343 226302 104352
rect 226156 100700 226208 100706
rect 226156 100642 226208 100648
rect 226064 100632 226116 100638
rect 226064 100574 226116 100580
rect 226260 99346 226288 104343
rect 227442 103864 227498 103873
rect 227442 103799 227498 103808
rect 227456 103698 227484 103799
rect 227444 103692 227496 103698
rect 227444 103634 227496 103640
rect 232148 100706 232176 115790
rect 258092 100706 258120 103564
rect 314212 102134 314240 103564
rect 338408 102134 338436 428567
rect 343638 428496 343694 428505
rect 343638 428431 343694 428440
rect 341524 310548 341576 310554
rect 341524 310490 341576 310496
rect 340144 309188 340196 309194
rect 340144 309130 340196 309136
rect 314200 102128 314252 102134
rect 314200 102070 314252 102076
rect 338396 102128 338448 102134
rect 338396 102070 338448 102076
rect 232136 100700 232188 100706
rect 232136 100642 232188 100648
rect 258080 100700 258132 100706
rect 258080 100642 258132 100648
rect 232148 99346 232176 100642
rect 226248 99340 226300 99346
rect 226248 99282 226300 99288
rect 232136 99340 232188 99346
rect 232136 99282 232188 99288
rect 232504 99340 232556 99346
rect 232504 99282 232556 99288
rect 224868 97980 224920 97986
rect 224868 97922 224920 97928
rect 215944 97640 215996 97646
rect 215944 97582 215996 97588
rect 215116 95192 215168 95198
rect 214746 95160 214802 95169
rect 215116 95134 215168 95140
rect 214746 95095 214802 95104
rect 116490 95024 116546 95033
rect 116490 94959 116546 94968
rect 116398 93936 116454 93945
rect 116398 93871 116400 93880
rect 116452 93871 116454 93880
rect 116400 93842 116452 93848
rect 116398 92712 116454 92721
rect 116398 92647 116454 92656
rect 116412 92546 116440 92647
rect 116400 92540 116452 92546
rect 116400 92482 116452 92488
rect 116398 91624 116454 91633
rect 116398 91559 116454 91568
rect 116412 91118 116440 91559
rect 116400 91112 116452 91118
rect 116400 91054 116452 91060
rect 116398 90400 116454 90409
rect 116504 90370 116532 94959
rect 215128 94353 215156 95134
rect 215114 94344 215170 94353
rect 215114 94279 215170 94288
rect 215208 93832 215260 93838
rect 215208 93774 215260 93780
rect 215116 93764 215168 93770
rect 215116 93706 215168 93712
rect 215128 93673 215156 93706
rect 215114 93664 215170 93673
rect 215114 93599 215170 93608
rect 215220 92857 215248 93774
rect 215206 92848 215262 92857
rect 215206 92783 215262 92792
rect 214838 92032 214894 92041
rect 214838 91967 214894 91976
rect 214562 90536 214618 90545
rect 214562 90471 214618 90480
rect 116398 90335 116454 90344
rect 116492 90364 116544 90370
rect 116412 89758 116440 90335
rect 116492 90306 116544 90312
rect 116400 89752 116452 89758
rect 116400 89694 116452 89700
rect 214286 89720 214342 89729
rect 214286 89655 214342 89664
rect 115938 89176 115994 89185
rect 115938 89111 115994 89120
rect 115952 88398 115980 89111
rect 115940 88392 115992 88398
rect 115940 88334 115992 88340
rect 116398 88088 116454 88097
rect 116398 88023 116454 88032
rect 214194 88088 214250 88097
rect 214194 88023 214250 88032
rect 116412 87038 116440 88023
rect 116400 87032 116452 87038
rect 116400 86974 116452 86980
rect 116306 86864 116362 86873
rect 116306 86799 116362 86808
rect 116320 85610 116348 86799
rect 116398 85776 116454 85785
rect 116398 85711 116454 85720
rect 116412 85678 116440 85711
rect 116400 85672 116452 85678
rect 116400 85614 116452 85620
rect 116308 85604 116360 85610
rect 116308 85546 116360 85552
rect 116398 84552 116454 84561
rect 116398 84487 116454 84496
rect 116412 84250 116440 84487
rect 116400 84244 116452 84250
rect 116400 84186 116452 84192
rect 105544 84176 105596 84182
rect 105544 84118 105596 84124
rect 214208 83722 214236 88023
rect 213932 83694 214236 83722
rect 116398 83328 116454 83337
rect 116398 83263 116454 83272
rect 116412 82890 116440 83263
rect 116400 82884 116452 82890
rect 116400 82826 116452 82832
rect 115938 82240 115994 82249
rect 115938 82175 115994 82184
rect 115952 81462 115980 82175
rect 115940 81456 115992 81462
rect 115940 81398 115992 81404
rect 116398 81016 116454 81025
rect 116398 80951 116454 80960
rect 116412 80102 116440 80951
rect 116400 80096 116452 80102
rect 116400 80038 116452 80044
rect 116214 79928 116270 79937
rect 116214 79863 116270 79872
rect 116228 78742 116256 79863
rect 213932 79642 213960 83694
rect 214012 83564 214064 83570
rect 214012 83506 214064 83512
rect 214024 80050 214052 83506
rect 214194 82648 214250 82657
rect 214194 82583 214250 82592
rect 214208 81462 214236 82583
rect 214196 81456 214248 81462
rect 214196 81398 214248 81404
rect 214024 80022 214236 80050
rect 214300 80034 214328 89655
rect 214470 86592 214526 86601
rect 214470 86527 214526 86536
rect 214378 84960 214434 84969
rect 214378 84895 214434 84904
rect 214392 83570 214420 84895
rect 214380 83564 214432 83570
rect 214380 83506 214432 83512
rect 214378 83464 214434 83473
rect 214378 83399 214434 83408
rect 213932 79614 214052 79642
rect 213918 79520 213974 79529
rect 213918 79455 213974 79464
rect 213932 78810 213960 79455
rect 116400 78804 116452 78810
rect 116400 78746 116452 78752
rect 213920 78804 213972 78810
rect 213920 78746 213972 78752
rect 116216 78736 116268 78742
rect 116412 78713 116440 78746
rect 116216 78678 116268 78684
rect 116398 78704 116454 78713
rect 214024 78674 214052 79614
rect 116398 78639 116454 78648
rect 214012 78668 214064 78674
rect 214012 78610 214064 78616
rect 213918 77888 213974 77897
rect 213918 77823 213974 77832
rect 116398 77480 116454 77489
rect 116398 77415 116454 77424
rect 116412 77314 116440 77415
rect 213932 77314 213960 77823
rect 116400 77308 116452 77314
rect 116400 77250 116452 77256
rect 213920 77308 213972 77314
rect 213920 77250 213972 77256
rect 116398 76392 116454 76401
rect 116398 76327 116454 76336
rect 213918 76392 213974 76401
rect 213918 76327 213974 76336
rect 116412 75954 116440 76327
rect 213932 76090 213960 76327
rect 213920 76084 213972 76090
rect 213920 76026 213972 76032
rect 116400 75948 116452 75954
rect 116400 75890 116452 75896
rect 214208 75750 214236 80022
rect 214288 80028 214340 80034
rect 214288 79970 214340 79976
rect 102876 75744 102928 75750
rect 102876 75686 102928 75692
rect 214196 75744 214248 75750
rect 214196 75686 214248 75692
rect 116398 75168 116454 75177
rect 116398 75103 116454 75112
rect 116412 74594 116440 75103
rect 213918 74760 213974 74769
rect 213918 74695 213974 74704
rect 213932 74662 213960 74695
rect 213920 74656 213972 74662
rect 213920 74598 213972 74604
rect 116400 74588 116452 74594
rect 116400 74530 116452 74536
rect 214392 74458 214420 83399
rect 214484 77178 214512 86527
rect 214576 79966 214604 90471
rect 214746 88904 214802 88913
rect 214746 88839 214802 88848
rect 214654 87408 214710 87417
rect 214654 87343 214710 87352
rect 214564 79960 214616 79966
rect 214564 79902 214616 79908
rect 214668 77246 214696 87343
rect 214760 78606 214788 88839
rect 214852 81326 214880 91967
rect 215022 91216 215078 91225
rect 215022 91151 215078 91160
rect 215036 81394 215064 91151
rect 232516 89706 232544 99282
rect 232424 89678 232544 89706
rect 215114 85776 215170 85785
rect 215114 85711 215170 85720
rect 215128 85610 215156 85711
rect 215116 85604 215168 85610
rect 215116 85546 215168 85552
rect 224224 85604 224276 85610
rect 224224 85546 224276 85552
rect 215114 84280 215170 84289
rect 215114 84215 215116 84224
rect 215168 84215 215170 84224
rect 215116 84186 215168 84192
rect 215944 82884 215996 82890
rect 215944 82826 215996 82832
rect 215206 81832 215262 81841
rect 215206 81767 215262 81776
rect 215024 81388 215076 81394
rect 215024 81330 215076 81336
rect 214840 81320 214892 81326
rect 214840 81262 214892 81268
rect 215114 81016 215170 81025
rect 215114 80951 215170 80960
rect 214930 80336 214986 80345
rect 214930 80271 214986 80280
rect 214838 78704 214894 78713
rect 214838 78639 214894 78648
rect 214748 78600 214800 78606
rect 214748 78542 214800 78548
rect 214656 77240 214708 77246
rect 214656 77182 214708 77188
rect 214472 77172 214524 77178
rect 214472 77114 214524 77120
rect 214746 75576 214802 75585
rect 214746 75511 214802 75520
rect 214380 74452 214432 74458
rect 214380 74394 214432 74400
rect 116398 74080 116454 74089
rect 116398 74015 116454 74024
rect 214102 74080 214158 74089
rect 214102 74015 214158 74024
rect 116412 73234 116440 74015
rect 213918 73264 213974 73273
rect 116400 73228 116452 73234
rect 213918 73199 213920 73208
rect 116400 73170 116452 73176
rect 213972 73199 213974 73208
rect 213920 73170 213972 73176
rect 101496 72956 101548 72962
rect 101496 72898 101548 72904
rect 116398 72856 116454 72865
rect 116398 72791 116454 72800
rect 116412 71806 116440 72791
rect 116400 71800 116452 71806
rect 116400 71742 116452 71748
rect 116582 71768 116638 71777
rect 116582 71703 116638 71712
rect 116398 70544 116454 70553
rect 116398 70479 116454 70488
rect 116412 70446 116440 70479
rect 116400 70440 116452 70446
rect 116400 70382 116452 70388
rect 116398 69320 116454 69329
rect 116398 69255 116454 69264
rect 116412 69086 116440 69255
rect 116400 69080 116452 69086
rect 116400 69022 116452 69028
rect 116398 68232 116454 68241
rect 116398 68167 116454 68176
rect 116412 67658 116440 68167
rect 116400 67652 116452 67658
rect 116400 67594 116452 67600
rect 116398 67008 116454 67017
rect 116398 66943 116454 66952
rect 100024 66904 100076 66910
rect 100024 66846 100076 66852
rect 116412 66298 116440 66943
rect 116400 66292 116452 66298
rect 116400 66234 116452 66240
rect 116398 65920 116454 65929
rect 116398 65855 116454 65864
rect 97356 65340 97408 65346
rect 97356 65282 97408 65288
rect 116412 64938 116440 65855
rect 116400 64932 116452 64938
rect 116400 64874 116452 64880
rect 115938 64696 115994 64705
rect 115938 64631 115994 64640
rect 115952 63578 115980 64631
rect 115940 63572 115992 63578
rect 115940 63514 115992 63520
rect 95976 63504 96028 63510
rect 95976 63446 96028 63452
rect 116214 63472 116270 63481
rect 116214 63407 116270 63416
rect 116228 62218 116256 63407
rect 116398 62384 116454 62393
rect 116398 62319 116454 62328
rect 116216 62212 116268 62218
rect 116216 62154 116268 62160
rect 116412 62150 116440 62319
rect 116400 62144 116452 62150
rect 116400 62086 116452 62092
rect 116596 62082 116624 71703
rect 214010 71632 214066 71641
rect 214010 71567 214066 71576
rect 213918 70952 213974 70961
rect 213918 70887 213974 70896
rect 213932 70446 213960 70887
rect 214024 70514 214052 71567
rect 214012 70508 214064 70514
rect 214012 70450 214064 70456
rect 213920 70440 213972 70446
rect 213920 70382 213972 70388
rect 214116 66230 214144 74015
rect 214562 72448 214618 72457
rect 214562 72383 214618 72392
rect 214470 68504 214526 68513
rect 214470 68439 214526 68448
rect 214484 67726 214512 68439
rect 214472 67720 214524 67726
rect 214472 67662 214524 67668
rect 214104 66224 214156 66230
rect 214104 66166 214156 66172
rect 214378 66192 214434 66201
rect 214378 66127 214434 66136
rect 214392 65550 214420 66127
rect 214380 65544 214432 65550
rect 214380 65486 214432 65492
rect 214010 65376 214066 65385
rect 214010 65311 214066 65320
rect 214024 64938 214052 65311
rect 214012 64932 214064 64938
rect 214012 64874 214064 64880
rect 214576 64870 214604 72383
rect 214654 70136 214710 70145
rect 214654 70071 214710 70080
rect 214668 69086 214696 70071
rect 214656 69080 214708 69086
rect 214656 69022 214708 69028
rect 214760 67590 214788 75511
rect 214852 70378 214880 78639
rect 214944 71738 214972 80271
rect 215128 80170 215156 80951
rect 215116 80164 215168 80170
rect 215116 80106 215168 80112
rect 215022 77208 215078 77217
rect 215022 77143 215078 77152
rect 214932 71732 214984 71738
rect 214932 71674 214984 71680
rect 214840 70372 214892 70378
rect 214840 70314 214892 70320
rect 215036 69018 215064 77143
rect 215220 73166 215248 81767
rect 215208 73160 215260 73166
rect 215208 73102 215260 73108
rect 215114 69320 215170 69329
rect 215114 69255 215170 69264
rect 215128 69154 215156 69255
rect 215116 69148 215168 69154
rect 215116 69090 215168 69096
rect 215024 69012 215076 69018
rect 215024 68954 215076 68960
rect 215114 67824 215170 67833
rect 215114 67759 215170 67768
rect 215128 67658 215156 67759
rect 215116 67652 215168 67658
rect 215116 67594 215168 67600
rect 214748 67584 214800 67590
rect 214748 67526 214800 67532
rect 215114 67008 215170 67017
rect 215114 66943 215170 66952
rect 215128 66298 215156 66943
rect 215116 66292 215168 66298
rect 215116 66234 215168 66240
rect 214564 64864 214616 64870
rect 214564 64806 214616 64812
rect 214562 64560 214618 64569
rect 214562 64495 214618 64504
rect 214576 63646 214604 64495
rect 215114 63880 215170 63889
rect 215114 63815 215170 63824
rect 214564 63640 214616 63646
rect 214564 63582 214616 63588
rect 215128 63578 215156 63815
rect 215116 63572 215168 63578
rect 215116 63514 215168 63520
rect 214654 63064 214710 63073
rect 214654 62999 214710 63008
rect 214668 62218 214696 62999
rect 215114 62248 215170 62257
rect 214656 62212 214708 62218
rect 215114 62183 215170 62192
rect 214656 62154 214708 62160
rect 215128 62150 215156 62183
rect 215116 62144 215168 62150
rect 215116 62086 215168 62092
rect 116584 62076 116636 62082
rect 116584 62018 116636 62024
rect 214562 61432 214618 61441
rect 214562 61367 214618 61376
rect 214576 61266 214604 61367
rect 214564 61260 214616 61266
rect 214564 61202 214616 61208
rect 116398 61160 116454 61169
rect 116398 61095 116454 61104
rect 116412 60790 116440 61095
rect 116400 60784 116452 60790
rect 215116 60784 215168 60790
rect 116400 60726 116452 60732
rect 215114 60752 215116 60761
rect 215168 60752 215170 60761
rect 215114 60687 215170 60696
rect 116398 60072 116454 60081
rect 116398 60007 116454 60016
rect 116412 59430 116440 60007
rect 214562 59936 214618 59945
rect 214562 59871 214618 59880
rect 214576 59430 214604 59871
rect 116400 59424 116452 59430
rect 116400 59366 116452 59372
rect 214564 59424 214616 59430
rect 214564 59366 214616 59372
rect 214102 59120 214158 59129
rect 214102 59055 214158 59064
rect 116398 58848 116454 58857
rect 116398 58783 116454 58792
rect 116412 58002 116440 58783
rect 214116 58070 214144 59055
rect 214194 58304 214250 58313
rect 214194 58239 214250 58248
rect 214104 58064 214156 58070
rect 214104 58006 214156 58012
rect 214208 58002 214236 58239
rect 116400 57996 116452 58002
rect 116400 57938 116452 57944
rect 214196 57996 214248 58002
rect 214196 57938 214248 57944
rect 116306 57624 116362 57633
rect 116306 57559 116362 57568
rect 213918 57624 213974 57633
rect 213918 57559 213974 57568
rect 116320 56642 116348 57559
rect 213932 56710 213960 57559
rect 214010 56808 214066 56817
rect 214010 56743 214066 56752
rect 213920 56704 213972 56710
rect 213920 56646 213972 56652
rect 214024 56642 214052 56743
rect 116308 56636 116360 56642
rect 116308 56578 116360 56584
rect 214012 56636 214064 56642
rect 214012 56578 214064 56584
rect 116306 56536 116362 56545
rect 116306 56471 116362 56480
rect 95146 55992 95202 56001
rect 95146 55927 95202 55936
rect 116320 55282 116348 56471
rect 215114 55992 215170 56001
rect 215114 55927 215170 55936
rect 116400 55344 116452 55350
rect 116398 55312 116400 55321
rect 116452 55312 116454 55321
rect 116308 55276 116360 55282
rect 215128 55282 215156 55927
rect 116398 55247 116454 55256
rect 215116 55276 215168 55282
rect 116308 55218 116360 55224
rect 215116 55218 215168 55224
rect 214746 55176 214802 55185
rect 214746 55111 214802 55120
rect 116398 54224 116454 54233
rect 116398 54159 116454 54168
rect 116412 53854 116440 54159
rect 214760 53854 214788 55111
rect 215114 54496 215170 54505
rect 215114 54431 215170 54440
rect 215128 53922 215156 54431
rect 215116 53916 215168 53922
rect 215116 53858 215168 53864
rect 116400 53848 116452 53854
rect 116400 53790 116452 53796
rect 214748 53848 214800 53854
rect 214748 53790 214800 53796
rect 214746 53680 214802 53689
rect 214746 53615 214802 53624
rect 116398 53000 116454 53009
rect 116398 52935 116454 52944
rect 116412 52494 116440 52935
rect 214760 52494 214788 53615
rect 215114 52864 215170 52873
rect 215114 52799 215170 52808
rect 215128 52562 215156 52799
rect 215116 52556 215168 52562
rect 215116 52498 215168 52504
rect 95148 52488 95200 52494
rect 95054 52456 95110 52465
rect 95148 52430 95200 52436
rect 116400 52488 116452 52494
rect 116400 52430 116452 52436
rect 214748 52488 214800 52494
rect 214748 52430 214800 52436
rect 95054 52391 95110 52400
rect 95056 49768 95108 49774
rect 95056 49710 95108 49716
rect 94778 47968 94834 47977
rect 94778 47903 94834 47912
rect 95068 45257 95096 49710
rect 95160 47025 95188 52430
rect 215114 52048 215170 52057
rect 215114 51983 215170 51992
rect 115938 51912 115994 51921
rect 115938 51847 115994 51856
rect 115952 51134 115980 51847
rect 214102 51368 214158 51377
rect 214102 51303 214158 51312
rect 214116 51134 214144 51303
rect 215128 51202 215156 51983
rect 215116 51196 215168 51202
rect 215116 51138 215168 51144
rect 115940 51128 115992 51134
rect 115940 51070 115992 51076
rect 214104 51128 214156 51134
rect 214104 51070 214156 51076
rect 116398 50688 116454 50697
rect 116398 50623 116454 50632
rect 116412 49774 116440 50623
rect 215206 50552 215262 50561
rect 215206 50487 215262 50496
rect 215116 49836 215168 49842
rect 215116 49778 215168 49784
rect 116400 49768 116452 49774
rect 215128 49745 215156 49778
rect 215220 49774 215248 50487
rect 215208 49768 215260 49774
rect 116400 49710 116452 49716
rect 215114 49736 215170 49745
rect 215208 49710 215260 49716
rect 215114 49671 215170 49680
rect 116398 49464 116454 49473
rect 116398 49399 116454 49408
rect 116124 48408 116176 48414
rect 116122 48376 116124 48385
rect 116176 48376 116178 48385
rect 116412 48346 116440 49399
rect 215114 48920 215170 48929
rect 215114 48855 215170 48864
rect 215128 48346 215156 48855
rect 116122 48311 116178 48320
rect 116400 48340 116452 48346
rect 116400 48282 116452 48288
rect 215116 48340 215168 48346
rect 215116 48282 215168 48288
rect 214746 48104 214802 48113
rect 214746 48039 214802 48048
rect 214010 47424 214066 47433
rect 214010 47359 214066 47368
rect 116398 47152 116454 47161
rect 116398 47087 116454 47096
rect 95146 47016 95202 47025
rect 116412 46986 116440 47087
rect 214024 46986 214052 47359
rect 214760 47054 214788 48039
rect 214748 47048 214800 47054
rect 214748 46990 214800 46996
rect 95146 46951 95202 46960
rect 116400 46980 116452 46986
rect 116400 46922 116452 46928
rect 214012 46980 214064 46986
rect 214012 46922 214064 46928
rect 215206 46608 215262 46617
rect 215206 46543 215262 46552
rect 116398 46064 116454 46073
rect 116398 45999 116454 46008
rect 116412 45626 116440 45999
rect 215114 45792 215170 45801
rect 215114 45727 215170 45736
rect 215128 45694 215156 45727
rect 215116 45688 215168 45694
rect 215116 45630 215168 45636
rect 215220 45626 215248 46543
rect 116400 45620 116452 45626
rect 116400 45562 116452 45568
rect 215208 45620 215260 45626
rect 215208 45562 215260 45568
rect 95054 45248 95110 45257
rect 95054 45183 95110 45192
rect 215206 44976 215262 44985
rect 215206 44911 215262 44920
rect 116398 44840 116454 44849
rect 116398 44775 116454 44784
rect 116412 44198 116440 44775
rect 215114 44296 215170 44305
rect 215220 44266 215248 44911
rect 215114 44231 215170 44240
rect 215208 44260 215260 44266
rect 215128 44198 215156 44231
rect 215208 44202 215260 44208
rect 94780 44192 94832 44198
rect 94780 44134 94832 44140
rect 116400 44192 116452 44198
rect 116400 44134 116452 44140
rect 215116 44192 215168 44198
rect 215116 44134 215168 44140
rect 94502 43480 94558 43489
rect 94502 43415 94558 43424
rect 94596 42832 94648 42838
rect 94596 42774 94648 42780
rect 94134 42528 94190 42537
rect 94134 42463 94190 42472
rect 93950 41712 94006 41721
rect 93950 41647 94006 41656
rect 94504 40180 94556 40186
rect 94504 40122 94556 40128
rect 94516 38185 94544 40122
rect 94608 39953 94636 42774
rect 94792 40769 94820 44134
rect 115938 43616 115994 43625
rect 115938 43551 115994 43560
rect 115952 42838 115980 43551
rect 214378 43480 214434 43489
rect 214378 43415 214434 43424
rect 214392 42838 214420 43415
rect 115940 42832 115992 42838
rect 115940 42774 115992 42780
rect 214380 42832 214432 42838
rect 214380 42774 214432 42780
rect 214102 42664 214158 42673
rect 214102 42599 214158 42608
rect 116398 42528 116454 42537
rect 116398 42463 116454 42472
rect 116412 41478 116440 42463
rect 214116 41478 214144 42599
rect 215114 41848 215170 41857
rect 215114 41783 215170 41792
rect 215128 41546 215156 41783
rect 215116 41540 215168 41546
rect 215116 41482 215168 41488
rect 95148 41472 95200 41478
rect 95148 41414 95200 41420
rect 116400 41472 116452 41478
rect 116400 41414 116452 41420
rect 214104 41472 214156 41478
rect 214104 41414 214156 41420
rect 94778 40760 94834 40769
rect 94778 40695 94834 40704
rect 95056 40112 95108 40118
rect 95056 40054 95108 40060
rect 94594 39944 94650 39953
rect 94594 39879 94650 39888
rect 94596 38684 94648 38690
rect 94596 38626 94648 38632
rect 94502 38176 94558 38185
rect 94502 38111 94558 38120
rect 93860 37324 93912 37330
rect 93860 37266 93912 37272
rect 93872 35465 93900 37266
rect 94608 36281 94636 38626
rect 95068 37233 95096 40054
rect 95160 39001 95188 41414
rect 116306 41304 116362 41313
rect 116306 41239 116362 41248
rect 116320 40186 116348 41239
rect 214654 41168 214710 41177
rect 214654 41103 214710 41112
rect 116398 40216 116454 40225
rect 116308 40180 116360 40186
rect 116398 40151 116454 40160
rect 116308 40122 116360 40128
rect 116412 40118 116440 40151
rect 214668 40118 214696 41103
rect 215114 40352 215170 40361
rect 215114 40287 215170 40296
rect 215128 40186 215156 40287
rect 215116 40180 215168 40186
rect 215116 40122 215168 40128
rect 116400 40112 116452 40118
rect 116400 40054 116452 40060
rect 214656 40112 214708 40118
rect 214656 40054 214708 40060
rect 214562 39536 214618 39545
rect 214562 39471 214618 39480
rect 95146 38992 95202 39001
rect 95146 38927 95202 38936
rect 116398 38992 116454 39001
rect 116398 38927 116454 38936
rect 116412 38690 116440 38927
rect 214576 38690 214604 39471
rect 215116 38752 215168 38758
rect 215114 38720 215116 38729
rect 215168 38720 215170 38729
rect 116400 38684 116452 38690
rect 116400 38626 116452 38632
rect 214564 38684 214616 38690
rect 215114 38655 215170 38664
rect 214564 38626 214616 38632
rect 215114 38040 215170 38049
rect 215114 37975 215170 37984
rect 116398 37768 116454 37777
rect 116398 37703 116454 37712
rect 116412 37330 116440 37703
rect 215128 37330 215156 37975
rect 116400 37324 116452 37330
rect 116400 37266 116452 37272
rect 215116 37324 215168 37330
rect 215116 37266 215168 37272
rect 95054 37224 95110 37233
rect 95054 37159 95110 37168
rect 214102 37224 214158 37233
rect 214102 37159 214158 37168
rect 116398 36680 116454 36689
rect 116398 36615 116454 36624
rect 94594 36272 94650 36281
rect 94594 36207 94650 36216
rect 116412 35970 116440 36615
rect 214116 36038 214144 37159
rect 215114 36408 215170 36417
rect 215114 36343 215170 36352
rect 214104 36032 214156 36038
rect 214104 35974 214156 35980
rect 215128 35970 215156 36343
rect 93952 35964 94004 35970
rect 93952 35906 94004 35912
rect 116400 35964 116452 35970
rect 116400 35906 116452 35912
rect 215116 35964 215168 35970
rect 215116 35906 215168 35912
rect 93858 35456 93914 35465
rect 93858 35391 93914 35400
rect 93964 34513 93992 35906
rect 214654 35592 214710 35601
rect 214654 35527 214710 35536
rect 116398 35456 116454 35465
rect 116398 35391 116454 35400
rect 116412 34542 116440 35391
rect 214668 34542 214696 35527
rect 215114 34912 215170 34921
rect 215114 34847 215170 34856
rect 215128 34610 215156 34847
rect 215116 34604 215168 34610
rect 215116 34546 215168 34552
rect 95148 34536 95200 34542
rect 93950 34504 94006 34513
rect 95148 34478 95200 34484
rect 116400 34536 116452 34542
rect 116400 34478 116452 34484
rect 214656 34536 214708 34542
rect 214656 34478 214708 34484
rect 93950 34439 94006 34448
rect 95160 33697 95188 34478
rect 116306 34368 116362 34377
rect 116306 34303 116362 34312
rect 95146 33688 95202 33697
rect 95146 33623 95202 33632
rect 116320 33182 116348 34303
rect 214562 34096 214618 34105
rect 214562 34031 214618 34040
rect 214576 33250 214604 34031
rect 215114 33280 215170 33289
rect 214564 33244 214616 33250
rect 215114 33215 215170 33224
rect 214564 33186 214616 33192
rect 215128 33182 215156 33215
rect 95148 33176 95200 33182
rect 95148 33118 95200 33124
rect 116308 33176 116360 33182
rect 215116 33176 215168 33182
rect 116308 33118 116360 33124
rect 116398 33144 116454 33153
rect 95160 32745 95188 33118
rect 215116 33118 215168 33124
rect 116398 33079 116454 33088
rect 95146 32736 95202 32745
rect 95146 32671 95202 32680
rect 116412 32434 116440 33079
rect 215956 32570 215984 82826
rect 220176 80164 220228 80170
rect 220176 80106 220228 80112
rect 218796 77308 218848 77314
rect 218796 77250 218848 77256
rect 216036 74656 216088 74662
rect 216036 74598 216088 74604
rect 216048 67522 216076 74598
rect 218060 73228 218112 73234
rect 218060 73170 218112 73176
rect 216036 67516 216088 67522
rect 216036 67458 216088 67464
rect 218072 66162 218100 73170
rect 218808 70310 218836 77250
rect 219440 76084 219492 76090
rect 219440 76026 219492 76032
rect 218796 70304 218848 70310
rect 218796 70246 218848 70252
rect 219452 68950 219480 76026
rect 220188 73098 220216 80106
rect 220820 78804 220872 78810
rect 220820 78746 220872 78752
rect 220176 73092 220228 73098
rect 220176 73034 220228 73040
rect 220832 71670 220860 78746
rect 224236 75886 224264 85546
rect 225604 84244 225656 84250
rect 225604 84186 225656 84192
rect 224224 75880 224276 75886
rect 224224 75822 224276 75828
rect 225616 74633 225644 84186
rect 226984 81456 227036 81462
rect 226984 81398 227036 81404
rect 225602 74624 225658 74633
rect 225602 74559 225658 74568
rect 226996 73273 227024 81398
rect 227352 81388 227404 81394
rect 227352 81330 227404 81336
rect 227364 80481 227392 81330
rect 227444 81320 227496 81326
rect 227444 81262 227496 81268
rect 227456 81161 227484 81262
rect 227442 81152 227498 81161
rect 227442 81087 227498 81096
rect 227350 80472 227406 80481
rect 227350 80407 227406 80416
rect 232424 80170 232452 89678
rect 340156 88330 340184 309130
rect 341536 135250 341564 310490
rect 341524 135244 341576 135250
rect 341524 135186 341576 135192
rect 343652 126721 343680 428431
rect 411904 227044 411956 227050
rect 411904 226986 411956 226992
rect 343638 126712 343694 126721
rect 343638 126647 343694 126656
rect 340144 88324 340196 88330
rect 340144 88266 340196 88272
rect 284484 83564 284536 83570
rect 284484 83506 284536 83512
rect 248144 82884 248196 82890
rect 248144 82826 248196 82832
rect 248156 81396 248184 82826
rect 284496 81396 284524 83506
rect 320824 83496 320876 83502
rect 320824 83438 320876 83444
rect 320836 81396 320864 83438
rect 232412 80164 232464 80170
rect 232412 80106 232464 80112
rect 227536 80028 227588 80034
rect 227536 79970 227588 79976
rect 232320 80028 232372 80034
rect 232320 79970 232372 79976
rect 227444 79960 227496 79966
rect 227444 79902 227496 79908
rect 227456 79801 227484 79902
rect 227442 79792 227498 79801
rect 227442 79727 227498 79736
rect 227548 79121 227576 79970
rect 227534 79112 227590 79121
rect 227534 79047 227590 79056
rect 227536 78668 227588 78674
rect 227536 78610 227588 78616
rect 227444 78600 227496 78606
rect 227442 78568 227444 78577
rect 227496 78568 227498 78577
rect 227442 78503 227498 78512
rect 227548 77897 227576 78610
rect 227534 77888 227590 77897
rect 227534 77823 227590 77832
rect 227444 77240 227496 77246
rect 227442 77208 227444 77217
rect 227496 77208 227498 77217
rect 227442 77143 227498 77152
rect 227536 77172 227588 77178
rect 227536 77114 227588 77120
rect 227548 76537 227576 77114
rect 227534 76528 227590 76537
rect 227534 76463 227590 76472
rect 227444 75880 227496 75886
rect 227442 75848 227444 75857
rect 227496 75848 227498 75857
rect 227442 75783 227498 75792
rect 227444 75744 227496 75750
rect 227444 75686 227496 75692
rect 227456 75313 227484 75686
rect 227442 75304 227498 75313
rect 227442 75239 227498 75248
rect 227444 74520 227496 74526
rect 227444 74462 227496 74468
rect 227456 73953 227484 74462
rect 227442 73944 227498 73953
rect 227442 73879 227498 73888
rect 226982 73264 227038 73273
rect 226982 73199 227038 73208
rect 227444 73160 227496 73166
rect 227444 73102 227496 73108
rect 227456 72729 227484 73102
rect 227536 73092 227588 73098
rect 227536 73034 227588 73040
rect 227442 72720 227498 72729
rect 227442 72655 227498 72664
rect 227548 72049 227576 73034
rect 227534 72040 227590 72049
rect 227534 71975 227590 71984
rect 227444 71732 227496 71738
rect 227444 71674 227496 71680
rect 220820 71664 220872 71670
rect 220820 71606 220872 71612
rect 227456 71369 227484 71674
rect 227536 71664 227588 71670
rect 227536 71606 227588 71612
rect 227442 71360 227498 71369
rect 227442 71295 227498 71304
rect 227548 70689 227576 71606
rect 227534 70680 227590 70689
rect 227534 70615 227590 70624
rect 224500 70508 224552 70514
rect 224500 70450 224552 70456
rect 224408 70440 224460 70446
rect 224408 70382 224460 70388
rect 224224 69148 224276 69154
rect 224224 69090 224276 69096
rect 224132 69080 224184 69086
rect 224132 69022 224184 69028
rect 219440 68944 219492 68950
rect 219440 68886 219492 68892
rect 218060 66156 218112 66162
rect 218060 66098 218112 66104
rect 216772 65544 216824 65550
rect 216772 65486 216824 65492
rect 216680 62212 216732 62218
rect 216680 62154 216732 62160
rect 216692 57934 216720 62154
rect 216784 60722 216812 65486
rect 216956 63640 217008 63646
rect 216956 63582 217008 63588
rect 216864 61260 216916 61266
rect 216864 61202 216916 61208
rect 216772 60716 216824 60722
rect 216772 60658 216824 60664
rect 216680 57928 216732 57934
rect 216680 57870 216732 57876
rect 216772 56704 216824 56710
rect 216772 56646 216824 56652
rect 216680 56636 216732 56642
rect 216680 56578 216732 56584
rect 216692 52426 216720 56578
rect 216680 52420 216732 52426
rect 216680 52362 216732 52368
rect 216784 52358 216812 56646
rect 216876 56574 216904 61202
rect 216968 59362 216996 63582
rect 224040 63572 224092 63578
rect 224040 63514 224092 63520
rect 217600 59424 217652 59430
rect 217600 59366 217652 59372
rect 216956 59356 217008 59362
rect 216956 59298 217008 59304
rect 217508 58064 217560 58070
rect 217508 58006 217560 58012
rect 217416 57996 217468 58002
rect 217416 57938 217468 57944
rect 216864 56568 216916 56574
rect 216864 56510 216916 56516
rect 217428 53718 217456 57938
rect 217520 53786 217548 58006
rect 217612 55214 217640 59366
rect 224052 57866 224080 63514
rect 224144 63510 224172 69022
rect 224132 63504 224184 63510
rect 224132 63446 224184 63452
rect 224236 63442 224264 69090
rect 224316 66292 224368 66298
rect 224316 66234 224368 66240
rect 224224 63436 224276 63442
rect 224224 63378 224276 63384
rect 224132 62144 224184 62150
rect 224132 62086 224184 62092
rect 224040 57860 224092 57866
rect 224040 57802 224092 57808
rect 224144 56506 224172 62086
rect 224224 60784 224276 60790
rect 224224 60726 224276 60732
rect 224132 56500 224184 56506
rect 224132 56442 224184 56448
rect 224236 55214 224264 60726
rect 224328 60654 224356 66234
rect 224420 64326 224448 70382
rect 224512 64530 224540 70450
rect 227444 70372 227496 70378
rect 227444 70314 227496 70320
rect 226524 70304 226576 70310
rect 226524 70246 226576 70252
rect 226536 69465 226564 70246
rect 227456 70009 227484 70314
rect 232332 70258 232360 79970
rect 232240 70230 232360 70258
rect 227442 70000 227498 70009
rect 227442 69935 227498 69944
rect 226522 69456 226578 69465
rect 226522 69391 226578 69400
rect 227444 69012 227496 69018
rect 227444 68954 227496 68960
rect 227456 68785 227484 68954
rect 227536 68944 227588 68950
rect 227536 68886 227588 68892
rect 227442 68776 227498 68785
rect 227442 68711 227498 68720
rect 227548 68105 227576 68886
rect 227534 68096 227590 68105
rect 227534 68031 227590 68040
rect 224684 67720 224736 67726
rect 224684 67662 224736 67668
rect 224592 64932 224644 64938
rect 224592 64874 224644 64880
rect 224500 64524 224552 64530
rect 224500 64466 224552 64472
rect 224408 64320 224460 64326
rect 224408 64262 224460 64268
rect 224316 60648 224368 60654
rect 224316 60590 224368 60596
rect 224604 59294 224632 64874
rect 224696 62082 224724 67662
rect 224868 67652 224920 67658
rect 224868 67594 224920 67600
rect 224684 62076 224736 62082
rect 224684 62018 224736 62024
rect 224880 62014 224908 67594
rect 227444 67584 227496 67590
rect 227444 67526 227496 67532
rect 227456 67425 227484 67526
rect 227536 67516 227588 67522
rect 227536 67458 227588 67464
rect 227442 67416 227498 67425
rect 227442 67351 227498 67360
rect 227548 66881 227576 67458
rect 227534 66872 227590 66881
rect 227534 66807 227590 66816
rect 227444 66224 227496 66230
rect 227442 66192 227444 66201
rect 227496 66192 227498 66201
rect 227442 66127 227498 66136
rect 227536 66156 227588 66162
rect 227536 66098 227588 66104
rect 227548 65521 227576 66098
rect 227534 65512 227590 65521
rect 227534 65447 227590 65456
rect 227444 64864 227496 64870
rect 227442 64832 227444 64841
rect 227496 64832 227498 64841
rect 227442 64767 227498 64776
rect 227444 64524 227496 64530
rect 227444 64466 227496 64472
rect 227456 64161 227484 64466
rect 227536 64320 227588 64326
rect 227536 64262 227588 64268
rect 227442 64152 227498 64161
rect 227442 64087 227498 64096
rect 227548 63617 227576 64262
rect 227534 63608 227590 63617
rect 227534 63543 227590 63552
rect 227444 63504 227496 63510
rect 227444 63446 227496 63452
rect 227456 62937 227484 63446
rect 227536 63436 227588 63442
rect 227536 63378 227588 63384
rect 227442 62928 227498 62937
rect 227442 62863 227498 62872
rect 227548 62257 227576 63378
rect 227534 62248 227590 62257
rect 227534 62183 227590 62192
rect 227536 62076 227588 62082
rect 227536 62018 227588 62024
rect 224868 62008 224920 62014
rect 224868 61950 224920 61956
rect 226708 62008 226760 62014
rect 226708 61950 226760 61956
rect 226720 61033 226748 61950
rect 227548 61577 227576 62018
rect 227534 61568 227590 61577
rect 227534 61503 227590 61512
rect 226706 61024 226762 61033
rect 226706 60959 226762 60968
rect 227444 60716 227496 60722
rect 227444 60658 227496 60664
rect 227076 60648 227128 60654
rect 227076 60590 227128 60596
rect 227088 60353 227116 60590
rect 227074 60344 227130 60353
rect 227074 60279 227130 60288
rect 227456 59673 227484 60658
rect 232240 60602 232268 70230
rect 232240 60574 232360 60602
rect 227442 59664 227498 59673
rect 227442 59599 227498 59608
rect 227536 59356 227588 59362
rect 227536 59298 227588 59304
rect 224592 59288 224644 59294
rect 224592 59230 224644 59236
rect 227444 59288 227496 59294
rect 227444 59230 227496 59236
rect 227456 58993 227484 59230
rect 227442 58984 227498 58993
rect 227442 58919 227498 58928
rect 227548 58313 227576 59298
rect 227534 58304 227590 58313
rect 227534 58239 227590 58248
rect 227444 57928 227496 57934
rect 232332 57882 232360 60574
rect 227444 57870 227496 57876
rect 227260 57860 227312 57866
rect 227260 57802 227312 57808
rect 227272 57769 227300 57802
rect 227258 57760 227314 57769
rect 227258 57695 227314 57704
rect 227456 57089 227484 57870
rect 232240 57854 232360 57882
rect 227442 57080 227498 57089
rect 227442 57015 227498 57024
rect 227444 56568 227496 56574
rect 227444 56510 227496 56516
rect 227260 56500 227312 56506
rect 227260 56442 227312 56448
rect 227272 56409 227300 56442
rect 227258 56400 227314 56409
rect 227258 56335 227314 56344
rect 227456 55729 227484 56510
rect 227442 55720 227498 55729
rect 227442 55655 227498 55664
rect 227536 55276 227588 55282
rect 227536 55218 227588 55224
rect 217600 55208 217652 55214
rect 217600 55150 217652 55156
rect 224224 55208 224276 55214
rect 227444 55208 227496 55214
rect 224224 55150 224276 55156
rect 227442 55176 227444 55185
rect 227496 55176 227498 55185
rect 227442 55111 227498 55120
rect 226524 55072 226576 55078
rect 226524 55014 226576 55020
rect 226536 54505 226564 55014
rect 226522 54496 226578 54505
rect 226522 54431 226578 54440
rect 226984 53916 227036 53922
rect 226984 53858 227036 53864
rect 226616 53848 226668 53854
rect 226616 53790 226668 53796
rect 217508 53780 217560 53786
rect 217508 53722 217560 53728
rect 217416 53712 217468 53718
rect 217416 53654 217468 53660
rect 226524 53712 226576 53718
rect 226524 53654 226576 53660
rect 226536 53145 226564 53654
rect 226522 53136 226578 53145
rect 226522 53071 226578 53080
rect 216772 52352 216824 52358
rect 216772 52294 216824 52300
rect 226340 51196 226392 51202
rect 226340 51138 226392 51144
rect 226352 47977 226380 51138
rect 226524 51128 226576 51134
rect 226524 51070 226576 51076
rect 226338 47968 226394 47977
rect 226338 47903 226394 47912
rect 226536 47297 226564 51070
rect 226628 50561 226656 53790
rect 226800 52556 226852 52562
rect 226800 52498 226852 52504
rect 226708 52488 226760 52494
rect 226708 52430 226760 52436
rect 226614 50552 226670 50561
rect 226614 50487 226670 50496
rect 226720 49337 226748 52430
rect 226706 49328 226762 49337
rect 226706 49263 226762 49272
rect 226812 48657 226840 52498
rect 226996 49881 227024 53858
rect 227442 53816 227498 53825
rect 227442 53751 227444 53760
rect 227496 53751 227498 53760
rect 227444 53722 227496 53728
rect 227258 52456 227314 52465
rect 227258 52391 227314 52400
rect 227444 52420 227496 52426
rect 227272 52358 227300 52391
rect 227444 52362 227496 52368
rect 227260 52352 227312 52358
rect 227260 52294 227312 52300
rect 227456 51921 227484 52362
rect 227442 51912 227498 51921
rect 227442 51847 227498 51856
rect 227548 51241 227576 55218
rect 227534 51232 227590 51241
rect 227534 51167 227590 51176
rect 232240 51082 232268 57854
rect 232240 51054 232360 51082
rect 226982 49872 227038 49881
rect 226982 49807 227038 49816
rect 227628 49836 227680 49842
rect 227628 49778 227680 49784
rect 227536 49768 227588 49774
rect 227536 49710 227588 49716
rect 226798 48648 226854 48657
rect 226798 48583 226854 48592
rect 227352 48340 227404 48346
rect 227352 48282 227404 48288
rect 226522 47288 226578 47297
rect 226522 47223 226578 47232
rect 226708 46980 226760 46986
rect 226708 46922 226760 46928
rect 226720 44033 226748 46922
rect 227260 45688 227312 45694
rect 227260 45630 227312 45636
rect 227076 45620 227128 45626
rect 227076 45562 227128 45568
rect 226706 44024 226762 44033
rect 226706 43959 226762 43968
rect 227088 43489 227116 45562
rect 227074 43480 227130 43489
rect 227074 43415 227130 43424
rect 226432 42832 226484 42838
rect 227272 42809 227300 45630
rect 227364 45393 227392 48282
rect 227444 47048 227496 47054
rect 227444 46990 227496 46996
rect 227350 45384 227406 45393
rect 227350 45319 227406 45328
rect 227456 44713 227484 46990
rect 227548 46617 227576 49710
rect 227534 46608 227590 46617
rect 227534 46543 227590 46552
rect 227640 46073 227668 49778
rect 232332 48362 232360 51054
rect 411916 49881 411944 226986
rect 413296 83570 413324 502930
rect 414032 502846 414184 502874
rect 414032 496126 414060 502846
rect 416148 500274 416176 502982
rect 420840 500954 420868 502982
rect 433444 502982 433596 503010
rect 435560 502982 435712 503010
rect 442000 502982 442152 503010
rect 446324 502982 446476 503010
rect 480824 502982 481312 503010
rect 422832 502846 423168 502874
rect 424948 502846 425008 502874
rect 427064 502846 427124 502874
rect 429272 502846 429332 502874
rect 431388 502846 431448 502874
rect 423140 500954 423168 502846
rect 424980 500954 425008 502846
rect 427096 500954 427124 502846
rect 429304 500954 429332 502846
rect 431420 500954 431448 502846
rect 433444 500954 433472 502982
rect 435560 500954 435588 502982
rect 437584 502846 437920 502874
rect 439700 502846 440036 502874
rect 437584 500954 437612 502846
rect 439700 500954 439728 502846
rect 442000 500954 442028 502982
rect 444360 502846 444420 502874
rect 444392 500954 444420 502846
rect 446324 500954 446352 502982
rect 448532 502846 448684 502874
rect 450464 502846 450800 502874
rect 453008 502846 453344 502874
rect 455124 502846 455368 502874
rect 457332 502846 457392 502874
rect 459448 502846 459508 502874
rect 448532 500954 448560 502846
rect 450464 500954 450492 502846
rect 453316 500954 453344 502846
rect 455340 500954 455368 502846
rect 457364 500954 457392 502846
rect 459480 502722 459508 502846
rect 461228 502846 461900 502874
rect 463772 502846 464108 502874
rect 465888 502846 465948 502874
rect 468096 502846 468156 502874
rect 470212 502846 470272 502874
rect 472420 502846 472756 502874
rect 474536 502846 474688 502874
rect 477756 502846 477816 502874
rect 461228 502722 461256 502846
rect 459468 502716 459520 502722
rect 459468 502658 459520 502664
rect 461216 502716 461268 502722
rect 461216 502658 461268 502664
rect 461872 500954 461900 502846
rect 464080 500954 464108 502846
rect 465920 500954 465948 502846
rect 468128 500954 468156 502846
rect 470244 500954 470272 502846
rect 472728 500954 472756 502846
rect 474660 500954 474688 502846
rect 477788 500954 477816 502846
rect 480824 500954 480852 502982
rect 481284 502926 481312 502982
rect 481272 502920 481324 502926
rect 484308 502920 484360 502926
rect 481272 502862 481324 502868
rect 484196 502868 484308 502874
rect 484196 502862 484360 502868
rect 487160 502920 487212 502926
rect 487212 502868 487508 502874
rect 487160 502862 487508 502868
rect 484196 502846 484348 502862
rect 487172 502846 487508 502862
rect 491740 502846 492076 502874
rect 492844 502846 493180 502874
rect 493948 502846 494008 502874
rect 495052 502846 495388 502874
rect 496064 502846 496768 502874
rect 497168 502846 497504 502874
rect 498272 502846 498608 502874
rect 492048 500954 492076 502846
rect 420828 500948 420880 500954
rect 420828 500890 420880 500896
rect 423128 500948 423180 500954
rect 423128 500890 423180 500896
rect 424968 500948 425020 500954
rect 424968 500890 425020 500896
rect 427084 500948 427136 500954
rect 427084 500890 427136 500896
rect 429292 500948 429344 500954
rect 429292 500890 429344 500896
rect 431408 500948 431460 500954
rect 431408 500890 431460 500896
rect 433432 500948 433484 500954
rect 433432 500890 433484 500896
rect 435548 500948 435600 500954
rect 435548 500890 435600 500896
rect 437572 500948 437624 500954
rect 437572 500890 437624 500896
rect 439688 500948 439740 500954
rect 439688 500890 439740 500896
rect 441988 500948 442040 500954
rect 441988 500890 442040 500896
rect 444380 500948 444432 500954
rect 444380 500890 444432 500896
rect 446312 500948 446364 500954
rect 446312 500890 446364 500896
rect 448520 500948 448572 500954
rect 448520 500890 448572 500896
rect 450452 500948 450504 500954
rect 450452 500890 450504 500896
rect 453304 500948 453356 500954
rect 453304 500890 453356 500896
rect 455328 500948 455380 500954
rect 455328 500890 455380 500896
rect 457352 500948 457404 500954
rect 457352 500890 457404 500896
rect 461860 500948 461912 500954
rect 461860 500890 461912 500896
rect 464068 500948 464120 500954
rect 464068 500890 464120 500896
rect 465908 500948 465960 500954
rect 465908 500890 465960 500896
rect 468116 500948 468168 500954
rect 468116 500890 468168 500896
rect 470232 500948 470284 500954
rect 470232 500890 470284 500896
rect 472716 500948 472768 500954
rect 472716 500890 472768 500896
rect 474648 500948 474700 500954
rect 474648 500890 474700 500896
rect 477776 500948 477828 500954
rect 477776 500890 477828 500896
rect 480812 500948 480864 500954
rect 480812 500890 480864 500896
rect 492036 500948 492088 500954
rect 492036 500890 492088 500896
rect 492588 500948 492640 500954
rect 492588 500890 492640 500896
rect 416136 500268 416188 500274
rect 416136 500210 416188 500216
rect 414020 496120 414072 496126
rect 414020 496062 414072 496068
rect 443644 494760 443696 494766
rect 443644 494702 443696 494708
rect 443656 450673 443684 494702
rect 492600 476814 492628 500890
rect 493152 499866 493180 502846
rect 493140 499860 493192 499866
rect 493140 499802 493192 499808
rect 492588 476808 492640 476814
rect 492588 476750 492640 476756
rect 493980 475425 494008 502846
rect 494704 499860 494756 499866
rect 494704 499802 494756 499808
rect 494716 479534 494744 499802
rect 495360 491978 495388 502846
rect 495348 491972 495400 491978
rect 495348 491914 495400 491920
rect 494704 479528 494756 479534
rect 494704 479470 494756 479476
rect 496740 478174 496768 502846
rect 497476 500177 497504 502846
rect 498384 500948 498436 500954
rect 498384 500890 498436 500896
rect 497462 500168 497518 500177
rect 497462 500103 497518 500112
rect 498396 497486 498424 500890
rect 498580 500274 498608 502846
rect 498948 502846 499284 502874
rect 500388 502846 500724 502874
rect 501492 502846 501828 502874
rect 502596 502846 502932 502874
rect 498948 500954 498976 502846
rect 498936 500948 498988 500954
rect 498936 500890 498988 500896
rect 500696 500313 500724 502846
rect 500682 500304 500738 500313
rect 498568 500268 498620 500274
rect 498568 500210 498620 500216
rect 499488 500268 499540 500274
rect 500682 500239 500738 500248
rect 499488 500210 499540 500216
rect 498384 497480 498436 497486
rect 498384 497422 498436 497428
rect 499500 490618 499528 500210
rect 501800 500070 501828 502846
rect 502432 500948 502484 500954
rect 502432 500890 502484 500896
rect 501788 500064 501840 500070
rect 501788 500006 501840 500012
rect 502248 500064 502300 500070
rect 502248 500006 502300 500012
rect 499488 490612 499540 490618
rect 499488 490554 499540 490560
rect 496728 478168 496780 478174
rect 496728 478110 496780 478116
rect 499304 475448 499356 475454
rect 493966 475416 494022 475425
rect 499304 475390 499356 475396
rect 493966 475351 494022 475360
rect 499316 473620 499344 475390
rect 502260 474026 502288 500006
rect 502444 494766 502472 500890
rect 502904 500274 502932 502846
rect 503272 502846 503608 502874
rect 504712 502846 505048 502874
rect 505816 502846 506152 502874
rect 506828 502846 507164 502874
rect 507932 502846 508268 502874
rect 509036 502846 509096 502874
rect 503272 500954 503300 502846
rect 503260 500948 503312 500954
rect 503260 500890 503312 500896
rect 502892 500268 502944 500274
rect 502892 500210 502944 500216
rect 502432 494760 502484 494766
rect 502432 494702 502484 494708
rect 505020 486470 505048 502846
rect 506124 500410 506152 502846
rect 507136 500682 507164 502846
rect 507124 500676 507176 500682
rect 507124 500618 507176 500624
rect 507768 500676 507820 500682
rect 507768 500618 507820 500624
rect 506112 500404 506164 500410
rect 506112 500346 506164 500352
rect 505008 486464 505060 486470
rect 505008 486406 505060 486412
rect 507780 475561 507808 500618
rect 508240 500449 508268 502846
rect 508226 500440 508282 500449
rect 508226 500375 508282 500384
rect 509068 500342 509096 502846
rect 509804 502846 510140 502874
rect 511152 502846 511488 502874
rect 512256 502846 512592 502874
rect 513360 502846 513696 502874
rect 514372 502846 514708 502874
rect 515476 502846 515812 502874
rect 516580 502846 516916 502874
rect 517684 502846 518020 502874
rect 518696 502846 518756 502874
rect 519800 502846 520228 502874
rect 520904 502846 521608 502874
rect 521916 502846 522252 502874
rect 523020 502846 523356 502874
rect 524124 502846 524368 502874
rect 525228 502846 525748 502874
rect 526240 502846 526576 502874
rect 527344 502846 527680 502874
rect 528448 502846 528508 502874
rect 529460 502846 529888 502874
rect 530564 502846 531268 502874
rect 531668 502846 532004 502874
rect 532772 502846 533108 502874
rect 533784 502846 533936 502874
rect 534888 502846 535408 502874
rect 535992 502846 536328 502874
rect 537004 502846 537340 502874
rect 509804 500954 509832 502846
rect 511460 500954 511488 502846
rect 509240 500948 509292 500954
rect 509240 500890 509292 500896
rect 509792 500948 509844 500954
rect 509792 500890 509844 500896
rect 511448 500948 511500 500954
rect 511448 500890 511500 500896
rect 511908 500948 511960 500954
rect 511908 500890 511960 500896
rect 509056 500336 509108 500342
rect 509056 500278 509108 500284
rect 509252 493338 509280 500890
rect 509240 493332 509292 493338
rect 509240 493274 509292 493280
rect 511920 483682 511948 500890
rect 512564 500721 512592 502846
rect 512550 500712 512606 500721
rect 512550 500647 512606 500656
rect 513668 500410 513696 502846
rect 514680 500585 514708 502846
rect 514666 500576 514722 500585
rect 514666 500511 514722 500520
rect 515784 500478 515812 502846
rect 515772 500472 515824 500478
rect 515772 500414 515824 500420
rect 512644 500404 512696 500410
rect 512644 500346 512696 500352
rect 513656 500404 513708 500410
rect 513656 500346 513708 500352
rect 511908 483676 511960 483682
rect 511908 483618 511960 483624
rect 507766 475552 507822 475561
rect 507766 475487 507822 475496
rect 512656 474094 512684 500346
rect 516888 500070 516916 502846
rect 516876 500064 516928 500070
rect 516876 500006 516928 500012
rect 517428 500064 517480 500070
rect 517428 500006 517480 500012
rect 517440 480962 517468 500006
rect 517992 499866 518020 502846
rect 517980 499860 518032 499866
rect 517980 499802 518032 499808
rect 517428 480956 517480 480962
rect 517428 480898 517480 480904
rect 518728 475386 518756 502846
rect 518808 499860 518860 499866
rect 518808 499802 518860 499808
rect 518716 475380 518768 475386
rect 518716 475322 518768 475328
rect 518820 474162 518848 499802
rect 520200 481030 520228 502846
rect 521580 483750 521608 502846
rect 522224 500954 522252 502846
rect 522212 500948 522264 500954
rect 522212 500890 522264 500896
rect 522948 500948 523000 500954
rect 522948 500890 523000 500896
rect 521568 483744 521620 483750
rect 521568 483686 521620 483692
rect 520188 481024 520240 481030
rect 520188 480966 520240 480972
rect 522960 478242 522988 500890
rect 523328 500546 523356 502846
rect 523316 500540 523368 500546
rect 523316 500482 523368 500488
rect 522948 478236 523000 478242
rect 522948 478178 523000 478184
rect 524340 476882 524368 502846
rect 525720 479670 525748 502846
rect 526548 500002 526576 502846
rect 527652 500954 527680 502846
rect 527640 500948 527692 500954
rect 527640 500890 527692 500896
rect 528376 500948 528428 500954
rect 528376 500890 528428 500896
rect 526536 499996 526588 500002
rect 526536 499938 526588 499944
rect 527088 499996 527140 500002
rect 527088 499938 527140 499944
rect 525708 479664 525760 479670
rect 525708 479606 525760 479612
rect 527100 479602 527128 499938
rect 527824 498840 527876 498846
rect 527824 498782 527876 498788
rect 527088 479596 527140 479602
rect 527088 479538 527140 479544
rect 524328 476876 524380 476882
rect 524328 476818 524380 476824
rect 527836 475454 527864 498782
rect 528388 482322 528416 500890
rect 528376 482316 528428 482322
rect 528376 482258 528428 482264
rect 528480 475454 528508 502846
rect 529860 481098 529888 502846
rect 529848 481092 529900 481098
rect 529848 481034 529900 481040
rect 531240 475522 531268 502846
rect 531976 500954 532004 502846
rect 533080 500954 533108 502846
rect 531964 500948 532016 500954
rect 531964 500890 532016 500896
rect 532608 500948 532660 500954
rect 532608 500890 532660 500896
rect 533068 500948 533120 500954
rect 533068 500890 533120 500896
rect 532620 478310 532648 500890
rect 533908 500614 533936 502846
rect 533988 500948 534040 500954
rect 533988 500890 534040 500896
rect 533896 500608 533948 500614
rect 533896 500550 533948 500556
rect 532608 478304 532660 478310
rect 532608 478246 532660 478252
rect 531228 475516 531280 475522
rect 531228 475458 531280 475464
rect 527824 475448 527876 475454
rect 527824 475390 527876 475396
rect 528468 475448 528520 475454
rect 528468 475390 528520 475396
rect 534000 474230 534028 500890
rect 535380 476950 535408 502846
rect 536300 500954 536328 502846
rect 536288 500948 536340 500954
rect 536288 500890 536340 500896
rect 536748 500948 536800 500954
rect 536748 500890 536800 500896
rect 536760 477018 536788 500890
rect 537312 500002 537340 502846
rect 538094 502602 538122 502860
rect 539212 502846 539548 502874
rect 540316 502846 540928 502874
rect 541328 502846 541664 502874
rect 542432 502846 542768 502874
rect 543536 502846 543688 502874
rect 544548 502846 544884 502874
rect 545652 502846 545988 502874
rect 546756 502846 547092 502874
rect 547860 502846 548196 502874
rect 548872 502846 549116 502874
rect 549976 502846 550588 502874
rect 551080 502846 551232 502874
rect 538048 502574 538122 502602
rect 537300 499996 537352 500002
rect 537300 499938 537352 499944
rect 536748 477012 536800 477018
rect 536748 476954 536800 476960
rect 535368 476944 535420 476950
rect 535368 476886 535420 476892
rect 538048 475590 538076 502574
rect 538128 499996 538180 500002
rect 538128 499938 538180 499944
rect 538036 475584 538088 475590
rect 538036 475526 538088 475532
rect 538140 474366 538168 499938
rect 538128 474360 538180 474366
rect 538128 474302 538180 474308
rect 539520 474298 539548 502846
rect 540900 478378 540928 502846
rect 541636 500954 541664 502846
rect 541624 500948 541676 500954
rect 541624 500890 541676 500896
rect 542268 500948 542320 500954
rect 542268 500890 542320 500896
rect 542280 478446 542308 500890
rect 542740 500750 542768 502846
rect 542728 500744 542780 500750
rect 542728 500686 542780 500692
rect 542268 478440 542320 478446
rect 542268 478382 542320 478388
rect 540888 478372 540940 478378
rect 540888 478314 540940 478320
rect 543660 475658 543688 502846
rect 544856 500682 544884 502846
rect 545960 500954 545988 502846
rect 547064 500954 547092 502846
rect 545948 500948 546000 500954
rect 545948 500890 546000 500896
rect 546408 500948 546460 500954
rect 546408 500890 546460 500896
rect 547052 500948 547104 500954
rect 547052 500890 547104 500896
rect 547788 500948 547840 500954
rect 547788 500890 547840 500896
rect 544844 500676 544896 500682
rect 544844 500618 544896 500624
rect 546420 477086 546448 500890
rect 546408 477080 546460 477086
rect 546408 477022 546460 477028
rect 543648 475652 543700 475658
rect 543648 475594 543700 475600
rect 539508 474292 539560 474298
rect 539508 474234 539560 474240
rect 533988 474224 534040 474230
rect 533988 474166 534040 474172
rect 518808 474156 518860 474162
rect 518808 474098 518860 474104
rect 512644 474088 512696 474094
rect 512644 474030 512696 474036
rect 502248 474020 502300 474026
rect 502248 473962 502300 473968
rect 546590 473512 546646 473521
rect 547800 473482 547828 500890
rect 548168 500546 548196 502846
rect 548156 500540 548208 500546
rect 548156 500482 548208 500488
rect 549088 499798 549116 502846
rect 549168 500540 549220 500546
rect 549168 500482 549220 500488
rect 549076 499792 549128 499798
rect 549076 499734 549128 499740
rect 549180 475726 549208 500482
rect 549904 500200 549956 500206
rect 549904 500142 549956 500148
rect 549168 475720 549220 475726
rect 549168 475662 549220 475668
rect 549916 474570 549944 500142
rect 550560 475862 550588 502846
rect 551204 481250 551232 502846
rect 552078 502602 552106 502860
rect 553196 502846 553348 502874
rect 554300 502846 554728 502874
rect 555404 502846 555556 502874
rect 552032 502574 552106 502602
rect 551376 500744 551428 500750
rect 551376 500686 551428 500692
rect 551284 499792 551336 499798
rect 551284 499734 551336 499740
rect 550928 481222 551232 481250
rect 550548 475856 550600 475862
rect 550548 475798 550600 475804
rect 550928 474638 550956 481222
rect 551008 480956 551060 480962
rect 551008 480898 551060 480904
rect 550916 474632 550968 474638
rect 550916 474574 550968 474580
rect 549904 474564 549956 474570
rect 549904 474506 549956 474512
rect 551020 473482 551048 480898
rect 551192 478236 551244 478242
rect 551192 478178 551244 478184
rect 551204 473550 551232 478178
rect 551192 473544 551244 473550
rect 551192 473486 551244 473492
rect 546590 473447 546592 473456
rect 546644 473447 546646 473456
rect 547788 473476 547840 473482
rect 546592 473418 546644 473424
rect 547788 473418 547840 473424
rect 551008 473476 551060 473482
rect 551008 473418 551060 473424
rect 443642 450664 443698 450673
rect 443642 450599 443698 450608
rect 551296 441674 551324 499734
rect 551388 445210 551416 500686
rect 551468 500472 551520 500478
rect 551468 500414 551520 500420
rect 551480 499526 551508 500414
rect 551560 500404 551612 500410
rect 551560 500346 551612 500352
rect 551468 499520 551520 499526
rect 551468 499462 551520 499468
rect 551468 489932 551520 489938
rect 551468 489874 551520 489880
rect 551480 480962 551508 489874
rect 551468 480956 551520 480962
rect 551468 480898 551520 480904
rect 551468 473476 551520 473482
rect 551468 473418 551520 473424
rect 551480 471782 551508 473418
rect 551468 471776 551520 471782
rect 551468 471718 551520 471724
rect 551572 468466 551600 500346
rect 551652 500336 551704 500342
rect 551652 500278 551704 500284
rect 551664 471918 551692 500278
rect 551744 500268 551796 500274
rect 551744 500210 551796 500216
rect 551652 471912 551704 471918
rect 551652 471854 551704 471860
rect 551756 471442 551784 500210
rect 551836 499520 551888 499526
rect 551836 499462 551888 499468
rect 551848 489938 551876 499462
rect 551836 489932 551888 489938
rect 551836 489874 551888 489880
rect 551836 476876 551888 476882
rect 551836 476818 551888 476824
rect 551744 471436 551796 471442
rect 551744 471378 551796 471384
rect 551572 468438 551784 468466
rect 551756 467922 551784 468438
rect 551572 467894 551784 467922
rect 551572 461428 551600 467894
rect 551652 467492 551704 467498
rect 551652 467434 551704 467440
rect 551664 463434 551692 467434
rect 551744 467356 551796 467362
rect 551744 467298 551796 467304
rect 551756 463622 551784 467298
rect 551744 463616 551796 463622
rect 551744 463558 551796 463564
rect 551664 463418 551784 463434
rect 551664 463412 551796 463418
rect 551664 463406 551744 463412
rect 551744 463354 551796 463360
rect 551744 461440 551796 461446
rect 551572 461400 551744 461428
rect 551744 461382 551796 461388
rect 551848 455326 551876 476818
rect 551928 474700 551980 474706
rect 551928 474642 551980 474648
rect 551940 473929 551968 474642
rect 551926 473920 551982 473929
rect 551926 473855 551982 473864
rect 551928 473544 551980 473550
rect 551928 473486 551980 473492
rect 551940 456550 551968 473486
rect 551928 456544 551980 456550
rect 551928 456486 551980 456492
rect 551836 455320 551888 455326
rect 551836 455262 551888 455268
rect 552032 446434 552060 502574
rect 553320 500954 553348 502846
rect 553308 500948 553360 500954
rect 553308 500890 553360 500896
rect 554044 500948 554096 500954
rect 554044 500890 554096 500896
rect 553308 497480 553360 497486
rect 553308 497422 553360 497428
rect 553216 494760 553268 494766
rect 553216 494702 553268 494708
rect 553124 493332 553176 493338
rect 553124 493274 553176 493280
rect 552664 483744 552716 483750
rect 552664 483686 552716 483692
rect 552388 482316 552440 482322
rect 552388 482258 552440 482264
rect 552112 476808 552164 476814
rect 552112 476750 552164 476756
rect 552124 473113 552152 476750
rect 552296 474360 552348 474366
rect 552296 474302 552348 474308
rect 552204 474156 552256 474162
rect 552204 474098 552256 474104
rect 552110 473104 552166 473113
rect 552110 473039 552166 473048
rect 552112 471436 552164 471442
rect 552112 471378 552164 471384
rect 552124 467265 552152 471378
rect 552110 467256 552166 467265
rect 552110 467191 552166 467200
rect 552216 467106 552244 474098
rect 552308 471442 552336 474302
rect 552296 471436 552348 471442
rect 552296 471378 552348 471384
rect 552294 471336 552350 471345
rect 552294 471271 552350 471280
rect 552124 467078 552244 467106
rect 552124 458969 552152 467078
rect 552204 467016 552256 467022
rect 552204 466958 552256 466964
rect 552110 458960 552166 458969
rect 552110 458895 552166 458904
rect 552112 456544 552164 456550
rect 552110 456512 552112 456521
rect 552164 456512 552166 456521
rect 552110 456447 552166 456456
rect 552112 455320 552164 455326
rect 552110 455288 552112 455297
rect 552164 455288 552166 455297
rect 552110 455223 552166 455232
rect 552216 448225 552244 466958
rect 552308 448769 552336 471271
rect 552400 453529 552428 482258
rect 552480 479664 552532 479670
rect 552480 479606 552532 479612
rect 552492 471442 552520 479606
rect 552572 477012 552624 477018
rect 552572 476954 552624 476960
rect 552480 471436 552532 471442
rect 552480 471378 552532 471384
rect 552584 471345 552612 476954
rect 552570 471336 552626 471345
rect 552570 471271 552626 471280
rect 552480 471232 552532 471238
rect 552480 471174 552532 471180
rect 552572 471232 552624 471238
rect 552572 471174 552624 471180
rect 552492 467022 552520 471174
rect 552480 467016 552532 467022
rect 552480 466958 552532 466964
rect 552480 466880 552532 466886
rect 552480 466822 552532 466828
rect 552386 453520 552442 453529
rect 552386 453455 552442 453464
rect 552492 450673 552520 466822
rect 552584 451217 552612 471174
rect 552676 459626 552704 483686
rect 553032 480820 553084 480826
rect 553032 480762 553084 480768
rect 552848 478304 552900 478310
rect 552848 478246 552900 478252
rect 552756 474224 552808 474230
rect 552756 474166 552808 474172
rect 552768 471578 552796 474166
rect 552756 471572 552808 471578
rect 552756 471514 552808 471520
rect 552756 471436 552808 471442
rect 552756 471378 552808 471384
rect 552768 471050 552796 471378
rect 552860 471238 552888 478246
rect 552940 475448 552992 475454
rect 552940 475390 552992 475396
rect 552952 471578 552980 475390
rect 552940 471572 552992 471578
rect 552940 471514 552992 471520
rect 552940 471436 552992 471442
rect 552940 471378 552992 471384
rect 552848 471232 552900 471238
rect 552848 471174 552900 471180
rect 552768 471022 552888 471050
rect 552756 470960 552808 470966
rect 552756 470902 552808 470908
rect 552768 466886 552796 470902
rect 552756 466880 552808 466886
rect 552756 466822 552808 466828
rect 552756 466744 552808 466750
rect 552756 466686 552808 466692
rect 552768 459746 552796 466686
rect 552860 461854 552888 471022
rect 552952 468625 552980 471378
rect 552938 468616 552994 468625
rect 552938 468551 552994 468560
rect 552940 468512 552992 468518
rect 552940 468454 552992 468460
rect 552848 461848 552900 461854
rect 552848 461790 552900 461796
rect 552952 461786 552980 468454
rect 553044 463706 553072 480762
rect 553136 471306 553164 493274
rect 553124 471300 553176 471306
rect 553124 471242 553176 471248
rect 553124 471164 553176 471170
rect 553124 471106 553176 471112
rect 553136 466750 553164 471106
rect 553124 466744 553176 466750
rect 553124 466686 553176 466692
rect 553228 466313 553256 494702
rect 553320 471442 553348 497422
rect 553676 478440 553728 478446
rect 553676 478382 553728 478388
rect 553584 477080 553636 477086
rect 553584 477022 553636 477028
rect 553400 475856 553452 475862
rect 553400 475798 553452 475804
rect 553308 471436 553360 471442
rect 553308 471378 553360 471384
rect 553308 471300 553360 471306
rect 553308 471242 553360 471248
rect 553214 466304 553270 466313
rect 553214 466239 553270 466248
rect 553044 463678 553164 463706
rect 553032 463616 553084 463622
rect 553030 463584 553032 463593
rect 553084 463584 553086 463593
rect 553030 463519 553086 463528
rect 553032 463412 553084 463418
rect 553032 463354 553084 463360
rect 552940 461780 552992 461786
rect 552940 461722 552992 461728
rect 552848 461440 552900 461446
rect 552848 461382 552900 461388
rect 552940 461440 552992 461446
rect 552940 461382 552992 461388
rect 552860 461009 552888 461382
rect 552846 461000 552902 461009
rect 552846 460935 552902 460944
rect 552756 459740 552808 459746
rect 552756 459682 552808 459688
rect 552676 459598 552888 459626
rect 552756 459536 552808 459542
rect 552756 459478 552808 459484
rect 552768 452985 552796 459478
rect 552860 456793 552888 459598
rect 552846 456784 552902 456793
rect 552846 456719 552902 456728
rect 552754 452976 552810 452985
rect 552754 452911 552810 452920
rect 552570 451208 552626 451217
rect 552570 451143 552626 451152
rect 552478 450664 552534 450673
rect 552478 450599 552534 450608
rect 552294 448760 552350 448769
rect 552294 448695 552350 448704
rect 552202 448216 552258 448225
rect 552202 448151 552258 448160
rect 552032 446406 552244 446434
rect 552018 445224 552074 445233
rect 551388 445182 552018 445210
rect 552018 445159 552074 445168
rect 552018 441688 552074 441697
rect 551296 441646 552018 441674
rect 552018 441623 552074 441632
rect 552216 439929 552244 446406
rect 552952 442513 552980 461382
rect 553044 459785 553072 463354
rect 553030 459776 553086 459785
rect 553030 459711 553086 459720
rect 553136 459241 553164 463678
rect 553320 462777 553348 471242
rect 553306 462768 553362 462777
rect 553306 462703 553362 462712
rect 553216 461848 553268 461854
rect 553216 461790 553268 461796
rect 553122 459232 553178 459241
rect 553122 459167 553178 459176
rect 553228 454481 553256 461790
rect 553214 454472 553270 454481
rect 553214 454407 553270 454416
rect 552938 442504 552994 442513
rect 552938 442439 552994 442448
rect 553412 440745 553440 475798
rect 553492 474632 553544 474638
rect 553492 474574 553544 474580
rect 553398 440736 553454 440745
rect 553398 440671 553454 440680
rect 553504 440201 553532 474574
rect 553596 443193 553624 477022
rect 553688 445505 553716 478382
rect 553768 475720 553820 475726
rect 553768 475662 553820 475668
rect 553674 445496 553730 445505
rect 553674 445431 553730 445440
rect 553582 443184 553638 443193
rect 553582 443119 553638 443128
rect 553780 441969 553808 475662
rect 553860 475652 553912 475658
rect 553860 475594 553912 475600
rect 553872 444417 553900 475594
rect 553952 474292 554004 474298
rect 553952 474234 554004 474240
rect 553964 446729 553992 474234
rect 554056 459610 554084 500890
rect 554136 500812 554188 500818
rect 554136 500754 554188 500760
rect 554148 467634 554176 500754
rect 554228 500608 554280 500614
rect 554228 500550 554280 500556
rect 554240 470422 554268 500550
rect 554596 481024 554648 481030
rect 554596 480966 554648 480972
rect 554504 479596 554556 479602
rect 554504 479538 554556 479544
rect 554320 476944 554372 476950
rect 554320 476886 554372 476892
rect 554228 470416 554280 470422
rect 554228 470358 554280 470364
rect 554136 467628 554188 467634
rect 554136 467570 554188 467576
rect 554044 459604 554096 459610
rect 554044 459546 554096 459552
rect 554332 449041 554360 476886
rect 554412 475516 554464 475522
rect 554412 475458 554464 475464
rect 554424 451489 554452 475458
rect 554516 453801 554544 479538
rect 554608 457337 554636 480966
rect 554700 465050 554728 502846
rect 555240 486464 555292 486470
rect 555240 486406 555292 486412
rect 555148 483676 555200 483682
rect 555148 483618 555200 483624
rect 554780 479528 554832 479534
rect 554780 479470 554832 479476
rect 554792 472161 554820 479470
rect 555056 475584 555108 475590
rect 555056 475526 555108 475532
rect 554964 474020 555016 474026
rect 554964 473962 555016 473968
rect 554778 472152 554834 472161
rect 554778 472087 554834 472096
rect 554780 472048 554832 472054
rect 554780 471990 554832 471996
rect 554688 465044 554740 465050
rect 554688 464986 554740 464992
rect 554792 463865 554820 471990
rect 554976 467537 555004 473962
rect 554962 467528 555018 467537
rect 554962 467463 555018 467472
rect 554778 463856 554834 463865
rect 554778 463791 554834 463800
rect 554964 459604 555016 459610
rect 554964 459546 555016 459552
rect 554594 457328 554650 457337
rect 554594 457263 554650 457272
rect 554502 453792 554558 453801
rect 554502 453727 554558 453736
rect 554410 451480 554466 451489
rect 554410 451415 554466 451424
rect 554318 449032 554374 449041
rect 554318 448967 554374 448976
rect 553950 446720 554006 446729
rect 553950 446655 554006 446664
rect 553858 444408 553914 444417
rect 553858 444343 553914 444352
rect 553766 441960 553822 441969
rect 553766 441895 553822 441904
rect 553490 440192 553546 440201
rect 553490 440127 553546 440136
rect 552202 439920 552258 439929
rect 552202 439855 552258 439864
rect 554976 438977 555004 459546
rect 555068 447273 555096 475526
rect 555160 462097 555188 483618
rect 555252 465633 555280 486406
rect 555424 475380 555476 475386
rect 555424 475322 555476 475328
rect 555332 474564 555384 474570
rect 555332 474506 555384 474512
rect 555238 465624 555294 465633
rect 555238 465559 555294 465568
rect 555146 462088 555202 462097
rect 555146 462023 555202 462032
rect 555344 455569 555372 474506
rect 555436 458017 555464 475322
rect 555422 458008 555478 458017
rect 555422 457943 555478 457952
rect 555330 455560 555386 455569
rect 555330 455495 555386 455504
rect 555054 447264 555110 447273
rect 555054 447199 555110 447208
rect 554962 438968 555018 438977
rect 554962 438903 555018 438912
rect 555528 437889 555556 502846
rect 556172 502846 556416 502874
rect 557520 502846 557672 502874
rect 555700 491972 555752 491978
rect 555700 491914 555752 491920
rect 555608 478372 555660 478378
rect 555608 478314 555660 478320
rect 555620 446185 555648 478314
rect 555712 471073 555740 491914
rect 555976 490612 556028 490618
rect 555976 490554 556028 490560
rect 555792 481092 555844 481098
rect 555792 481034 555844 481040
rect 555698 471064 555754 471073
rect 555698 470999 555754 471008
rect 555700 470416 555752 470422
rect 555700 470358 555752 470364
rect 555712 449721 555740 470358
rect 555804 452033 555832 481034
rect 555884 478168 555936 478174
rect 555884 478110 555936 478116
rect 555896 470393 555924 478110
rect 555882 470384 555938 470393
rect 555882 470319 555938 470328
rect 555988 469305 556016 490554
rect 556068 474088 556120 474094
rect 556068 474030 556120 474036
rect 555974 469296 556030 469305
rect 555974 469231 556030 469240
rect 555976 467628 556028 467634
rect 555976 467570 556028 467576
rect 555884 465044 555936 465050
rect 555884 464986 555936 464992
rect 555790 452024 555846 452033
rect 555790 451959 555846 451968
rect 555698 449712 555754 449721
rect 555698 449647 555754 449656
rect 555606 446176 555662 446185
rect 555606 446111 555662 446120
rect 555896 438433 555924 464986
rect 555988 443737 556016 467570
rect 556080 465089 556108 474030
rect 556066 465080 556122 465089
rect 556066 465015 556122 465024
rect 555974 443728 556030 443737
rect 555974 443663 556030 443672
rect 555882 438424 555938 438433
rect 555882 438359 555938 438368
rect 555514 437880 555570 437889
rect 555514 437815 555570 437824
rect 554964 437368 555016 437374
rect 554964 437310 555016 437316
rect 554780 437164 554832 437170
rect 554780 437106 554832 437112
rect 554792 436665 554820 437106
rect 554778 436656 554834 436665
rect 554778 436591 554834 436600
rect 554976 436121 555004 437310
rect 556066 437200 556122 437209
rect 556172 437186 556200 502846
rect 556804 500268 556856 500274
rect 556804 500210 556856 500216
rect 556122 437158 556200 437186
rect 556066 437135 556122 437144
rect 554962 436112 555018 436121
rect 554872 436076 554924 436082
rect 554962 436047 555018 436056
rect 554872 436018 554924 436024
rect 554780 436008 554832 436014
rect 554780 435950 554832 435956
rect 554792 435441 554820 435950
rect 554778 435432 554834 435441
rect 554778 435367 554834 435376
rect 554884 434897 554912 436018
rect 554870 434888 554926 434897
rect 554870 434823 554926 434832
rect 554780 434716 554832 434722
rect 554780 434658 554832 434664
rect 554792 434217 554820 434658
rect 554872 434648 554924 434654
rect 554872 434590 554924 434596
rect 554778 434208 554834 434217
rect 554778 434143 554834 434152
rect 554884 433673 554912 434590
rect 554870 433664 554926 433673
rect 554870 433599 554926 433608
rect 554872 433288 554924 433294
rect 554872 433230 554924 433236
rect 554780 433220 554832 433226
rect 554780 433162 554832 433168
rect 554792 433129 554820 433162
rect 554778 433120 554834 433129
rect 554778 433055 554834 433064
rect 554884 432449 554912 433230
rect 554870 432440 554926 432449
rect 554870 432375 554926 432384
rect 554964 431928 555016 431934
rect 554778 431896 554834 431905
rect 554964 431870 555016 431876
rect 554778 431831 554780 431840
rect 554832 431831 554834 431840
rect 554780 431802 554832 431808
rect 554872 431792 554924 431798
rect 554872 431734 554924 431740
rect 554884 431361 554912 431734
rect 554870 431352 554926 431361
rect 554870 431287 554926 431296
rect 554976 430681 555004 431870
rect 554962 430672 555018 430681
rect 554962 430607 555018 430616
rect 554872 430568 554924 430574
rect 554872 430510 554924 430516
rect 554780 430500 554832 430506
rect 554780 430442 554832 430448
rect 554792 430137 554820 430442
rect 554778 430128 554834 430137
rect 554778 430063 554834 430072
rect 554884 429593 554912 430510
rect 554870 429584 554926 429593
rect 554870 429519 554926 429528
rect 554780 429140 554832 429146
rect 554780 429082 554832 429088
rect 554792 428369 554820 429082
rect 556816 428942 556844 500210
rect 557644 437170 557672 502846
rect 557736 502846 558624 502874
rect 559300 502846 559636 502874
rect 560312 502846 560740 502874
rect 561692 502846 561844 502874
rect 561968 502846 562948 502874
rect 563072 502846 563960 502874
rect 564452 502846 565064 502874
rect 565832 502846 566168 502874
rect 567180 502846 567240 502874
rect 557736 437374 557764 502846
rect 559300 500954 559328 502846
rect 558184 500948 558236 500954
rect 558184 500890 558236 500896
rect 559288 500948 559340 500954
rect 559288 500890 559340 500896
rect 557724 437368 557776 437374
rect 557724 437310 557776 437316
rect 557632 437164 557684 437170
rect 557632 437106 557684 437112
rect 558196 436014 558224 500890
rect 560312 436082 560340 502846
rect 560944 499588 560996 499594
rect 560944 499530 560996 499536
rect 560300 436076 560352 436082
rect 560300 436018 560352 436024
rect 558184 436008 558236 436014
rect 558184 435950 558236 435956
rect 560956 431798 560984 499530
rect 561692 434722 561720 502846
rect 561680 434716 561732 434722
rect 561680 434658 561732 434664
rect 561968 434654 561996 502846
rect 561956 434648 562008 434654
rect 561956 434590 562008 434596
rect 563072 433226 563100 502846
rect 563704 462392 563756 462398
rect 563704 462334 563756 462340
rect 563060 433220 563112 433226
rect 563060 433162 563112 433168
rect 560944 431792 560996 431798
rect 560944 431734 560996 431740
rect 554872 428936 554924 428942
rect 554870 428904 554872 428913
rect 556804 428936 556856 428942
rect 554924 428904 554926 428913
rect 556804 428878 556856 428884
rect 554870 428839 554926 428848
rect 554778 428360 554834 428369
rect 554778 428295 554834 428304
rect 554778 427816 554834 427825
rect 554778 427751 554780 427760
rect 554832 427751 554834 427760
rect 554780 427722 554832 427728
rect 499316 426426 499344 427516
rect 499304 426420 499356 426426
rect 499304 426362 499356 426368
rect 563716 325650 563744 462334
rect 564452 433294 564480 502846
rect 564440 433288 564492 433294
rect 564440 433230 564492 433236
rect 565832 431866 565860 502846
rect 567212 499594 567240 502846
rect 567304 502846 568284 502874
rect 568592 502846 569388 502874
rect 569972 502846 570492 502874
rect 571352 502846 571504 502874
rect 571628 502846 572608 502874
rect 572732 502846 573712 502874
rect 574112 502846 574724 502874
rect 567200 499588 567252 499594
rect 567200 499530 567252 499536
rect 567304 431934 567332 502846
rect 567292 431928 567344 431934
rect 567292 431870 567344 431876
rect 565820 431860 565872 431866
rect 565820 431802 565872 431808
rect 568592 430506 568620 502846
rect 569972 430574 570000 502846
rect 571352 500274 571380 502846
rect 571340 500268 571392 500274
rect 571340 500210 571392 500216
rect 569960 430568 570012 430574
rect 569960 430510 570012 430516
rect 568580 430500 568632 430506
rect 568580 430442 568632 430448
rect 571628 429146 571656 502846
rect 571616 429140 571668 429146
rect 571616 429082 571668 429088
rect 572732 427786 572760 502846
rect 574112 498846 574140 502846
rect 574100 498840 574152 498846
rect 574100 498782 574152 498788
rect 572720 427780 572772 427786
rect 572720 427722 572772 427728
rect 563704 325644 563756 325650
rect 563704 325586 563756 325592
rect 560944 306400 560996 306406
rect 560944 306342 560996 306348
rect 413284 83564 413336 83570
rect 413284 83506 413336 83512
rect 487620 62824 487672 62830
rect 487620 62766 487672 62772
rect 487632 60860 487660 62766
rect 411902 49872 411958 49881
rect 411902 49807 411958 49816
rect 232240 48334 232360 48362
rect 227626 46064 227682 46073
rect 227626 45999 227682 46008
rect 227442 44704 227498 44713
rect 227442 44639 227498 44648
rect 227444 44260 227496 44266
rect 227444 44202 227496 44208
rect 226432 42774 226484 42780
rect 227258 42800 227314 42809
rect 226340 41472 226392 41478
rect 226340 41414 226392 41420
rect 226352 40225 226380 41414
rect 226444 40769 226472 42774
rect 227258 42735 227314 42744
rect 227456 42129 227484 44202
rect 227536 44192 227588 44198
rect 227536 44134 227588 44140
rect 227442 42120 227498 42129
rect 227442 42055 227498 42064
rect 226616 41540 226668 41546
rect 226616 41482 226668 41488
rect 226430 40760 226486 40769
rect 226430 40695 226486 40704
rect 226338 40216 226394 40225
rect 226338 40151 226394 40160
rect 226628 39545 226656 41482
rect 227548 41449 227576 44134
rect 227534 41440 227590 41449
rect 227534 41375 227590 41384
rect 232240 41290 232268 48334
rect 560956 41410 560984 306342
rect 576136 95198 576164 696934
rect 580262 686352 580318 686361
rect 580262 686287 580318 686296
rect 579618 651128 579674 651137
rect 579618 651063 579674 651072
rect 579632 650078 579660 651063
rect 577504 650072 577556 650078
rect 577504 650014 577556 650020
rect 579620 650072 579672 650078
rect 579620 650014 579672 650020
rect 576216 579692 576268 579698
rect 576216 579634 576268 579640
rect 576124 95192 576176 95198
rect 576124 95134 576176 95140
rect 576228 62830 576256 579634
rect 577516 93770 577544 650014
rect 578882 604208 578938 604217
rect 578882 604143 578938 604152
rect 577596 509652 577648 509658
rect 577596 509594 577648 509600
rect 577608 327078 577636 509594
rect 577596 327072 577648 327078
rect 577596 327014 577648 327020
rect 578896 93838 578924 604143
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 579698 580212 580751
rect 580172 579692 580224 579698
rect 580172 579634 580224 579640
rect 580170 557288 580226 557297
rect 580170 557223 580226 557232
rect 580184 556238 580212 557223
rect 580172 556232 580224 556238
rect 580172 556174 580224 556180
rect 579618 510368 579674 510377
rect 579618 510303 579674 510312
rect 579632 509658 579660 510303
rect 579620 509652 579672 509658
rect 579620 509594 579672 509600
rect 580170 463448 580226 463457
rect 580170 463383 580226 463392
rect 580184 462398 580212 463383
rect 580172 462392 580224 462398
rect 580172 462334 580224 462340
rect 580170 416528 580226 416537
rect 580170 416463 580226 416472
rect 580184 415478 580212 416463
rect 580172 415472 580224 415478
rect 580172 415414 580224 415420
rect 580170 369608 580226 369617
rect 580170 369543 580226 369552
rect 580184 368558 580212 369543
rect 580172 368552 580224 368558
rect 580172 368494 580224 368500
rect 580170 322688 580226 322697
rect 580170 322623 580226 322632
rect 580184 321638 580212 322623
rect 580172 321632 580224 321638
rect 580172 321574 580224 321580
rect 580172 276004 580224 276010
rect 580172 275946 580224 275952
rect 580184 275777 580212 275946
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 579988 229084 580040 229090
rect 579988 229026 580040 229032
rect 580000 228857 580028 229026
rect 579986 228848 580042 228857
rect 579986 228783 580042 228792
rect 579988 182164 580040 182170
rect 579988 182106 580040 182112
rect 580000 181937 580028 182106
rect 579986 181928 580042 181937
rect 579986 181863 580042 181872
rect 580172 135244 580224 135250
rect 580172 135186 580224 135192
rect 580184 134881 580212 135186
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 578884 93832 578936 93838
rect 578884 93774 578936 93780
rect 577504 93764 577556 93770
rect 577504 93706 577556 93712
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 87961 580212 88266
rect 580170 87952 580226 87961
rect 580170 87887 580226 87896
rect 580276 83502 580304 686287
rect 580354 639432 580410 639441
rect 580354 639367 580410 639376
rect 580368 502994 580396 639367
rect 580446 592512 580502 592521
rect 580446 592447 580502 592456
rect 580460 569226 580488 592447
rect 580448 569220 580500 569226
rect 580448 569162 580500 569168
rect 580906 545592 580962 545601
rect 580906 545527 580962 545536
rect 580356 502988 580408 502994
rect 580356 502930 580408 502936
rect 580920 498681 580948 545527
rect 580906 498672 580962 498681
rect 580906 498607 580962 498616
rect 580920 451761 580948 498607
rect 580906 451752 580962 451761
rect 580906 451687 580962 451696
rect 580920 404841 580948 451687
rect 580906 404832 580962 404841
rect 580906 404767 580962 404776
rect 580920 357921 580948 404767
rect 580906 357912 580962 357921
rect 580906 357847 580962 357856
rect 580920 310865 580948 357847
rect 580354 310856 580410 310865
rect 580354 310791 580410 310800
rect 580906 310856 580962 310865
rect 580906 310791 580962 310800
rect 580368 303618 580396 310791
rect 580356 303612 580408 303618
rect 580356 303554 580408 303560
rect 580368 263945 580396 303554
rect 580354 263936 580410 263945
rect 580354 263871 580410 263880
rect 580906 263936 580962 263945
rect 580906 263871 580962 263880
rect 580920 217025 580948 263871
rect 580906 217016 580962 217025
rect 580906 216951 580962 216960
rect 580920 170105 580948 216951
rect 580906 170096 580962 170105
rect 580906 170031 580962 170040
rect 580920 123185 580948 170031
rect 580906 123176 580962 123185
rect 580906 123111 580962 123120
rect 580264 83496 580316 83502
rect 580264 83438 580316 83444
rect 580920 76265 580948 123111
rect 580906 76256 580962 76265
rect 580906 76191 580962 76200
rect 576216 62824 576268 62830
rect 576216 62766 576268 62772
rect 560944 41404 560996 41410
rect 560944 41346 560996 41352
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 232240 41262 232360 41290
rect 227444 40180 227496 40186
rect 227444 40122 227496 40128
rect 227076 40112 227128 40118
rect 227076 40054 227128 40060
rect 226614 39536 226670 39545
rect 226614 39471 226670 39480
rect 227088 38865 227116 40054
rect 227074 38856 227130 38865
rect 227074 38791 227130 38800
rect 226708 38684 226760 38690
rect 226708 38626 226760 38632
rect 226720 37641 226748 38626
rect 227456 38185 227484 40122
rect 227536 38752 227588 38758
rect 227536 38694 227588 38700
rect 227442 38176 227498 38185
rect 227442 38111 227498 38120
rect 226706 37632 226762 37641
rect 226706 37567 226762 37576
rect 227444 37324 227496 37330
rect 227444 37266 227496 37272
rect 227456 36281 227484 37266
rect 227548 36961 227576 38694
rect 232332 38570 232360 41262
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 563702 38720 563758 38729
rect 563702 38655 563758 38664
rect 231964 38542 232360 38570
rect 227534 36952 227590 36961
rect 227534 36887 227590 36896
rect 227442 36272 227498 36281
rect 227442 36207 227498 36216
rect 226708 36032 226760 36038
rect 226708 35974 226760 35980
rect 226720 35601 226748 35974
rect 227444 35964 227496 35970
rect 227444 35906 227496 35912
rect 226706 35592 226762 35601
rect 226706 35527 226762 35536
rect 227456 34921 227484 35906
rect 227442 34912 227498 34921
rect 227442 34847 227498 34856
rect 227352 34604 227404 34610
rect 227352 34546 227404 34552
rect 227364 33697 227392 34546
rect 227444 34536 227496 34542
rect 227444 34478 227496 34484
rect 227456 34377 227484 34478
rect 227442 34368 227498 34377
rect 227442 34303 227498 34312
rect 227350 33688 227406 33697
rect 227350 33623 227406 33632
rect 227444 33244 227496 33250
rect 227444 33186 227496 33192
rect 227456 33017 227484 33186
rect 227536 33176 227588 33182
rect 227536 33118 227588 33124
rect 227442 33008 227498 33017
rect 227442 32943 227498 32952
rect 213920 32564 213972 32570
rect 213920 32506 213972 32512
rect 215944 32564 215996 32570
rect 215944 32506 215996 32512
rect 95148 32428 95200 32434
rect 95148 32370 95200 32376
rect 116400 32428 116452 32434
rect 116400 32370 116452 32376
rect 95160 31929 95188 32370
rect 116398 32056 116454 32065
rect 116398 31991 116454 32000
rect 95146 31920 95202 31929
rect 95146 31855 95202 31864
rect 116412 31822 116440 31991
rect 71688 31816 71740 31822
rect 32310 31784 32366 31793
rect 71346 31764 71688 31770
rect 71346 31758 71740 31764
rect 116400 31816 116452 31822
rect 213932 31793 213960 32506
rect 215114 32464 215170 32473
rect 215114 32399 215116 32408
rect 215168 32399 215170 32408
rect 227444 32428 227496 32434
rect 215116 32370 215168 32376
rect 227444 32370 227496 32376
rect 227456 31793 227484 32370
rect 227548 32337 227576 33118
rect 227534 32328 227590 32337
rect 227534 32263 227590 32272
rect 116400 31758 116452 31764
rect 213918 31784 213974 31793
rect 71346 31742 71728 31758
rect 32310 31719 32366 31728
rect 213918 31719 213974 31728
rect 227442 31784 227498 31793
rect 227442 31719 227498 31728
rect 29932 31346 29960 31484
rect 32324 31346 32352 31719
rect 159100 31606 159850 31634
rect 161676 31606 162518 31634
rect 178236 31606 178986 31634
rect 179892 31606 180734 31634
rect 182560 31606 183310 31634
rect 208688 31606 209346 31634
rect 29920 31340 29972 31346
rect 29920 31282 29972 31288
rect 32312 31340 32364 31346
rect 32312 31282 32364 31288
rect 105544 30320 105596 30326
rect 120000 30297 120028 31484
rect 120092 31470 120842 31498
rect 105544 30262 105596 30268
rect 119986 30288 120042 30297
rect 95884 30252 95936 30258
rect 95884 30194 95936 30200
rect 50344 30184 50396 30190
rect 50344 30126 50396 30132
rect 31024 29912 31076 29918
rect 31024 29854 31076 29860
rect 25504 29776 25556 29782
rect 25504 29718 25556 29724
rect 10324 28280 10376 28286
rect 10324 28222 10376 28228
rect 10336 3738 10364 28222
rect 11704 25560 11756 25566
rect 11704 25502 11756 25508
rect 10416 10328 10468 10334
rect 10416 10270 10468 10276
rect 10324 3732 10376 3738
rect 10324 3674 10376 3680
rect 10048 3664 10100 3670
rect 10048 3606 10100 3612
rect 9128 3460 9180 3466
rect 9128 3402 9180 3408
rect 10060 480 10088 3606
rect 10428 3534 10456 10270
rect 11244 3800 11296 3806
rect 11244 3742 11296 3748
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 11256 480 11284 3742
rect 11716 3398 11744 25502
rect 13728 14476 13780 14482
rect 13728 14418 13780 14424
rect 12438 4856 12494 4865
rect 12438 4791 12494 4800
rect 11704 3392 11756 3398
rect 11704 3334 11756 3340
rect 12452 480 12480 4791
rect 13740 3482 13768 14418
rect 18328 8968 18380 8974
rect 18328 8910 18380 8916
rect 17224 4888 17276 4894
rect 17224 4830 17276 4836
rect 14832 3732 14884 3738
rect 14832 3674 14884 3680
rect 13648 3454 13768 3482
rect 13648 480 13676 3454
rect 14844 480 14872 3674
rect 16028 3324 16080 3330
rect 16028 3266 16080 3272
rect 16040 480 16068 3266
rect 17236 480 17264 4830
rect 18340 480 18368 8910
rect 21916 4820 21968 4826
rect 21916 4762 21968 4768
rect 19524 4072 19576 4078
rect 19524 4014 19576 4020
rect 19536 480 19564 4014
rect 20720 3256 20772 3262
rect 20720 3198 20772 3204
rect 20732 480 20760 3198
rect 21928 480 21956 4762
rect 25516 3670 25544 29718
rect 28264 29640 28316 29646
rect 28264 29582 28316 29588
rect 26700 4956 26752 4962
rect 26700 4898 26752 4904
rect 25504 3664 25556 3670
rect 25504 3606 25556 3612
rect 24308 3528 24360 3534
rect 24308 3470 24360 3476
rect 23112 3460 23164 3466
rect 23112 3402 23164 3408
rect 23124 480 23152 3402
rect 24320 480 24348 3470
rect 25502 3360 25558 3369
rect 25502 3295 25558 3304
rect 25516 480 25544 3295
rect 26712 480 26740 4898
rect 28276 3738 28304 29582
rect 30288 5024 30340 5030
rect 30288 4966 30340 4972
rect 28264 3732 28316 3738
rect 28264 3674 28316 3680
rect 29092 3732 29144 3738
rect 29092 3674 29144 3680
rect 27896 3664 27948 3670
rect 27896 3606 27948 3612
rect 27908 480 27936 3606
rect 29104 480 29132 3674
rect 30300 480 30328 4966
rect 31036 3806 31064 29854
rect 46204 29436 46256 29442
rect 46204 29378 46256 29384
rect 38568 11824 38620 11830
rect 38568 11766 38620 11772
rect 31484 7608 31536 7614
rect 31484 7550 31536 7556
rect 31024 3800 31076 3806
rect 31024 3742 31076 3748
rect 31496 480 31524 7550
rect 37372 6384 37424 6390
rect 37372 6326 37424 6332
rect 33876 6316 33928 6322
rect 33876 6258 33928 6264
rect 32680 3392 32732 3398
rect 32680 3334 32732 3340
rect 32692 480 32720 3334
rect 33888 480 33916 6258
rect 36176 3868 36228 3874
rect 36176 3810 36228 3816
rect 34980 3800 35032 3806
rect 34980 3742 35032 3748
rect 34992 480 35020 3742
rect 36188 480 36216 3810
rect 37384 480 37412 6326
rect 38580 480 38608 11766
rect 44548 6520 44600 6526
rect 44548 6462 44600 6468
rect 40960 6452 41012 6458
rect 40960 6394 41012 6400
rect 39764 3120 39816 3126
rect 39764 3062 39816 3068
rect 39776 480 39804 3062
rect 40972 480 41000 6394
rect 43352 4004 43404 4010
rect 43352 3946 43404 3952
rect 42156 3936 42208 3942
rect 42156 3878 42208 3884
rect 42168 480 42196 3878
rect 43364 480 43392 3946
rect 44560 480 44588 6462
rect 45468 4140 45520 4146
rect 45468 4082 45520 4088
rect 45480 3738 45508 4082
rect 46216 4078 46244 29378
rect 48228 15904 48280 15910
rect 48228 15846 48280 15852
rect 46848 13184 46900 13190
rect 46848 13126 46900 13132
rect 46204 4072 46256 4078
rect 46204 4014 46256 4020
rect 45468 3732 45520 3738
rect 45468 3674 45520 3680
rect 46860 3398 46888 13126
rect 46940 4072 46992 4078
rect 46940 4014 46992 4020
rect 45744 3392 45796 3398
rect 45744 3334 45796 3340
rect 46848 3392 46900 3398
rect 46848 3334 46900 3340
rect 45756 480 45784 3334
rect 46952 480 46980 4014
rect 48240 3482 48268 15846
rect 49332 6588 49384 6594
rect 49332 6530 49384 6536
rect 48148 3454 48268 3482
rect 48148 480 48176 3454
rect 49344 480 49372 6530
rect 50356 4146 50384 30126
rect 82084 30116 82136 30122
rect 82084 30058 82136 30064
rect 53104 30048 53156 30054
rect 53104 29990 53156 29996
rect 52368 24132 52420 24138
rect 52368 24074 52420 24080
rect 50344 4140 50396 4146
rect 50344 4082 50396 4088
rect 52380 3398 52408 24074
rect 51632 3392 51684 3398
rect 51632 3334 51684 3340
rect 52368 3392 52420 3398
rect 52368 3334 52420 3340
rect 52828 3392 52880 3398
rect 52828 3334 52880 3340
rect 50528 3324 50580 3330
rect 50528 3266 50580 3272
rect 50540 480 50568 3266
rect 51644 480 51672 3334
rect 52840 480 52868 3334
rect 53116 3126 53144 29990
rect 75184 29980 75236 29986
rect 75184 29922 75236 29928
rect 66904 29844 66956 29850
rect 66904 29786 66956 29792
rect 60004 29708 60056 29714
rect 60004 29650 60056 29656
rect 57244 29164 57296 29170
rect 57244 29106 57296 29112
rect 53748 18624 53800 18630
rect 53748 18566 53800 18572
rect 53760 3398 53788 18566
rect 56508 17264 56560 17270
rect 56508 17206 56560 17212
rect 56416 6656 56468 6662
rect 56416 6598 56468 6604
rect 53748 3392 53800 3398
rect 53748 3334 53800 3340
rect 54024 3392 54076 3398
rect 54024 3334 54076 3340
rect 53104 3120 53156 3126
rect 53104 3062 53156 3068
rect 54036 480 54064 3334
rect 55220 3120 55272 3126
rect 55220 3062 55272 3068
rect 55232 480 55260 3062
rect 56428 480 56456 6598
rect 56520 3126 56548 17206
rect 56508 3120 56560 3126
rect 56508 3062 56560 3068
rect 57256 3058 57284 29106
rect 59268 21412 59320 21418
rect 59268 21354 59320 21360
rect 57612 4140 57664 4146
rect 57612 4082 57664 4088
rect 57244 3052 57296 3058
rect 57244 2994 57296 3000
rect 57624 480 57652 4082
rect 59280 3330 59308 21354
rect 60016 4146 60044 29650
rect 61384 29096 61436 29102
rect 61384 29038 61436 29044
rect 60648 28348 60700 28354
rect 60648 28290 60700 28296
rect 60004 4140 60056 4146
rect 60004 4082 60056 4088
rect 60660 3330 60688 28290
rect 58808 3324 58860 3330
rect 58808 3266 58860 3272
rect 59268 3324 59320 3330
rect 59268 3266 59320 3272
rect 60004 3324 60056 3330
rect 60004 3266 60056 3272
rect 60648 3324 60700 3330
rect 60648 3266 60700 3272
rect 61200 3324 61252 3330
rect 61200 3266 61252 3272
rect 58820 480 58848 3266
rect 60016 480 60044 3266
rect 61212 480 61240 3266
rect 61396 3126 61424 29038
rect 63408 22772 63460 22778
rect 63408 22714 63460 22720
rect 61384 3120 61436 3126
rect 61384 3062 61436 3068
rect 63420 2990 63448 22714
rect 66168 19984 66220 19990
rect 66168 19926 66220 19932
rect 66180 19310 66208 19926
rect 66168 19304 66220 19310
rect 66168 19246 66220 19252
rect 65984 9716 66036 9722
rect 65984 9658 66036 9664
rect 65996 9602 66024 9658
rect 65904 9574 66024 9602
rect 63592 6724 63644 6730
rect 63592 6666 63644 6672
rect 62396 2984 62448 2990
rect 62396 2926 62448 2932
rect 63408 2984 63460 2990
rect 63408 2926 63460 2932
rect 62408 480 62436 2926
rect 63604 480 63632 6666
rect 64788 3868 64840 3874
rect 64788 3810 64840 3816
rect 64800 480 64828 3810
rect 65904 610 65932 9574
rect 66916 3874 66944 29786
rect 68008 29232 68060 29238
rect 68008 29174 68060 29180
rect 68020 28966 68048 29174
rect 68008 28960 68060 28966
rect 68008 28902 68060 28908
rect 67548 25628 67600 25634
rect 67548 25570 67600 25576
rect 67560 12510 67588 25570
rect 74448 24200 74500 24206
rect 74448 24142 74500 24148
rect 68100 19372 68152 19378
rect 68100 19314 68152 19320
rect 67548 12504 67600 12510
rect 67548 12446 67600 12452
rect 67180 9716 67232 9722
rect 67180 9658 67232 9664
rect 66904 3868 66956 3874
rect 66904 3810 66956 3816
rect 65892 604 65944 610
rect 65892 546 65944 552
rect 65984 604 66036 610
rect 65984 546 66036 552
rect 65996 480 66024 546
rect 67192 480 67220 9658
rect 68112 3194 68140 19314
rect 70676 6792 70728 6798
rect 70676 6734 70728 6740
rect 69480 5160 69532 5166
rect 69480 5102 69532 5108
rect 68284 3256 68336 3262
rect 68284 3198 68336 3204
rect 68100 3188 68152 3194
rect 68100 3130 68152 3136
rect 68296 480 68324 3198
rect 69492 480 69520 5102
rect 70688 480 70716 6734
rect 73068 5092 73120 5098
rect 73068 5034 73120 5040
rect 71872 2984 71924 2990
rect 71872 2926 71924 2932
rect 71884 480 71912 2926
rect 73080 480 73108 5034
rect 74460 3482 74488 24142
rect 74276 3454 74488 3482
rect 74276 480 74304 3454
rect 75196 2990 75224 29922
rect 77852 6860 77904 6866
rect 77852 6802 77904 6808
rect 76656 5228 76708 5234
rect 76656 5170 76708 5176
rect 75460 3052 75512 3058
rect 75460 2994 75512 3000
rect 75184 2984 75236 2990
rect 75184 2926 75236 2932
rect 75472 480 75500 2994
rect 76668 480 76696 5170
rect 77864 480 77892 6802
rect 80244 5296 80296 5302
rect 80244 5238 80296 5244
rect 79048 3120 79100 3126
rect 79048 3062 79100 3068
rect 79060 480 79088 3062
rect 80256 480 80284 5238
rect 81440 3188 81492 3194
rect 81440 3130 81492 3136
rect 81452 480 81480 3130
rect 82096 3126 82124 30058
rect 85488 22840 85540 22846
rect 85488 22782 85540 22788
rect 82728 15972 82780 15978
rect 82728 15914 82780 15920
rect 82740 3194 82768 15914
rect 83832 5364 83884 5370
rect 83832 5306 83884 5312
rect 82728 3188 82780 3194
rect 82728 3130 82780 3136
rect 82084 3120 82136 3126
rect 82084 3062 82136 3068
rect 82636 3052 82688 3058
rect 82636 2994 82688 3000
rect 82648 480 82676 2994
rect 83844 480 83872 5306
rect 85500 3126 85528 22782
rect 89628 18692 89680 18698
rect 89628 18634 89680 18640
rect 87328 5432 87380 5438
rect 87328 5374 87380 5380
rect 84936 3120 84988 3126
rect 84936 3062 84988 3068
rect 85488 3120 85540 3126
rect 85488 3062 85540 3068
rect 84948 480 84976 3062
rect 86132 2984 86184 2990
rect 86132 2926 86184 2932
rect 86144 480 86172 2926
rect 87340 480 87368 5374
rect 89640 3126 89668 18634
rect 92388 17332 92440 17338
rect 92388 17274 92440 17280
rect 90916 5500 90968 5506
rect 90916 5442 90968 5448
rect 88524 3120 88576 3126
rect 88524 3062 88576 3068
rect 89628 3120 89680 3126
rect 89628 3062 89680 3068
rect 88536 480 88564 3062
rect 89720 2848 89772 2854
rect 89720 2790 89772 2796
rect 89732 480 89760 2790
rect 90928 480 90956 5442
rect 92400 3482 92428 17274
rect 94504 4752 94556 4758
rect 94504 4694 94556 4700
rect 92124 3454 92428 3482
rect 92124 480 92152 3454
rect 93308 2984 93360 2990
rect 93308 2926 93360 2932
rect 93320 480 93348 2926
rect 94516 480 94544 4694
rect 95896 3074 95924 30194
rect 102784 29368 102836 29374
rect 102784 29310 102836 29316
rect 96528 21480 96580 21486
rect 96528 21422 96580 21428
rect 95620 3046 95924 3074
rect 95424 2848 95476 2854
rect 95620 2802 95648 3046
rect 96540 2922 96568 21422
rect 99196 20052 99248 20058
rect 99196 19994 99248 20000
rect 98092 4684 98144 4690
rect 98092 4626 98144 4632
rect 95700 2916 95752 2922
rect 95700 2858 95752 2864
rect 96528 2916 96580 2922
rect 96528 2858 96580 2864
rect 96896 2916 96948 2922
rect 96896 2858 96948 2864
rect 95476 2796 95648 2802
rect 95424 2790 95648 2796
rect 95436 2774 95648 2790
rect 95712 480 95740 2858
rect 96908 480 96936 2858
rect 98104 480 98132 4626
rect 99208 3482 99236 19994
rect 101588 4616 101640 4622
rect 101588 4558 101640 4564
rect 99208 3454 99328 3482
rect 99300 480 99328 3454
rect 100484 2848 100536 2854
rect 100484 2790 100536 2796
rect 100496 480 100524 2790
rect 101600 480 101628 4558
rect 102796 3074 102824 29310
rect 103428 28416 103480 28422
rect 103428 28358 103480 28364
rect 102704 3046 102824 3074
rect 102704 2922 102732 3046
rect 103440 2922 103468 28358
rect 105176 4480 105228 4486
rect 105176 4422 105228 4428
rect 102692 2916 102744 2922
rect 102692 2858 102744 2864
rect 102784 2916 102836 2922
rect 102784 2858 102836 2864
rect 103428 2916 103480 2922
rect 103428 2858 103480 2864
rect 103980 2916 104032 2922
rect 103980 2858 104032 2864
rect 102796 480 102824 2858
rect 103992 480 104020 2858
rect 105188 480 105216 4422
rect 105556 2922 105584 30262
rect 119986 30223 120042 30232
rect 111708 29572 111760 29578
rect 111708 29514 111760 29520
rect 110328 26920 110380 26926
rect 110328 26862 110380 26868
rect 107568 20732 107620 20738
rect 107568 20674 107620 20680
rect 107580 2922 107608 20674
rect 108764 4548 108816 4554
rect 108764 4490 108816 4496
rect 105544 2916 105596 2922
rect 105544 2858 105596 2864
rect 106372 2916 106424 2922
rect 106372 2858 106424 2864
rect 107568 2916 107620 2922
rect 107568 2858 107620 2864
rect 107660 2916 107712 2922
rect 107660 2858 107712 2864
rect 106384 480 106412 2858
rect 107672 2802 107700 2858
rect 107580 2774 107700 2802
rect 107580 480 107608 2774
rect 108776 480 108804 4490
rect 110340 3346 110368 26862
rect 109972 3318 110368 3346
rect 109972 480 110000 3318
rect 111720 2922 111748 29514
rect 115848 29504 115900 29510
rect 115848 29446 115900 29452
rect 114468 24268 114520 24274
rect 114468 24210 114520 24216
rect 112352 4412 112404 4418
rect 112352 4354 112404 4360
rect 111156 2916 111208 2922
rect 111156 2858 111208 2864
rect 111708 2916 111760 2922
rect 111708 2858 111760 2864
rect 111168 480 111196 2858
rect 112364 480 112392 4354
rect 113178 3904 113234 3913
rect 113178 3839 113180 3848
rect 113232 3839 113234 3848
rect 113180 3810 113232 3816
rect 113454 3632 113510 3641
rect 114480 3602 114508 24210
rect 115860 3602 115888 29446
rect 117964 29300 118016 29306
rect 117964 29242 118016 29248
rect 117136 18760 117188 18766
rect 117136 18702 117188 18708
rect 115940 4276 115992 4282
rect 115940 4218 115992 4224
rect 113454 3567 113456 3576
rect 113508 3567 113510 3576
rect 113548 3596 113600 3602
rect 113456 3538 113508 3544
rect 113548 3538 113600 3544
rect 114468 3596 114520 3602
rect 114468 3538 114520 3544
rect 114744 3596 114796 3602
rect 114744 3538 114796 3544
rect 115848 3596 115900 3602
rect 115848 3538 115900 3544
rect 113560 480 113588 3538
rect 114756 480 114784 3538
rect 115952 480 115980 4218
rect 116030 3632 116086 3641
rect 116030 3567 116032 3576
rect 116084 3567 116086 3576
rect 116032 3538 116084 3544
rect 117148 480 117176 18702
rect 117976 3602 118004 29242
rect 120000 29034 120028 30223
rect 119988 29028 120040 29034
rect 119988 28970 120040 28976
rect 120092 10334 120120 31470
rect 121656 28286 121684 31484
rect 122208 31470 122590 31498
rect 121644 28280 121696 28286
rect 121644 28222 121696 28228
rect 122208 22506 122236 31470
rect 122748 29300 122800 29306
rect 122748 29242 122800 29248
rect 121460 22500 121512 22506
rect 121460 22442 121512 22448
rect 122196 22500 122248 22506
rect 122196 22442 122248 22448
rect 121472 22098 121500 22442
rect 121460 22092 121512 22098
rect 121460 22034 121512 22040
rect 121644 22092 121696 22098
rect 121644 22034 121696 22040
rect 121656 19310 121684 22034
rect 121644 19304 121696 19310
rect 121644 19246 121696 19252
rect 121368 17400 121420 17406
rect 121368 17342 121420 17348
rect 120080 10328 120132 10334
rect 120080 10270 120132 10276
rect 119436 4344 119488 4350
rect 119436 4286 119488 4292
rect 118698 3904 118754 3913
rect 118698 3839 118700 3848
rect 118752 3839 118754 3848
rect 118700 3810 118752 3816
rect 117964 3596 118016 3602
rect 117964 3538 118016 3544
rect 118240 3596 118292 3602
rect 118240 3538 118292 3544
rect 118252 480 118280 3538
rect 119448 480 119476 4286
rect 121380 3738 121408 17342
rect 121644 12436 121696 12442
rect 121644 12378 121696 12384
rect 121656 6186 121684 12378
rect 121644 6180 121696 6186
rect 121644 6122 121696 6128
rect 122760 3738 122788 29242
rect 123404 29238 123432 31484
rect 123392 29232 123444 29238
rect 123392 29174 123444 29180
rect 124324 29034 124352 31484
rect 124312 29028 124364 29034
rect 124312 28970 124364 28976
rect 125152 25566 125180 31484
rect 125704 31470 126086 31498
rect 125508 29232 125560 29238
rect 125508 29174 125560 29180
rect 125140 25560 125192 25566
rect 125140 25502 125192 25508
rect 125416 22908 125468 22914
rect 125416 22850 125468 22856
rect 122932 4344 122984 4350
rect 122930 4312 122932 4321
rect 123024 4344 123076 4350
rect 122984 4312 122986 4321
rect 123024 4286 123076 4292
rect 122930 4247 122986 4256
rect 120632 3732 120684 3738
rect 120632 3674 120684 3680
rect 121368 3732 121420 3738
rect 121368 3674 121420 3680
rect 121828 3732 121880 3738
rect 121828 3674 121880 3680
rect 122748 3732 122800 3738
rect 122748 3674 122800 3680
rect 120644 480 120672 3674
rect 121840 480 121868 3674
rect 123036 480 123064 4286
rect 125428 3738 125456 22850
rect 124220 3732 124272 3738
rect 124220 3674 124272 3680
rect 125416 3732 125468 3738
rect 125416 3674 125468 3680
rect 124232 480 124260 3674
rect 125520 3618 125548 29174
rect 125704 6254 125732 31470
rect 126900 29782 126928 31484
rect 127728 29918 127756 31484
rect 128372 31470 128662 31498
rect 129200 31470 129490 31498
rect 127716 29912 127768 29918
rect 127716 29854 127768 29860
rect 126888 29776 126940 29782
rect 126888 29718 126940 29724
rect 126888 13116 126940 13122
rect 126888 13058 126940 13064
rect 126900 9654 126928 13058
rect 126888 9648 126940 9654
rect 126888 9590 126940 9596
rect 127806 7576 127862 7585
rect 127806 7511 127862 7520
rect 125692 6248 125744 6254
rect 125692 6190 125744 6196
rect 125692 4344 125744 4350
rect 125690 4312 125692 4321
rect 125744 4312 125746 4321
rect 125690 4247 125746 4256
rect 125428 3590 125548 3618
rect 125428 480 125456 3590
rect 126612 604 126664 610
rect 126612 546 126664 552
rect 126624 480 126652 546
rect 127820 480 127848 7511
rect 128372 4865 128400 31470
rect 129200 26874 129228 31470
rect 130396 29646 130424 31484
rect 130384 29640 130436 29646
rect 130384 29582 130436 29588
rect 131224 29170 131252 31484
rect 131316 31470 132158 31498
rect 132604 31470 132986 31498
rect 131212 29164 131264 29170
rect 131212 29106 131264 29112
rect 128556 26846 129228 26874
rect 128556 14482 128584 26846
rect 128544 14476 128596 14482
rect 128544 14418 128596 14424
rect 131028 13252 131080 13258
rect 131028 13194 131080 13200
rect 129002 11656 129058 11665
rect 129002 11591 129058 11600
rect 128358 4856 128414 4865
rect 128358 4791 128414 4800
rect 129016 480 129044 11591
rect 131040 3874 131068 13194
rect 131316 12594 131344 31470
rect 131224 12566 131344 12594
rect 131224 4894 131252 12566
rect 132500 11756 132552 11762
rect 132500 11698 132552 11704
rect 131394 7712 131450 7721
rect 131394 7647 131450 7656
rect 131212 4888 131264 4894
rect 131212 4830 131264 4836
rect 130200 3868 130252 3874
rect 130200 3810 130252 3816
rect 131028 3868 131080 3874
rect 131028 3810 131080 3816
rect 129830 3632 129886 3641
rect 129830 3567 129886 3576
rect 129844 3534 129872 3567
rect 129832 3528 129884 3534
rect 129832 3470 129884 3476
rect 130212 480 130240 3810
rect 131408 480 131436 7647
rect 132512 7290 132540 11698
rect 132604 8974 132632 31470
rect 133800 29442 133828 31484
rect 133788 29436 133840 29442
rect 133788 29378 133840 29384
rect 134720 29102 134748 31484
rect 135364 31470 135562 31498
rect 135640 31470 136482 31498
rect 136652 31470 137310 31498
rect 134708 29096 134760 29102
rect 134708 29038 134760 29044
rect 132592 8968 132644 8974
rect 132592 8910 132644 8916
rect 134890 8936 134946 8945
rect 134890 8871 134946 8880
rect 132512 7262 132632 7290
rect 132604 480 132632 7262
rect 133236 3664 133288 3670
rect 133234 3632 133236 3641
rect 133288 3632 133290 3641
rect 133234 3567 133290 3576
rect 133788 2100 133840 2106
rect 133788 2042 133840 2048
rect 133800 480 133828 2042
rect 134904 480 134932 8871
rect 135364 4826 135392 31470
rect 135640 12594 135668 31470
rect 135548 12566 135668 12594
rect 135548 12458 135576 12566
rect 135456 12430 135576 12458
rect 135352 4820 135404 4826
rect 135352 4762 135404 4768
rect 135456 3534 135484 12430
rect 136086 10296 136142 10305
rect 136086 10231 136142 10240
rect 135444 3528 135496 3534
rect 135444 3470 135496 3476
rect 136100 480 136128 10231
rect 136652 3670 136680 31470
rect 138112 26784 138164 26790
rect 138112 26726 138164 26732
rect 138124 4962 138152 26726
rect 138112 4956 138164 4962
rect 138112 4898 138164 4904
rect 136640 3664 136692 3670
rect 136640 3606 136692 3612
rect 137284 3664 137336 3670
rect 137284 3606 137336 3612
rect 137296 480 137324 3606
rect 138216 3369 138244 31484
rect 138768 31470 139058 31498
rect 139412 31470 139886 31498
rect 138768 26790 138796 31470
rect 138756 26784 138808 26790
rect 138756 26726 138808 26732
rect 138478 9072 138534 9081
rect 138478 9007 138534 9016
rect 138202 3360 138258 3369
rect 138202 3295 138258 3304
rect 138492 480 138520 9007
rect 139412 3806 139440 31470
rect 140686 14512 140742 14521
rect 140686 14447 140742 14456
rect 140700 4146 140728 14447
rect 139676 4140 139728 4146
rect 139676 4082 139728 4088
rect 140688 4140 140740 4146
rect 140688 4082 140740 4088
rect 139400 3800 139452 3806
rect 139400 3742 139452 3748
rect 139688 480 139716 4082
rect 140792 3466 140820 31484
rect 140884 31470 141634 31498
rect 142264 31470 142554 31498
rect 140884 5030 140912 31470
rect 142066 10432 142122 10441
rect 142066 10367 142122 10376
rect 140962 6216 141018 6225
rect 140962 6151 141018 6160
rect 140872 5024 140924 5030
rect 140872 4966 140924 4972
rect 140780 3460 140832 3466
rect 140780 3402 140832 3408
rect 140976 2802 141004 6151
rect 140884 2774 141004 2802
rect 140884 480 140912 2774
rect 142080 480 142108 10367
rect 142264 7614 142292 31470
rect 143368 29918 143396 31484
rect 143552 31470 144302 31498
rect 145024 31470 145130 31498
rect 145760 31470 146050 31498
rect 146312 31470 146878 31498
rect 147706 31470 147812 31498
rect 143356 29912 143408 29918
rect 143356 29854 143408 29860
rect 142252 7608 142304 7614
rect 142252 7550 142304 7556
rect 143264 7608 143316 7614
rect 143264 7550 143316 7556
rect 143276 480 143304 7550
rect 143552 6322 143580 31470
rect 144920 26784 144972 26790
rect 144920 26726 144972 26732
rect 144182 14648 144238 14657
rect 144182 14583 144238 14592
rect 144196 7614 144224 14583
rect 144184 7608 144236 7614
rect 144184 7550 144236 7556
rect 143540 6316 143592 6322
rect 143540 6258 143592 6264
rect 144460 6180 144512 6186
rect 144460 6122 144512 6128
rect 144472 480 144500 6122
rect 144932 3738 144960 26726
rect 144920 3732 144972 3738
rect 144920 3674 144972 3680
rect 145024 3534 145052 31470
rect 145760 26790 145788 31470
rect 145748 26784 145800 26790
rect 145748 26726 145800 26732
rect 145654 10568 145710 10577
rect 145654 10503 145710 10512
rect 145012 3528 145064 3534
rect 145012 3470 145064 3476
rect 145668 480 145696 10503
rect 146312 6390 146340 31470
rect 147784 11830 147812 31470
rect 148612 30054 148640 31484
rect 149164 31470 149454 31498
rect 149992 31470 150374 31498
rect 150452 31470 151202 31498
rect 151832 31470 152122 31498
rect 152476 31470 152950 31498
rect 153212 31470 153778 31498
rect 148600 30048 148652 30054
rect 148600 29990 148652 29996
rect 149060 26784 149112 26790
rect 149060 26726 149112 26732
rect 147772 11824 147824 11830
rect 147772 11766 147824 11772
rect 146852 10464 146904 10470
rect 146852 10406 146904 10412
rect 146300 6384 146352 6390
rect 146300 6326 146352 6332
rect 146864 480 146892 10406
rect 148046 7848 148102 7857
rect 148046 7783 148102 7792
rect 148060 480 148088 7783
rect 149072 3942 149100 26726
rect 149164 6458 149192 31470
rect 149992 26790 150020 31470
rect 149980 26784 150032 26790
rect 149980 26726 150032 26732
rect 149152 6452 149204 6458
rect 149152 6394 149204 6400
rect 149244 6248 149296 6254
rect 149244 6190 149296 6196
rect 149060 3936 149112 3942
rect 149060 3878 149112 3884
rect 149256 480 149284 6190
rect 150452 4010 150480 31470
rect 150624 9036 150676 9042
rect 150624 8978 150676 8984
rect 150440 4004 150492 4010
rect 150440 3946 150492 3952
rect 150636 2802 150664 8978
rect 151542 7984 151598 7993
rect 151542 7919 151598 7928
rect 150452 2774 150664 2802
rect 150452 480 150480 2774
rect 151556 480 151584 7919
rect 151832 6526 151860 31470
rect 152476 29186 152504 31470
rect 152108 29158 152504 29186
rect 152108 13190 152136 29158
rect 152464 29028 152516 29034
rect 152464 28970 152516 28976
rect 152096 13184 152148 13190
rect 152096 13126 152148 13132
rect 151820 6520 151872 6526
rect 151820 6462 151872 6468
rect 152476 4078 152504 28970
rect 152464 4072 152516 4078
rect 152464 4014 152516 4020
rect 153212 3806 153240 31470
rect 154580 26784 154632 26790
rect 154580 26726 154632 26732
rect 153936 8968 153988 8974
rect 153936 8910 153988 8916
rect 153200 3800 153252 3806
rect 153200 3742 153252 3748
rect 152740 3528 152792 3534
rect 152740 3470 152792 3476
rect 152752 480 152780 3470
rect 153948 480 153976 8910
rect 154592 6594 154620 26726
rect 154684 15910 154712 31484
rect 155144 31470 155526 31498
rect 155144 26790 155172 31470
rect 156432 29034 156460 31484
rect 156420 29028 156472 29034
rect 156420 28970 156472 28976
rect 156604 29028 156656 29034
rect 156604 28970 156656 28976
rect 155132 26784 155184 26790
rect 155132 26726 155184 26732
rect 154672 15904 154724 15910
rect 154672 15846 154724 15852
rect 156326 11792 156382 11801
rect 156326 11727 156382 11736
rect 155130 8120 155186 8129
rect 155130 8055 155186 8064
rect 154580 6588 154632 6594
rect 154580 6530 154632 6536
rect 155144 480 155172 8055
rect 156340 480 156368 11727
rect 156616 3398 156644 28970
rect 157260 24138 157288 31484
rect 157352 31470 158194 31498
rect 157248 24132 157300 24138
rect 157248 24074 157300 24080
rect 157352 18630 157380 31470
rect 159008 29034 159036 31484
rect 158996 29028 159048 29034
rect 158996 28970 159048 28976
rect 159100 26738 159128 31606
rect 160112 31470 160770 31498
rect 159364 29028 159416 29034
rect 159364 28970 159416 28976
rect 158824 26710 159128 26738
rect 157340 18624 157392 18630
rect 157340 18566 157392 18572
rect 158824 17270 158852 26710
rect 158812 17264 158864 17270
rect 158812 17206 158864 17212
rect 158718 8256 158774 8265
rect 158718 8191 158774 8200
rect 157524 4072 157576 4078
rect 157524 4014 157576 4020
rect 156604 3392 156656 3398
rect 156604 3334 156656 3340
rect 157536 480 157564 4014
rect 158732 480 158760 8191
rect 159376 3330 159404 28970
rect 160008 11824 160060 11830
rect 160008 11766 160060 11772
rect 159364 3324 159416 3330
rect 159364 3266 159416 3272
rect 160020 626 160048 11766
rect 160112 6662 160140 31470
rect 161584 29714 161612 31484
rect 161572 29708 161624 29714
rect 161572 29650 161624 29656
rect 161676 22114 161704 31606
rect 162124 29096 162176 29102
rect 162124 29038 162176 29044
rect 161584 22086 161704 22114
rect 161584 21418 161612 22086
rect 161572 21412 161624 21418
rect 161572 21354 161624 21360
rect 161388 10328 161440 10334
rect 161388 10270 161440 10276
rect 160100 6656 160152 6662
rect 160100 6598 160152 6604
rect 159928 598 160048 626
rect 161400 610 161428 10270
rect 162136 3262 162164 29038
rect 163332 28354 163360 31484
rect 163504 30184 163556 30190
rect 163504 30126 163556 30132
rect 163320 28348 163372 28354
rect 163320 28290 163372 28296
rect 163516 7698 163544 30126
rect 164252 29034 164280 31484
rect 164884 30048 164936 30054
rect 164884 29990 164936 29996
rect 164240 29028 164292 29034
rect 164240 28970 164292 28976
rect 164698 11928 164754 11937
rect 164698 11863 164754 11872
rect 163424 7670 163544 7698
rect 162308 3528 162360 3534
rect 162308 3470 162360 3476
rect 162124 3256 162176 3262
rect 162124 3198 162176 3204
rect 161112 604 161164 610
rect 159928 480 159956 598
rect 161112 546 161164 552
rect 161388 604 161440 610
rect 161388 546 161440 552
rect 161124 480 161152 546
rect 162320 480 162348 3470
rect 163424 3194 163452 7670
rect 163504 7608 163556 7614
rect 163504 7550 163556 7556
rect 163412 3188 163464 3194
rect 163412 3130 163464 3136
rect 163516 480 163544 7550
rect 164712 480 164740 11863
rect 164896 3126 164924 29990
rect 165080 22778 165108 31484
rect 165724 31470 166014 31498
rect 165068 22772 165120 22778
rect 165068 22714 165120 22720
rect 165724 6730 165752 31470
rect 166264 29912 166316 29918
rect 166264 29854 166316 29860
rect 165712 6724 165764 6730
rect 165712 6666 165764 6672
rect 164884 3120 164936 3126
rect 164884 3062 164936 3068
rect 166276 3058 166304 29854
rect 166828 29850 166856 31484
rect 167012 31470 167670 31498
rect 166816 29844 166868 29850
rect 166816 29786 166868 29792
rect 167012 19990 167040 31470
rect 168576 25634 168604 31484
rect 169116 29844 169168 29850
rect 169116 29786 169168 29792
rect 169024 29776 169076 29782
rect 169024 29718 169076 29724
rect 168564 25628 168616 25634
rect 168564 25570 168616 25576
rect 167000 19984 167052 19990
rect 167000 19926 167052 19932
rect 167092 7676 167144 7682
rect 167092 7618 167144 7624
rect 166264 3052 166316 3058
rect 166264 2994 166316 3000
rect 165896 1012 165948 1018
rect 165896 954 165948 960
rect 165908 480 165936 954
rect 167104 480 167132 7618
rect 168196 4004 168248 4010
rect 168196 3946 168248 3952
rect 168208 480 168236 3946
rect 169036 2922 169064 29718
rect 169128 2990 169156 29786
rect 169404 29034 169432 31484
rect 169772 31470 170338 31498
rect 171166 31470 171272 31498
rect 169392 29028 169444 29034
rect 169392 28970 169444 28976
rect 169772 5166 169800 31470
rect 171244 6798 171272 31470
rect 172072 29986 172100 31484
rect 172532 31470 172914 31498
rect 172060 29980 172112 29986
rect 172060 29922 172112 29928
rect 171784 29708 171836 29714
rect 171784 29650 171836 29656
rect 171796 12186 171824 29650
rect 171612 12158 171824 12186
rect 171232 6792 171284 6798
rect 171232 6734 171284 6740
rect 169760 5160 169812 5166
rect 169760 5102 169812 5108
rect 169392 3664 169444 3670
rect 169392 3606 169444 3612
rect 169116 2984 169168 2990
rect 169116 2926 169168 2932
rect 169024 2916 169076 2922
rect 169024 2858 169076 2864
rect 169404 480 169432 3606
rect 170588 3392 170640 3398
rect 170588 3334 170640 3340
rect 170600 480 170628 3334
rect 171612 2854 171640 12158
rect 171782 12064 171838 12073
rect 171782 11999 171838 12008
rect 171600 2848 171652 2854
rect 171600 2790 171652 2796
rect 171796 480 171824 11999
rect 172532 5098 172560 31470
rect 173164 29640 173216 29646
rect 173164 29582 173216 29588
rect 172520 5092 172572 5098
rect 172520 5034 172572 5040
rect 172980 4140 173032 4146
rect 172980 4082 173032 4088
rect 172992 480 173020 4082
rect 173176 3602 173204 29582
rect 173728 24206 173756 31484
rect 174648 30190 174676 31484
rect 175292 31470 175490 31498
rect 175568 31470 176410 31498
rect 174636 30184 174688 30190
rect 174636 30126 174688 30132
rect 173716 24200 173768 24206
rect 173716 24142 173768 24148
rect 174176 14476 174228 14482
rect 174176 14418 174228 14424
rect 173808 13184 173860 13190
rect 173808 13126 173860 13132
rect 173820 4146 173848 13126
rect 174188 9042 174216 14418
rect 174176 9036 174228 9042
rect 174176 8978 174228 8984
rect 174176 7744 174228 7750
rect 174176 7686 174228 7692
rect 173808 4140 173860 4146
rect 173808 4082 173860 4088
rect 173164 3596 173216 3602
rect 173164 3538 173216 3544
rect 174188 480 174216 7686
rect 175292 5234 175320 31470
rect 175568 12458 175596 31470
rect 177224 30122 177252 31484
rect 178052 31470 178158 31498
rect 177212 30116 177264 30122
rect 177212 30058 177264 30064
rect 175384 12430 175596 12458
rect 175384 6866 175412 12430
rect 175464 11892 175516 11898
rect 175464 11834 175516 11840
rect 175372 6860 175424 6866
rect 175372 6802 175424 6808
rect 175476 6746 175504 11834
rect 177764 7812 177816 7818
rect 177764 7754 177816 7760
rect 175384 6718 175504 6746
rect 175280 5228 175332 5234
rect 175280 5170 175332 5176
rect 175384 480 175412 6718
rect 176476 3732 176528 3738
rect 176476 3674 176528 3680
rect 176488 1850 176516 3674
rect 176488 1822 176608 1850
rect 176580 480 176608 1822
rect 177776 480 177804 7754
rect 178052 5302 178080 31470
rect 178236 22114 178264 31606
rect 179800 30054 179828 31484
rect 179788 30048 179840 30054
rect 179788 29990 179840 29996
rect 179892 26738 179920 31606
rect 178144 22086 178264 22114
rect 179524 26710 179920 26738
rect 178144 15978 178172 22086
rect 178132 15972 178184 15978
rect 178132 15914 178184 15920
rect 179524 12510 179552 26710
rect 181548 22846 181576 31484
rect 182468 29918 182496 31484
rect 182456 29912 182508 29918
rect 182456 29854 182508 29860
rect 181536 22840 181588 22846
rect 181536 22782 181588 22788
rect 182560 22114 182588 31606
rect 182284 22086 182588 22114
rect 183572 31470 184230 31498
rect 182284 19310 182312 22086
rect 182272 19304 182324 19310
rect 182272 19246 182324 19252
rect 183572 18698 183600 31470
rect 185044 30258 185072 31484
rect 185136 31470 185886 31498
rect 186424 31470 186806 31498
rect 185032 30252 185084 30258
rect 185032 30194 185084 30200
rect 185136 20074 185164 31470
rect 184952 20046 185164 20074
rect 184952 19394 184980 20046
rect 184952 19366 185072 19394
rect 185044 19310 185072 19366
rect 184572 19304 184624 19310
rect 184572 19246 184624 19252
rect 185032 19304 185084 19310
rect 185032 19246 185084 19252
rect 183560 18692 183612 18698
rect 183560 18634 183612 18640
rect 179512 12504 179564 12510
rect 179512 12446 179564 12452
rect 182548 12028 182600 12034
rect 182548 11970 182600 11976
rect 179328 11960 179380 11966
rect 179328 11902 179380 11908
rect 178040 5296 178092 5302
rect 178040 5238 178092 5244
rect 179340 610 179368 11902
rect 179420 9716 179472 9722
rect 179420 9658 179472 9664
rect 182180 9716 182232 9722
rect 182180 9658 182232 9664
rect 179432 5370 179460 9658
rect 182192 5438 182220 9658
rect 182180 5432 182232 5438
rect 182180 5374 182232 5380
rect 179420 5364 179472 5370
rect 179420 5306 179472 5312
rect 182178 3632 182234 3641
rect 180156 3596 180208 3602
rect 182178 3567 182180 3576
rect 180156 3538 180208 3544
rect 182232 3567 182234 3576
rect 182180 3538 182232 3544
rect 178960 604 179012 610
rect 178960 546 179012 552
rect 179328 604 179380 610
rect 179328 546 179380 552
rect 178972 480 179000 546
rect 180168 480 180196 3538
rect 181352 3256 181404 3262
rect 181352 3198 181404 3204
rect 181364 480 181392 3198
rect 182560 480 182588 11970
rect 184584 9761 184612 19246
rect 186424 17338 186452 31470
rect 187620 29850 187648 31484
rect 187712 31470 188554 31498
rect 189184 31470 189382 31498
rect 187608 29844 187660 29850
rect 187608 29786 187660 29792
rect 186412 17332 186464 17338
rect 186412 17274 186464 17280
rect 186228 12096 186280 12102
rect 186228 12038 186280 12044
rect 184570 9752 184626 9761
rect 184570 9687 184626 9696
rect 184754 9752 184810 9761
rect 184754 9687 184810 9696
rect 184848 9716 184900 9722
rect 184768 5506 184796 9687
rect 184848 9658 184900 9664
rect 184756 5500 184808 5506
rect 184756 5442 184808 5448
rect 184756 3868 184808 3874
rect 184756 3810 184808 3816
rect 182638 3632 182694 3641
rect 182638 3567 182640 3576
rect 182692 3567 182694 3576
rect 182640 3538 182692 3544
rect 183744 2508 183796 2514
rect 183744 2450 183796 2456
rect 183756 480 183784 2450
rect 184768 1986 184796 3810
rect 184860 2514 184888 9658
rect 184848 2508 184900 2514
rect 184848 2450 184900 2456
rect 184768 1958 184888 1986
rect 184860 480 184888 1958
rect 186240 626 186268 12038
rect 187712 4758 187740 31470
rect 189184 21486 189212 31470
rect 190288 29374 190316 31484
rect 190472 31470 191130 31498
rect 191944 31470 192050 31498
rect 190276 29368 190328 29374
rect 190276 29310 190328 29316
rect 189172 21480 189224 21486
rect 189172 21422 189224 21428
rect 188988 15224 189040 15230
rect 188988 15166 189040 15172
rect 187700 4752 187752 4758
rect 187700 4694 187752 4700
rect 187240 3800 187292 3806
rect 187240 3742 187292 3748
rect 186056 598 186268 626
rect 186056 480 186084 598
rect 187252 480 187280 3742
rect 189000 3330 189028 15166
rect 190368 12164 190420 12170
rect 190368 12106 190420 12112
rect 190380 3398 190408 12106
rect 190472 4690 190500 31470
rect 191944 20058 191972 31470
rect 192864 29782 192892 31484
rect 193232 31470 193706 31498
rect 192852 29776 192904 29782
rect 192852 29718 192904 29724
rect 191932 20052 191984 20058
rect 191932 19994 191984 20000
rect 191748 13388 191800 13394
rect 191748 13330 191800 13336
rect 190460 4684 190512 4690
rect 190460 4626 190512 4632
rect 191760 3398 191788 13330
rect 193232 4622 193260 31470
rect 194612 28422 194640 31484
rect 195440 30326 195468 31484
rect 195992 31470 196374 31498
rect 195428 30320 195480 30326
rect 195428 30262 195480 30268
rect 194600 28416 194652 28422
rect 194600 28358 194652 28364
rect 195888 15292 195940 15298
rect 195888 15234 195940 15240
rect 194508 12232 194560 12238
rect 194508 12174 194560 12180
rect 193220 4616 193272 4622
rect 193220 4558 193272 4564
rect 189632 3392 189684 3398
rect 189632 3334 189684 3340
rect 190368 3392 190420 3398
rect 190368 3334 190420 3340
rect 190828 3392 190880 3398
rect 190828 3334 190880 3340
rect 191748 3392 191800 3398
rect 191748 3334 191800 3340
rect 194416 3392 194468 3398
rect 194416 3334 194468 3340
rect 188436 3324 188488 3330
rect 188436 3266 188488 3272
rect 188988 3324 189040 3330
rect 188988 3266 189040 3272
rect 188448 480 188476 3266
rect 189644 480 189672 3334
rect 190840 480 190868 3334
rect 193220 3120 193272 3126
rect 193220 3062 193272 3068
rect 192024 2168 192076 2174
rect 192024 2110 192076 2116
rect 192036 480 192064 2110
rect 193232 480 193260 3062
rect 194428 480 194456 3334
rect 194520 3126 194548 12174
rect 195520 7948 195572 7954
rect 195520 7890 195572 7896
rect 195532 3330 195560 7890
rect 195520 3324 195572 3330
rect 195520 3266 195572 3272
rect 194508 3120 194560 3126
rect 194508 3062 194560 3068
rect 195900 626 195928 15234
rect 195992 4486 196020 31470
rect 197188 26246 197216 31484
rect 198108 29714 198136 31484
rect 198752 31470 198950 31498
rect 198096 29708 198148 29714
rect 198096 29650 198148 29656
rect 197176 26240 197228 26246
rect 197176 26182 197228 26188
rect 196808 12300 196860 12306
rect 196808 12242 196860 12248
rect 195980 4480 196032 4486
rect 195980 4422 196032 4428
rect 195624 598 195928 626
rect 195624 480 195652 598
rect 196820 480 196848 12242
rect 198004 4820 198056 4826
rect 198004 4762 198056 4768
rect 198016 480 198044 4762
rect 198752 4554 198780 31470
rect 199764 26926 199792 31484
rect 200684 29578 200712 31484
rect 200672 29572 200724 29578
rect 200672 29514 200724 29520
rect 199752 26920 199804 26926
rect 199752 26862 199804 26868
rect 201512 4978 201540 31484
rect 202432 24274 202460 31484
rect 203260 29510 203288 31484
rect 203904 31470 204194 31498
rect 204272 31470 205022 31498
rect 203248 29504 203300 29510
rect 203248 29446 203300 29452
rect 202420 24268 202472 24274
rect 202420 24210 202472 24216
rect 203904 22166 203932 31470
rect 203064 22160 203116 22166
rect 203064 22102 203116 22108
rect 203892 22160 203944 22166
rect 203892 22102 203944 22108
rect 202788 15428 202840 15434
rect 202788 15370 202840 15376
rect 202800 9654 202828 15370
rect 202788 9648 202840 9654
rect 202788 9590 202840 9596
rect 201420 4950 201540 4978
rect 198740 4548 198792 4554
rect 198740 4490 198792 4496
rect 201420 4418 201448 4950
rect 201498 4856 201554 4865
rect 201498 4791 201554 4800
rect 201408 4412 201460 4418
rect 201408 4354 201460 4360
rect 200396 2304 200448 2310
rect 200396 2246 200448 2252
rect 199200 2236 199252 2242
rect 199200 2178 199252 2184
rect 199212 480 199240 2178
rect 200408 480 200436 2246
rect 201512 480 201540 4791
rect 203076 4282 203104 22102
rect 204272 18766 204300 31470
rect 205836 29646 205864 31484
rect 206020 31470 206770 31498
rect 207032 31470 207598 31498
rect 205824 29640 205876 29646
rect 205824 29582 205876 29588
rect 206020 26874 206048 31470
rect 205836 26846 206048 26874
rect 204260 18760 204312 18766
rect 204260 18702 204312 18708
rect 204168 15360 204220 15366
rect 204168 15302 204220 15308
rect 203064 4276 203116 4282
rect 203064 4218 203116 4224
rect 204180 2530 204208 15302
rect 204904 14544 204956 14550
rect 205836 14498 205864 26846
rect 207032 17406 207060 31470
rect 208504 29306 208532 31484
rect 208492 29300 208544 29306
rect 208492 29242 208544 29248
rect 208688 26738 208716 31606
rect 208596 26710 208716 26738
rect 207020 17400 207072 17406
rect 207020 17342 207072 17348
rect 208596 14498 208624 26710
rect 210252 22914 210280 31484
rect 211080 29238 211108 31484
rect 231964 30297 231992 38542
rect 284588 30297 284616 31484
rect 231950 30288 232006 30297
rect 231950 30223 232006 30232
rect 284574 30288 284630 30297
rect 284574 30223 284630 30232
rect 211068 29232 211120 29238
rect 211068 29174 211120 29180
rect 411260 27600 411312 27606
rect 411258 27568 411260 27577
rect 411312 27568 411314 27577
rect 411258 27503 411314 27512
rect 210240 22908 210292 22914
rect 210240 22850 210292 22856
rect 437598 16510 437888 16538
rect 378048 16380 378100 16386
rect 378048 16322 378100 16328
rect 318064 16312 318116 16318
rect 318064 16254 318116 16260
rect 300124 16244 300176 16250
rect 300124 16186 300176 16192
rect 286324 16176 286376 16182
rect 286324 16118 286376 16124
rect 285588 16040 285640 16046
rect 285588 15982 285640 15988
rect 280068 15972 280120 15978
rect 280068 15914 280120 15920
rect 278688 15904 278740 15910
rect 278688 15846 278740 15852
rect 273168 15836 273220 15842
rect 273168 15778 273220 15784
rect 266268 15768 266320 15774
rect 266268 15710 266320 15716
rect 259368 15700 259420 15706
rect 259368 15642 259420 15648
rect 240048 15632 240100 15638
rect 240048 15574 240100 15580
rect 233148 15564 233200 15570
rect 233148 15506 233200 15512
rect 222108 15496 222160 15502
rect 222108 15438 222160 15444
rect 214564 14612 214616 14618
rect 214564 14554 214616 14560
rect 204904 14486 204956 14492
rect 204916 8974 204944 14486
rect 205744 14470 205864 14498
rect 208504 14470 208624 14498
rect 205744 9722 205772 14470
rect 208308 13456 208360 13462
rect 208308 13398 208360 13404
rect 205732 9716 205784 9722
rect 205732 9658 205784 9664
rect 206008 9716 206060 9722
rect 206008 9658 206060 9664
rect 204904 8968 204956 8974
rect 204904 8910 204956 8916
rect 205086 4992 205142 5001
rect 205086 4927 205142 4936
rect 203904 2502 204208 2530
rect 202696 604 202748 610
rect 202696 546 202748 552
rect 202708 480 202736 546
rect 203904 480 203932 2502
rect 205100 480 205128 4927
rect 206020 4350 206048 9658
rect 206282 9208 206338 9217
rect 206282 9143 206338 9152
rect 206008 4344 206060 4350
rect 206008 4286 206060 4292
rect 206296 480 206324 9143
rect 208320 4078 208348 13398
rect 208504 9722 208532 14470
rect 211068 13592 211120 13598
rect 211068 13534 211120 13540
rect 208492 9716 208544 9722
rect 208492 9658 208544 9664
rect 208860 9716 208912 9722
rect 208860 9658 208912 9664
rect 208676 4888 208728 4894
rect 208676 4830 208728 4836
rect 207480 4072 207532 4078
rect 207480 4014 207532 4020
rect 208308 4072 208360 4078
rect 208308 4014 208360 4020
rect 207492 480 207520 4014
rect 208688 480 208716 4830
rect 208872 4214 208900 9658
rect 209872 8968 209924 8974
rect 209872 8910 209924 8916
rect 208860 4208 208912 4214
rect 208860 4150 208912 4156
rect 209884 480 209912 8910
rect 211080 480 211108 13534
rect 213460 9036 213512 9042
rect 213460 8978 213512 8984
rect 212262 5128 212318 5137
rect 212262 5063 212318 5072
rect 212276 480 212304 5063
rect 213472 480 213500 8978
rect 214576 3398 214604 14554
rect 219256 13524 219308 13530
rect 219256 13466 219308 13472
rect 217048 9104 217100 9110
rect 217048 9046 217100 9052
rect 215852 5024 215904 5030
rect 215852 4966 215904 4972
rect 214564 3392 214616 3398
rect 214564 3334 214616 3340
rect 214656 2372 214708 2378
rect 214656 2314 214708 2320
rect 214668 480 214696 2314
rect 215864 480 215892 4966
rect 217060 480 217088 9046
rect 219268 3398 219296 13466
rect 220544 9172 220596 9178
rect 220544 9114 220596 9120
rect 219348 5092 219400 5098
rect 219348 5034 219400 5040
rect 218152 3392 218204 3398
rect 218152 3334 218204 3340
rect 219256 3392 219308 3398
rect 219256 3334 219308 3340
rect 218164 480 218192 3334
rect 219360 480 219388 5034
rect 220556 480 220584 9114
rect 220820 8016 220872 8022
rect 220820 7958 220872 7964
rect 220832 4146 220860 7958
rect 220820 4140 220872 4146
rect 220820 4082 220872 4088
rect 222120 3482 222148 15438
rect 232502 13016 232558 13025
rect 232502 12951 232558 12960
rect 225604 12368 225656 12374
rect 225604 12310 225656 12316
rect 224132 9240 224184 9246
rect 224132 9182 224184 9188
rect 222936 5160 222988 5166
rect 222936 5102 222988 5108
rect 221752 3454 222148 3482
rect 221752 480 221780 3454
rect 222948 480 222976 5102
rect 224144 480 224172 9182
rect 225328 4072 225380 4078
rect 225328 4014 225380 4020
rect 225340 480 225368 4014
rect 225616 4010 225644 12310
rect 229100 12164 229152 12170
rect 229100 12106 229152 12112
rect 229112 11558 229140 12106
rect 229100 11552 229152 11558
rect 229100 11494 229152 11500
rect 231308 9376 231360 9382
rect 231308 9318 231360 9324
rect 227720 9308 227772 9314
rect 227720 9250 227772 9256
rect 226524 5228 226576 5234
rect 226524 5170 226576 5176
rect 225604 4004 225656 4010
rect 225604 3946 225656 3952
rect 226536 480 226564 5170
rect 227732 480 227760 9250
rect 230112 5296 230164 5302
rect 230112 5238 230164 5244
rect 228916 2440 228968 2446
rect 228916 2382 228968 2388
rect 228928 480 228956 2382
rect 230124 480 230152 5238
rect 231320 480 231348 9318
rect 232516 3942 232544 12951
rect 232504 3936 232556 3942
rect 232504 3878 232556 3884
rect 233160 3398 233188 15506
rect 239402 13152 239458 13161
rect 239402 13087 239458 13096
rect 238668 12164 238720 12170
rect 238668 12106 238720 12112
rect 238680 11558 238708 12106
rect 238668 11552 238720 11558
rect 238668 11494 238720 11500
rect 238392 9512 238444 9518
rect 238392 9454 238444 9460
rect 234804 9444 234856 9450
rect 234804 9386 234856 9392
rect 233700 5364 233752 5370
rect 233700 5306 233752 5312
rect 232504 3392 232556 3398
rect 232504 3334 232556 3340
rect 233148 3392 233200 3398
rect 233148 3334 233200 3340
rect 232516 480 232544 3334
rect 233712 480 233740 5306
rect 234816 480 234844 9386
rect 237196 5432 237248 5438
rect 237196 5374 237248 5380
rect 236000 2508 236052 2514
rect 236000 2450 236052 2456
rect 236012 480 236040 2450
rect 237208 480 237236 5374
rect 238404 480 238432 9454
rect 239416 3534 239444 13087
rect 240060 3534 240088 15574
rect 257344 13660 257396 13666
rect 257344 13602 257396 13608
rect 250442 13424 250498 13433
rect 250442 13359 250498 13368
rect 243542 13288 243598 13297
rect 243542 13223 243598 13232
rect 241980 9580 242032 9586
rect 241980 9522 242032 9528
rect 240784 5500 240836 5506
rect 240784 5442 240836 5448
rect 239404 3528 239456 3534
rect 239404 3470 239456 3476
rect 239588 3528 239640 3534
rect 239588 3470 239640 3476
rect 240048 3528 240100 3534
rect 240048 3470 240100 3476
rect 239600 480 239628 3470
rect 240796 480 240824 5442
rect 241992 480 242020 9522
rect 243556 3670 243584 13223
rect 246302 12200 246358 12209
rect 246302 12135 246358 12144
rect 248420 12164 248472 12170
rect 245568 9648 245620 9654
rect 245568 9590 245620 9596
rect 244372 4752 244424 4758
rect 244372 4694 244424 4700
rect 243544 3664 243596 3670
rect 243544 3606 243596 3612
rect 243176 2576 243228 2582
rect 243176 2518 243228 2524
rect 243188 480 243216 2518
rect 244384 480 244412 4694
rect 245580 480 245608 9590
rect 246316 3466 246344 12135
rect 248420 12106 248472 12112
rect 248432 11558 248460 12106
rect 248420 11552 248472 11558
rect 248420 11494 248472 11500
rect 249156 8900 249208 8906
rect 249156 8842 249208 8848
rect 247960 4684 248012 4690
rect 247960 4626 248012 4632
rect 246764 4004 246816 4010
rect 246764 3946 246816 3952
rect 246304 3460 246356 3466
rect 246304 3402 246356 3408
rect 246776 480 246804 3946
rect 247972 480 248000 4626
rect 249168 480 249196 8842
rect 250456 3738 250484 13359
rect 252652 8832 252704 8838
rect 252652 8774 252704 8780
rect 251456 4616 251508 4622
rect 251456 4558 251508 4564
rect 250444 3732 250496 3738
rect 250444 3674 250496 3680
rect 250352 3664 250404 3670
rect 250352 3606 250404 3612
rect 250364 480 250392 3606
rect 251468 480 251496 4558
rect 252664 480 252692 8774
rect 256240 8764 256292 8770
rect 256240 8706 256292 8712
rect 255044 4548 255096 4554
rect 255044 4490 255096 4496
rect 253848 2916 253900 2922
rect 253848 2858 253900 2864
rect 253860 480 253888 2858
rect 255056 480 255084 4490
rect 256252 480 256280 8706
rect 257356 3602 257384 13602
rect 257988 12164 258040 12170
rect 257988 12106 258040 12112
rect 258000 11558 258028 12106
rect 257988 11552 258040 11558
rect 257988 11494 258040 11500
rect 257436 3936 257488 3942
rect 257436 3878 257488 3884
rect 257344 3596 257396 3602
rect 257344 3538 257396 3544
rect 257448 480 257476 3878
rect 259380 3534 259408 15642
rect 261484 13728 261536 13734
rect 261484 13670 261536 13676
rect 259828 8696 259880 8702
rect 259828 8638 259880 8644
rect 258632 3528 258684 3534
rect 258632 3470 258684 3476
rect 259368 3528 259420 3534
rect 259368 3470 259420 3476
rect 258644 480 258672 3470
rect 259840 480 259868 8638
rect 261496 3806 261524 13670
rect 263416 8628 263468 8634
rect 263416 8570 263468 8576
rect 261484 3800 261536 3806
rect 261484 3742 261536 3748
rect 261024 2848 261076 2854
rect 261024 2790 261076 2796
rect 261036 480 261064 2790
rect 262220 2644 262272 2650
rect 262220 2586 262272 2592
rect 262232 480 262260 2586
rect 263428 480 263456 8570
rect 264612 3732 264664 3738
rect 264612 3674 264664 3680
rect 264624 480 264652 3674
rect 266280 3534 266308 15710
rect 268384 13796 268436 13802
rect 268384 13738 268436 13744
rect 267740 12164 267792 12170
rect 267740 12106 267792 12112
rect 267752 11558 267780 12106
rect 267740 11552 267792 11558
rect 267740 11494 267792 11500
rect 267004 8560 267056 8566
rect 267004 8502 267056 8508
rect 265808 3528 265860 3534
rect 265808 3470 265860 3476
rect 266268 3528 266320 3534
rect 266268 3470 266320 3476
rect 265820 480 265848 3470
rect 267016 480 267044 8502
rect 268396 3874 268424 13738
rect 270500 8492 270552 8498
rect 270500 8434 270552 8440
rect 268384 3868 268436 3874
rect 268384 3810 268436 3816
rect 268108 3596 268160 3602
rect 268108 3538 268160 3544
rect 268120 480 268148 3538
rect 269304 2712 269356 2718
rect 269304 2654 269356 2660
rect 269316 480 269344 2654
rect 270512 480 270540 8434
rect 271696 3528 271748 3534
rect 273180 3482 273208 15778
rect 275284 12436 275336 12442
rect 275284 12378 275336 12384
rect 275296 4078 275324 12378
rect 277308 12164 277360 12170
rect 277308 12106 277360 12112
rect 277320 11558 277348 12106
rect 277308 11552 277360 11558
rect 277308 11494 277360 11500
rect 275284 4072 275336 4078
rect 275284 4014 275336 4020
rect 271696 3470 271748 3476
rect 271708 480 271736 3470
rect 272904 3454 273208 3482
rect 272904 480 272932 3454
rect 278700 3398 278728 15846
rect 275284 3392 275336 3398
rect 275284 3334 275336 3340
rect 277676 3392 277728 3398
rect 277676 3334 277728 3340
rect 278688 3392 278740 3398
rect 278688 3334 278740 3340
rect 278870 3360 278926 3369
rect 274088 2780 274140 2786
rect 274088 2722 274140 2728
rect 274100 480 274128 2722
rect 275296 480 275324 3334
rect 276480 2032 276532 2038
rect 276480 1974 276532 1980
rect 276492 480 276520 1974
rect 277688 480 277716 3334
rect 278870 3295 278926 3304
rect 278884 480 278912 3295
rect 280080 480 280108 15914
rect 283654 6352 283710 6361
rect 283654 6287 283710 6296
rect 282460 3324 282512 3330
rect 282460 3266 282512 3272
rect 281264 1964 281316 1970
rect 281264 1906 281316 1912
rect 281276 480 281304 1906
rect 282472 480 282500 3266
rect 283668 480 283696 6287
rect 285600 3398 285628 15982
rect 286336 4010 286364 16118
rect 296628 16108 296680 16114
rect 296628 16050 296680 16056
rect 287060 12164 287112 12170
rect 287060 12106 287112 12112
rect 287072 11558 287100 12106
rect 287060 11552 287112 11558
rect 287060 11494 287112 11500
rect 289728 10396 289780 10402
rect 289728 10338 289780 10344
rect 287152 6316 287204 6322
rect 287152 6258 287204 6264
rect 286324 4004 286376 4010
rect 286324 3946 286376 3952
rect 285954 3496 286010 3505
rect 285954 3431 286010 3440
rect 284760 3392 284812 3398
rect 284760 3334 284812 3340
rect 285588 3392 285640 3398
rect 285588 3334 285640 3340
rect 284772 480 284800 3334
rect 285968 480 285996 3431
rect 287164 480 287192 6258
rect 289740 3346 289768 10338
rect 292304 8084 292356 8090
rect 292304 8026 292356 8032
rect 290740 6384 290792 6390
rect 290740 6326 290792 6332
rect 289556 3318 289768 3346
rect 288348 1896 288400 1902
rect 288348 1838 288400 1844
rect 288360 480 288388 1838
rect 289556 480 289584 3318
rect 290752 480 290780 6326
rect 291936 4480 291988 4486
rect 291936 4422 291988 4428
rect 291948 480 291976 4422
rect 292316 3602 292344 8026
rect 294328 6452 294380 6458
rect 294328 6394 294380 6400
rect 293130 3632 293186 3641
rect 292304 3596 292356 3602
rect 293130 3567 293186 3576
rect 292304 3538 292356 3544
rect 292580 2916 292632 2922
rect 292580 2858 292632 2864
rect 292592 1766 292620 2858
rect 292580 1760 292632 1766
rect 292580 1702 292632 1708
rect 293144 480 293172 3567
rect 294340 480 294368 6394
rect 296640 3602 296668 16050
rect 298008 10668 298060 10674
rect 298008 10610 298060 10616
rect 297916 6520 297968 6526
rect 297916 6462 297968 6468
rect 295524 3596 295576 3602
rect 295524 3538 295576 3544
rect 296628 3596 296680 3602
rect 296628 3538 296680 3544
rect 296720 3596 296772 3602
rect 296720 3538 296772 3544
rect 295536 480 295564 3538
rect 296732 480 296760 3538
rect 297928 480 297956 6462
rect 298020 3602 298048 10610
rect 300136 3942 300164 16186
rect 311808 14816 311860 14822
rect 311808 14758 311860 14764
rect 305000 14748 305052 14754
rect 305000 14690 305052 14696
rect 302240 14680 302292 14686
rect 302240 14622 302292 14628
rect 302252 10402 302280 14622
rect 304264 13048 304316 13054
rect 304264 12990 304316 12996
rect 302240 10396 302292 10402
rect 302240 10338 302292 10344
rect 303528 10396 303580 10402
rect 303528 10338 303580 10344
rect 301412 6588 301464 6594
rect 301412 6530 301464 6536
rect 300124 3936 300176 3942
rect 300124 3878 300176 3884
rect 298008 3596 298060 3602
rect 298008 3538 298060 3544
rect 300308 3392 300360 3398
rect 300308 3334 300360 3340
rect 299112 1828 299164 1834
rect 299112 1770 299164 1776
rect 299124 480 299152 1770
rect 300320 480 300348 3334
rect 301424 480 301452 6530
rect 303540 3602 303568 10338
rect 304276 3670 304304 12990
rect 305012 10674 305040 14690
rect 306380 12164 306432 12170
rect 306380 12106 306432 12112
rect 306392 11558 306420 12106
rect 306380 11552 306432 11558
rect 306380 11494 306432 11500
rect 305000 10668 305052 10674
rect 305000 10610 305052 10616
rect 310428 10600 310480 10606
rect 310428 10542 310480 10548
rect 306288 10532 306340 10538
rect 306288 10474 306340 10480
rect 305000 6656 305052 6662
rect 305000 6598 305052 6604
rect 304264 3664 304316 3670
rect 304264 3606 304316 3612
rect 302608 3596 302660 3602
rect 302608 3538 302660 3544
rect 303528 3596 303580 3602
rect 303528 3538 303580 3544
rect 302620 480 302648 3538
rect 303804 3120 303856 3126
rect 303804 3062 303856 3068
rect 303816 480 303844 3062
rect 305012 480 305040 6598
rect 306300 3482 306328 10474
rect 308588 6724 308640 6730
rect 308588 6666 308640 6672
rect 307392 3664 307444 3670
rect 307392 3606 307444 3612
rect 306208 3454 306328 3482
rect 306208 480 306236 3454
rect 307404 480 307432 3606
rect 308600 480 308628 6666
rect 310440 3398 310468 10542
rect 311820 3398 311848 14758
rect 313280 14068 313332 14074
rect 313280 14010 313332 14016
rect 313292 10470 313320 14010
rect 315948 12164 316000 12170
rect 315948 12106 316000 12112
rect 315960 11558 315988 12106
rect 315948 11552 316000 11558
rect 315948 11494 316000 11500
rect 317328 10668 317380 10674
rect 317328 10610 317380 10616
rect 313280 10464 313332 10470
rect 313280 10406 313332 10412
rect 314568 10464 314620 10470
rect 314568 10406 314620 10412
rect 312176 6792 312228 6798
rect 312176 6734 312228 6740
rect 309784 3392 309836 3398
rect 309784 3334 309836 3340
rect 310428 3392 310480 3398
rect 310428 3334 310480 3340
rect 310980 3392 311032 3398
rect 310980 3334 311032 3340
rect 311808 3392 311860 3398
rect 311808 3334 311860 3340
rect 309796 480 309824 3334
rect 310992 480 311020 3334
rect 311164 2848 311216 2854
rect 311164 2790 311216 2796
rect 311176 1698 311204 2790
rect 311164 1692 311216 1698
rect 311164 1634 311216 1640
rect 312188 480 312216 6734
rect 314476 3800 314528 3806
rect 314476 3742 314528 3748
rect 313372 3392 313424 3398
rect 313372 3334 313424 3340
rect 313384 480 313412 3334
rect 314488 1986 314516 3742
rect 314580 3398 314608 10406
rect 315764 6860 315816 6866
rect 315764 6802 315816 6808
rect 314568 3392 314620 3398
rect 314568 3334 314620 3340
rect 314488 1958 314608 1986
rect 314580 480 314608 1958
rect 315776 480 315804 6802
rect 317340 3482 317368 10610
rect 318076 3738 318104 16254
rect 354588 15156 354640 15162
rect 354588 15098 354640 15104
rect 340788 15088 340840 15094
rect 340788 15030 340840 15036
rect 332508 15020 332560 15026
rect 332508 14962 332560 14968
rect 325608 14952 325660 14958
rect 325608 14894 325660 14900
rect 318708 14884 318760 14890
rect 318708 14826 318760 14832
rect 318064 3732 318116 3738
rect 318064 3674 318116 3680
rect 316972 3454 317368 3482
rect 316972 480 317000 3454
rect 318720 3398 318748 14826
rect 324228 10804 324280 10810
rect 324228 10746 324280 10752
rect 321468 10736 321520 10742
rect 321468 10678 321520 10684
rect 319260 6112 319312 6118
rect 319260 6054 319312 6060
rect 318064 3392 318116 3398
rect 318064 3334 318116 3340
rect 318708 3392 318760 3398
rect 318708 3334 318760 3340
rect 318076 480 318104 3334
rect 319272 480 319300 6054
rect 321480 3398 321508 10678
rect 322848 6044 322900 6050
rect 322848 5986 322900 5992
rect 321652 3732 321704 3738
rect 321652 3674 321704 3680
rect 320456 3392 320508 3398
rect 320456 3334 320508 3340
rect 321468 3392 321520 3398
rect 321468 3334 321520 3340
rect 320468 480 320496 3334
rect 321664 480 321692 3674
rect 322860 480 322888 5986
rect 324240 3482 324268 10746
rect 325620 3482 325648 14894
rect 330300 13864 330352 13870
rect 330300 13806 330352 13812
rect 325700 12164 325752 12170
rect 325700 12106 325752 12112
rect 325712 11558 325740 12106
rect 325700 11552 325752 11558
rect 325700 11494 325752 11500
rect 328368 10872 328420 10878
rect 328368 10814 328420 10820
rect 326436 5976 326488 5982
rect 326436 5918 326488 5924
rect 324056 3454 324268 3482
rect 325252 3454 325648 3482
rect 324056 480 324084 3454
rect 325252 480 325280 3454
rect 326448 480 326476 5918
rect 328380 3194 328408 10814
rect 330312 10334 330340 13806
rect 330300 10328 330352 10334
rect 330300 10270 330352 10276
rect 332416 10328 332468 10334
rect 332416 10270 332468 10276
rect 330024 5908 330076 5914
rect 330024 5850 330076 5856
rect 328828 3936 328880 3942
rect 328828 3878 328880 3884
rect 327632 3188 327684 3194
rect 327632 3130 327684 3136
rect 328368 3188 328420 3194
rect 328368 3130 328420 3136
rect 327644 480 327672 3130
rect 328840 480 328868 3878
rect 330036 480 330064 5850
rect 332428 3874 332456 10270
rect 331220 3868 331272 3874
rect 331220 3810 331272 3816
rect 332416 3868 332468 3874
rect 332416 3810 332468 3816
rect 331232 480 331260 3810
rect 332520 3482 332548 14962
rect 335268 12164 335320 12170
rect 335268 12106 335320 12112
rect 335280 11558 335308 12106
rect 335268 11552 335320 11558
rect 335268 11494 335320 11500
rect 339408 11008 339460 11014
rect 339408 10950 339460 10956
rect 335268 10940 335320 10946
rect 335268 10882 335320 10888
rect 333612 5840 333664 5846
rect 333612 5782 333664 5788
rect 332428 3454 332548 3482
rect 332428 480 332456 3454
rect 333624 480 333652 5782
rect 335280 3398 335308 10882
rect 337108 5772 337160 5778
rect 337108 5714 337160 5720
rect 335912 3868 335964 3874
rect 335912 3810 335964 3816
rect 334716 3392 334768 3398
rect 334716 3334 334768 3340
rect 335268 3392 335320 3398
rect 335268 3334 335320 3340
rect 334728 480 334756 3334
rect 335924 480 335952 3810
rect 337120 480 337148 5714
rect 339420 3398 339448 10950
rect 340696 5704 340748 5710
rect 340696 5646 340748 5652
rect 338304 3392 338356 3398
rect 338304 3334 338356 3340
rect 339408 3392 339460 3398
rect 339408 3334 339460 3340
rect 339500 3392 339552 3398
rect 339500 3334 339552 3340
rect 338316 480 338344 3334
rect 339512 480 339540 3334
rect 340708 480 340736 5646
rect 340800 3398 340828 15030
rect 349068 12980 349120 12986
rect 349068 12922 349120 12928
rect 342168 10260 342220 10266
rect 342168 10202 342220 10208
rect 342180 3482 342208 10202
rect 346308 10192 346360 10198
rect 346308 10134 346360 10140
rect 344284 5636 344336 5642
rect 344284 5578 344336 5584
rect 343088 4004 343140 4010
rect 343088 3946 343140 3952
rect 341904 3454 342208 3482
rect 340788 3392 340840 3398
rect 340788 3334 340840 3340
rect 341904 480 341932 3454
rect 342902 2408 342958 2417
rect 342902 2343 342904 2352
rect 342956 2343 342958 2352
rect 342904 2314 342956 2320
rect 343100 480 343128 3946
rect 344296 480 344324 5578
rect 346320 3398 346348 10134
rect 348976 10124 349028 10130
rect 348976 10066 349028 10072
rect 345480 3392 345532 3398
rect 345480 3334 345532 3340
rect 346308 3392 346360 3398
rect 346308 3334 346360 3340
rect 347872 3392 347924 3398
rect 347872 3334 347924 3340
rect 345492 480 345520 3334
rect 346676 2848 346728 2854
rect 346676 2790 346728 2796
rect 346688 480 346716 2790
rect 347686 2408 347742 2417
rect 347686 2343 347688 2352
rect 347740 2343 347742 2352
rect 347688 2314 347740 2320
rect 347412 2304 347464 2310
rect 347412 2246 347464 2252
rect 347424 2122 347452 2246
rect 347688 2236 347740 2242
rect 347688 2178 347740 2184
rect 347700 2122 347728 2178
rect 347424 2094 347728 2122
rect 347884 480 347912 3334
rect 348988 1578 349016 10066
rect 349080 3398 349108 12922
rect 351828 12912 351880 12918
rect 351828 12854 351880 12860
rect 350264 4072 350316 4078
rect 350264 4014 350316 4020
rect 349068 3392 349120 3398
rect 349068 3334 349120 3340
rect 348988 1550 349108 1578
rect 349080 480 349108 1550
rect 350276 480 350304 4014
rect 351840 3398 351868 12854
rect 353208 10056 353260 10062
rect 353208 9998 353260 10004
rect 353220 3398 353248 9998
rect 354600 3398 354628 15098
rect 361488 14408 361540 14414
rect 361488 14350 361540 14356
rect 358728 12708 358780 12714
rect 358728 12650 358780 12656
rect 357348 9988 357400 9994
rect 357348 9930 357400 9936
rect 354956 4412 355008 4418
rect 354956 4354 355008 4360
rect 351368 3392 351420 3398
rect 351368 3334 351420 3340
rect 351828 3392 351880 3398
rect 351828 3334 351880 3340
rect 352564 3392 352616 3398
rect 352564 3334 352616 3340
rect 353208 3392 353260 3398
rect 353208 3334 353260 3340
rect 353760 3392 353812 3398
rect 353760 3334 353812 3340
rect 354588 3392 354640 3398
rect 354588 3334 354640 3340
rect 351380 480 351408 3334
rect 352576 480 352604 3334
rect 353772 480 353800 3334
rect 354968 480 354996 4354
rect 357360 3398 357388 9930
rect 358740 3482 358768 12650
rect 360108 9920 360160 9926
rect 360108 9862 360160 9868
rect 360120 3482 360148 9862
rect 361500 4146 361528 14350
rect 368388 14340 368440 14346
rect 368388 14282 368440 14288
rect 364984 12708 365036 12714
rect 364984 12650 365036 12656
rect 363328 9852 363380 9858
rect 363328 9794 363380 9800
rect 360936 4140 360988 4146
rect 360936 4082 360988 4088
rect 361488 4140 361540 4146
rect 361488 4082 361540 4088
rect 358556 3454 358768 3482
rect 359752 3454 360148 3482
rect 356152 3392 356204 3398
rect 356152 3334 356204 3340
rect 357348 3392 357400 3398
rect 357348 3334 357400 3340
rect 356164 480 356192 3334
rect 357348 3256 357400 3262
rect 357348 3198 357400 3204
rect 357360 480 357388 3198
rect 358556 480 358584 3454
rect 359752 480 359780 3454
rect 360948 480 360976 4082
rect 362132 1624 362184 1630
rect 362132 1566 362184 1572
rect 362144 480 362172 1566
rect 363340 480 363368 9794
rect 364524 4140 364576 4146
rect 364524 4082 364576 4088
rect 364536 480 364564 4082
rect 364996 3330 365024 12650
rect 367008 9784 367060 9790
rect 367008 9726 367060 9732
rect 365720 8152 365772 8158
rect 365720 8094 365772 8100
rect 364984 3324 365036 3330
rect 364984 3266 365036 3272
rect 365732 480 365760 8094
rect 367020 626 367048 9726
rect 368400 626 368428 14282
rect 375196 14272 375248 14278
rect 375196 14214 375248 14220
rect 370412 8424 370464 8430
rect 370412 8366 370464 8372
rect 369216 8220 369268 8226
rect 369216 8162 369268 8168
rect 366928 598 367048 626
rect 368032 598 368428 626
rect 366928 480 366956 598
rect 368032 480 368060 598
rect 369228 480 369256 8162
rect 370424 480 370452 8366
rect 372804 8288 372856 8294
rect 372804 8230 372856 8236
rect 371608 3188 371660 3194
rect 371608 3130 371660 3136
rect 371620 480 371648 3130
rect 372816 480 372844 8230
rect 374000 4344 374052 4350
rect 374000 4286 374052 4292
rect 374012 480 374040 4286
rect 375208 480 375236 14214
rect 376392 7540 376444 7546
rect 376392 7482 376444 7488
rect 376404 480 376432 7482
rect 378060 3330 378088 16322
rect 383568 14204 383620 14210
rect 383568 14146 383620 14152
rect 382188 11688 382240 11694
rect 382188 11630 382240 11636
rect 379980 7472 380032 7478
rect 379980 7414 380032 7420
rect 377588 3324 377640 3330
rect 377588 3266 377640 3272
rect 378048 3324 378100 3330
rect 378048 3266 378100 3272
rect 377600 480 377628 3266
rect 378784 3052 378836 3058
rect 378784 2994 378836 3000
rect 378796 480 378824 2994
rect 379992 480 380020 7414
rect 382200 3330 382228 11630
rect 383476 7404 383528 7410
rect 383476 7346 383528 7352
rect 383292 4208 383344 4214
rect 383292 4150 383344 4156
rect 383304 3330 383332 4150
rect 383488 3482 383516 7346
rect 383580 4214 383608 14146
rect 390468 14136 390520 14142
rect 390468 14078 390520 14084
rect 387708 12776 387760 12782
rect 387708 12718 387760 12724
rect 384948 11620 385000 11626
rect 384948 11562 385000 11568
rect 383568 4208 383620 4214
rect 383568 4150 383620 4156
rect 384960 3482 384988 11562
rect 385776 5568 385828 5574
rect 385776 5510 385828 5516
rect 383488 3454 383608 3482
rect 381176 3324 381228 3330
rect 381176 3266 381228 3272
rect 382188 3324 382240 3330
rect 382188 3266 382240 3272
rect 382372 3324 382424 3330
rect 382372 3266 382424 3272
rect 383292 3324 383344 3330
rect 383292 3266 383344 3272
rect 381188 480 381216 3266
rect 381542 2136 381598 2145
rect 381542 2071 381544 2080
rect 381596 2071 381598 2080
rect 381544 2042 381596 2048
rect 382384 480 382412 3266
rect 383580 480 383608 3454
rect 384684 3454 384988 3482
rect 384684 480 384712 3454
rect 385788 3126 385816 5510
rect 387720 3262 387748 12718
rect 389088 11552 389140 11558
rect 389088 11494 389140 11500
rect 389100 3262 389128 11494
rect 390480 3262 390508 14078
rect 397368 14000 397420 14006
rect 397368 13942 397420 13948
rect 393228 12912 393280 12918
rect 393228 12854 393280 12860
rect 393240 12510 393268 12854
rect 393228 12504 393280 12510
rect 393228 12446 393280 12452
rect 391848 11484 391900 11490
rect 391848 11426 391900 11432
rect 390652 7336 390704 7342
rect 390652 7278 390704 7284
rect 387064 3256 387116 3262
rect 387064 3198 387116 3204
rect 387708 3256 387760 3262
rect 387708 3198 387760 3204
rect 388260 3256 388312 3262
rect 388260 3198 388312 3204
rect 389088 3256 389140 3262
rect 389088 3198 389140 3204
rect 389456 3256 389508 3262
rect 389456 3198 389508 3204
rect 390468 3256 390520 3262
rect 390468 3198 390520 3204
rect 385776 3120 385828 3126
rect 385776 3062 385828 3068
rect 385868 3052 385920 3058
rect 385868 2994 385920 3000
rect 385880 480 385908 2994
rect 386326 2136 386382 2145
rect 386326 2071 386328 2080
rect 386380 2071 386382 2080
rect 386328 2042 386380 2048
rect 385960 1828 386012 1834
rect 385960 1770 386012 1776
rect 386328 1828 386380 1834
rect 386328 1770 386380 1776
rect 385972 1714 386000 1770
rect 386340 1714 386368 1770
rect 385972 1686 386368 1714
rect 387076 480 387104 3198
rect 388272 480 388300 3198
rect 389468 480 389496 3198
rect 390664 480 390692 7278
rect 391860 480 391888 11426
rect 395988 11416 396040 11422
rect 395988 11358 396040 11364
rect 394240 7268 394292 7274
rect 394240 7210 394292 7216
rect 393044 2984 393096 2990
rect 393044 2926 393096 2932
rect 393056 480 393084 2926
rect 394252 480 394280 7210
rect 396000 3126 396028 11358
rect 397380 3126 397408 13942
rect 408408 13932 408460 13938
rect 408408 13874 408460 13880
rect 402980 12912 403032 12918
rect 403032 12860 403112 12866
rect 402980 12854 403112 12860
rect 402992 12838 403112 12854
rect 403084 12510 403112 12838
rect 403072 12504 403124 12510
rect 403072 12446 403124 12452
rect 400128 11348 400180 11354
rect 400128 11290 400180 11296
rect 397828 7200 397880 7206
rect 397828 7142 397880 7148
rect 395436 3120 395488 3126
rect 395436 3062 395488 3068
rect 395988 3120 396040 3126
rect 395988 3062 396040 3068
rect 396632 3120 396684 3126
rect 396632 3062 396684 3068
rect 397368 3120 397420 3126
rect 397368 3062 397420 3068
rect 395448 480 395476 3062
rect 396644 480 396672 3062
rect 397840 480 397868 7142
rect 400140 3126 400168 11290
rect 407028 11280 407080 11286
rect 407028 11222 407080 11228
rect 403624 9716 403676 9722
rect 403624 9658 403676 9664
rect 402520 8356 402572 8362
rect 402520 8298 402572 8304
rect 401324 7132 401376 7138
rect 401324 7074 401376 7080
rect 399024 3120 399076 3126
rect 399024 3062 399076 3068
rect 400128 3120 400180 3126
rect 400128 3062 400180 3068
rect 400220 3120 400272 3126
rect 400220 3062 400272 3068
rect 399036 480 399064 3062
rect 400232 480 400260 3062
rect 401336 480 401364 7074
rect 402532 480 402560 8298
rect 403636 3126 403664 9658
rect 404912 7064 404964 7070
rect 404912 7006 404964 7012
rect 403624 3120 403676 3126
rect 403624 3062 403676 3068
rect 403716 3120 403768 3126
rect 403716 3062 403768 3068
rect 403728 480 403756 3062
rect 404924 480 404952 7006
rect 407040 3534 407068 11222
rect 408420 3534 408448 13874
rect 414216 13122 414244 16388
rect 414204 13116 414256 13122
rect 414204 13058 414256 13064
rect 412548 12912 412600 12918
rect 410430 12880 410486 12889
rect 410430 12815 410486 12824
rect 412546 12880 412548 12889
rect 412600 12880 412602 12889
rect 412546 12815 412602 12824
rect 409788 12640 409840 12646
rect 409788 12582 409840 12588
rect 409696 11212 409748 11218
rect 409696 11154 409748 11160
rect 406108 3528 406160 3534
rect 406108 3470 406160 3476
rect 407028 3528 407080 3534
rect 407028 3470 407080 3476
rect 407304 3528 407356 3534
rect 407304 3470 407356 3476
rect 408408 3528 408460 3534
rect 408408 3470 408460 3476
rect 408500 3528 408552 3534
rect 408500 3470 408552 3476
rect 406120 480 406148 3470
rect 407316 480 407344 3470
rect 408512 480 408540 3470
rect 409708 480 409736 11154
rect 409800 3534 409828 12582
rect 410444 12510 410472 12815
rect 410432 12504 410484 12510
rect 410432 12446 410484 12452
rect 410524 12504 410576 12510
rect 410524 12446 410576 12452
rect 409788 3528 409840 3534
rect 409788 3470 409840 3476
rect 410536 3058 410564 12446
rect 413928 11144 413980 11150
rect 413928 11086 413980 11092
rect 412088 6996 412140 7002
rect 412088 6938 412140 6944
rect 410524 3052 410576 3058
rect 410524 2994 410576 3000
rect 410892 2916 410944 2922
rect 410892 2858 410944 2864
rect 410904 480 410932 2858
rect 412100 480 412128 6938
rect 413940 3534 413968 11086
rect 414584 7585 414612 16388
rect 414952 11665 414980 16388
rect 415320 13258 415348 16388
rect 415308 13252 415360 13258
rect 415308 13194 415360 13200
rect 414938 11656 414994 11665
rect 414938 11591 414994 11600
rect 415492 11076 415544 11082
rect 415492 11018 415544 11024
rect 414570 7576 414626 7585
rect 414570 7511 414626 7520
rect 413284 3528 413336 3534
rect 413284 3470 413336 3476
rect 413928 3528 413980 3534
rect 413928 3470 413980 3476
rect 413296 480 413324 3470
rect 414480 3052 414532 3058
rect 414480 2994 414532 3000
rect 414492 480 414520 2994
rect 415400 2440 415452 2446
rect 415398 2408 415400 2417
rect 415452 2408 415454 2417
rect 415398 2343 415454 2352
rect 415504 2106 415532 11018
rect 415688 7721 415716 16388
rect 416056 11762 416084 16388
rect 416332 16374 416530 16402
rect 416044 11756 416096 11762
rect 416044 11698 416096 11704
rect 416332 11082 416360 16374
rect 416688 13116 416740 13122
rect 416688 13058 416740 13064
rect 416320 11076 416372 11082
rect 416320 11018 416372 11024
rect 415674 7712 415730 7721
rect 415674 7647 415730 7656
rect 416700 3534 416728 13058
rect 416884 8945 416912 16388
rect 417252 10305 417280 16388
rect 417436 16374 417634 16402
rect 417712 16374 418002 16402
rect 417238 10296 417294 10305
rect 417238 10231 417294 10240
rect 416870 8936 416926 8945
rect 416870 8871 416926 8880
rect 417436 8786 417464 16374
rect 417712 9081 417740 16374
rect 418356 14521 418384 16388
rect 418540 16374 418830 16402
rect 418342 14512 418398 14521
rect 418342 14447 418398 14456
rect 417976 11756 418028 11762
rect 417976 11698 418028 11704
rect 417698 9072 417754 9081
rect 417698 9007 417754 9016
rect 416792 8758 417464 8786
rect 416792 4962 416820 8758
rect 416780 4956 416832 4962
rect 416780 4898 416832 4904
rect 417988 3534 418016 11698
rect 418540 6225 418568 16374
rect 419184 10441 419212 16388
rect 419552 14657 419580 16388
rect 419736 16374 419934 16402
rect 419538 14648 419594 14657
rect 419538 14583 419594 14592
rect 419448 13252 419500 13258
rect 419448 13194 419500 13200
rect 419170 10432 419226 10441
rect 419170 10367 419226 10376
rect 418526 6216 418582 6225
rect 418526 6151 418582 6160
rect 418068 4208 418120 4214
rect 418068 4150 418120 4156
rect 415676 3528 415728 3534
rect 415676 3470 415728 3476
rect 416688 3528 416740 3534
rect 416688 3470 416740 3476
rect 416872 3528 416924 3534
rect 416872 3470 416924 3476
rect 417976 3528 418028 3534
rect 417976 3470 418028 3476
rect 415492 2100 415544 2106
rect 415492 2042 415544 2048
rect 415688 480 415716 3470
rect 416884 480 416912 3470
rect 418080 3346 418108 4150
rect 417988 3318 418108 3346
rect 417988 480 418016 3318
rect 419460 626 419488 13194
rect 419736 6186 419764 16374
rect 420288 10577 420316 16388
rect 420656 14074 420684 16388
rect 420644 14068 420696 14074
rect 420644 14010 420696 14016
rect 420828 14068 420880 14074
rect 420828 14010 420880 14016
rect 420274 10568 420330 10577
rect 420274 10503 420330 10512
rect 419724 6180 419776 6186
rect 419724 6122 419776 6128
rect 420368 6180 420420 6186
rect 420368 6122 420420 6128
rect 419184 598 419488 626
rect 419184 480 419212 598
rect 420380 480 420408 6122
rect 420840 4214 420868 14010
rect 421116 7857 421144 16388
rect 421208 16374 421498 16402
rect 421102 7848 421158 7857
rect 421102 7783 421158 7792
rect 421208 6254 421236 16374
rect 421852 14482 421880 16388
rect 421840 14476 421892 14482
rect 421840 14418 421892 14424
rect 422220 7993 422248 16388
rect 422298 13832 422354 13841
rect 422298 13767 422300 13776
rect 422352 13767 422354 13776
rect 422300 13738 422352 13744
rect 422300 12912 422352 12918
rect 422298 12880 422300 12889
rect 422352 12880 422354 12889
rect 422298 12815 422354 12824
rect 422588 12209 422616 16388
rect 422956 14550 422984 16388
rect 422944 14544 422996 14550
rect 422944 14486 422996 14492
rect 422574 12200 422630 12209
rect 422574 12135 422630 12144
rect 423416 8129 423444 16388
rect 423588 12572 423640 12578
rect 423588 12514 423640 12520
rect 423402 8120 423458 8129
rect 423402 8055 423458 8064
rect 422206 7984 422262 7993
rect 422206 7919 422262 7928
rect 421196 6248 421248 6254
rect 421196 6190 421248 6196
rect 420828 4208 420880 4214
rect 420828 4150 420880 4156
rect 421378 3768 421434 3777
rect 421378 3703 421434 3712
rect 421392 3534 421420 3703
rect 423600 3534 423628 12514
rect 423784 11801 423812 16388
rect 424152 14618 424180 16388
rect 424140 14612 424192 14618
rect 424140 14554 424192 14560
rect 423770 11792 423826 11801
rect 423770 11727 423826 11736
rect 424520 8265 424548 16388
rect 424888 11082 424916 16388
rect 425256 13870 425284 16388
rect 425244 13864 425296 13870
rect 425428 13864 425480 13870
rect 425244 13806 425296 13812
rect 425426 13832 425428 13841
rect 425480 13832 425482 13841
rect 425426 13767 425482 13776
rect 425716 13161 425744 16388
rect 425702 13152 425758 13161
rect 425702 13087 425758 13096
rect 424876 11076 424928 11082
rect 424876 11018 424928 11024
rect 425060 11076 425112 11082
rect 425060 11018 425112 11024
rect 424506 8256 424562 8265
rect 424506 8191 424562 8200
rect 423956 6248 424008 6254
rect 423956 6190 424008 6196
rect 421380 3528 421432 3534
rect 421380 3470 421432 3476
rect 422760 3528 422812 3534
rect 422760 3470 422812 3476
rect 423588 3528 423640 3534
rect 423588 3470 423640 3476
rect 421564 3052 421616 3058
rect 421564 2994 421616 3000
rect 421576 480 421604 2994
rect 422772 480 422800 3470
rect 423968 480 423996 6190
rect 425072 2854 425100 11018
rect 426084 7614 426112 16388
rect 426452 11937 426480 16388
rect 426820 13025 426848 16388
rect 426806 13016 426862 13025
rect 426806 12951 426862 12960
rect 426438 11928 426494 11937
rect 426438 11863 426494 11872
rect 426440 11824 426492 11830
rect 426440 11766 426492 11772
rect 426072 7608 426124 7614
rect 426072 7550 426124 7556
rect 426348 4956 426400 4962
rect 426348 4898 426400 4904
rect 425060 2848 425112 2854
rect 425060 2790 425112 2796
rect 425152 2848 425204 2854
rect 425152 2790 425204 2796
rect 424968 2440 425020 2446
rect 424966 2408 424968 2417
rect 425020 2408 425022 2417
rect 424966 2343 425022 2352
rect 425164 480 425192 2790
rect 426360 480 426388 4898
rect 426452 3534 426480 11766
rect 427188 7682 427216 16388
rect 427556 12374 427584 16388
rect 428016 13297 428044 16388
rect 428002 13288 428058 13297
rect 428002 13223 428058 13232
rect 427544 12368 427596 12374
rect 427544 12310 427596 12316
rect 428384 7886 428412 16388
rect 428752 12073 428780 16388
rect 429120 13190 429148 16388
rect 429108 13184 429160 13190
rect 429108 13126 429160 13132
rect 429200 13184 429252 13190
rect 429200 13126 429252 13132
rect 428924 12368 428976 12374
rect 428924 12310 428976 12316
rect 428738 12064 428794 12073
rect 428738 11999 428794 12008
rect 428936 9738 428964 12310
rect 429212 9738 429240 13126
rect 428936 9710 429056 9738
rect 428372 7880 428424 7886
rect 428372 7822 428424 7828
rect 427176 7676 427228 7682
rect 427176 7618 427228 7624
rect 427544 7608 427596 7614
rect 427544 7550 427596 7556
rect 426530 3768 426586 3777
rect 426530 3703 426586 3712
rect 426544 3534 426572 3703
rect 426440 3528 426492 3534
rect 426440 3470 426492 3476
rect 426532 3528 426584 3534
rect 426532 3470 426584 3476
rect 427556 480 427584 7550
rect 429028 3210 429056 9710
rect 429120 9710 429240 9738
rect 429120 3369 429148 9710
rect 429488 7750 429516 16388
rect 429580 16374 429870 16402
rect 429580 11966 429608 16374
rect 430316 13433 430344 16388
rect 430302 13424 430358 13433
rect 430302 13359 430358 13368
rect 429568 11960 429620 11966
rect 429568 11902 429620 11908
rect 430488 11960 430540 11966
rect 430488 11902 430540 11908
rect 429476 7744 429528 7750
rect 429476 7686 429528 7692
rect 429936 4276 429988 4282
rect 429936 4218 429988 4224
rect 429106 3360 429162 3369
rect 429106 3295 429162 3304
rect 429028 3182 429148 3210
rect 429120 626 429148 3182
rect 428752 598 429148 626
rect 428752 480 428780 598
rect 429948 480 429976 4218
rect 430500 3505 430528 11902
rect 430684 7818 430712 16388
rect 431052 12034 431080 16388
rect 431420 13666 431448 16388
rect 431408 13660 431460 13666
rect 431408 13602 431460 13608
rect 431684 12368 431736 12374
rect 431684 12310 431736 12316
rect 431040 12028 431092 12034
rect 431040 11970 431092 11976
rect 430672 7812 430724 7818
rect 430672 7754 430724 7760
rect 431132 7676 431184 7682
rect 431132 7618 431184 7624
rect 430486 3496 430542 3505
rect 430486 3431 430542 3440
rect 431144 480 431172 7618
rect 431696 3641 431724 12310
rect 431788 7954 431816 16388
rect 431868 12912 431920 12918
rect 431866 12880 431868 12889
rect 431920 12880 431922 12889
rect 431866 12815 431922 12824
rect 432156 12102 432184 16388
rect 432616 13326 432644 16388
rect 432604 13320 432656 13326
rect 432604 13262 432656 13268
rect 432144 12096 432196 12102
rect 432144 12038 432196 12044
rect 432984 8022 433012 16388
rect 433352 12170 433380 16388
rect 433720 13734 433748 16388
rect 434088 15230 434116 16388
rect 434076 15224 434128 15230
rect 434076 15166 434128 15172
rect 433708 13728 433760 13734
rect 433708 13670 433760 13676
rect 433984 13728 434036 13734
rect 433984 13670 434036 13676
rect 433340 12164 433392 12170
rect 433340 12106 433392 12112
rect 433432 12096 433484 12102
rect 433432 12038 433484 12044
rect 432972 8016 433024 8022
rect 432972 7958 433024 7964
rect 431776 7948 431828 7954
rect 431776 7890 431828 7896
rect 431682 3632 431738 3641
rect 431682 3567 431738 3576
rect 433444 3534 433472 12038
rect 433524 4208 433576 4214
rect 433524 4150 433576 4156
rect 433432 3528 433484 3534
rect 433432 3470 433484 3476
rect 432328 3460 432380 3466
rect 432328 3402 432380 3408
rect 432340 480 432368 3402
rect 433536 480 433564 4150
rect 433996 3670 434024 13670
rect 434456 11898 434484 16388
rect 434916 13394 434944 16388
rect 435298 16374 435496 16402
rect 434904 13388 434956 13394
rect 434904 13330 434956 13336
rect 435364 13388 435416 13394
rect 435364 13330 435416 13336
rect 434444 11892 434496 11898
rect 434444 11834 434496 11840
rect 434810 9752 434866 9761
rect 434810 9687 434866 9696
rect 434824 9602 434852 9687
rect 434824 9574 434944 9602
rect 434628 7744 434680 7750
rect 434628 7686 434680 7692
rect 433984 3664 434036 3670
rect 433984 3606 434036 3612
rect 434640 480 434668 7686
rect 434720 2440 434772 2446
rect 434718 2408 434720 2417
rect 434772 2408 434774 2417
rect 434718 2343 434774 2352
rect 434916 2174 434944 9574
rect 435376 3806 435404 13330
rect 435468 9897 435496 16374
rect 435652 12238 435680 16388
rect 436020 13666 436048 16388
rect 436388 15298 436416 16388
rect 436376 15292 436428 15298
rect 436376 15234 436428 15240
rect 436008 13660 436060 13666
rect 436008 13602 436060 13608
rect 436756 12306 436784 16388
rect 436848 16374 437230 16402
rect 436744 12300 436796 12306
rect 436744 12242 436796 12248
rect 435640 12232 435692 12238
rect 435640 12174 435692 12180
rect 436100 11960 436152 11966
rect 436100 11902 436152 11908
rect 435454 9888 435510 9897
rect 435454 9823 435510 9832
rect 436112 3942 436140 11902
rect 436848 4826 436876 16374
rect 437572 13184 437624 13190
rect 437572 13126 437624 13132
rect 437480 11892 437532 11898
rect 437480 11834 437532 11840
rect 437492 4865 437520 11834
rect 437478 4856 437534 4865
rect 436836 4820 436888 4826
rect 436836 4762 436888 4768
rect 437020 4820 437072 4826
rect 437478 4791 437534 4800
rect 437020 4762 437072 4768
rect 436100 3936 436152 3942
rect 436100 3878 436152 3884
rect 435364 3800 435416 3806
rect 435364 3742 435416 3748
rect 435824 3528 435876 3534
rect 435824 3470 435876 3476
rect 434904 2168 434956 2174
rect 434904 2110 434956 2116
rect 435836 480 435864 3470
rect 437032 480 437060 4762
rect 437584 2310 437612 13126
rect 437860 11234 437888 16510
rect 446968 16510 447166 16538
rect 447336 16510 447534 16538
rect 480548 16510 480930 16538
rect 493612 16510 493902 16538
rect 512748 16510 513130 16538
rect 516336 16510 516534 16538
rect 437952 13190 437980 16388
rect 438044 16374 438334 16402
rect 437940 13184 437992 13190
rect 437940 13126 437992 13132
rect 438044 11898 438072 16374
rect 438688 15434 438716 16388
rect 438676 15428 438728 15434
rect 438676 15370 438728 15376
rect 439056 15366 439084 16388
rect 439332 16374 439530 16402
rect 439044 15360 439096 15366
rect 439044 15302 439096 15308
rect 439332 13666 439360 16374
rect 438860 13660 438912 13666
rect 438860 13602 438912 13608
rect 439320 13660 439372 13666
rect 439320 13602 439372 13608
rect 438032 11892 438084 11898
rect 438032 11834 438084 11840
rect 437768 11206 437888 11234
rect 437572 2304 437624 2310
rect 437572 2246 437624 2252
rect 437768 2242 437796 11206
rect 438216 7812 438268 7818
rect 438216 7754 438268 7760
rect 437756 2236 437808 2242
rect 437756 2178 437808 2184
rect 438228 480 438256 7754
rect 438872 5001 438900 13602
rect 439320 13320 439372 13326
rect 439320 13262 439372 13268
rect 438858 4992 438914 5001
rect 438858 4927 438914 4936
rect 439332 3602 439360 13262
rect 439884 9217 439912 16388
rect 440252 13462 440280 16388
rect 440436 16374 440634 16402
rect 440240 13456 440292 13462
rect 440240 13398 440292 13404
rect 439870 9208 439926 9217
rect 439870 9143 439926 9152
rect 440436 4894 440464 16374
rect 440988 8974 441016 16388
rect 441356 13598 441384 16388
rect 441344 13592 441396 13598
rect 441344 13534 441396 13540
rect 441712 12096 441764 12102
rect 441712 12038 441764 12044
rect 440976 8968 441028 8974
rect 440976 8910 441028 8916
rect 441724 5030 441752 12038
rect 441816 5137 441844 16388
rect 442184 9042 442212 16388
rect 442368 16374 442566 16402
rect 442644 16374 442934 16402
rect 443012 16374 443302 16402
rect 442172 9036 442224 9042
rect 442172 8978 442224 8984
rect 442368 8922 442396 16374
rect 442644 12102 442672 16374
rect 442632 12096 442684 12102
rect 442632 12038 442684 12044
rect 443012 9110 443040 16374
rect 443656 13530 443684 16388
rect 443748 16374 444130 16402
rect 443644 13524 443696 13530
rect 443644 13466 443696 13472
rect 443748 11642 443776 16374
rect 443828 14544 443880 14550
rect 443828 14486 443880 14492
rect 443196 11614 443776 11642
rect 443000 9104 443052 9110
rect 443000 9046 443052 9052
rect 442000 8894 442396 8922
rect 441896 7880 441948 7886
rect 441896 7822 441948 7828
rect 441802 5128 441858 5137
rect 441802 5063 441858 5072
rect 441712 5024 441764 5030
rect 441712 4966 441764 4972
rect 440424 4888 440476 4894
rect 440424 4830 440476 4836
rect 440608 4888 440660 4894
rect 440608 4830 440660 4836
rect 439412 3936 439464 3942
rect 439412 3878 439464 3884
rect 439320 3596 439372 3602
rect 439320 3538 439372 3544
rect 439424 480 439452 3878
rect 440620 480 440648 4830
rect 441908 3482 441936 7822
rect 441816 3454 441936 3482
rect 441816 480 441844 3454
rect 442000 2378 442028 8894
rect 443196 5098 443224 11614
rect 443840 10690 443868 14486
rect 443564 10662 443868 10690
rect 443184 5092 443236 5098
rect 443184 5034 443236 5040
rect 443564 3942 443592 10662
rect 444484 9178 444512 16388
rect 444852 15502 444880 16388
rect 445036 16374 445234 16402
rect 444840 15496 444892 15502
rect 444840 15438 444892 15444
rect 444472 9172 444524 9178
rect 444472 9114 444524 9120
rect 445036 9058 445064 16374
rect 445588 9314 445616 16388
rect 445668 13456 445720 13462
rect 445668 13398 445720 13404
rect 445576 9308 445628 9314
rect 445576 9250 445628 9256
rect 445300 9240 445352 9246
rect 445300 9182 445352 9188
rect 444484 9030 445064 9058
rect 444484 5166 444512 9030
rect 444472 5160 444524 5166
rect 444472 5102 444524 5108
rect 444196 5024 444248 5030
rect 444196 4966 444248 4972
rect 443552 3936 443604 3942
rect 443552 3878 443604 3884
rect 443000 3664 443052 3670
rect 443000 3606 443052 3612
rect 442078 2408 442134 2417
rect 441988 2372 442040 2378
rect 442078 2343 442080 2352
rect 441988 2314 442040 2320
rect 442132 2343 442134 2352
rect 442080 2314 442132 2320
rect 443012 480 443040 3606
rect 444208 480 444236 4966
rect 445312 3738 445340 9182
rect 445300 3732 445352 3738
rect 445300 3674 445352 3680
rect 445680 610 445708 13398
rect 445956 12442 445984 16388
rect 446140 16374 446430 16402
rect 445944 12436 445996 12442
rect 445944 12378 445996 12384
rect 446140 11642 446168 16374
rect 445864 11614 446168 11642
rect 445864 5234 445892 11614
rect 446784 9382 446812 16388
rect 446968 9897 446996 16510
rect 446954 9888 447010 9897
rect 446954 9823 447010 9832
rect 447230 9752 447286 9761
rect 447230 9687 447286 9696
rect 446772 9376 446824 9382
rect 446772 9318 446824 9324
rect 446220 9308 446272 9314
rect 446220 9250 446272 9256
rect 445852 5228 445904 5234
rect 445852 5170 445904 5176
rect 446232 3874 446260 9250
rect 446220 3868 446272 3874
rect 446220 3810 446272 3816
rect 446588 3596 446640 3602
rect 446588 3538 446640 3544
rect 445392 604 445444 610
rect 445392 546 445444 552
rect 445668 604 445720 610
rect 445668 546 445720 552
rect 445404 480 445432 546
rect 446600 480 446628 3538
rect 447244 2378 447272 9687
rect 447336 5302 447364 16510
rect 447784 14612 447836 14618
rect 447784 14554 447836 14560
rect 447324 5296 447376 5302
rect 447324 5238 447376 5244
rect 447796 3602 447824 14554
rect 447888 9450 447916 16388
rect 448256 15570 448284 16388
rect 448244 15564 448296 15570
rect 448244 15506 448296 15512
rect 447876 9444 447928 9450
rect 447876 9386 447928 9392
rect 448716 5370 448744 16388
rect 448808 16374 449098 16402
rect 449176 16374 449466 16402
rect 449544 16374 449834 16402
rect 448808 9518 448836 16374
rect 448796 9512 448848 9518
rect 448796 9454 448848 9460
rect 448704 5364 448756 5370
rect 448704 5306 448756 5312
rect 447876 5092 447928 5098
rect 447876 5034 447928 5040
rect 447784 3596 447836 3602
rect 447784 3538 447836 3544
rect 447888 2564 447916 5034
rect 449176 2802 449204 16374
rect 449544 5438 449572 16374
rect 450188 9110 450216 16388
rect 450556 15638 450584 16388
rect 450648 16374 451030 16402
rect 451292 16374 451398 16402
rect 451568 16374 451766 16402
rect 451844 16374 452134 16402
rect 450544 15632 450596 15638
rect 450544 15574 450596 15580
rect 450176 9104 450228 9110
rect 450176 9046 450228 9052
rect 450648 5506 450676 16374
rect 451292 9586 451320 16374
rect 451280 9580 451332 9586
rect 451280 9522 451332 9528
rect 451188 9512 451240 9518
rect 451188 9454 451240 9460
rect 450636 5500 450688 5506
rect 450636 5442 450688 5448
rect 449532 5432 449584 5438
rect 449532 5374 449584 5380
rect 451200 4010 451228 9454
rect 451280 5160 451332 5166
rect 451280 5102 451332 5108
rect 451188 4004 451240 4010
rect 451188 3946 451240 3952
rect 447796 2536 447916 2564
rect 449084 2774 449204 2802
rect 447232 2372 447284 2378
rect 447232 2314 447284 2320
rect 447796 480 447824 2536
rect 448980 2508 449032 2514
rect 448980 2450 449032 2456
rect 448992 480 449020 2450
rect 449084 2446 449112 2774
rect 449072 2440 449124 2446
rect 449072 2382 449124 2388
rect 450176 2100 450228 2106
rect 450176 2042 450228 2048
rect 450188 480 450216 2042
rect 451292 480 451320 5102
rect 451568 2582 451596 16374
rect 451844 4758 451872 16374
rect 452488 9586 452516 16388
rect 452856 16182 452884 16388
rect 452948 16374 453330 16402
rect 452844 16176 452896 16182
rect 452844 16118 452896 16124
rect 452476 9580 452528 9586
rect 452476 9522 452528 9528
rect 452660 9580 452712 9586
rect 452660 9522 452712 9528
rect 452476 9036 452528 9042
rect 452476 8978 452528 8984
rect 451832 4752 451884 4758
rect 451832 4694 451884 4700
rect 451556 2576 451608 2582
rect 451556 2518 451608 2524
rect 452488 480 452516 8978
rect 452672 3806 452700 9522
rect 452752 9376 452804 9382
rect 452752 9318 452804 9324
rect 452660 3800 452712 3806
rect 452660 3742 452712 3748
rect 452764 3398 452792 9318
rect 452948 4690 452976 16374
rect 453684 8906 453712 16388
rect 454052 13054 454080 16388
rect 454144 16374 454434 16402
rect 454040 13048 454092 13054
rect 454040 12990 454092 12996
rect 453672 8900 453724 8906
rect 453672 8842 453724 8848
rect 452936 4684 452988 4690
rect 452936 4626 452988 4632
rect 454144 4622 454172 16374
rect 454788 8838 454816 16388
rect 454972 16374 455170 16402
rect 455432 16374 455630 16402
rect 454776 8832 454828 8838
rect 454776 8774 454828 8780
rect 454972 7426 455000 16374
rect 454236 7398 455000 7426
rect 454132 4616 454184 4622
rect 454132 4558 454184 4564
rect 452752 3392 452804 3398
rect 452752 3334 452804 3340
rect 453672 3392 453724 3398
rect 453672 3334 453724 3340
rect 453684 480 453712 3334
rect 454236 1766 454264 7398
rect 454868 5228 454920 5234
rect 454868 5170 454920 5176
rect 454224 1760 454276 1766
rect 454224 1702 454276 1708
rect 454880 480 454908 5170
rect 455432 4554 455460 16374
rect 455984 8770 456012 16388
rect 456352 16250 456380 16388
rect 456340 16244 456392 16250
rect 456340 16186 456392 16192
rect 456720 15706 456748 16388
rect 456708 15700 456760 15706
rect 456708 15642 456760 15648
rect 456984 15224 457036 15230
rect 456984 15166 457036 15172
rect 456892 12096 456944 12102
rect 456892 12038 456944 12044
rect 456064 9104 456116 9110
rect 456064 9046 456116 9052
rect 455972 8764 456024 8770
rect 455972 8706 456024 8712
rect 455420 4548 455472 4554
rect 455420 4490 455472 4496
rect 456076 480 456104 9046
rect 456904 2650 456932 12038
rect 456892 2644 456944 2650
rect 456892 2586 456944 2592
rect 456996 1698 457024 15166
rect 457088 8702 457116 16388
rect 457456 15230 457484 16388
rect 457640 16374 457930 16402
rect 457444 15224 457496 15230
rect 457444 15166 457496 15172
rect 457444 13864 457496 13870
rect 457444 13806 457496 13812
rect 457076 8696 457128 8702
rect 457076 8638 457128 8644
rect 457260 3732 457312 3738
rect 457260 3674 457312 3680
rect 456984 1692 457036 1698
rect 456984 1634 457036 1640
rect 457272 480 457300 3674
rect 457456 3398 457484 13806
rect 457640 12102 457668 16374
rect 457628 12096 457680 12102
rect 457628 12038 457680 12044
rect 458284 8634 458312 16388
rect 458376 16374 458666 16402
rect 458376 16318 458404 16374
rect 458364 16312 458416 16318
rect 458364 16254 458416 16260
rect 459020 15774 459048 16388
rect 459008 15768 459060 15774
rect 459008 15710 459060 15716
rect 458548 9444 458600 9450
rect 458548 9386 458600 9392
rect 458272 8628 458324 8634
rect 458272 8570 458324 8576
rect 458456 5296 458508 5302
rect 458456 5238 458508 5244
rect 457444 3392 457496 3398
rect 457444 3334 457496 3340
rect 458468 480 458496 5238
rect 458560 3194 458588 9386
rect 459388 8566 459416 16388
rect 459572 16374 459770 16402
rect 459848 16374 460230 16402
rect 459376 8560 459428 8566
rect 459376 8502 459428 8508
rect 459572 8090 459600 16374
rect 459744 9172 459796 9178
rect 459744 9114 459796 9120
rect 459560 8084 459612 8090
rect 459560 8026 459612 8032
rect 458548 3188 458600 3194
rect 458548 3130 458600 3136
rect 459756 626 459784 9114
rect 459848 2718 459876 16374
rect 460584 8498 460612 16388
rect 460952 12510 460980 16388
rect 461320 15842 461348 16388
rect 461308 15836 461360 15842
rect 461308 15778 461360 15784
rect 461584 13456 461636 13462
rect 461584 13398 461636 13404
rect 461032 13388 461084 13394
rect 461032 13330 461084 13336
rect 460940 12504 460992 12510
rect 460940 12446 460992 12452
rect 460572 8492 460624 8498
rect 460572 8434 460624 8440
rect 460848 3868 460900 3874
rect 460848 3810 460900 3816
rect 459836 2712 459888 2718
rect 459836 2654 459888 2660
rect 459664 598 459784 626
rect 459664 480 459692 598
rect 460860 480 460888 3810
rect 461044 2786 461072 13330
rect 461596 4146 461624 13398
rect 461688 13394 461716 16388
rect 461676 13388 461728 13394
rect 461676 13330 461728 13336
rect 462056 11082 462084 16388
rect 462424 16374 462530 16402
rect 462044 11076 462096 11082
rect 462044 11018 462096 11024
rect 462044 5364 462096 5370
rect 462044 5306 462096 5312
rect 461584 4140 461636 4146
rect 461584 4082 461636 4088
rect 461032 2780 461084 2786
rect 461032 2722 461084 2728
rect 462056 480 462084 5306
rect 462424 2038 462452 16374
rect 462884 15910 462912 16388
rect 462872 15904 462924 15910
rect 462872 15846 462924 15852
rect 463252 13802 463280 16388
rect 463620 15978 463648 16388
rect 463896 16374 464002 16402
rect 463608 15972 463660 15978
rect 463608 15914 463660 15920
rect 463240 13796 463292 13802
rect 463240 13738 463292 13744
rect 463792 12028 463844 12034
rect 463792 11970 463844 11976
rect 463240 9240 463292 9246
rect 463240 9182 463292 9188
rect 462412 2032 462464 2038
rect 462412 1974 462464 1980
rect 463252 480 463280 9182
rect 463804 6361 463832 11970
rect 463790 6352 463846 6361
rect 463790 6287 463846 6296
rect 463896 1970 463924 16374
rect 464252 13524 464304 13530
rect 464252 13466 464304 13472
rect 464264 2990 464292 13466
rect 464356 12714 464384 16388
rect 464448 16374 464830 16402
rect 464344 12708 464396 12714
rect 464344 12650 464396 12656
rect 464448 12034 464476 16374
rect 465184 16046 465212 16388
rect 465172 16040 465224 16046
rect 465172 15982 465224 15988
rect 465552 12170 465580 16388
rect 465644 16374 465934 16402
rect 466196 16374 466302 16402
rect 465540 12164 465592 12170
rect 465540 12106 465592 12112
rect 464436 12028 464488 12034
rect 464436 11970 464488 11976
rect 465644 11642 465672 16374
rect 465184 11614 465672 11642
rect 465184 6322 465212 11614
rect 466196 11082 466224 16374
rect 466656 14686 466684 16388
rect 466748 16374 467130 16402
rect 467300 16374 467498 16402
rect 466644 14680 466696 14686
rect 466644 14622 466696 14628
rect 466748 11642 466776 16374
rect 466564 11614 466776 11642
rect 465356 11076 465408 11082
rect 465356 11018 465408 11024
rect 466184 11076 466236 11082
rect 466184 11018 466236 11024
rect 465172 6316 465224 6322
rect 465172 6258 465224 6264
rect 464436 3800 464488 3806
rect 464436 3742 464488 3748
rect 464252 2984 464304 2990
rect 464252 2926 464304 2932
rect 463884 1964 463936 1970
rect 463884 1906 463936 1912
rect 464448 480 464476 3742
rect 465368 1902 465396 11018
rect 466564 6390 466592 11614
rect 467300 11506 467328 16374
rect 467748 13388 467800 13394
rect 467748 13330 467800 13336
rect 466748 11478 467328 11506
rect 466552 6384 466604 6390
rect 466552 6326 466604 6332
rect 465632 5432 465684 5438
rect 465632 5374 465684 5380
rect 465356 1896 465408 1902
rect 465356 1838 465408 1844
rect 465644 480 465672 5374
rect 466748 4486 466776 11478
rect 466736 4480 466788 4486
rect 466736 4422 466788 4428
rect 467760 2990 467788 13330
rect 467852 12374 467880 16388
rect 468036 16374 468234 16402
rect 467840 12368 467892 12374
rect 467840 12310 467892 12316
rect 468036 6458 468064 16374
rect 468588 16114 468616 16388
rect 468576 16108 468628 16114
rect 468576 16050 468628 16056
rect 468956 14754 468984 16388
rect 469324 16374 469430 16402
rect 469508 16374 469798 16402
rect 468944 14748 468996 14754
rect 468944 14690 468996 14696
rect 469036 14680 469088 14686
rect 469036 14622 469088 14628
rect 468024 6452 468076 6458
rect 468024 6394 468076 6400
rect 469048 3398 469076 14622
rect 469324 6526 469352 16374
rect 469404 12028 469456 12034
rect 469404 11970 469456 11976
rect 469416 6594 469444 11970
rect 469404 6588 469456 6594
rect 469404 6530 469456 6536
rect 469312 6520 469364 6526
rect 469312 6462 469364 6468
rect 469128 5500 469180 5506
rect 469128 5442 469180 5448
rect 467932 3392 467984 3398
rect 467932 3334 467984 3340
rect 469036 3392 469088 3398
rect 469036 3334 469088 3340
rect 466828 2984 466880 2990
rect 466828 2926 466880 2932
rect 467748 2984 467800 2990
rect 467748 2926 467800 2932
rect 466840 480 466868 2926
rect 467944 480 467972 3334
rect 469140 480 469168 5442
rect 469508 1834 469536 16374
rect 470152 13734 470180 16388
rect 470244 16374 470534 16402
rect 470140 13728 470192 13734
rect 470140 13670 470192 13676
rect 470244 12034 470272 16374
rect 470232 12028 470284 12034
rect 470232 11970 470284 11976
rect 470692 11892 470744 11898
rect 470692 11834 470744 11840
rect 470704 6662 470732 11834
rect 470888 10402 470916 16388
rect 471072 16374 471270 16402
rect 471440 16374 471730 16402
rect 470876 10396 470928 10402
rect 470876 10338 470928 10344
rect 471072 10282 471100 16374
rect 471440 11898 471468 16374
rect 471428 11892 471480 11898
rect 471428 11834 471480 11840
rect 472084 10538 472112 16388
rect 472452 11966 472480 16388
rect 472636 16374 472834 16402
rect 472440 11960 472492 11966
rect 472440 11902 472492 11908
rect 472636 11642 472664 16374
rect 472176 11614 472664 11642
rect 472072 10532 472124 10538
rect 472072 10474 472124 10480
rect 470888 10254 471100 10282
rect 470692 6656 470744 6662
rect 470692 6598 470744 6604
rect 470324 6316 470376 6322
rect 470324 6258 470376 6264
rect 469496 1828 469548 1834
rect 469496 1770 469548 1776
rect 470336 480 470364 6258
rect 470888 5574 470916 10254
rect 472176 6730 472204 11614
rect 473188 10606 473216 16388
rect 473556 14822 473584 16388
rect 473740 16374 474030 16402
rect 473544 14816 473596 14822
rect 473544 14758 473596 14764
rect 473740 11642 473768 16374
rect 473464 11614 473768 11642
rect 473176 10600 473228 10606
rect 473176 10542 473228 10548
rect 473464 6798 473492 11614
rect 474384 10470 474412 16388
rect 474752 13666 474780 16388
rect 474936 16374 475134 16402
rect 474740 13660 474792 13666
rect 474740 13602 474792 13608
rect 474372 10464 474424 10470
rect 474372 10406 474424 10412
rect 474936 6866 474964 16374
rect 475488 10674 475516 16388
rect 475856 14890 475884 16388
rect 476224 16374 476330 16402
rect 475844 14884 475896 14890
rect 475844 14826 475896 14832
rect 476028 14748 476080 14754
rect 476028 14690 476080 14696
rect 475476 10668 475528 10674
rect 475476 10610 475528 10616
rect 474924 6860 474976 6866
rect 474924 6802 474976 6808
rect 473452 6792 473504 6798
rect 473452 6734 473504 6740
rect 472164 6724 472216 6730
rect 472164 6666 472216 6672
rect 471888 6520 471940 6526
rect 471888 6462 471940 6468
rect 470876 5568 470928 5574
rect 470876 5510 470928 5516
rect 471520 3936 471572 3942
rect 471520 3878 471572 3884
rect 471532 480 471560 3878
rect 471900 3330 471928 6462
rect 473912 6384 473964 6390
rect 473912 6326 473964 6332
rect 472716 4752 472768 4758
rect 472716 4694 472768 4700
rect 471888 3324 471940 3330
rect 471888 3266 471940 3272
rect 472728 480 472756 4694
rect 473360 3596 473412 3602
rect 473360 3538 473412 3544
rect 473452 3596 473504 3602
rect 473452 3538 473504 3544
rect 473372 3482 473400 3538
rect 473464 3482 473492 3538
rect 473372 3454 473492 3482
rect 473924 480 473952 6326
rect 476040 3398 476068 14690
rect 476120 6656 476172 6662
rect 476120 6598 476172 6604
rect 475108 3392 475160 3398
rect 475108 3334 475160 3340
rect 476028 3392 476080 3398
rect 476028 3334 476080 3340
rect 475120 480 475148 3334
rect 476132 3262 476160 6598
rect 476224 6118 476252 16374
rect 476684 10742 476712 16388
rect 476672 10736 476724 10742
rect 476672 10678 476724 10684
rect 477052 9654 477080 16388
rect 477236 16374 477434 16402
rect 477040 9648 477092 9654
rect 477040 9590 477092 9596
rect 477236 9466 477264 16374
rect 477788 10810 477816 16388
rect 478156 14958 478184 16388
rect 478340 16374 478630 16402
rect 478144 14952 478196 14958
rect 478144 14894 478196 14900
rect 477776 10804 477828 10810
rect 477776 10746 477828 10752
rect 478340 10690 478368 16374
rect 478788 14816 478840 14822
rect 478788 14758 478840 14764
rect 476316 9438 477264 9466
rect 477512 10662 478368 10690
rect 476212 6112 476264 6118
rect 476212 6054 476264 6060
rect 476316 6050 476344 9438
rect 476304 6044 476356 6050
rect 476304 5986 476356 5992
rect 477512 5982 477540 10662
rect 477592 6452 477644 6458
rect 477592 6394 477644 6400
rect 477500 5976 477552 5982
rect 477500 5918 477552 5924
rect 476304 4684 476356 4690
rect 476304 4626 476356 4632
rect 476120 3256 476172 3262
rect 476120 3198 476172 3204
rect 476316 480 476344 4626
rect 477500 3392 477552 3398
rect 477500 3334 477552 3340
rect 477512 480 477540 3334
rect 477604 3126 477632 6394
rect 478696 4004 478748 4010
rect 478696 3946 478748 3952
rect 477592 3120 477644 3126
rect 477592 3062 477644 3068
rect 478708 480 478736 3946
rect 478800 3398 478828 14758
rect 478984 10878 479012 16388
rect 479352 12034 479380 16388
rect 479536 16374 479734 16402
rect 479340 12028 479392 12034
rect 479340 11970 479392 11976
rect 479536 11642 479564 16374
rect 479076 11614 479564 11642
rect 478972 10872 479024 10878
rect 478972 10814 479024 10820
rect 479076 5914 479104 11614
rect 479524 10600 479576 10606
rect 479524 10542 479576 10548
rect 479064 5908 479116 5914
rect 479064 5850 479116 5856
rect 478788 3392 478840 3398
rect 478788 3334 478840 3340
rect 479536 2922 479564 10542
rect 480088 10334 480116 16388
rect 480456 15026 480484 16388
rect 480444 15020 480496 15026
rect 480444 14962 480496 14968
rect 480548 12458 480576 16510
rect 493612 16454 493640 16510
rect 492864 16448 492916 16454
rect 480364 12430 480576 12458
rect 480076 10328 480128 10334
rect 480076 10270 480128 10276
rect 480364 5846 480392 12430
rect 481284 10946 481312 16388
rect 481272 10940 481324 10946
rect 481272 10882 481324 10888
rect 481548 10328 481600 10334
rect 481548 10270 481600 10276
rect 480720 6588 480772 6594
rect 480720 6530 480772 6536
rect 480352 5840 480404 5846
rect 480352 5782 480404 5788
rect 479892 4616 479944 4622
rect 479892 4558 479944 4564
rect 479524 2916 479576 2922
rect 479524 2858 479576 2864
rect 479904 480 479932 4558
rect 480732 3058 480760 6530
rect 481560 3398 481588 10270
rect 481652 9314 481680 16388
rect 481836 16374 482034 16402
rect 481640 9308 481692 9314
rect 481640 9250 481692 9256
rect 481836 5778 481864 16374
rect 482388 11014 482416 16388
rect 482756 15094 482784 16388
rect 483230 16374 483336 16402
rect 482744 15088 482796 15094
rect 482744 15030 482796 15036
rect 482928 14884 482980 14890
rect 482928 14826 482980 14832
rect 482376 11008 482428 11014
rect 482376 10950 482428 10956
rect 481824 5772 481876 5778
rect 481824 5714 481876 5720
rect 482940 3398 482968 14826
rect 483112 11824 483164 11830
rect 483112 11766 483164 11772
rect 483124 5642 483152 11766
rect 483308 5710 483336 16374
rect 483584 10266 483612 16388
rect 483572 10260 483624 10266
rect 483572 10202 483624 10208
rect 483952 9518 483980 16388
rect 484044 16374 484334 16402
rect 484044 11830 484072 16374
rect 484032 11824 484084 11830
rect 484032 11766 484084 11772
rect 484688 10198 484716 16388
rect 485056 11966 485084 16388
rect 485516 12986 485544 16388
rect 485504 12980 485556 12986
rect 485504 12922 485556 12928
rect 485044 11960 485096 11966
rect 485044 11902 485096 11908
rect 485044 10668 485096 10674
rect 485044 10610 485096 10616
rect 484676 10192 484728 10198
rect 484676 10134 484728 10140
rect 483940 9512 483992 9518
rect 483940 9454 483992 9460
rect 483480 9308 483532 9314
rect 483480 9250 483532 9256
rect 483296 5704 483348 5710
rect 483296 5646 483348 5652
rect 483112 5636 483164 5642
rect 483112 5578 483164 5584
rect 481088 3392 481140 3398
rect 481088 3334 481140 3340
rect 481548 3392 481600 3398
rect 481548 3334 481600 3340
rect 482284 3392 482336 3398
rect 482284 3334 482336 3340
rect 482928 3392 482980 3398
rect 482928 3334 482980 3340
rect 480720 3052 480772 3058
rect 480720 2994 480772 3000
rect 481100 480 481128 3334
rect 482296 480 482324 3334
rect 483492 480 483520 9250
rect 484584 4548 484636 4554
rect 484584 4490 484636 4496
rect 484596 480 484624 4490
rect 485056 2854 485084 10610
rect 485884 10130 485912 16388
rect 485872 10124 485924 10130
rect 485872 10066 485924 10072
rect 486252 9586 486280 16388
rect 486620 12918 486648 16388
rect 486712 16374 487002 16402
rect 486608 12912 486660 12918
rect 486608 12854 486660 12860
rect 486712 10062 486740 16374
rect 487356 15162 487384 16388
rect 487540 16374 487830 16402
rect 487344 15156 487396 15162
rect 487344 15098 487396 15104
rect 487068 14952 487120 14958
rect 487068 14894 487120 14900
rect 486976 10396 487028 10402
rect 486976 10338 487028 10344
rect 486700 10056 486752 10062
rect 486700 9998 486752 10004
rect 486240 9580 486292 9586
rect 486240 9522 486292 9528
rect 485780 3392 485832 3398
rect 485780 3334 485832 3340
rect 485044 2848 485096 2854
rect 485044 2790 485096 2796
rect 485792 480 485820 3334
rect 486988 480 487016 10338
rect 487080 3398 487108 14894
rect 487540 11642 487568 16374
rect 487264 11614 487568 11642
rect 487264 4418 487292 11614
rect 488184 9994 488212 16388
rect 488172 9988 488224 9994
rect 488172 9930 488224 9936
rect 488552 9382 488580 16388
rect 488920 12850 488948 16388
rect 488908 12844 488960 12850
rect 488908 12786 488960 12792
rect 489288 9926 489316 16388
rect 489656 14414 489684 16388
rect 489828 15088 489880 15094
rect 489828 15030 489880 15036
rect 489644 14408 489696 14414
rect 489644 14350 489696 14356
rect 489276 9920 489328 9926
rect 489276 9862 489328 9868
rect 488540 9376 488592 9382
rect 488540 9318 488592 9324
rect 488172 4480 488224 4486
rect 488172 4422 488224 4428
rect 487252 4412 487304 4418
rect 487252 4354 487304 4360
rect 487068 3392 487120 3398
rect 487068 3334 487120 3340
rect 488184 480 488212 4422
rect 489840 3398 489868 15030
rect 489368 3392 489420 3398
rect 489368 3334 489420 3340
rect 489828 3392 489880 3398
rect 489828 3334 489880 3340
rect 489380 480 489408 3334
rect 490116 1630 490144 16388
rect 490484 9858 490512 16388
rect 490852 13462 490880 16388
rect 490944 16374 491234 16402
rect 492864 16390 492916 16396
rect 493600 16448 493652 16454
rect 493600 16390 493652 16396
rect 490840 13456 490892 13462
rect 490840 13398 490892 13404
rect 490472 9852 490524 9858
rect 490472 9794 490524 9800
rect 490944 8158 490972 16374
rect 491208 13456 491260 13462
rect 491208 13398 491260 13404
rect 490932 8152 490984 8158
rect 490932 8094 490984 8100
rect 491220 3398 491248 13398
rect 491588 9790 491616 16388
rect 491956 14346 491984 16388
rect 491944 14340 491996 14346
rect 491944 14282 491996 14288
rect 491576 9784 491628 9790
rect 491576 9726 491628 9732
rect 492416 8226 492444 16388
rect 492784 8430 492812 16388
rect 492772 8424 492824 8430
rect 492772 8366 492824 8372
rect 492404 8220 492456 8226
rect 492404 8162 492456 8168
rect 491760 4412 491812 4418
rect 491760 4354 491812 4360
rect 490564 3392 490616 3398
rect 490564 3334 490616 3340
rect 491208 3392 491260 3398
rect 491208 3334 491260 3340
rect 490104 1624 490156 1630
rect 490104 1566 490156 1572
rect 490576 480 490604 3334
rect 491772 480 491800 4354
rect 492876 4350 492904 16390
rect 493152 9450 493180 16388
rect 493140 9444 493192 9450
rect 493140 9386 493192 9392
rect 493520 8294 493548 16388
rect 494256 14278 494284 16388
rect 494244 14272 494296 14278
rect 494244 14214 494296 14220
rect 494244 9444 494296 9450
rect 494244 9386 494296 9392
rect 493508 8288 493560 8294
rect 493508 8230 493560 8236
rect 492864 4344 492916 4350
rect 492864 4286 492916 4292
rect 492956 4072 493008 4078
rect 492956 4014 493008 4020
rect 492968 480 492996 4014
rect 494256 626 494284 9386
rect 494716 7546 494744 16388
rect 494808 16386 495098 16402
rect 494796 16380 495098 16386
rect 494848 16374 495098 16380
rect 495466 16374 495664 16402
rect 494796 16322 494848 16328
rect 495348 9376 495400 9382
rect 495348 9318 495400 9324
rect 494704 7540 494756 7546
rect 494704 7482 494756 7488
rect 494164 598 494284 626
rect 494164 480 494192 598
rect 495360 480 495388 9318
rect 495636 6526 495664 16374
rect 495820 7478 495848 16388
rect 496188 11694 496216 16388
rect 496556 14210 496584 16388
rect 496728 15020 496780 15026
rect 496728 14962 496780 14968
rect 496544 14204 496596 14210
rect 496544 14146 496596 14152
rect 496176 11688 496228 11694
rect 496176 11630 496228 11636
rect 495808 7472 495860 7478
rect 495808 7414 495860 7420
rect 495624 6520 495676 6526
rect 495624 6462 495676 6468
rect 496740 610 496768 14962
rect 497016 7410 497044 16388
rect 497096 12436 497148 12442
rect 497096 12378 497148 12384
rect 497004 7404 497056 7410
rect 497004 7346 497056 7352
rect 497108 7290 497136 12378
rect 497384 11626 497412 16388
rect 497752 12442 497780 16388
rect 498120 12782 498148 16388
rect 498108 12776 498160 12782
rect 498108 12718 498160 12724
rect 497740 12436 497792 12442
rect 497740 12378 497792 12384
rect 497372 11620 497424 11626
rect 497372 11562 497424 11568
rect 498488 11558 498516 16388
rect 498856 14142 498884 16388
rect 498844 14136 498896 14142
rect 498844 14078 498896 14084
rect 498476 11552 498528 11558
rect 498476 11494 498528 11500
rect 498108 10464 498160 10470
rect 498108 10406 498160 10412
rect 496924 7262 497136 7290
rect 496924 6662 496952 7262
rect 496912 6656 496964 6662
rect 496912 6598 496964 6604
rect 498120 626 498148 10406
rect 499316 7342 499344 16388
rect 499684 11490 499712 16388
rect 500052 13530 500080 16388
rect 500040 13524 500092 13530
rect 500040 13466 500092 13472
rect 499672 11484 499724 11490
rect 499672 11426 499724 11432
rect 499488 10532 499540 10538
rect 499488 10474 499540 10480
rect 499304 7336 499356 7342
rect 499304 7278 499356 7284
rect 499500 3398 499528 10474
rect 500420 7274 500448 16388
rect 500788 11422 500816 16388
rect 501156 14006 501184 16388
rect 501144 14000 501196 14006
rect 501144 13942 501196 13948
rect 500776 11416 500828 11422
rect 500776 11358 500828 11364
rect 500408 7268 500460 7274
rect 500408 7210 500460 7216
rect 501616 7206 501644 16388
rect 501984 11354 502012 16388
rect 502248 11824 502300 11830
rect 502248 11766 502300 11772
rect 501972 11348 502024 11354
rect 501972 11290 502024 11296
rect 501604 7200 501656 7206
rect 501604 7142 501656 7148
rect 500132 4140 500184 4146
rect 500132 4082 500184 4088
rect 498936 3392 498988 3398
rect 498936 3334 498988 3340
rect 499488 3392 499540 3398
rect 499488 3334 499540 3340
rect 496544 604 496596 610
rect 496544 546 496596 552
rect 496728 604 496780 610
rect 496728 546 496780 552
rect 497752 598 498148 626
rect 496556 480 496584 546
rect 497752 480 497780 598
rect 498948 480 498976 3334
rect 500144 480 500172 4082
rect 502260 3534 502288 11766
rect 502352 9722 502380 16388
rect 502524 14408 502576 14414
rect 502524 14350 502576 14356
rect 502340 9716 502392 9722
rect 502340 9658 502392 9664
rect 502536 6458 502564 14350
rect 502720 7138 502748 16388
rect 503088 8362 503116 16388
rect 503180 16374 503470 16402
rect 503180 14414 503208 16374
rect 503628 15156 503680 15162
rect 503628 15098 503680 15104
rect 503168 14408 503220 14414
rect 503168 14350 503220 14356
rect 503536 11892 503588 11898
rect 503536 11834 503588 11840
rect 503076 8356 503128 8362
rect 503076 8298 503128 8304
rect 502708 7132 502760 7138
rect 502708 7074 502760 7080
rect 502524 6452 502576 6458
rect 502524 6394 502576 6400
rect 502352 4146 502564 4162
rect 502340 4140 502576 4146
rect 502392 4134 502524 4140
rect 502340 4082 502392 4088
rect 502524 4082 502576 4088
rect 503548 3534 503576 11834
rect 501236 3528 501288 3534
rect 501236 3470 501288 3476
rect 502248 3528 502300 3534
rect 502248 3470 502300 3476
rect 502432 3528 502484 3534
rect 502432 3470 502484 3476
rect 503536 3528 503588 3534
rect 503536 3470 503588 3476
rect 501248 480 501276 3470
rect 502444 480 502472 3470
rect 503640 480 503668 15098
rect 503916 7070 503944 16388
rect 504284 11286 504312 16388
rect 504652 13938 504680 16388
rect 504640 13932 504692 13938
rect 504640 13874 504692 13880
rect 505020 12646 505048 16388
rect 505008 12640 505060 12646
rect 505008 12582 505060 12588
rect 504272 11280 504324 11286
rect 504272 11222 504324 11228
rect 505388 11218 505416 16388
rect 505376 11212 505428 11218
rect 505376 11154 505428 11160
rect 505756 10606 505784 16388
rect 505744 10600 505796 10606
rect 505744 10542 505796 10548
rect 503904 7064 503956 7070
rect 503904 7006 503956 7012
rect 506216 7002 506244 16388
rect 506584 11150 506612 16388
rect 506952 13326 506980 16388
rect 506940 13320 506992 13326
rect 506940 13262 506992 13268
rect 507320 13122 507348 16388
rect 507308 13116 507360 13122
rect 507308 13058 507360 13064
rect 507688 11762 507716 16388
rect 507768 14408 507820 14414
rect 507768 14350 507820 14356
rect 507676 11756 507728 11762
rect 507676 11698 507728 11704
rect 506572 11144 506624 11150
rect 506572 11086 506624 11092
rect 506204 6996 506256 7002
rect 506204 6938 506256 6944
rect 506020 6520 506072 6526
rect 506020 6462 506072 6468
rect 504824 6452 504876 6458
rect 504824 6394 504876 6400
rect 504836 480 504864 6394
rect 506032 480 506060 6462
rect 507780 3534 507808 14350
rect 508056 14074 508084 16388
rect 508044 14068 508096 14074
rect 508044 14010 508096 14016
rect 508516 13258 508544 16388
rect 508700 16374 508898 16402
rect 509266 16374 509372 16402
rect 508504 13252 508556 13258
rect 508504 13194 508556 13200
rect 508700 11694 508728 16374
rect 507860 11688 507912 11694
rect 507860 11630 507912 11636
rect 508688 11688 508740 11694
rect 508688 11630 508740 11636
rect 507872 6186 507900 11630
rect 509344 6594 509372 16374
rect 509620 12578 509648 16388
rect 509804 16374 510002 16402
rect 509608 12572 509660 12578
rect 509608 12514 509660 12520
rect 509804 11642 509832 16374
rect 509884 14000 509936 14006
rect 509884 13942 509936 13948
rect 509528 11614 509832 11642
rect 509332 6588 509384 6594
rect 509332 6530 509384 6536
rect 509528 6254 509556 11614
rect 509516 6248 509568 6254
rect 509516 6190 509568 6196
rect 507860 6180 507912 6186
rect 507860 6122 507912 6128
rect 508412 4344 508464 4350
rect 508412 4286 508464 4292
rect 507216 3528 507268 3534
rect 507216 3470 507268 3476
rect 507768 3528 507820 3534
rect 507768 3470 507820 3476
rect 507228 480 507256 3470
rect 508424 480 508452 4286
rect 509608 3528 509660 3534
rect 509608 3470 509660 3476
rect 509620 480 509648 3470
rect 509896 3466 509924 13942
rect 510356 10674 510384 16388
rect 510830 16374 510936 16402
rect 510528 13116 510580 13122
rect 510528 13058 510580 13064
rect 510344 10668 510396 10674
rect 510344 10610 510396 10616
rect 510540 3534 510568 13058
rect 510712 11688 510764 11694
rect 510712 11630 510764 11636
rect 510724 4282 510752 11630
rect 510908 4962 510936 16374
rect 511184 7614 511212 16388
rect 511552 14482 511580 16388
rect 511644 16374 511934 16402
rect 511540 14476 511592 14482
rect 511540 14418 511592 14424
rect 511264 13932 511316 13938
rect 511264 13874 511316 13880
rect 511172 7608 511224 7614
rect 511172 7550 511224 7556
rect 510896 4956 510948 4962
rect 510896 4898 510948 4904
rect 510712 4276 510764 4282
rect 510712 4218 510764 4224
rect 510528 3528 510580 3534
rect 510528 3470 510580 3476
rect 509884 3460 509936 3466
rect 509884 3402 509936 3408
rect 510804 3460 510856 3466
rect 510804 3402 510856 3408
rect 510816 480 510844 3402
rect 511276 3398 511304 13874
rect 511644 11694 511672 16374
rect 511632 11688 511684 11694
rect 511632 11630 511684 11636
rect 512288 7682 512316 16388
rect 512656 14006 512684 16388
rect 512644 14000 512696 14006
rect 512644 13942 512696 13948
rect 512276 7676 512328 7682
rect 512276 7618 512328 7624
rect 512000 7608 512052 7614
rect 512748 7562 512776 16510
rect 513484 7750 513512 16388
rect 513564 14476 513616 14482
rect 513564 14418 513616 14424
rect 513472 7744 513524 7750
rect 513472 7686 513524 7692
rect 513196 7676 513248 7682
rect 513196 7618 513248 7624
rect 512000 7550 512052 7556
rect 511264 3392 511316 3398
rect 511264 3334 511316 3340
rect 512012 480 512040 7550
rect 512104 7534 512776 7562
rect 512104 4214 512132 7534
rect 512092 4208 512144 4214
rect 512092 4150 512144 4156
rect 513208 480 513236 7618
rect 513576 4826 513604 14418
rect 513852 13938 513880 16388
rect 514036 16374 514234 16402
rect 514036 14482 514064 16374
rect 514024 14476 514076 14482
rect 514024 14418 514076 14424
rect 514024 14340 514076 14346
rect 514024 14282 514076 14288
rect 513840 13932 513892 13938
rect 513840 13874 513892 13880
rect 513564 4820 513616 4826
rect 513564 4762 513616 4768
rect 514036 3874 514064 14282
rect 514588 7818 514616 16388
rect 514956 14550 514984 16388
rect 515140 16374 515430 16402
rect 514944 14544 514996 14550
rect 514944 14486 514996 14492
rect 514576 7812 514628 7818
rect 514576 7754 514628 7760
rect 515140 4894 515168 16374
rect 515784 7886 515812 16388
rect 516166 16374 516272 16402
rect 516048 13252 516100 13258
rect 516048 13194 516100 13200
rect 515772 7880 515824 7886
rect 515772 7822 515824 7828
rect 515128 4888 515180 4894
rect 515128 4830 515180 4836
rect 516060 4146 516088 13194
rect 515588 4140 515640 4146
rect 515588 4082 515640 4088
rect 516048 4140 516100 4146
rect 516048 4082 516100 4088
rect 514024 3868 514076 3874
rect 514024 3810 514076 3816
rect 514392 3392 514444 3398
rect 514392 3334 514444 3340
rect 514404 480 514432 3334
rect 515600 480 515628 4082
rect 516244 3602 516272 16374
rect 516336 5030 516364 16510
rect 516888 13190 516916 16388
rect 517256 14618 517284 16388
rect 517244 14612 517296 14618
rect 517244 14554 517296 14560
rect 517428 14476 517480 14482
rect 517428 14418 517480 14424
rect 516876 13184 516928 13190
rect 516876 13126 516928 13132
rect 516324 5024 516376 5030
rect 516324 4966 516376 4972
rect 517440 4146 517468 14418
rect 517716 5098 517744 16388
rect 518084 8974 518112 16388
rect 518176 16374 518466 16402
rect 518544 16374 518834 16402
rect 519004 16374 519202 16402
rect 518072 8968 518124 8974
rect 518072 8910 518124 8916
rect 517704 5092 517756 5098
rect 517704 5034 517756 5040
rect 516784 4140 516836 4146
rect 516784 4082 516836 4088
rect 517428 4140 517480 4146
rect 517428 4082 517480 4088
rect 516232 3596 516284 3602
rect 516232 3538 516284 3544
rect 516796 480 516824 4082
rect 517888 4072 517940 4078
rect 517888 4014 517940 4020
rect 517900 480 517928 4014
rect 518176 3670 518204 16374
rect 518348 14000 518400 14006
rect 518348 13942 518400 13948
rect 518360 4146 518388 13942
rect 518544 5166 518572 16374
rect 519004 9042 519032 16374
rect 519556 13870 519584 16388
rect 519648 16374 520030 16402
rect 520292 16374 520398 16402
rect 520568 16374 520766 16402
rect 520844 16374 521134 16402
rect 519544 13864 519596 13870
rect 519544 13806 519596 13812
rect 518992 9036 519044 9042
rect 518992 8978 519044 8984
rect 519084 6180 519136 6186
rect 519084 6122 519136 6128
rect 518532 5160 518584 5166
rect 518532 5102 518584 5108
rect 518348 4140 518400 4146
rect 518348 4082 518400 4088
rect 518164 3664 518216 3670
rect 518164 3606 518216 3612
rect 519096 480 519124 6122
rect 519648 5234 519676 16374
rect 519728 14136 519780 14142
rect 519728 14078 519780 14084
rect 519636 5228 519688 5234
rect 519636 5170 519688 5176
rect 519740 3874 519768 14078
rect 520292 9110 520320 16374
rect 520280 9104 520332 9110
rect 520280 9046 520332 9052
rect 520280 4140 520332 4146
rect 520280 4082 520332 4088
rect 519728 3868 519780 3874
rect 519728 3810 519780 3816
rect 520292 480 520320 4082
rect 520568 3738 520596 16374
rect 520844 5302 520872 16374
rect 520924 14272 520976 14278
rect 520924 14214 520976 14220
rect 520832 5296 520884 5302
rect 520832 5238 520884 5244
rect 520556 3732 520608 3738
rect 520556 3674 520608 3680
rect 520936 3466 520964 14214
rect 521488 9178 521516 16388
rect 521568 14544 521620 14550
rect 521568 14486 521620 14492
rect 521476 9172 521528 9178
rect 521476 9114 521528 9120
rect 521580 4146 521608 14486
rect 521856 14346 521884 16388
rect 521948 16374 522330 16402
rect 521844 14340 521896 14346
rect 521844 14282 521896 14288
rect 521948 5370 521976 16374
rect 522304 14340 522356 14346
rect 522304 14282 522356 14288
rect 521936 5364 521988 5370
rect 521936 5306 521988 5312
rect 521568 4140 521620 4146
rect 521568 4082 521620 4088
rect 520924 3460 520976 3466
rect 520924 3402 520976 3408
rect 522316 3398 522344 14282
rect 522684 9246 522712 16388
rect 523066 16374 523264 16402
rect 522672 9240 522724 9246
rect 522672 9182 522724 9188
rect 523236 3806 523264 16374
rect 523328 16374 523434 16402
rect 523328 5438 523356 16374
rect 523684 14680 523736 14686
rect 523684 14622 523736 14628
rect 523316 5432 523368 5438
rect 523316 5374 523368 5380
rect 523696 4078 523724 14622
rect 523788 13394 523816 16388
rect 524156 14618 524184 16388
rect 524524 16374 524630 16402
rect 524708 16374 524998 16402
rect 525076 16374 525366 16402
rect 525444 16374 525734 16402
rect 525904 16374 526102 16402
rect 524144 14612 524196 14618
rect 524144 14554 524196 14560
rect 524328 14612 524380 14618
rect 524328 14554 524380 14560
rect 523776 13388 523828 13394
rect 523776 13330 523828 13336
rect 524340 4146 524368 14554
rect 524420 11756 524472 11762
rect 524420 11698 524472 11704
rect 524432 6322 524460 11698
rect 524420 6316 524472 6322
rect 524420 6258 524472 6264
rect 524524 5506 524552 16374
rect 524708 11762 524736 16374
rect 524696 11756 524748 11762
rect 524696 11698 524748 11704
rect 524604 11688 524656 11694
rect 525076 11642 525104 16374
rect 525156 14204 525208 14210
rect 525156 14146 525208 14152
rect 524604 11630 524656 11636
rect 524512 5500 524564 5506
rect 524512 5442 524564 5448
rect 524616 4758 524644 11630
rect 524708 11614 525104 11642
rect 524604 4752 524656 4758
rect 524604 4694 524656 4700
rect 523868 4140 523920 4146
rect 523868 4082 523920 4088
rect 524328 4140 524380 4146
rect 524328 4082 524380 4088
rect 523684 4072 523736 4078
rect 523684 4014 523736 4020
rect 523224 3800 523276 3806
rect 523224 3742 523276 3748
rect 522672 3460 522724 3466
rect 522672 3402 522724 3408
rect 522304 3392 522356 3398
rect 522304 3334 522356 3340
rect 521476 3324 521528 3330
rect 521476 3266 521528 3272
rect 521488 480 521516 3266
rect 522684 480 522712 3402
rect 523880 480 523908 4082
rect 524708 3942 524736 11614
rect 525168 10554 525196 14146
rect 525444 11694 525472 16374
rect 525432 11688 525484 11694
rect 525432 11630 525484 11636
rect 524984 10526 525196 10554
rect 524696 3936 524748 3942
rect 524696 3878 524748 3884
rect 524984 3330 525012 10526
rect 525904 6390 525932 16374
rect 526456 14754 526484 16388
rect 526548 16374 526930 16402
rect 526444 14748 526496 14754
rect 526444 14690 526496 14696
rect 526548 11642 526576 16374
rect 527284 14822 527312 16388
rect 527376 16374 527666 16402
rect 527744 16374 528034 16402
rect 527272 14816 527324 14822
rect 527272 14758 527324 14764
rect 526628 14748 526680 14754
rect 526628 14690 526680 14696
rect 525996 11614 526576 11642
rect 525892 6384 525944 6390
rect 525892 6326 525944 6332
rect 525996 4690 526024 11614
rect 526640 10826 526668 14690
rect 527272 11688 527324 11694
rect 527272 11630 527324 11636
rect 526364 10798 526668 10826
rect 525984 4684 526036 4690
rect 525984 4626 526036 4632
rect 526260 3596 526312 3602
rect 526260 3538 526312 3544
rect 525064 3528 525116 3534
rect 525064 3470 525116 3476
rect 524972 3324 525024 3330
rect 524972 3266 525024 3272
rect 525076 480 525104 3470
rect 526272 480 526300 3538
rect 526364 3534 526392 10798
rect 527284 4622 527312 11630
rect 527272 4616 527324 4622
rect 527272 4558 527324 4564
rect 527376 4010 527404 16374
rect 527744 11694 527772 16374
rect 527732 11688 527784 11694
rect 527732 11630 527784 11636
rect 528388 10334 528416 16388
rect 528756 14890 528784 16388
rect 528744 14884 528796 14890
rect 528744 14826 528796 14832
rect 528468 14068 528520 14074
rect 528468 14010 528520 14016
rect 528376 10328 528428 10334
rect 528376 10270 528428 10276
rect 527364 4004 527416 4010
rect 527364 3946 527416 3952
rect 526352 3528 526404 3534
rect 526352 3470 526404 3476
rect 528480 3466 528508 14010
rect 528836 12572 528888 12578
rect 528836 12514 528888 12520
rect 528848 11642 528876 12514
rect 528756 11614 528876 11642
rect 528756 4554 528784 11614
rect 529216 9314 529244 16388
rect 529308 16374 529598 16402
rect 529308 12578 529336 16374
rect 529952 14958 529980 16388
rect 529940 14952 529992 14958
rect 529940 14894 529992 14900
rect 529848 14816 529900 14822
rect 529848 14758 529900 14764
rect 529296 12572 529348 12578
rect 529296 12514 529348 12520
rect 529204 9308 529256 9314
rect 529204 9250 529256 9256
rect 528744 4548 528796 4554
rect 528744 4490 528796 4496
rect 529860 3534 529888 14758
rect 530320 10402 530348 16388
rect 530308 10396 530360 10402
rect 530308 10338 530360 10344
rect 530688 9722 530716 16388
rect 531056 15094 531084 16388
rect 531044 15088 531096 15094
rect 531044 15030 531096 15036
rect 531228 14952 531280 14958
rect 531228 14894 531280 14900
rect 530124 9716 530176 9722
rect 530124 9658 530176 9664
rect 530676 9716 530728 9722
rect 530676 9658 530728 9664
rect 530136 4486 530164 9658
rect 530124 4480 530176 4486
rect 530124 4422 530176 4428
rect 528652 3528 528704 3534
rect 528652 3470 528704 3476
rect 529848 3528 529900 3534
rect 531240 3482 531268 14894
rect 531516 13462 531544 16388
rect 531700 16374 531898 16402
rect 531504 13456 531556 13462
rect 531504 13398 531556 13404
rect 531700 11642 531728 16374
rect 532252 14006 532280 16388
rect 532344 16374 532634 16402
rect 532240 14000 532292 14006
rect 532240 13942 532292 13948
rect 531516 11614 531728 11642
rect 531516 4418 531544 11614
rect 532344 9450 532372 16374
rect 532608 14884 532660 14890
rect 532608 14826 532660 14832
rect 532332 9444 532384 9450
rect 532332 9386 532384 9392
rect 531504 4412 531556 4418
rect 531504 4354 531556 4360
rect 532620 3482 532648 14826
rect 532988 9382 533016 16388
rect 533356 15026 533384 16388
rect 533344 15020 533396 15026
rect 533344 14962 533396 14968
rect 533816 10470 533844 16388
rect 533988 15020 534040 15026
rect 533988 14962 534040 14968
rect 533804 10464 533856 10470
rect 533804 10406 533856 10412
rect 532976 9376 533028 9382
rect 532976 9318 533028 9324
rect 533252 8968 533304 8974
rect 533252 8910 533304 8916
rect 533264 3602 533292 8910
rect 533252 3596 533304 3602
rect 533252 3538 533304 3544
rect 534000 3534 534028 14962
rect 534184 10538 534212 16388
rect 534552 14142 534580 16388
rect 534540 14136 534592 14142
rect 534540 14078 534592 14084
rect 534920 11830 534948 16388
rect 535288 11898 535316 16388
rect 535656 15162 535684 16388
rect 535748 16374 536130 16402
rect 536300 16374 536498 16402
rect 535644 15156 535696 15162
rect 535644 15098 535696 15104
rect 535368 15088 535420 15094
rect 535368 15030 535420 15036
rect 535276 11892 535328 11898
rect 535276 11834 535328 11840
rect 534908 11824 534960 11830
rect 534908 11766 534960 11772
rect 534724 11756 534776 11762
rect 534724 11698 534776 11704
rect 534172 10532 534224 10538
rect 534172 10474 534224 10480
rect 529848 3470 529900 3476
rect 527456 3460 527508 3466
rect 527456 3402 527508 3408
rect 528468 3460 528520 3466
rect 528468 3402 528520 3408
rect 527468 480 527496 3402
rect 528664 480 528692 3470
rect 531056 3454 531268 3482
rect 532252 3454 532648 3482
rect 533436 3528 533488 3534
rect 533436 3470 533488 3476
rect 533988 3528 534040 3534
rect 533988 3470 534040 3476
rect 534540 3528 534592 3534
rect 534540 3470 534592 3476
rect 529848 3392 529900 3398
rect 529848 3334 529900 3340
rect 529860 480 529888 3334
rect 531056 480 531084 3454
rect 532252 480 532280 3454
rect 533448 480 533476 3470
rect 534552 480 534580 3470
rect 534736 3330 534764 11698
rect 535380 3534 535408 15030
rect 535748 11642 535776 16374
rect 535564 11614 535776 11642
rect 535564 6458 535592 11614
rect 536300 11506 536328 16374
rect 536852 14414 536880 16388
rect 537036 16374 537234 16402
rect 536840 14408 536892 14414
rect 536840 14350 536892 14356
rect 536748 14136 536800 14142
rect 536748 14078 536800 14084
rect 535656 11478 536328 11506
rect 535656 6526 535684 11478
rect 535644 6520 535696 6526
rect 535644 6462 535696 6468
rect 535552 6452 535604 6458
rect 535552 6394 535604 6400
rect 535368 3528 535420 3534
rect 535368 3470 535420 3476
rect 536760 3330 536788 14078
rect 537036 4350 537064 16374
rect 537588 13122 537616 16388
rect 537956 14278 537984 16388
rect 538128 15156 538180 15162
rect 538128 15098 538180 15104
rect 537944 14272 537996 14278
rect 537944 14214 537996 14220
rect 537576 13116 537628 13122
rect 537576 13058 537628 13064
rect 537024 4344 537076 4350
rect 537024 4286 537076 4292
rect 536932 3596 536984 3602
rect 536932 3538 536984 3544
rect 534724 3324 534776 3330
rect 534724 3266 534776 3272
rect 535736 3324 535788 3330
rect 535736 3266 535788 3272
rect 536748 3324 536800 3330
rect 536748 3266 536800 3272
rect 535748 480 535776 3266
rect 536944 480 536972 3538
rect 538140 480 538168 15098
rect 538416 7614 538444 16388
rect 538784 7682 538812 16388
rect 539152 14346 539180 16388
rect 539140 14340 539192 14346
rect 539140 14282 539192 14288
rect 539520 13258 539548 16388
rect 539888 14482 539916 16388
rect 540256 14686 540284 16388
rect 540532 16374 540730 16402
rect 540244 14680 540296 14686
rect 540244 14622 540296 14628
rect 539876 14476 539928 14482
rect 539876 14418 539928 14424
rect 539508 13252 539560 13258
rect 539508 13194 539560 13200
rect 538772 7676 538824 7682
rect 538772 7618 538824 7624
rect 538404 7608 538456 7614
rect 538404 7550 538456 7556
rect 540532 6934 540560 16374
rect 541084 14550 541112 16388
rect 541072 14544 541124 14550
rect 541072 14486 541124 14492
rect 541452 14210 541480 16388
rect 541440 14204 541492 14210
rect 541440 14146 541492 14152
rect 541820 11762 541848 16388
rect 542188 14618 542216 16388
rect 542556 14754 542584 16388
rect 542544 14748 542596 14754
rect 542544 14690 542596 14696
rect 542176 14612 542228 14618
rect 542176 14554 542228 14560
rect 541808 11756 541860 11762
rect 541808 11698 541860 11704
rect 543016 8974 543044 16388
rect 543384 14074 543412 16388
rect 543752 14822 543780 16388
rect 543936 16374 544134 16402
rect 543740 14816 543792 14822
rect 543740 14758 543792 14764
rect 543648 14204 543700 14210
rect 543648 14146 543700 14152
rect 543372 14068 543424 14074
rect 543372 14010 543424 14016
rect 543004 8968 543056 8974
rect 543004 8910 543056 8916
rect 539600 6928 539652 6934
rect 539600 6870 539652 6876
rect 540520 6928 540572 6934
rect 540520 6870 540572 6876
rect 539612 6186 539640 6870
rect 539600 6180 539652 6186
rect 539600 6122 539652 6128
rect 543660 3466 543688 14146
rect 543936 3534 543964 16374
rect 544488 14958 544516 16388
rect 544476 14952 544528 14958
rect 544476 14894 544528 14900
rect 544856 14890 544884 16388
rect 545316 15026 545344 16388
rect 545684 15094 545712 16388
rect 545672 15088 545724 15094
rect 545672 15030 545724 15036
rect 545304 15020 545356 15026
rect 545304 14962 545356 14968
rect 544844 14884 544896 14890
rect 544844 14826 544896 14832
rect 544384 14408 544436 14414
rect 544384 14350 544436 14356
rect 544108 3732 544160 3738
rect 544108 3674 544160 3680
rect 543924 3528 543976 3534
rect 543924 3470 543976 3476
rect 542912 3460 542964 3466
rect 542912 3402 542964 3408
rect 543648 3460 543700 3466
rect 543648 3402 543700 3408
rect 539324 3392 539376 3398
rect 539324 3334 539376 3340
rect 539336 480 539364 3334
rect 541716 3256 541768 3262
rect 541716 3198 541768 3204
rect 540520 2916 540572 2922
rect 540520 2858 540572 2864
rect 540532 480 540560 2858
rect 541728 480 541756 3198
rect 542924 480 542952 3402
rect 544120 480 544148 3674
rect 544396 3602 544424 14350
rect 546052 14278 546080 16388
rect 546316 14544 546368 14550
rect 546316 14486 546368 14492
rect 546040 14272 546092 14278
rect 546040 14214 546092 14220
rect 545764 14204 545816 14210
rect 545764 14146 545816 14152
rect 545028 14068 545080 14074
rect 545028 14010 545080 14016
rect 545040 3738 545068 14010
rect 545304 3868 545356 3874
rect 545304 3810 545356 3816
rect 545028 3732 545080 3738
rect 545028 3674 545080 3680
rect 544384 3596 544436 3602
rect 544384 3538 544436 3544
rect 545316 480 545344 3810
rect 545776 3398 545804 14146
rect 546328 3874 546356 14486
rect 546420 14414 546448 16388
rect 546788 15162 546816 16388
rect 546776 15156 546828 15162
rect 546776 15098 546828 15104
rect 546408 14408 546460 14414
rect 546408 14350 546460 14356
rect 547156 14210 547184 16388
rect 547340 16374 547630 16402
rect 547998 16374 548104 16402
rect 547144 14204 547196 14210
rect 547144 14146 547196 14152
rect 546316 3868 546368 3874
rect 546316 3810 546368 3816
rect 545764 3392 545816 3398
rect 545764 3334 545816 3340
rect 546500 3392 546552 3398
rect 546500 3334 546552 3340
rect 546512 480 546540 3334
rect 547340 2922 547368 16374
rect 547788 14476 547840 14482
rect 547788 14418 547840 14424
rect 547696 14408 547748 14414
rect 547696 14350 547748 14356
rect 547708 3398 547736 14350
rect 547696 3392 547748 3398
rect 547696 3334 547748 3340
rect 547800 3210 547828 14418
rect 548076 3262 548104 16374
rect 548352 14346 548380 16388
rect 548340 14340 548392 14346
rect 548340 14282 548392 14288
rect 548720 14074 548748 16388
rect 549088 14550 549116 16388
rect 549076 14544 549128 14550
rect 549076 14486 549128 14492
rect 549456 14414 549484 16388
rect 549916 14482 549944 16388
rect 549904 14476 549956 14482
rect 549904 14418 549956 14424
rect 549444 14408 549496 14414
rect 549444 14350 549496 14356
rect 548708 14068 548760 14074
rect 548708 14010 548760 14016
rect 550284 9722 550312 16388
rect 550652 13954 550680 16388
rect 550560 13926 550680 13954
rect 550836 16374 551034 16402
rect 548892 9716 548944 9722
rect 548892 9658 548944 9664
rect 550272 9716 550324 9722
rect 550272 9658 550324 9664
rect 547708 3182 547828 3210
rect 548064 3256 548116 3262
rect 548064 3198 548116 3204
rect 547328 2916 547380 2922
rect 547328 2858 547380 2864
rect 547708 480 547736 3182
rect 548904 480 548932 9658
rect 550560 4146 550588 13926
rect 550088 4140 550140 4146
rect 550088 4082 550140 4088
rect 550548 4140 550600 4146
rect 550548 4082 550600 4088
rect 550100 480 550128 4082
rect 550836 2854 550864 16374
rect 551388 14414 551416 16388
rect 551376 14408 551428 14414
rect 551376 14350 551428 14356
rect 551756 13870 551784 16388
rect 551928 14408 551980 14414
rect 551928 14350 551980 14356
rect 551744 13864 551796 13870
rect 551744 13806 551796 13812
rect 551940 4146 551968 14350
rect 552216 11354 552244 16388
rect 552584 14142 552612 16388
rect 552572 14136 552624 14142
rect 552572 14078 552624 14084
rect 552952 14074 552980 16388
rect 552940 14068 552992 14074
rect 552940 14010 552992 14016
rect 553320 14006 553348 16388
rect 553688 14278 553716 16388
rect 553676 14272 553728 14278
rect 553676 14214 553728 14220
rect 554056 14210 554084 16388
rect 554044 14204 554096 14210
rect 554044 14146 554096 14152
rect 553308 14000 553360 14006
rect 553308 13942 553360 13948
rect 554516 13870 554544 16388
rect 554884 14550 554912 16388
rect 555252 14958 555280 16388
rect 555240 14952 555292 14958
rect 555240 14894 555292 14900
rect 554872 14544 554924 14550
rect 554872 14486 554924 14492
rect 555240 14136 555292 14142
rect 555240 14078 555292 14084
rect 553400 13864 553452 13870
rect 553400 13806 553452 13812
rect 554504 13864 554556 13870
rect 554504 13806 554556 13812
rect 552204 11348 552256 11354
rect 552204 11290 552256 11296
rect 551928 4140 551980 4146
rect 551928 4082 551980 4088
rect 552388 4140 552440 4146
rect 552388 4082 552440 4088
rect 550824 2848 550876 2854
rect 550824 2790 550876 2796
rect 551192 2780 551244 2786
rect 551192 2722 551244 2728
rect 551204 480 551232 2722
rect 552400 480 552428 4082
rect 553412 2854 553440 13806
rect 555252 12442 555280 14078
rect 555424 14068 555476 14074
rect 555424 14010 555476 14016
rect 555240 12436 555292 12442
rect 555240 12378 555292 12384
rect 554964 11348 555016 11354
rect 554964 11290 555016 11296
rect 553400 2848 553452 2854
rect 553400 2790 553452 2796
rect 553584 2780 553636 2786
rect 553584 2722 553636 2728
rect 553596 480 553624 2722
rect 554976 610 555004 11290
rect 555436 4146 555464 14010
rect 555516 14000 555568 14006
rect 555516 13942 555568 13948
rect 555424 4140 555476 4146
rect 555424 4082 555476 4088
rect 555528 4010 555556 13942
rect 555620 13938 555648 16388
rect 556002 16374 556108 16402
rect 555608 13932 555660 13938
rect 555608 13874 555660 13880
rect 555976 13932 556028 13938
rect 555976 13874 556028 13880
rect 555884 12436 555936 12442
rect 555884 12378 555936 12384
rect 555516 4004 555568 4010
rect 555516 3946 555568 3952
rect 555896 2938 555924 12378
rect 555988 3126 556016 13874
rect 556080 3194 556108 16374
rect 556356 13938 556384 16388
rect 556344 13932 556396 13938
rect 556344 13874 556396 13880
rect 556816 13870 556844 16388
rect 557198 16374 557304 16402
rect 556988 14272 557040 14278
rect 556988 14214 557040 14220
rect 556896 14204 556948 14210
rect 556896 14146 556948 14152
rect 556712 13864 556764 13870
rect 556712 13806 556764 13812
rect 556804 13864 556856 13870
rect 556804 13806 556856 13812
rect 556724 3602 556752 13806
rect 556908 3670 556936 14146
rect 557000 4078 557028 14214
rect 557172 4140 557224 4146
rect 557172 4082 557224 4088
rect 556988 4072 557040 4078
rect 556988 4014 557040 4020
rect 556896 3664 556948 3670
rect 556896 3606 556948 3612
rect 556712 3596 556764 3602
rect 556712 3538 556764 3544
rect 556068 3188 556120 3194
rect 556068 3130 556120 3136
rect 555976 3120 556028 3126
rect 555976 3062 556028 3068
rect 555896 2910 556016 2938
rect 554780 604 554832 610
rect 554780 546 554832 552
rect 554964 604 555016 610
rect 554964 546 555016 552
rect 554792 480 554820 546
rect 555988 480 556016 2910
rect 557184 480 557212 4082
rect 557276 3942 557304 16374
rect 557552 13938 557580 16388
rect 557356 13932 557408 13938
rect 557356 13874 557408 13880
rect 557540 13932 557592 13938
rect 557540 13874 557592 13880
rect 557264 3936 557316 3942
rect 557264 3878 557316 3884
rect 557368 3262 557396 13874
rect 557920 13870 557948 16388
rect 558302 16374 558592 16402
rect 558670 16374 558776 16402
rect 557448 13864 557500 13870
rect 557448 13806 557500 13812
rect 557908 13864 557960 13870
rect 557908 13806 557960 13812
rect 557460 3330 557488 13806
rect 558368 4004 558420 4010
rect 558368 3946 558420 3952
rect 557448 3324 557500 3330
rect 557448 3266 557500 3272
rect 557356 3256 557408 3262
rect 557356 3198 557408 3204
rect 558380 480 558408 3946
rect 558564 3738 558592 16374
rect 558644 13864 558696 13870
rect 558644 13806 558696 13812
rect 558656 4146 558684 13806
rect 558644 4140 558696 4146
rect 558644 4082 558696 4088
rect 558748 3874 558776 16374
rect 559116 13938 559144 16388
rect 559498 16374 559788 16402
rect 558828 13932 558880 13938
rect 558828 13874 558880 13880
rect 559104 13932 559156 13938
rect 559104 13874 559156 13880
rect 558736 3868 558788 3874
rect 558736 3810 558788 3816
rect 558552 3732 558604 3738
rect 558552 3674 558604 3680
rect 558840 3058 558868 13874
rect 559564 4072 559616 4078
rect 559564 4014 559616 4020
rect 558828 3052 558880 3058
rect 558828 2994 558880 3000
rect 559576 480 559604 4014
rect 559760 3806 559788 16374
rect 559852 13870 559880 16388
rect 560036 16374 560234 16402
rect 559840 13864 559892 13870
rect 559840 13806 559892 13812
rect 559748 3800 559800 3806
rect 559748 3742 559800 3748
rect 560036 3398 560064 16374
rect 560116 13932 560168 13938
rect 560116 13874 560168 13880
rect 560128 3942 560156 13874
rect 560588 13870 560616 16388
rect 560970 16374 561628 16402
rect 560208 13864 560260 13870
rect 560208 13806 560260 13812
rect 560576 13864 560628 13870
rect 560576 13806 560628 13812
rect 561496 13864 561548 13870
rect 561496 13806 561548 13812
rect 560116 3936 560168 3942
rect 560116 3878 560168 3884
rect 560220 3738 560248 13806
rect 560208 3732 560260 3738
rect 560208 3674 560260 3680
rect 560760 3664 560812 3670
rect 560760 3606 560812 3612
rect 560024 3392 560076 3398
rect 560024 3334 560076 3340
rect 560772 480 560800 3606
rect 561508 3466 561536 13806
rect 561600 3670 561628 16374
rect 563060 14952 563112 14958
rect 563060 14894 563112 14900
rect 561588 3664 561640 3670
rect 561588 3606 561640 3612
rect 561956 3596 562008 3602
rect 561956 3538 562008 3544
rect 561496 3460 561548 3466
rect 561496 3402 561548 3408
rect 561968 480 561996 3538
rect 563072 3534 563100 14894
rect 563152 14544 563204 14550
rect 563152 14486 563204 14492
rect 563060 3528 563112 3534
rect 563060 3470 563112 3476
rect 563164 480 563192 14486
rect 563716 3602 563744 38655
rect 580920 29345 580948 76191
rect 580906 29336 580962 29345
rect 580906 29271 580962 29280
rect 572628 4140 572680 4146
rect 572628 4082 572680 4088
rect 570236 4072 570288 4078
rect 570236 4014 570288 4020
rect 563704 3596 563756 3602
rect 563704 3538 563756 3544
rect 564348 3528 564400 3534
rect 564348 3470 564400 3476
rect 564360 480 564388 3470
rect 569040 3324 569092 3330
rect 569040 3266 569092 3272
rect 567844 3256 567896 3262
rect 567844 3198 567896 3204
rect 566740 3188 566792 3194
rect 566740 3130 566792 3136
rect 565544 3120 565596 3126
rect 565544 3062 565596 3068
rect 565556 480 565584 3062
rect 566752 480 566780 3130
rect 567856 480 567884 3198
rect 569052 480 569080 3266
rect 570248 480 570276 4014
rect 571432 3392 571484 3398
rect 571432 3334 571484 3340
rect 571444 480 571472 3334
rect 572640 480 572668 4082
rect 573824 4004 573876 4010
rect 573824 3946 573876 3952
rect 573836 480 573864 3946
rect 576216 3936 576268 3942
rect 576216 3878 576268 3884
rect 575020 3868 575072 3874
rect 575020 3810 575072 3816
rect 575032 480 575060 3810
rect 576228 480 576256 3878
rect 577412 3800 577464 3806
rect 577412 3742 577464 3748
rect 577424 480 577452 3742
rect 578608 3732 578660 3738
rect 578608 3674 578660 3680
rect 578620 480 578648 3674
rect 582196 3664 582248 3670
rect 582196 3606 582248 3612
rect 581000 3528 581052 3534
rect 581000 3470 581052 3476
rect 579804 3460 579856 3466
rect 579804 3402 579856 3408
rect 579816 480 579844 3402
rect 581012 480 581040 3470
rect 582208 480 582236 3606
rect 583392 3596 583444 3602
rect 583392 3538 583444 3544
rect 583404 480 583432 3538
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3514 682216 3570 682272
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 3054 653520 3110 653576
rect 3422 624824 3478 624880
rect 3330 610408 3386 610464
rect 3146 553016 3202 553072
rect 2870 509904 2926 509960
rect 3514 595992 3570 596048
rect 3514 567296 3570 567352
rect 3514 538600 3570 538656
rect 3514 495508 3570 495544
rect 3514 495488 3516 495508
rect 3516 495488 3568 495508
rect 3568 495488 3570 495508
rect 3146 481072 3202 481128
rect 3422 452376 3478 452432
rect 3422 437960 3478 438016
rect 2778 380568 2834 380624
rect 2778 366152 2834 366208
rect 3146 337456 3202 337512
rect 2778 323040 2834 323096
rect 2778 309032 2834 309088
rect 2778 308760 2834 308816
rect 2778 280064 2834 280120
rect 2778 265648 2834 265704
rect 2778 236952 2834 237008
rect 2778 222536 2834 222592
rect 2778 193840 2834 193896
rect 2778 179424 2834 179480
rect 2778 150728 2834 150784
rect 2778 136312 2834 136368
rect 2778 107616 2834 107672
rect 2778 93200 2834 93256
rect 2778 64504 2834 64560
rect 2778 50088 2834 50144
rect 3514 423700 3570 423736
rect 3514 423680 3516 423700
rect 3516 423680 3568 423700
rect 3568 423680 3570 423700
rect 4802 394984 4858 395040
rect 3514 309032 3570 309088
rect 3606 294344 3662 294400
rect 4802 173712 4858 173768
rect 6182 65456 6238 65512
rect 3514 35808 3570 35864
rect 2778 21392 2834 21448
rect 2778 7112 2834 7168
rect 12530 443536 12586 443592
rect 116582 622376 116638 622432
rect 28630 611496 28686 611552
rect 27710 609592 27766 609648
rect 27526 608912 27582 608968
rect 27158 607144 27214 607200
rect 27066 601160 27122 601216
rect 26974 598712 27030 598768
rect 24950 593952 25006 594008
rect 24858 572872 24914 572928
rect 24766 572328 24822 572384
rect 24674 571804 24730 571840
rect 24674 571784 24676 571804
rect 24676 571784 24728 571804
rect 24728 571784 24730 571804
rect 26054 592728 26110 592784
rect 25870 591504 25926 591560
rect 25778 587968 25834 588024
rect 25686 585520 25742 585576
rect 25502 584296 25558 584352
rect 25318 583072 25374 583128
rect 25226 581984 25282 582040
rect 25134 580760 25190 580816
rect 25042 579536 25098 579592
rect 25410 581304 25466 581360
rect 25594 583752 25650 583808
rect 25962 589736 26018 589792
rect 26790 596400 26846 596456
rect 26698 592184 26754 592240
rect 26606 584976 26662 585032
rect 26514 582528 26570 582584
rect 26422 578856 26478 578912
rect 26146 578312 26202 578368
rect 26238 574096 26294 574152
rect 26330 573552 26386 573608
rect 26882 595176 26938 595232
rect 27434 606600 27490 606656
rect 27250 605920 27306 605976
rect 27342 604152 27398 604208
rect 27618 608368 27674 608424
rect 28630 607280 28686 607336
rect 27802 605376 27858 605432
rect 28538 602520 28594 602576
rect 27894 601976 27950 602032
rect 28078 601840 28134 601896
rect 27986 597624 28042 597680
rect 28630 600208 28686 600264
rect 28538 598848 28594 598904
rect 28170 597080 28226 597136
rect 28630 597080 28686 597136
rect 28446 595312 28502 595368
rect 28262 594088 28318 594144
rect 28354 592864 28410 592920
rect 28538 590416 28594 590472
rect 28446 588648 28502 588704
rect 28630 590008 28686 590064
rect 28262 588104 28318 588160
rect 28354 586880 28410 586936
rect 28630 586880 28686 586936
rect 28630 585656 28686 585712
rect 28630 579672 28686 579728
rect 28630 577224 28686 577280
rect 28630 576680 28686 576736
rect 28630 576000 28686 576056
rect 28630 575084 28632 575104
rect 28632 575084 28684 575104
rect 28684 575084 28686 575104
rect 28630 575048 28686 575084
rect 28630 574948 28632 574968
rect 28632 574948 28684 574968
rect 28684 574948 28686 574968
rect 28630 574912 28686 574948
rect 29182 571512 29238 571568
rect 73802 532616 73858 532672
rect 279146 618296 279202 618352
rect 139582 594768 139638 594824
rect 80242 533568 80298 533624
rect 82450 533432 82506 533488
rect 100758 559544 100814 559600
rect 90546 554104 90602 554160
rect 90362 553968 90418 554024
rect 92110 530848 92166 530904
rect 93214 530712 93270 530768
rect 94226 530576 94282 530632
rect 97538 533296 97594 533352
rect 96434 532480 96490 532536
rect 98550 532344 98606 532400
rect 100758 532208 100814 532264
rect 102874 532072 102930 532128
rect 103978 531936 104034 531992
rect 106094 529896 106150 529952
rect 119066 530168 119122 530224
rect 115846 530032 115902 530088
rect 141698 531392 141754 531448
rect 154670 532752 154726 532808
rect 153566 531528 153622 531584
rect 155682 531664 155738 531720
rect 166446 532888 166502 532944
rect 162214 531800 162270 531856
rect 175094 533160 175150 533216
rect 170770 533024 170826 533080
rect 188066 531936 188122 531992
rect 280158 563760 280214 563816
rect 280158 553152 280214 553208
rect 107566 528536 107622 528592
rect 115110 528264 115166 528320
rect 115938 528284 115994 528320
rect 115938 528264 115940 528284
rect 115940 528264 115992 528284
rect 115992 528264 115994 528284
rect 125322 528162 125378 528218
rect 21362 492496 21418 492552
rect 104898 497392 104954 497448
rect 107198 499976 107254 500032
rect 110418 497936 110474 497992
rect 113178 500384 113234 500440
rect 112626 500248 112682 500304
rect 110602 497800 110658 497856
rect 109038 497664 109094 497720
rect 107658 497528 107714 497584
rect 106186 489096 106242 489152
rect 115938 500656 115994 500712
rect 114742 500520 114798 500576
rect 118698 500792 118754 500848
rect 120078 500792 120134 500848
rect 114558 500112 114614 500168
rect 132590 500792 132646 500848
rect 134154 499976 134210 500032
rect 136270 499840 136326 499896
rect 142066 500792 142122 500848
rect 138478 499704 138534 499760
rect 144642 500792 144698 500848
rect 132590 499568 132646 499624
rect 142066 499568 142122 499624
rect 144642 499568 144698 499624
rect 147034 500792 147090 500848
rect 148138 500792 148194 500848
rect 149242 500792 149298 500848
rect 150346 500792 150402 500848
rect 151358 500792 151414 500848
rect 152462 500792 152518 500848
rect 146022 500656 146078 500712
rect 151910 486512 151966 486568
rect 153014 489096 153070 489152
rect 152002 486376 152058 486432
rect 121366 401512 121422 401568
rect 115754 401376 115810 401432
rect 114466 401240 114522 401296
rect 111706 400968 111762 401024
rect 111614 400832 111670 400888
rect 77942 363704 77998 363760
rect 21362 357584 21418 357640
rect 75826 351056 75882 351112
rect 109590 351464 109646 351520
rect 107566 351328 107622 351384
rect 104898 351056 104954 351112
rect 106186 351056 106242 351112
rect 108670 351192 108726 351248
rect 112902 351600 112958 351656
rect 115846 401104 115902 401160
rect 119342 351736 119398 351792
rect 117134 350920 117190 350976
rect 122470 351736 122526 351792
rect 124678 350512 124734 350568
rect 126886 350648 126942 350704
rect 129094 350784 129150 350840
rect 129738 350784 129794 350840
rect 129738 350512 129794 350568
rect 135166 400696 135222 400752
rect 136546 400560 136602 400616
rect 139306 400424 139362 400480
rect 146206 400288 146262 400344
rect 144918 350920 144974 350976
rect 144918 350512 144974 350568
rect 145562 351192 145618 351248
rect 145562 350920 145618 350976
rect 146298 351464 146354 351520
rect 146942 351464 146998 351520
rect 148046 351464 148102 351520
rect 149426 351464 149482 351520
rect 150070 351464 150126 351520
rect 151174 351464 151230 351520
rect 152370 351464 152426 351520
rect 146298 351192 146354 351248
rect 153382 500828 153384 500848
rect 153384 500828 153436 500848
rect 153436 500828 153438 500848
rect 153382 500792 153438 500828
rect 153474 500520 153530 500576
rect 156050 465296 156106 465352
rect 185582 450880 185638 450936
rect 190182 500792 190238 500848
rect 191286 500792 191342 500848
rect 189078 500656 189134 500712
rect 194506 500112 194562 500168
rect 280526 528400 280582 528456
rect 280526 518880 280582 518936
rect 281538 515888 281594 515944
rect 280342 495488 280398 495544
rect 280342 489912 280398 489968
rect 280158 479984 280214 480040
rect 279606 471824 279662 471880
rect 280158 470600 280214 470656
rect 280250 451152 280306 451208
rect 280250 445712 280306 445768
rect 280342 439456 280398 439512
rect 280342 434696 280398 434752
rect 281538 430480 281594 430536
rect 281630 421232 281686 421288
rect 189446 351736 189502 351792
rect 191194 351736 191250 351792
rect 189906 351600 189962 351656
rect 194138 357448 194194 357504
rect 280342 347520 280398 347576
rect 280342 338136 280398 338192
rect 280342 326984 280398 327040
rect 17130 274896 17186 274952
rect 67178 236000 67234 236056
rect 113362 295296 113418 295352
rect 116398 221176 116454 221232
rect 116122 219952 116178 220008
rect 104806 219272 104862 219328
rect 116398 218864 116454 218920
rect 104806 217948 104808 217968
rect 104808 217948 104860 217968
rect 104860 217948 104862 217968
rect 104806 217912 104862 217948
rect 116398 217640 116454 217696
rect 104806 216588 104808 216608
rect 104808 216588 104860 216608
rect 104860 216588 104862 216608
rect 104806 216552 104862 216588
rect 115938 216552 115994 216608
rect 104806 215600 104862 215656
rect 116398 215348 116454 215384
rect 116398 215328 116400 215348
rect 116400 215328 116452 215348
rect 116452 215328 116454 215348
rect 104806 214648 104862 214704
rect 116398 214104 116454 214160
rect 104806 213424 104862 213480
rect 115938 213016 115994 213072
rect 104438 212064 104494 212120
rect 116306 211792 116362 211848
rect 104806 210840 104862 210896
rect 116306 210704 116362 210760
rect 104806 209480 104862 209536
rect 116030 209480 116086 209536
rect 116398 208256 116454 208312
rect 104806 208120 104862 208176
rect 116306 207168 116362 207224
rect 104806 206916 104862 206952
rect 104806 206896 104808 206916
rect 104808 206896 104860 206916
rect 104860 206896 104862 206916
rect 104714 206216 104770 206272
rect 115938 205944 115994 206000
rect 104806 204992 104862 205048
rect 116398 204856 116454 204912
rect 104806 203632 104862 203688
rect 116306 203632 116362 203688
rect 104806 202408 104862 202464
rect 116122 202408 116178 202464
rect 116122 201320 116178 201376
rect 104806 201048 104862 201104
rect 115938 200132 115940 200152
rect 115940 200132 115992 200152
rect 115992 200132 115994 200152
rect 104806 199824 104862 199880
rect 115938 200096 115994 200132
rect 115938 199008 115994 199064
rect 104806 198464 104862 198520
rect 104806 197260 104862 197296
rect 116122 197784 116178 197840
rect 104806 197240 104808 197260
rect 104808 197240 104860 197260
rect 104860 197240 104862 197260
rect 116398 196696 116454 196752
rect 104714 196560 104770 196616
rect 115938 195472 115994 195528
rect 104806 195336 104862 195392
rect 116122 194248 116178 194304
rect 104806 193976 104862 194032
rect 116398 193160 116454 193216
rect 104438 192752 104494 192808
rect 104438 191392 104494 191448
rect 116030 191956 116086 191992
rect 116030 191936 116032 191956
rect 116032 191936 116084 191956
rect 116084 191936 116086 191956
rect 116490 190848 116546 190904
rect 104714 190168 104770 190224
rect 116398 189624 116454 189680
rect 104806 188808 104862 188864
rect 104806 187448 104862 187504
rect 104806 186244 104862 186280
rect 116398 188400 116454 188456
rect 115938 187312 115994 187368
rect 104806 186224 104808 186244
rect 104808 186224 104860 186244
rect 104860 186224 104862 186244
rect 116030 186088 116086 186144
rect 104714 185544 104770 185600
rect 104806 184320 104862 184376
rect 104806 182960 104862 183016
rect 104806 181736 104862 181792
rect 116398 185020 116454 185056
rect 116398 185000 116400 185020
rect 116400 185000 116452 185020
rect 116452 185000 116454 185020
rect 116398 183776 116454 183832
rect 115938 182552 115994 182608
rect 115938 181464 115994 181520
rect 104806 180376 104862 180432
rect 116398 180240 116454 180296
rect 104806 179016 104862 179072
rect 115938 179152 115994 179208
rect 104162 177792 104218 177848
rect 104162 176432 104218 176488
rect 104806 175228 104862 175264
rect 115938 177928 115994 177984
rect 116398 176840 116454 176896
rect 104806 175208 104808 175228
rect 104808 175208 104860 175228
rect 104860 175208 104862 175228
rect 104530 174528 104586 174584
rect 116398 175616 116454 175672
rect 115938 174392 115994 174448
rect 104806 173304 104862 173360
rect 104438 172080 104494 172136
rect 116398 173304 116454 173360
rect 116122 172080 116178 172136
rect 104806 170720 104862 170776
rect 104162 168136 104218 168192
rect 116306 170992 116362 171048
rect 104806 169360 104862 169416
rect 104254 166912 104310 166968
rect 116398 169788 116454 169824
rect 116398 169768 116400 169788
rect 116400 169768 116452 169788
rect 116452 169768 116454 169788
rect 116398 168544 116454 168600
rect 115938 167456 115994 167512
rect 104806 165552 104862 165608
rect 104622 164872 104678 164928
rect 115938 166232 115994 166288
rect 116122 165144 116178 165200
rect 104806 163648 104862 163704
rect 104806 162288 104862 162344
rect 116398 163920 116454 163976
rect 116214 162696 116270 162752
rect 104806 160928 104862 160984
rect 103702 158616 103758 158672
rect 116398 161608 116454 161664
rect 116398 160384 116454 160440
rect 104806 159704 104862 159760
rect 116398 159296 116454 159352
rect 104254 157256 104310 157312
rect 116398 158072 116454 158128
rect 116030 156984 116086 157040
rect 104806 155896 104862 155952
rect 104346 154400 104402 154456
rect 104622 153856 104678 153912
rect 116030 155760 116086 155816
rect 116398 154572 116400 154592
rect 116400 154572 116452 154592
rect 116452 154572 116454 154592
rect 116398 154536 116454 154572
rect 115938 153448 115994 153504
rect 104806 152632 104862 152688
rect 116398 152224 116454 152280
rect 104254 151544 104310 151600
rect 116398 151136 116454 151192
rect 103794 150320 103850 150376
rect 103702 148960 103758 149016
rect 116398 149912 116454 149968
rect 104346 147600 104402 147656
rect 103518 140528 103574 140584
rect 116398 148688 116454 148744
rect 115938 147600 115994 147656
rect 116398 146376 116454 146432
rect 104806 146240 104862 146296
rect 116030 145288 116086 145344
rect 104714 144744 104770 144800
rect 104622 144200 104678 144256
rect 116398 144064 116454 144120
rect 104530 142976 104586 143032
rect 116398 142840 116454 142896
rect 104162 141752 104218 141808
rect 116398 141752 116454 141808
rect 103702 139304 103758 139360
rect 116398 140528 116454 140584
rect 116306 139476 116308 139496
rect 116308 139476 116360 139496
rect 116360 139476 116362 139496
rect 104346 137944 104402 138000
rect 104806 136584 104862 136640
rect 116306 139440 116362 139476
rect 115846 138216 115902 138272
rect 104806 135088 104862 135144
rect 104806 133728 104862 133784
rect 104714 133184 104770 133240
rect 104346 131960 104402 132016
rect 116398 137128 116454 137184
rect 115938 135904 115994 135960
rect 116398 134680 116454 134736
rect 103978 130600 104034 130656
rect 104806 129240 104862 129296
rect 116398 132368 116454 132424
rect 115938 131280 115994 131336
rect 116398 128832 116454 128888
rect 104806 128016 104862 128072
rect 116398 127744 116454 127800
rect 32218 125024 32274 125080
rect 116398 126520 116454 126576
rect 116398 125432 116454 125488
rect 116306 124208 116362 124264
rect 146022 254124 146024 254144
rect 146024 254124 146076 254144
rect 146076 254124 146078 254144
rect 146022 254088 146078 254124
rect 149518 254124 149520 254144
rect 149520 254124 149572 254144
rect 149572 254124 149574 254144
rect 149518 254088 149574 254124
rect 185582 274896 185638 274952
rect 189078 320456 189134 320512
rect 192390 320320 192446 320376
rect 190182 320184 190238 320240
rect 191286 320184 191342 320240
rect 194506 320184 194562 320240
rect 193402 319368 193458 319424
rect 282274 586064 282330 586120
rect 282274 430480 282330 430536
rect 348790 700576 348846 700632
rect 282918 683168 282974 683224
rect 283286 683168 283342 683224
rect 284298 608776 284354 608832
rect 283102 578176 283158 578232
rect 283286 578176 283342 578232
rect 282918 550568 282974 550624
rect 283102 550568 283158 550624
rect 282826 527312 282882 527368
rect 283010 527176 283066 527232
rect 282918 518880 282974 518936
rect 283194 518880 283250 518936
rect 282918 482976 282974 483032
rect 283102 482976 283158 483032
rect 284298 392672 284354 392728
rect 282458 369824 282514 369880
rect 282550 360032 282606 360088
rect 282274 335960 282330 336016
rect 282182 322088 282238 322144
rect 280342 317600 280398 317656
rect 280342 317328 280398 317384
rect 280342 309576 280398 309632
rect 279514 295840 279570 295896
rect 280710 295024 280766 295080
rect 280710 277616 280766 277672
rect 282182 255040 282238 255096
rect 280526 251096 280582 251152
rect 280526 241576 280582 241632
rect 209778 235184 209834 235240
rect 250442 235184 250498 235240
rect 205822 233824 205878 233880
rect 205730 229744 205786 229800
rect 204534 228248 204590 228304
rect 207018 232464 207074 232520
rect 208858 223624 208914 223680
rect 213918 221312 213974 221368
rect 214010 220496 214066 220552
rect 213918 219680 213974 219736
rect 213918 218864 213974 218920
rect 214010 218184 214066 218240
rect 213918 217368 213974 217424
rect 213918 216588 213920 216608
rect 213920 216588 213972 216608
rect 213972 216588 213974 216608
rect 213918 216552 213974 216588
rect 213918 215736 213974 215792
rect 213918 215056 213974 215112
rect 214010 214240 214066 214296
rect 213918 213424 213974 213480
rect 214010 212608 214066 212664
rect 213918 211928 213974 211984
rect 214010 211112 214066 211168
rect 213918 210296 213974 210352
rect 213918 209480 213974 209536
rect 214010 208800 214066 208856
rect 213918 207984 213974 208040
rect 214010 207168 214066 207224
rect 213918 206352 213974 206408
rect 214010 205672 214066 205728
rect 213918 204856 213974 204912
rect 213918 204040 213974 204096
rect 214010 203224 214066 203280
rect 213918 202408 213974 202464
rect 214010 201728 214066 201784
rect 213918 200912 213974 200968
rect 214010 200096 214066 200152
rect 213918 199280 213974 199336
rect 213918 198620 213974 198656
rect 213918 198600 213920 198620
rect 213920 198600 213972 198620
rect 213972 198600 213974 198620
rect 214010 197784 214066 197840
rect 213918 196968 213974 197024
rect 214010 196152 214066 196208
rect 213918 195472 213974 195528
rect 214010 194656 214066 194712
rect 213918 193840 213974 193896
rect 213918 193024 213974 193080
rect 214010 192344 214066 192400
rect 213918 191528 213974 191584
rect 214010 190712 214066 190768
rect 213918 189896 213974 189952
rect 214010 189216 214066 189272
rect 213918 188400 213974 188456
rect 213918 186768 213974 186824
rect 213918 185272 213974 185328
rect 214194 187584 214250 187640
rect 214102 184456 214158 184512
rect 214286 181872 214342 181928
rect 213918 180548 213920 180568
rect 213920 180548 213972 180568
rect 213972 180548 213974 180568
rect 213918 180512 213974 180548
rect 213918 179052 213920 179072
rect 213920 179052 213972 179072
rect 213972 179052 213974 179072
rect 213918 179016 213974 179052
rect 214010 178200 214066 178256
rect 213918 177384 213974 177440
rect 214010 175888 214066 175944
rect 214470 185952 214526 186008
rect 214378 179696 214434 179752
rect 214286 176568 214342 176624
rect 214194 175072 214250 175128
rect 213918 174256 213974 174312
rect 214194 173848 214250 173904
rect 214010 173440 214066 173496
rect 213918 172760 213974 172816
rect 213918 171128 213974 171184
rect 213918 169496 213974 169552
rect 213918 168000 213974 168056
rect 214470 173884 214472 173904
rect 214472 173884 214524 173904
rect 214524 173884 214526 173904
rect 214470 173848 214526 173884
rect 214378 171944 214434 172000
rect 213918 166368 213974 166424
rect 214010 165688 214066 165744
rect 213918 164872 213974 164928
rect 213918 164092 213920 164112
rect 213920 164092 213972 164112
rect 213972 164092 213974 164112
rect 213918 164056 213974 164092
rect 213918 163240 213974 163296
rect 213918 162560 213974 162616
rect 213918 161744 213974 161800
rect 213918 160928 213974 160984
rect 213918 160112 213974 160168
rect 213918 156984 213974 157040
rect 214102 156304 214158 156360
rect 213918 155488 213974 155544
rect 214010 153856 214066 153912
rect 213918 153176 213974 153232
rect 213918 152360 213974 152416
rect 213918 151544 213974 151600
rect 213918 150728 213974 150784
rect 213918 149912 213974 149968
rect 213918 149232 213974 149288
rect 213918 148416 213974 148472
rect 214010 147600 214066 147656
rect 213918 146784 213974 146840
rect 214010 146104 214066 146160
rect 213918 145288 213974 145344
rect 214010 144472 214066 144528
rect 213918 143676 213974 143712
rect 213918 143656 213920 143676
rect 213920 143656 213972 143676
rect 213972 143656 213974 143676
rect 214562 143520 214618 143576
rect 214010 142976 214066 143032
rect 213918 142196 213920 142216
rect 213920 142196 213972 142216
rect 213972 142196 213974 142216
rect 213918 142160 213974 142196
rect 213918 141344 213974 141400
rect 214010 140528 214066 140584
rect 213918 139848 213974 139904
rect 214010 139032 214066 139088
rect 213918 138216 213974 138272
rect 214010 137400 214066 137456
rect 213918 136740 213974 136776
rect 213918 136720 213920 136740
rect 213920 136720 213972 136740
rect 213972 136720 213974 136740
rect 213918 135904 213974 135960
rect 214010 135088 214066 135144
rect 213918 134272 213974 134328
rect 117134 133592 117190 133648
rect 214010 133456 214066 133512
rect 213918 132776 213974 132832
rect 214010 131960 214066 132016
rect 213918 131180 213920 131200
rect 213920 131180 213972 131200
rect 213972 131180 213974 131200
rect 213918 131144 213974 131180
rect 213918 130328 213974 130384
rect 116674 130056 116730 130112
rect 213918 129648 213974 129704
rect 213918 128832 213974 128888
rect 213918 128016 213974 128072
rect 213918 127200 213974 127256
rect 213918 126520 213974 126576
rect 213918 125704 213974 125760
rect 213918 124908 213974 124944
rect 213918 124888 213920 124908
rect 213920 124888 213972 124908
rect 213972 124888 213974 124908
rect 213918 124108 213920 124128
rect 213920 124108 213972 124128
rect 213972 124108 213974 124128
rect 213918 124072 213974 124108
rect 213918 123428 213920 123448
rect 213920 123428 213972 123448
rect 213972 123428 213974 123448
rect 213918 123392 213974 123428
rect 116582 122984 116638 123040
rect 213918 122576 213974 122632
rect 116398 121896 116454 121952
rect 213918 121760 213974 121816
rect 213918 120944 213974 121000
rect 116398 120672 116454 120728
rect 213918 120264 213974 120320
rect 116398 119584 116454 119640
rect 213918 119448 213974 119504
rect 94502 98912 94558 98968
rect 213918 118652 213974 118688
rect 213918 118632 213920 118652
rect 213920 118632 213972 118652
rect 213972 118632 213974 118652
rect 116398 118360 116454 118416
rect 214010 117816 214066 117872
rect 116398 117136 116454 117192
rect 116122 116068 116178 116104
rect 116122 116048 116124 116068
rect 116124 116048 116176 116068
rect 116176 116048 116178 116068
rect 94686 97960 94742 98016
rect 94594 97144 94650 97200
rect 94778 96192 94834 96248
rect 94410 92656 94466 92712
rect 94318 87216 94374 87272
rect 94410 86400 94466 86456
rect 94226 85448 94282 85504
rect 94226 82864 94282 82920
rect 94134 81912 94190 81968
rect 94410 80960 94466 81016
rect 94410 79192 94466 79248
rect 94594 91704 94650 91760
rect 94502 78376 94558 78432
rect 94226 77424 94282 77480
rect 213918 117000 213974 117056
rect 214010 116320 214066 116376
rect 213918 115504 213974 115560
rect 116398 114824 116454 114880
rect 214010 114688 214066 114744
rect 213918 113872 213974 113928
rect 116398 113736 116454 113792
rect 214010 113192 214066 113248
rect 94962 95376 95018 95432
rect 94870 94424 94926 94480
rect 94778 89936 94834 89992
rect 95146 93508 95148 93528
rect 95148 93508 95200 93528
rect 95200 93508 95202 93528
rect 95146 93472 95202 93508
rect 116398 112512 116454 112568
rect 213918 112376 213974 112432
rect 213918 111560 213974 111616
rect 116398 111424 116454 111480
rect 214010 110744 214066 110800
rect 116398 110200 116454 110256
rect 213918 110064 213974 110120
rect 214010 109248 214066 109304
rect 116306 108976 116362 109032
rect 214470 108976 214526 109032
rect 213918 108432 213974 108488
rect 116398 107888 116454 107944
rect 95054 90888 95110 90944
rect 94962 89120 95018 89176
rect 94686 80144 94742 80200
rect 94594 76472 94650 76528
rect 94594 75692 94596 75712
rect 94596 75692 94648 75712
rect 94648 75692 94650 75712
rect 94594 75656 94650 75692
rect 94410 72120 94466 72176
rect 93858 68484 93860 68504
rect 93860 68484 93912 68504
rect 93912 68484 93914 68504
rect 93858 68448 93914 68484
rect 93950 61376 94006 61432
rect 94226 57704 94282 57760
rect 94594 73888 94650 73944
rect 94502 63960 94558 64016
rect 94410 59472 94466 59528
rect 94318 56888 94374 56944
rect 93858 50632 93914 50688
rect 93950 49680 94006 49736
rect 94778 72936 94834 72992
rect 95146 88204 95148 88224
rect 95148 88204 95200 88224
rect 95200 88204 95202 88224
rect 95146 88168 95202 88204
rect 95146 84632 95202 84688
rect 95146 83680 95202 83736
rect 94962 74704 95018 74760
rect 94870 71168 94926 71224
rect 94870 70252 94872 70272
rect 94872 70252 94924 70272
rect 94924 70252 94926 70272
rect 94870 70216 94926 70252
rect 94686 65864 94742 65920
rect 94686 64912 94742 64968
rect 94594 60424 94650 60480
rect 94870 63144 94926 63200
rect 95054 69400 95110 69456
rect 95146 67632 95202 67688
rect 95146 66680 95202 66736
rect 94962 62192 95018 62248
rect 94778 58656 94834 58712
rect 94686 55120 94742 55176
rect 94502 54168 94558 54224
rect 94410 51448 94466 51504
rect 94042 48864 94098 48920
rect 94226 46144 94282 46200
rect 94410 44376 94466 44432
rect 94962 53216 95018 53272
rect 214010 107616 214066 107672
rect 213918 106936 213974 106992
rect 116398 106664 116454 106720
rect 213918 106120 213974 106176
rect 116398 105576 116454 105632
rect 214010 105304 214066 105360
rect 213918 104488 213974 104544
rect 116398 104352 116454 104408
rect 214838 167184 214894 167240
rect 214746 158616 214802 158672
rect 229006 221312 229062 221368
rect 226338 220804 226340 220824
rect 226340 220804 226392 220824
rect 226392 220804 226394 220824
rect 226338 220768 226394 220804
rect 226338 220124 226340 220144
rect 226340 220124 226392 220144
rect 226392 220124 226394 220144
rect 226338 220088 226394 220124
rect 226430 219544 226486 219600
rect 226338 219000 226394 219056
rect 226430 218320 226486 218376
rect 226338 217776 226394 217832
rect 226430 217232 226486 217288
rect 226338 216552 226394 216608
rect 226430 216008 226486 216064
rect 226338 215464 226394 215520
rect 226430 214784 226486 214840
rect 226338 214240 226394 214296
rect 226430 213560 226486 213616
rect 226338 213016 226394 213072
rect 226522 212472 226578 212528
rect 226062 211792 226118 211848
rect 225970 210704 226026 210760
rect 226246 211248 226302 211304
rect 226154 210024 226210 210080
rect 226062 209480 226118 209536
rect 225786 207712 225842 207768
rect 225602 205264 225658 205320
rect 225694 204720 225750 204776
rect 225970 207168 226026 207224
rect 225878 206488 225934 206544
rect 226246 208936 226302 208992
rect 226154 207984 226210 208040
rect 226246 205944 226302 206000
rect 226062 203496 226118 203552
rect 225970 202952 226026 203008
rect 225786 202408 225842 202464
rect 225694 199960 225750 200016
rect 215206 183640 215262 183696
rect 215022 182824 215078 182880
rect 215206 182144 215262 182200
rect 215022 170312 215078 170368
rect 225878 200640 225934 200696
rect 226246 204176 226302 204232
rect 226154 201728 226210 201784
rect 226338 201184 226394 201240
rect 226430 199416 226486 199472
rect 226338 198872 226394 198928
rect 226430 198192 226486 198248
rect 226338 197648 226394 197704
rect 226338 196968 226394 197024
rect 226706 196424 226762 196480
rect 226522 195880 226578 195936
rect 226338 195200 226394 195256
rect 226430 194676 226486 194712
rect 226430 194656 226432 194676
rect 226432 194656 226484 194676
rect 226484 194656 226486 194676
rect 226338 194112 226394 194168
rect 226430 193432 226486 193488
rect 226430 192888 226486 192944
rect 226338 192344 226394 192400
rect 226430 191664 226486 191720
rect 226522 191120 226578 191176
rect 226338 190440 226394 190496
rect 226430 189896 226486 189952
rect 226338 189352 226394 189408
rect 226338 188672 226394 188728
rect 215114 168816 215170 168872
rect 226430 188128 226486 188184
rect 226338 186904 226394 186960
rect 226430 186396 226432 186416
rect 226432 186396 226484 186416
rect 226484 186396 226486 186416
rect 226430 186360 226486 186396
rect 226338 185816 226394 185872
rect 226430 185136 226486 185192
rect 226338 184592 226394 184648
rect 227074 187584 227130 187640
rect 226982 184048 227038 184104
rect 226430 183368 226486 183424
rect 225694 182824 225750 182880
rect 225602 178064 225658 178120
rect 226338 182144 226394 182200
rect 226338 181600 226394 181656
rect 226338 181056 226394 181112
rect 226430 180376 226486 180432
rect 226338 179832 226394 179888
rect 226338 179288 226394 179344
rect 226430 178608 226486 178664
rect 226338 177520 226394 177576
rect 226430 176840 226486 176896
rect 226890 176296 226946 176352
rect 227442 175752 227498 175808
rect 296626 527448 296682 527504
rect 298098 527468 298154 527504
rect 298098 527448 298100 527468
rect 298100 527448 298152 527468
rect 298152 527448 298154 527468
rect 288530 527212 288532 527232
rect 288532 527212 288584 527232
rect 288584 527212 288586 527232
rect 288530 527176 288586 527212
rect 288898 317056 288954 317112
rect 289726 325216 289782 325272
rect 289634 308896 289690 308952
rect 300858 305496 300914 305552
rect 292578 302776 292634 302832
rect 302974 527176 303030 527232
rect 304262 328208 304318 328264
rect 303618 326304 303674 326360
rect 303618 324400 303674 324456
rect 304354 322496 304410 322552
rect 304446 320592 304502 320648
rect 303618 318688 303674 318744
rect 304354 316920 304410 316976
rect 304262 315016 304318 315072
rect 303618 313112 303674 313168
rect 303618 311208 303674 311264
rect 303618 309304 303674 309360
rect 303618 307400 303674 307456
rect 313278 613400 313334 613456
rect 313278 462712 313334 462768
rect 478510 700440 478566 700496
rect 543462 700304 543518 700360
rect 314658 515752 314714 515808
rect 314658 439592 314714 439648
rect 580170 697992 580226 698048
rect 506018 663856 506074 663912
rect 552018 641688 552074 641744
rect 551650 639512 551706 639568
rect 456062 635160 456118 635216
rect 455418 591640 455474 591696
rect 326894 567840 326950 567896
rect 325054 532072 325110 532128
rect 408590 531936 408646 531992
rect 421378 533160 421434 533216
rect 425702 533024 425758 533080
rect 430026 532888 430082 532944
rect 434258 531800 434314 531856
rect 440514 567840 440570 567896
rect 441802 532752 441858 532808
rect 441618 532072 441674 532128
rect 440790 531664 440846 531720
rect 442998 531528 443054 531584
rect 456798 616256 456854 616312
rect 550822 569744 550878 569800
rect 551006 569744 551062 569800
rect 550822 569472 550878 569528
rect 454774 531392 454830 531448
rect 493966 560904 494022 560960
rect 477498 530168 477554 530224
rect 480626 530032 480682 530088
rect 493782 534656 493838 534712
rect 492034 531120 492090 531176
rect 490378 529896 490434 529952
rect 499486 545672 499542 545728
rect 498566 532344 498622 532400
rect 495346 532208 495402 532264
rect 497462 532072 497518 532128
rect 496358 531936 496414 531992
rect 508226 533568 508282 533624
rect 506110 533432 506166 533488
rect 501786 533296 501842 533352
rect 500682 530712 500738 530768
rect 505006 532616 505062 532672
rect 503626 532480 503682 532536
rect 502890 530576 502946 530632
rect 507122 530984 507178 531040
rect 509054 530848 509110 530904
rect 551006 563216 551062 563272
rect 551006 560224 551062 560280
rect 551006 555464 551062 555520
rect 516874 531800 516930 531856
rect 515770 531120 515826 531176
rect 545946 531256 546002 531312
rect 551374 632168 551430 632224
rect 551558 628360 551614 628416
rect 551374 627952 551430 628008
rect 551466 622376 551522 622432
rect 551374 621288 551430 621344
rect 551374 618568 551430 618624
rect 551374 617480 551430 617536
rect 551650 627952 551706 628008
rect 551558 618432 551614 618488
rect 551650 616392 551706 616448
rect 551374 601568 551430 601624
rect 551374 599936 551430 599992
rect 551374 595176 551430 595232
rect 551374 595076 551376 595096
rect 551376 595076 551428 595096
rect 551428 595076 551430 595096
rect 551374 595040 551430 595076
rect 551374 592340 551430 592376
rect 551374 592320 551376 592340
rect 551376 592320 551428 592340
rect 551428 592320 551430 592340
rect 551374 592204 551430 592240
rect 551374 592184 551376 592204
rect 551376 592184 551428 592204
rect 551428 592184 551430 592204
rect 551374 586916 551376 586936
rect 551376 586916 551428 586936
rect 551428 586916 551430 586936
rect 551374 586880 551430 586916
rect 551374 586236 551376 586256
rect 551376 586236 551428 586256
rect 551428 586236 551430 586256
rect 551374 586200 551430 586236
rect 551374 581984 551430 582040
rect 551374 577496 551430 577552
rect 551650 613808 551706 613864
rect 551558 612720 551614 612776
rect 551742 613672 551798 613728
rect 551650 612176 551706 612232
rect 551650 611632 551706 611688
rect 551742 601160 551798 601216
rect 551742 600344 551798 600400
rect 551834 597896 551890 597952
rect 553398 641008 553454 641064
rect 552202 639920 552258 639976
rect 552110 638696 552166 638752
rect 552294 637472 552350 637528
rect 552386 631352 552442 631408
rect 552478 624008 552534 624064
rect 552570 614352 552626 614408
rect 553030 608232 553086 608288
rect 552662 604560 552718 604616
rect 552754 599664 552810 599720
rect 552846 597216 552902 597272
rect 552938 594768 552994 594824
rect 553122 605784 553178 605840
rect 553214 603336 553270 603392
rect 553306 595992 553362 596048
rect 553306 576000 553362 576056
rect 553306 574776 553362 574832
rect 553306 574116 553362 574152
rect 553306 574096 553308 574116
rect 553308 574096 553360 574116
rect 553360 574096 553362 574116
rect 553306 572872 553362 572928
rect 553306 571668 553362 571704
rect 553306 571648 553308 571668
rect 553308 571648 553360 571668
rect 553360 571648 553362 571668
rect 553306 570016 553362 570072
rect 553490 633800 553546 633856
rect 553582 630128 553638 630184
rect 553766 627680 553822 627736
rect 553674 626456 553730 626512
rect 553858 625232 553914 625288
rect 553950 620336 554006 620392
rect 554134 617888 554190 617944
rect 554042 615576 554098 615632
rect 554226 616800 554282 616856
rect 554318 610680 554374 610736
rect 554410 609456 554466 609512
rect 554502 607008 554558 607064
rect 554594 593680 554650 593736
rect 554686 592456 554742 592512
rect 554594 590008 554650 590064
rect 554594 588804 554650 588840
rect 554594 588784 554596 588804
rect 554596 588784 554648 588804
rect 554648 588784 554650 588804
rect 554594 587560 554650 587616
rect 554778 591232 554834 591288
rect 554870 586356 554926 586392
rect 554870 586336 554872 586356
rect 554872 586336 554924 586356
rect 554924 586336 554926 586356
rect 554870 585148 554872 585168
rect 554872 585148 554924 585168
rect 554924 585148 554926 585168
rect 554870 585112 554926 585148
rect 554870 583772 554926 583808
rect 554870 583752 554872 583772
rect 554872 583752 554924 583772
rect 554924 583752 554926 583772
rect 555422 582664 555478 582720
rect 554870 581052 554926 581088
rect 554870 581032 554872 581052
rect 554872 581032 554924 581052
rect 554924 581032 554926 581052
rect 554870 579692 554926 579728
rect 554870 579672 554872 579692
rect 554872 579672 554924 579692
rect 554924 579672 554926 579692
rect 554870 578448 554926 578504
rect 554870 577224 554926 577280
rect 489274 528536 489330 528592
rect 471702 528264 471758 528320
rect 317418 527176 317474 527232
rect 317418 526904 317474 526960
rect 315946 515752 316002 515808
rect 320546 482976 320602 483032
rect 320730 482976 320786 483032
rect 338118 428712 338174 428768
rect 338394 428576 338450 428632
rect 338118 198600 338174 198656
rect 283378 173848 283434 173904
rect 232226 173168 232282 173224
rect 283378 173168 283434 173224
rect 214930 157800 214986 157856
rect 214930 154672 214986 154728
rect 214746 143520 214802 143576
rect 214746 108976 214802 109032
rect 214010 103808 214066 103864
rect 116306 103128 116362 103184
rect 213918 102992 213974 103048
rect 214010 102176 214066 102232
rect 116306 102040 116362 102096
rect 213918 101360 213974 101416
rect 116398 100836 116454 100872
rect 116398 100816 116400 100836
rect 116400 100816 116452 100836
rect 116452 100816 116454 100836
rect 213918 100544 213974 100600
rect 214010 99864 214066 99920
rect 116398 99728 116454 99784
rect 116398 98504 116454 98560
rect 116398 97280 116454 97336
rect 214102 97416 214158 97472
rect 213918 96736 213974 96792
rect 116306 96192 116362 96248
rect 214654 98232 214710 98288
rect 214562 95920 214618 95976
rect 215114 99048 215170 99104
rect 232318 154536 232374 154592
rect 232502 154536 232558 154592
rect 227442 149368 227498 149424
rect 227442 148824 227498 148880
rect 227534 148144 227590 148200
rect 227442 147620 227498 147656
rect 227442 147600 227444 147620
rect 227444 147600 227496 147620
rect 227496 147600 227498 147620
rect 226982 146920 227038 146976
rect 227534 146376 227590 146432
rect 227442 145832 227498 145888
rect 226706 145152 226762 145208
rect 226522 143928 226578 143984
rect 226890 142840 226946 142896
rect 226706 141616 226762 141672
rect 227442 144608 227498 144664
rect 227442 143420 227444 143440
rect 227444 143420 227496 143440
rect 227496 143420 227498 143440
rect 227442 143384 227498 143420
rect 227258 140936 227314 140992
rect 226522 136720 226578 136776
rect 227074 140392 227130 140448
rect 227626 142160 227682 142216
rect 227534 139712 227590 139768
rect 227442 139168 227498 139224
rect 227350 138624 227406 138680
rect 226706 137400 226762 137456
rect 226614 136176 226670 136232
rect 226430 135632 226486 135688
rect 227442 137964 227498 138000
rect 227442 137944 227444 137964
rect 227444 137944 227496 137964
rect 227496 137944 227498 137964
rect 226798 134952 226854 135008
rect 227442 134408 227498 134464
rect 227074 133728 227130 133784
rect 227626 133184 227682 133240
rect 227534 132504 227590 132560
rect 227350 131960 227406 132016
rect 227442 131416 227498 131472
rect 226706 130736 226762 130792
rect 227074 130192 227130 130248
rect 226522 129512 226578 129568
rect 227534 128968 227590 129024
rect 227442 128424 227498 128480
rect 226338 127744 226394 127800
rect 227442 127200 227498 127256
rect 227442 126520 227498 126576
rect 227442 125976 227498 126032
rect 227442 125296 227498 125352
rect 227258 124752 227314 124808
rect 227258 124208 227314 124264
rect 227258 123528 227314 123584
rect 227442 122984 227498 123040
rect 227442 122304 227498 122360
rect 227442 121760 227498 121816
rect 227442 121216 227498 121272
rect 227442 120536 227498 120592
rect 226430 119992 226486 120048
rect 226338 119312 226394 119368
rect 226246 118768 226302 118824
rect 226154 117544 226210 117600
rect 227442 118088 227498 118144
rect 227442 117000 227498 117056
rect 226246 116320 226302 116376
rect 226154 115096 226210 115152
rect 226062 114552 226118 114608
rect 225970 113328 226026 113384
rect 225878 112104 225934 112160
rect 225786 110336 225842 110392
rect 225602 109112 225658 109168
rect 225694 107888 225750 107944
rect 227074 115776 227130 115832
rect 226246 114008 226302 114064
rect 226154 112784 226210 112840
rect 226062 110880 226118 110936
rect 226246 111560 226302 111616
rect 226338 109792 226394 109848
rect 226154 108568 226210 108624
rect 225970 107344 226026 107400
rect 225878 106800 225934 106856
rect 226062 105576 226118 105632
rect 226246 105712 226302 105768
rect 227442 104916 227498 104952
rect 227442 104896 227444 104916
rect 227444 104896 227496 104916
rect 227496 104896 227498 104916
rect 226246 104352 226302 104408
rect 227442 103808 227498 103864
rect 343638 428440 343694 428496
rect 214746 95104 214802 95160
rect 116490 94968 116546 95024
rect 116398 93900 116454 93936
rect 116398 93880 116400 93900
rect 116400 93880 116452 93900
rect 116452 93880 116454 93900
rect 116398 92656 116454 92712
rect 116398 91568 116454 91624
rect 116398 90344 116454 90400
rect 215114 94288 215170 94344
rect 215114 93608 215170 93664
rect 215206 92792 215262 92848
rect 214838 91976 214894 92032
rect 214562 90480 214618 90536
rect 214286 89664 214342 89720
rect 115938 89120 115994 89176
rect 116398 88032 116454 88088
rect 214194 88032 214250 88088
rect 116306 86808 116362 86864
rect 116398 85720 116454 85776
rect 116398 84496 116454 84552
rect 116398 83272 116454 83328
rect 115938 82184 115994 82240
rect 116398 80960 116454 81016
rect 116214 79872 116270 79928
rect 214194 82592 214250 82648
rect 214470 86536 214526 86592
rect 214378 84904 214434 84960
rect 214378 83408 214434 83464
rect 213918 79464 213974 79520
rect 116398 78648 116454 78704
rect 213918 77832 213974 77888
rect 116398 77424 116454 77480
rect 116398 76336 116454 76392
rect 213918 76336 213974 76392
rect 116398 75112 116454 75168
rect 213918 74704 213974 74760
rect 214746 88848 214802 88904
rect 214654 87352 214710 87408
rect 215022 91160 215078 91216
rect 215114 85720 215170 85776
rect 215114 84244 215170 84280
rect 215114 84224 215116 84244
rect 215116 84224 215168 84244
rect 215168 84224 215170 84244
rect 215206 81776 215262 81832
rect 215114 80960 215170 81016
rect 214930 80280 214986 80336
rect 214838 78648 214894 78704
rect 214746 75520 214802 75576
rect 116398 74024 116454 74080
rect 214102 74024 214158 74080
rect 213918 73228 213974 73264
rect 213918 73208 213920 73228
rect 213920 73208 213972 73228
rect 213972 73208 213974 73228
rect 116398 72800 116454 72856
rect 116582 71712 116638 71768
rect 116398 70488 116454 70544
rect 116398 69264 116454 69320
rect 116398 68176 116454 68232
rect 116398 66952 116454 67008
rect 116398 65864 116454 65920
rect 115938 64640 115994 64696
rect 116214 63416 116270 63472
rect 116398 62328 116454 62384
rect 214010 71576 214066 71632
rect 213918 70896 213974 70952
rect 214562 72392 214618 72448
rect 214470 68448 214526 68504
rect 214378 66136 214434 66192
rect 214010 65320 214066 65376
rect 214654 70080 214710 70136
rect 215022 77152 215078 77208
rect 215114 69264 215170 69320
rect 215114 67768 215170 67824
rect 215114 66952 215170 67008
rect 214562 64504 214618 64560
rect 215114 63824 215170 63880
rect 214654 63008 214710 63064
rect 215114 62192 215170 62248
rect 214562 61376 214618 61432
rect 116398 61104 116454 61160
rect 215114 60732 215116 60752
rect 215116 60732 215168 60752
rect 215168 60732 215170 60752
rect 215114 60696 215170 60732
rect 116398 60016 116454 60072
rect 214562 59880 214618 59936
rect 214102 59064 214158 59120
rect 116398 58792 116454 58848
rect 214194 58248 214250 58304
rect 116306 57568 116362 57624
rect 213918 57568 213974 57624
rect 214010 56752 214066 56808
rect 116306 56480 116362 56536
rect 95146 55936 95202 55992
rect 215114 55936 215170 55992
rect 116398 55292 116400 55312
rect 116400 55292 116452 55312
rect 116452 55292 116454 55312
rect 116398 55256 116454 55292
rect 214746 55120 214802 55176
rect 116398 54168 116454 54224
rect 215114 54440 215170 54496
rect 214746 53624 214802 53680
rect 116398 52944 116454 53000
rect 215114 52808 215170 52864
rect 95054 52400 95110 52456
rect 94778 47912 94834 47968
rect 215114 51992 215170 52048
rect 115938 51856 115994 51912
rect 214102 51312 214158 51368
rect 116398 50632 116454 50688
rect 215206 50496 215262 50552
rect 215114 49680 215170 49736
rect 116398 49408 116454 49464
rect 116122 48356 116124 48376
rect 116124 48356 116176 48376
rect 116176 48356 116178 48376
rect 116122 48320 116178 48356
rect 215114 48864 215170 48920
rect 214746 48048 214802 48104
rect 214010 47368 214066 47424
rect 116398 47096 116454 47152
rect 95146 46960 95202 47016
rect 215206 46552 215262 46608
rect 116398 46008 116454 46064
rect 215114 45736 215170 45792
rect 95054 45192 95110 45248
rect 215206 44920 215262 44976
rect 116398 44784 116454 44840
rect 215114 44240 215170 44296
rect 94502 43424 94558 43480
rect 94134 42472 94190 42528
rect 93950 41656 94006 41712
rect 115938 43560 115994 43616
rect 214378 43424 214434 43480
rect 214102 42608 214158 42664
rect 116398 42472 116454 42528
rect 215114 41792 215170 41848
rect 94778 40704 94834 40760
rect 94594 39888 94650 39944
rect 94502 38120 94558 38176
rect 116306 41248 116362 41304
rect 214654 41112 214710 41168
rect 116398 40160 116454 40216
rect 215114 40296 215170 40352
rect 214562 39480 214618 39536
rect 95146 38936 95202 38992
rect 116398 38936 116454 38992
rect 215114 38700 215116 38720
rect 215116 38700 215168 38720
rect 215168 38700 215170 38720
rect 215114 38664 215170 38700
rect 215114 37984 215170 38040
rect 116398 37712 116454 37768
rect 95054 37168 95110 37224
rect 214102 37168 214158 37224
rect 116398 36624 116454 36680
rect 94594 36216 94650 36272
rect 215114 36352 215170 36408
rect 93858 35400 93914 35456
rect 214654 35536 214710 35592
rect 116398 35400 116454 35456
rect 215114 34856 215170 34912
rect 93950 34448 94006 34504
rect 116306 34312 116362 34368
rect 95146 33632 95202 33688
rect 214562 34040 214618 34096
rect 215114 33224 215170 33280
rect 116398 33088 116454 33144
rect 95146 32680 95202 32736
rect 225602 74568 225658 74624
rect 227442 81096 227498 81152
rect 227350 80416 227406 80472
rect 343638 126656 343694 126712
rect 227442 79736 227498 79792
rect 227534 79056 227590 79112
rect 227442 78548 227444 78568
rect 227444 78548 227496 78568
rect 227496 78548 227498 78568
rect 227442 78512 227498 78548
rect 227534 77832 227590 77888
rect 227442 77188 227444 77208
rect 227444 77188 227496 77208
rect 227496 77188 227498 77208
rect 227442 77152 227498 77188
rect 227534 76472 227590 76528
rect 227442 75828 227444 75848
rect 227444 75828 227496 75848
rect 227496 75828 227498 75848
rect 227442 75792 227498 75828
rect 227442 75248 227498 75304
rect 227442 73888 227498 73944
rect 226982 73208 227038 73264
rect 227442 72664 227498 72720
rect 227534 71984 227590 72040
rect 227442 71304 227498 71360
rect 227534 70624 227590 70680
rect 227442 69944 227498 70000
rect 226522 69400 226578 69456
rect 227442 68720 227498 68776
rect 227534 68040 227590 68096
rect 227442 67360 227498 67416
rect 227534 66816 227590 66872
rect 227442 66172 227444 66192
rect 227444 66172 227496 66192
rect 227496 66172 227498 66192
rect 227442 66136 227498 66172
rect 227534 65456 227590 65512
rect 227442 64812 227444 64832
rect 227444 64812 227496 64832
rect 227496 64812 227498 64832
rect 227442 64776 227498 64812
rect 227442 64096 227498 64152
rect 227534 63552 227590 63608
rect 227442 62872 227498 62928
rect 227534 62192 227590 62248
rect 227534 61512 227590 61568
rect 226706 60968 226762 61024
rect 227074 60288 227130 60344
rect 227442 59608 227498 59664
rect 227442 58928 227498 58984
rect 227534 58248 227590 58304
rect 227258 57704 227314 57760
rect 227442 57024 227498 57080
rect 227258 56344 227314 56400
rect 227442 55664 227498 55720
rect 227442 55156 227444 55176
rect 227444 55156 227496 55176
rect 227496 55156 227498 55176
rect 227442 55120 227498 55156
rect 226522 54440 226578 54496
rect 226522 53080 226578 53136
rect 226338 47912 226394 47968
rect 226614 50496 226670 50552
rect 226706 49272 226762 49328
rect 227442 53780 227498 53816
rect 227442 53760 227444 53780
rect 227444 53760 227496 53780
rect 227496 53760 227498 53780
rect 227258 52400 227314 52456
rect 227442 51856 227498 51912
rect 227534 51176 227590 51232
rect 226982 49816 227038 49872
rect 226798 48592 226854 48648
rect 226522 47232 226578 47288
rect 226706 43968 226762 44024
rect 227074 43424 227130 43480
rect 227350 45328 227406 45384
rect 227534 46552 227590 46608
rect 497462 500112 497518 500168
rect 500682 500248 500738 500304
rect 493966 475360 494022 475416
rect 508226 500384 508282 500440
rect 512550 500656 512606 500712
rect 514666 500520 514722 500576
rect 507766 475496 507822 475552
rect 546590 473476 546646 473512
rect 546590 473456 546592 473476
rect 546592 473456 546644 473476
rect 546644 473456 546646 473476
rect 443642 450608 443698 450664
rect 551926 473864 551982 473920
rect 552110 473048 552166 473104
rect 552110 467200 552166 467256
rect 552294 471280 552350 471336
rect 552110 458904 552166 458960
rect 552110 456492 552112 456512
rect 552112 456492 552164 456512
rect 552164 456492 552166 456512
rect 552110 456456 552166 456492
rect 552110 455268 552112 455288
rect 552112 455268 552164 455288
rect 552164 455268 552166 455288
rect 552110 455232 552166 455268
rect 552570 471280 552626 471336
rect 552386 453464 552442 453520
rect 552938 468560 552994 468616
rect 553214 466248 553270 466304
rect 553030 463564 553032 463584
rect 553032 463564 553084 463584
rect 553084 463564 553086 463584
rect 553030 463528 553086 463564
rect 552846 460944 552902 461000
rect 552846 456728 552902 456784
rect 552754 452920 552810 452976
rect 552570 451152 552626 451208
rect 552478 450608 552534 450664
rect 552294 448704 552350 448760
rect 552202 448160 552258 448216
rect 552018 445168 552074 445224
rect 552018 441632 552074 441688
rect 553030 459720 553086 459776
rect 553306 462712 553362 462768
rect 553122 459176 553178 459232
rect 553214 454416 553270 454472
rect 552938 442448 552994 442504
rect 553398 440680 553454 440736
rect 553674 445440 553730 445496
rect 553582 443128 553638 443184
rect 554778 472096 554834 472152
rect 554962 467472 555018 467528
rect 554778 463800 554834 463856
rect 554594 457272 554650 457328
rect 554502 453736 554558 453792
rect 554410 451424 554466 451480
rect 554318 448976 554374 449032
rect 553950 446664 554006 446720
rect 553858 444352 553914 444408
rect 553766 441904 553822 441960
rect 553490 440136 553546 440192
rect 552202 439864 552258 439920
rect 555238 465568 555294 465624
rect 555146 462032 555202 462088
rect 555422 457952 555478 458008
rect 555330 455504 555386 455560
rect 555054 447208 555110 447264
rect 554962 438912 555018 438968
rect 555698 471008 555754 471064
rect 555882 470328 555938 470384
rect 555974 469240 556030 469296
rect 555790 451968 555846 452024
rect 555698 449656 555754 449712
rect 555606 446120 555662 446176
rect 556066 465024 556122 465080
rect 555974 443672 556030 443728
rect 555882 438368 555938 438424
rect 555514 437824 555570 437880
rect 554778 436600 554834 436656
rect 556066 437144 556122 437200
rect 554962 436056 555018 436112
rect 554778 435376 554834 435432
rect 554870 434832 554926 434888
rect 554778 434152 554834 434208
rect 554870 433608 554926 433664
rect 554778 433064 554834 433120
rect 554870 432384 554926 432440
rect 554778 431860 554834 431896
rect 554778 431840 554780 431860
rect 554780 431840 554832 431860
rect 554832 431840 554834 431860
rect 554870 431296 554926 431352
rect 554962 430616 555018 430672
rect 554778 430072 554834 430128
rect 554870 429528 554926 429584
rect 554870 428884 554872 428904
rect 554872 428884 554924 428904
rect 554924 428884 554926 428904
rect 554870 428848 554926 428884
rect 554778 428304 554834 428360
rect 554778 427780 554834 427816
rect 554778 427760 554780 427780
rect 554780 427760 554832 427780
rect 554832 427760 554834 427780
rect 411902 49816 411958 49872
rect 227626 46008 227682 46064
rect 227442 44648 227498 44704
rect 227258 42744 227314 42800
rect 227442 42064 227498 42120
rect 226430 40704 226486 40760
rect 226338 40160 226394 40216
rect 227534 41384 227590 41440
rect 580262 686296 580318 686352
rect 579618 651072 579674 651128
rect 578882 604152 578938 604208
rect 580170 580760 580226 580816
rect 580170 557232 580226 557288
rect 579618 510312 579674 510368
rect 580170 463392 580226 463448
rect 580170 416472 580226 416528
rect 580170 369552 580226 369608
rect 580170 322632 580226 322688
rect 580170 275712 580226 275768
rect 579986 228792 580042 228848
rect 579986 181872 580042 181928
rect 580170 134816 580226 134872
rect 580170 87896 580226 87952
rect 580354 639376 580410 639432
rect 580446 592456 580502 592512
rect 580906 545536 580962 545592
rect 580906 498616 580962 498672
rect 580906 451696 580962 451752
rect 580906 404776 580962 404832
rect 580906 357856 580962 357912
rect 580354 310800 580410 310856
rect 580906 310800 580962 310856
rect 580354 263880 580410 263936
rect 580906 263880 580962 263936
rect 580906 216960 580962 217016
rect 580906 170040 580962 170096
rect 580906 123120 580962 123176
rect 580906 76200 580962 76256
rect 226614 39480 226670 39536
rect 227074 38800 227130 38856
rect 227442 38120 227498 38176
rect 226706 37576 226762 37632
rect 580170 40976 580226 41032
rect 563702 38664 563758 38720
rect 227534 36896 227590 36952
rect 227442 36216 227498 36272
rect 226706 35536 226762 35592
rect 227442 34856 227498 34912
rect 227442 34312 227498 34368
rect 227350 33632 227406 33688
rect 227442 32952 227498 33008
rect 116398 32000 116454 32056
rect 95146 31864 95202 31920
rect 32310 31728 32366 31784
rect 215114 32428 215170 32464
rect 215114 32408 215116 32428
rect 215116 32408 215168 32428
rect 215168 32408 215170 32428
rect 227534 32272 227590 32328
rect 213918 31728 213974 31784
rect 227442 31728 227498 31784
rect 12438 4800 12494 4856
rect 25502 3304 25558 3360
rect 119986 30232 120042 30288
rect 113178 3868 113234 3904
rect 113178 3848 113180 3868
rect 113180 3848 113232 3868
rect 113232 3848 113234 3868
rect 113454 3596 113510 3632
rect 113454 3576 113456 3596
rect 113456 3576 113508 3596
rect 113508 3576 113510 3596
rect 116030 3596 116086 3632
rect 116030 3576 116032 3596
rect 116032 3576 116084 3596
rect 116084 3576 116086 3596
rect 118698 3868 118754 3904
rect 118698 3848 118700 3868
rect 118700 3848 118752 3868
rect 118752 3848 118754 3868
rect 122930 4292 122932 4312
rect 122932 4292 122984 4312
rect 122984 4292 122986 4312
rect 122930 4256 122986 4292
rect 127806 7520 127862 7576
rect 125690 4292 125692 4312
rect 125692 4292 125744 4312
rect 125744 4292 125746 4312
rect 125690 4256 125746 4292
rect 129002 11600 129058 11656
rect 128358 4800 128414 4856
rect 131394 7656 131450 7712
rect 129830 3576 129886 3632
rect 134890 8880 134946 8936
rect 133234 3612 133236 3632
rect 133236 3612 133288 3632
rect 133288 3612 133290 3632
rect 133234 3576 133290 3612
rect 136086 10240 136142 10296
rect 138478 9016 138534 9072
rect 138202 3304 138258 3360
rect 140686 14456 140742 14512
rect 142066 10376 142122 10432
rect 140962 6160 141018 6216
rect 144182 14592 144238 14648
rect 145654 10512 145710 10568
rect 148046 7792 148102 7848
rect 151542 7928 151598 7984
rect 156326 11736 156382 11792
rect 155130 8064 155186 8120
rect 158718 8200 158774 8256
rect 164698 11872 164754 11928
rect 171782 12008 171838 12064
rect 182178 3596 182234 3632
rect 182178 3576 182180 3596
rect 182180 3576 182232 3596
rect 182232 3576 182234 3596
rect 184570 9696 184626 9752
rect 184754 9696 184810 9752
rect 182638 3596 182694 3632
rect 182638 3576 182640 3596
rect 182640 3576 182692 3596
rect 182692 3576 182694 3596
rect 201498 4800 201554 4856
rect 231950 30232 232006 30288
rect 284574 30232 284630 30288
rect 411258 27548 411260 27568
rect 411260 27548 411312 27568
rect 411312 27548 411314 27568
rect 411258 27512 411314 27548
rect 205086 4936 205142 4992
rect 206282 9152 206338 9208
rect 212262 5072 212318 5128
rect 232502 12960 232558 13016
rect 239402 13096 239458 13152
rect 250442 13368 250498 13424
rect 243542 13232 243598 13288
rect 246302 12144 246358 12200
rect 278870 3304 278926 3360
rect 283654 6296 283710 6352
rect 285954 3440 286010 3496
rect 293130 3576 293186 3632
rect 342902 2372 342958 2408
rect 342902 2352 342904 2372
rect 342904 2352 342956 2372
rect 342956 2352 342958 2372
rect 347686 2372 347742 2408
rect 347686 2352 347688 2372
rect 347688 2352 347740 2372
rect 347740 2352 347742 2372
rect 381542 2100 381598 2136
rect 381542 2080 381544 2100
rect 381544 2080 381596 2100
rect 381596 2080 381598 2100
rect 386326 2100 386382 2136
rect 386326 2080 386328 2100
rect 386328 2080 386380 2100
rect 386380 2080 386382 2100
rect 410430 12824 410486 12880
rect 412546 12860 412548 12880
rect 412548 12860 412600 12880
rect 412600 12860 412602 12880
rect 412546 12824 412602 12860
rect 414938 11600 414994 11656
rect 414570 7520 414626 7576
rect 415398 2388 415400 2408
rect 415400 2388 415452 2408
rect 415452 2388 415454 2408
rect 415398 2352 415454 2388
rect 415674 7656 415730 7712
rect 417238 10240 417294 10296
rect 416870 8880 416926 8936
rect 418342 14456 418398 14512
rect 417698 9016 417754 9072
rect 419538 14592 419594 14648
rect 419170 10376 419226 10432
rect 418526 6160 418582 6216
rect 420274 10512 420330 10568
rect 421102 7792 421158 7848
rect 422298 13796 422354 13832
rect 422298 13776 422300 13796
rect 422300 13776 422352 13796
rect 422352 13776 422354 13796
rect 422298 12860 422300 12880
rect 422300 12860 422352 12880
rect 422352 12860 422354 12880
rect 422298 12824 422354 12860
rect 422574 12144 422630 12200
rect 423402 8064 423458 8120
rect 422206 7928 422262 7984
rect 421378 3712 421434 3768
rect 423770 11736 423826 11792
rect 425426 13812 425428 13832
rect 425428 13812 425480 13832
rect 425480 13812 425482 13832
rect 425426 13776 425482 13812
rect 425702 13096 425758 13152
rect 424506 8200 424562 8256
rect 426806 12960 426862 13016
rect 426438 11872 426494 11928
rect 424966 2388 424968 2408
rect 424968 2388 425020 2408
rect 425020 2388 425022 2408
rect 424966 2352 425022 2388
rect 428002 13232 428058 13288
rect 428738 12008 428794 12064
rect 426530 3712 426586 3768
rect 430302 13368 430358 13424
rect 429106 3304 429162 3360
rect 430486 3440 430542 3496
rect 431866 12860 431868 12880
rect 431868 12860 431920 12880
rect 431920 12860 431922 12880
rect 431866 12824 431922 12860
rect 431682 3576 431738 3632
rect 434810 9696 434866 9752
rect 434718 2388 434720 2408
rect 434720 2388 434772 2408
rect 434772 2388 434774 2408
rect 434718 2352 434774 2388
rect 435454 9832 435510 9888
rect 437478 4800 437534 4856
rect 438858 4936 438914 4992
rect 439870 9152 439926 9208
rect 441802 5072 441858 5128
rect 442078 2372 442134 2408
rect 442078 2352 442080 2372
rect 442080 2352 442132 2372
rect 442132 2352 442134 2372
rect 446954 9832 447010 9888
rect 447230 9696 447286 9752
rect 463790 6296 463846 6352
rect 580906 29280 580962 29336
<< metal3 >>
rect 317086 700572 317092 700636
rect 317156 700634 317162 700636
rect 348785 700634 348851 700637
rect 317156 700632 348851 700634
rect 317156 700576 348790 700632
rect 348846 700576 348851 700632
rect 317156 700574 348851 700576
rect 317156 700572 317162 700574
rect 348785 700571 348851 700574
rect 317270 700436 317276 700500
rect 317340 700498 317346 700500
rect 478505 700498 478571 700501
rect 317340 700496 478571 700498
rect 317340 700440 478510 700496
rect 478566 700440 478571 700496
rect 317340 700438 478571 700440
rect 317340 700436 317346 700438
rect 478505 700435 478571 700438
rect 316902 700300 316908 700364
rect 316972 700362 316978 700364
rect 543457 700362 543523 700365
rect 316972 700360 543523 700362
rect 316972 700304 543462 700360
rect 543518 700304 543523 700360
rect 316972 700302 543523 700304
rect 316972 700300 316978 700302
rect 543457 700299 543523 700302
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 580257 686354 580323 686357
rect 583520 686354 584960 686444
rect 580257 686352 584960 686354
rect 580257 686296 580262 686352
rect 580318 686296 584960 686352
rect 580257 686294 584960 686296
rect 580257 686291 580323 686294
rect 583520 686204 584960 686294
rect 282913 683226 282979 683229
rect 283281 683226 283347 683229
rect 282913 683224 283347 683226
rect 282913 683168 282918 683224
rect 282974 683168 283286 683224
rect 283342 683168 283347 683224
rect 282913 683166 283347 683168
rect 282913 683163 282979 683166
rect 283281 683163 283347 683166
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 583520 674508 584960 674748
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 492438 663852 492444 663916
rect 492508 663914 492514 663916
rect 506013 663914 506079 663917
rect 492508 663912 506079 663914
rect 492508 663856 506018 663912
rect 506074 663856 506079 663912
rect 492508 663854 506079 663856
rect 492508 663852 492514 663854
rect 506013 663851 506079 663854
rect 583520 662676 584960 662916
rect 548374 662084 548380 662148
rect 548444 662146 548450 662148
rect 548444 662086 551386 662146
rect 548444 662084 548450 662086
rect 551326 661844 551386 662086
rect 551326 660108 551386 660620
rect 551318 660044 551324 660108
rect 551388 660044 551394 660108
rect 551510 658884 551570 659396
rect 551502 658820 551508 658884
rect 551572 658820 551578 658884
rect 553342 658202 553348 658204
rect 551908 658142 553348 658202
rect 553342 658140 553348 658142
rect 553412 658140 553418 658204
rect 553526 656978 553532 656980
rect 551908 656918 553532 656978
rect 553526 656916 553532 656918
rect 553596 656916 553602 656980
rect 553710 655754 553716 655756
rect 551908 655694 553716 655754
rect 553710 655692 553716 655694
rect 553780 655692 553786 655756
rect 552790 654530 552796 654532
rect 551908 654470 552796 654530
rect 552790 654468 552796 654470
rect 552860 654468 552866 654532
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 551326 653172 551386 653276
rect 551318 653108 551324 653172
rect 551388 653108 551394 653172
rect 551878 651538 551938 652052
rect 552054 651538 552060 651540
rect 551878 651478 552060 651538
rect 552054 651476 552060 651478
rect 552124 651476 552130 651540
rect 579613 651130 579679 651133
rect 583520 651130 584960 651220
rect 579613 651128 584960 651130
rect 579613 651072 579618 651128
rect 579674 651072 584960 651128
rect 579613 651070 584960 651072
rect 579613 651067 579679 651070
rect 583520 650980 584960 651070
rect 553894 650858 553900 650860
rect 551908 650798 553900 650858
rect 553894 650796 553900 650798
rect 553964 650796 553970 650860
rect 551326 649092 551386 649604
rect 551318 649028 551324 649092
rect 551388 649028 551394 649092
rect 552238 648410 552244 648412
rect 551908 648350 552244 648410
rect 552238 648348 552244 648350
rect 552308 648348 552314 648412
rect 552422 647186 552428 647188
rect 551908 647126 552428 647186
rect 552422 647124 552428 647126
rect 552492 647124 552498 647188
rect 551326 645828 551386 645932
rect 551318 645764 551324 645828
rect 551388 645764 551394 645828
rect 552606 644738 552612 644740
rect 551908 644678 552612 644738
rect 552606 644676 552612 644678
rect 552676 644676 552682 644740
rect 554078 643514 554084 643516
rect 551908 643454 554084 643514
rect 554078 643452 554084 643454
rect 554148 643452 554154 643516
rect 551878 641746 551938 642260
rect 552013 641746 552079 641749
rect 551878 641744 552079 641746
rect 551878 641688 552018 641744
rect 552074 641688 552079 641744
rect 551878 641686 552079 641688
rect 552013 641683 552079 641686
rect 553393 641066 553459 641069
rect 551908 641064 553459 641066
rect 551908 641008 553398 641064
rect 553454 641008 553459 641064
rect 551908 641006 553459 641008
rect 553393 641003 553459 641006
rect 552197 639978 552263 639981
rect 551908 639976 552263 639978
rect 551908 639920 552202 639976
rect 552258 639920 552263 639976
rect 551908 639918 552263 639920
rect 552197 639915 552263 639918
rect 551318 639644 551324 639708
rect 551388 639644 551394 639708
rect 551326 639436 551386 639644
rect 551502 639508 551508 639572
rect 551572 639570 551578 639572
rect 551645 639570 551711 639573
rect 551572 639568 551711 639570
rect 551572 639512 551650 639568
rect 551706 639512 551711 639568
rect 551572 639510 551711 639512
rect 551572 639508 551578 639510
rect 551645 639507 551711 639510
rect 551318 639372 551324 639436
rect 551388 639372 551394 639436
rect 580349 639434 580415 639437
rect 583520 639434 584960 639524
rect 580349 639432 584960 639434
rect 580349 639376 580354 639432
rect 580410 639376 584960 639432
rect 580349 639374 584960 639376
rect 580349 639371 580415 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 552105 638754 552171 638757
rect 551908 638752 552171 638754
rect 551908 638696 552110 638752
rect 552166 638696 552171 638752
rect 551908 638694 552171 638696
rect 552105 638691 552171 638694
rect 552289 637530 552355 637533
rect 551908 637528 552355 637530
rect 551908 637472 552294 637528
rect 552350 637472 552355 637528
rect 551908 637470 552355 637472
rect 552289 637467 552355 637470
rect 551326 636036 551386 636276
rect 551318 635972 551324 636036
rect 551388 635972 551394 636036
rect 456057 635218 456123 635221
rect 454020 635216 456123 635218
rect 454020 635160 456062 635216
rect 456118 635160 456123 635216
rect 454020 635158 456123 635160
rect 456057 635155 456123 635158
rect 551878 634948 551938 635052
rect 551870 634884 551876 634948
rect 551940 634884 551946 634948
rect 553485 633858 553551 633861
rect 551908 633856 553551 633858
rect 551908 633800 553490 633856
rect 553546 633800 553551 633856
rect 551908 633798 553551 633800
rect 553485 633795 553551 633798
rect 551326 632229 551386 632604
rect 551326 632224 551435 632229
rect 551326 632168 551374 632224
rect 551430 632168 551435 632224
rect 551326 632166 551435 632168
rect 551369 632163 551435 632166
rect 552381 631410 552447 631413
rect 551908 631408 552447 631410
rect 551908 631352 552386 631408
rect 552442 631352 552447 631408
rect 551908 631350 552447 631352
rect 552381 631347 552447 631350
rect 553577 630186 553643 630189
rect 551908 630184 553643 630186
rect 551908 630128 553582 630184
rect 553638 630128 553643 630184
rect 551908 630126 553643 630128
rect 553577 630123 553643 630126
rect 551510 628421 551570 628932
rect 551510 628416 551619 628421
rect 551510 628360 551558 628416
rect 551614 628360 551619 628416
rect 551510 628358 551619 628360
rect 551553 628355 551619 628358
rect 551369 628012 551435 628013
rect 551318 628010 551324 628012
rect 551278 627950 551324 628010
rect 551388 628008 551435 628012
rect 551645 628012 551711 628013
rect 551645 628010 551692 628012
rect 551430 627952 551435 628008
rect 551318 627948 551324 627950
rect 551388 627948 551435 627952
rect 551600 628008 551692 628010
rect 551600 627952 551650 628008
rect 551600 627950 551692 627952
rect 551369 627947 551435 627948
rect 551645 627948 551692 627950
rect 551756 627948 551762 628012
rect 551645 627947 551711 627948
rect 553761 627738 553827 627741
rect 551908 627736 553827 627738
rect 551908 627680 553766 627736
rect 553822 627680 553827 627736
rect 551908 627678 553827 627680
rect 553761 627675 553827 627678
rect 583520 627588 584960 627828
rect 553669 626514 553735 626517
rect 551908 626512 553735 626514
rect 551908 626456 553674 626512
rect 553730 626456 553735 626512
rect 551908 626454 553735 626456
rect 553669 626451 553735 626454
rect 553853 625290 553919 625293
rect 551908 625288 553919 625290
rect 551908 625232 553858 625288
rect 553914 625232 553919 625288
rect 551908 625230 553919 625232
rect 553853 625227 553919 625230
rect -960 624882 480 624972
rect 3417 624882 3483 624885
rect -960 624880 3483 624882
rect -960 624824 3422 624880
rect 3478 624824 3483 624880
rect -960 624822 3483 624824
rect -960 624732 480 624822
rect 3417 624819 3483 624822
rect 552473 624066 552539 624069
rect 551908 624064 552539 624066
rect 551908 624008 552478 624064
rect 552534 624008 552539 624064
rect 551908 624006 552539 624008
rect 552473 624003 552539 624006
rect 551510 622437 551570 622812
rect 113398 622372 113404 622436
rect 113468 622434 113474 622436
rect 116577 622434 116643 622437
rect 113468 622432 116643 622434
rect 113468 622376 116582 622432
rect 116638 622376 116643 622432
rect 113468 622374 116643 622376
rect 113468 622372 113474 622374
rect 116577 622371 116643 622374
rect 551461 622432 551570 622437
rect 551461 622376 551466 622432
rect 551522 622376 551570 622432
rect 551461 622374 551570 622376
rect 551461 622371 551527 622374
rect 551326 621349 551386 621588
rect 551326 621344 551435 621349
rect 551326 621288 551374 621344
rect 551430 621288 551435 621344
rect 551326 621286 551435 621288
rect 551369 621283 551435 621286
rect 553945 620394 554011 620397
rect 551908 620392 554011 620394
rect 551908 620336 553950 620392
rect 554006 620336 554011 620392
rect 551908 620334 554011 620336
rect 553945 620331 554011 620334
rect 551369 618628 551435 618629
rect 551318 618564 551324 618628
rect 551388 618626 551435 618628
rect 551388 618624 551480 618626
rect 551430 618568 551480 618624
rect 551388 618566 551480 618568
rect 551388 618564 551435 618566
rect 551369 618563 551435 618564
rect 551553 618490 551619 618493
rect 551694 618490 551754 619140
rect 551553 618488 551754 618490
rect 551553 618432 551558 618488
rect 551614 618432 551754 618488
rect 551553 618430 551754 618432
rect 551553 618427 551619 618430
rect 279141 618354 279207 618357
rect 280654 618354 280660 618356
rect 279141 618352 280660 618354
rect 279141 618296 279146 618352
rect 279202 618296 280660 618352
rect 279141 618294 280660 618296
rect 279141 618291 279207 618294
rect 280654 618292 280660 618294
rect 280724 618292 280730 618356
rect 551318 618292 551324 618356
rect 551388 618354 551394 618356
rect 551686 618354 551692 618356
rect 551388 618294 551692 618354
rect 551388 618292 551394 618294
rect 551686 618292 551692 618294
rect 551756 618292 551762 618356
rect 554129 617946 554195 617949
rect 551908 617944 554195 617946
rect 551908 617888 554134 617944
rect 554190 617888 554195 617944
rect 551908 617886 554195 617888
rect 554129 617883 554195 617886
rect 106222 617612 106228 617676
rect 106292 617674 106298 617676
rect 113398 617674 113404 617676
rect 106292 617614 113404 617674
rect 106292 617612 106298 617614
rect 113398 617612 113404 617614
rect 113468 617612 113474 617676
rect 551369 617540 551435 617541
rect 551318 617538 551324 617540
rect 551278 617478 551324 617538
rect 551388 617536 551435 617540
rect 551430 617480 551435 617536
rect 551318 617476 551324 617478
rect 551388 617476 551435 617480
rect 551369 617475 551435 617476
rect 25446 617340 25452 617404
rect 25516 617402 25522 617404
rect 25516 617342 28060 617402
rect 25516 617340 25522 617342
rect 27654 616796 27660 616860
rect 27724 616858 27730 616860
rect 554221 616858 554287 616861
rect 27724 616798 28060 616858
rect 551908 616856 554287 616858
rect 551908 616800 554226 616856
rect 554282 616800 554287 616856
rect 551908 616798 554287 616800
rect 27724 616796 27730 616798
rect 554221 616795 554287 616798
rect 551318 616388 551324 616452
rect 551388 616450 551394 616452
rect 551645 616450 551711 616453
rect 551388 616448 551711 616450
rect 551388 616392 551650 616448
rect 551706 616392 551711 616448
rect 551388 616390 551711 616392
rect 551388 616388 551394 616390
rect 551645 616387 551711 616390
rect 456793 616314 456859 616317
rect 456793 616312 460092 616314
rect 456793 616256 456798 616312
rect 456854 616256 460092 616312
rect 456793 616254 460092 616256
rect 456793 616251 456859 616254
rect 27470 616116 27476 616180
rect 27540 616178 27546 616180
rect 27540 616118 28060 616178
rect 27540 616116 27546 616118
rect 21214 615708 21220 615772
rect 21284 615770 21290 615772
rect 22134 615770 22140 615772
rect 21284 615710 22140 615770
rect 21284 615708 21290 615710
rect 22134 615708 22140 615710
rect 22204 615708 22210 615772
rect 28574 615708 28580 615772
rect 28644 615708 28650 615772
rect 583520 615756 584960 615996
rect 28582 615604 28642 615708
rect 554037 615634 554103 615637
rect 551908 615632 554103 615634
rect 551908 615576 554042 615632
rect 554098 615576 554103 615632
rect 551908 615574 554103 615576
rect 554037 615571 554103 615574
rect 27286 614892 27292 614956
rect 27356 614954 27362 614956
rect 27356 614894 28060 614954
rect 27356 614892 27362 614894
rect 25262 614348 25268 614412
rect 25332 614410 25338 614412
rect 552565 614410 552631 614413
rect 25332 614350 28060 614410
rect 551908 614408 552631 614410
rect 551908 614352 552570 614408
rect 552626 614352 552631 614408
rect 551908 614350 552631 614352
rect 25332 614348 25338 614350
rect 552565 614347 552631 614350
rect 27102 613804 27108 613868
rect 27172 613866 27178 613868
rect 27172 613806 28060 613866
rect 27172 613804 27178 613806
rect 551318 613804 551324 613868
rect 551388 613866 551394 613868
rect 551645 613866 551711 613869
rect 551388 613864 551711 613866
rect 551388 613808 551650 613864
rect 551706 613808 551711 613864
rect 551388 613806 551711 613808
rect 551388 613804 551394 613806
rect 551645 613803 551711 613806
rect 551318 613668 551324 613732
rect 551388 613730 551394 613732
rect 551737 613730 551803 613733
rect 551388 613728 551803 613730
rect 551388 613672 551742 613728
rect 551798 613672 551803 613728
rect 551388 613670 551803 613672
rect 551388 613668 551394 613670
rect 551737 613667 551803 613670
rect 313273 613458 313339 613461
rect 313273 613456 316204 613458
rect 313273 613400 313278 613456
rect 313334 613400 316204 613456
rect 313273 613398 316204 613400
rect 313273 613395 313339 613398
rect 28214 612780 28274 613156
rect 551510 612781 551570 613156
rect 28206 612716 28212 612780
rect 28276 612716 28282 612780
rect 551510 612776 551619 612781
rect 551510 612720 551558 612776
rect 551614 612720 551619 612776
rect 551510 612718 551619 612720
rect 551553 612715 551619 612718
rect 28030 612100 28090 612612
rect 551502 612308 551508 612372
rect 551572 612370 551578 612372
rect 551686 612370 551692 612372
rect 551572 612310 551692 612370
rect 551572 612308 551578 612310
rect 551686 612308 551692 612310
rect 551756 612308 551762 612372
rect 551318 612172 551324 612236
rect 551388 612234 551394 612236
rect 551645 612234 551711 612237
rect 551388 612232 551711 612234
rect 551388 612176 551650 612232
rect 551706 612176 551711 612232
rect 551388 612174 551711 612176
rect 551388 612172 551394 612174
rect 551645 612171 551711 612174
rect 28022 612036 28028 612100
rect 28092 612036 28098 612100
rect 28582 611557 28642 611932
rect 551694 611693 551754 611932
rect 551645 611688 551754 611693
rect 551645 611632 551650 611688
rect 551706 611632 551754 611688
rect 551645 611630 551754 611632
rect 551645 611627 551711 611630
rect 28582 611552 28691 611557
rect 28582 611496 28630 611552
rect 28686 611496 28691 611552
rect 28582 611494 28691 611496
rect 28625 611491 28691 611494
rect 26918 611356 26924 611420
rect 26988 611418 26994 611420
rect 26988 611358 28060 611418
rect 26988 611356 26994 611358
rect 27838 610812 27844 610876
rect 27908 610874 27914 610876
rect 27908 610814 28060 610874
rect 27908 610812 27914 610814
rect 554313 610738 554379 610741
rect 551908 610736 554379 610738
rect 551908 610680 554318 610736
rect 554374 610680 554379 610736
rect 551908 610678 554379 610680
rect 554313 610675 554379 610678
rect -960 610466 480 610556
rect 3325 610466 3391 610469
rect -960 610464 3391 610466
rect -960 610408 3330 610464
rect 3386 610408 3391 610464
rect -960 610406 3391 610408
rect -960 610316 480 610406
rect 3325 610403 3391 610406
rect 26734 610132 26740 610196
rect 26804 610194 26810 610196
rect 26804 610134 28060 610194
rect 26804 610132 26810 610134
rect 27705 609650 27771 609653
rect 27705 609648 28060 609650
rect 27705 609592 27710 609648
rect 27766 609592 28060 609648
rect 27705 609590 28060 609592
rect 27705 609587 27771 609590
rect 554405 609514 554471 609517
rect 551908 609512 554471 609514
rect 551908 609456 554410 609512
rect 554466 609456 554471 609512
rect 551908 609454 554471 609456
rect 554405 609451 554471 609454
rect 27521 608970 27587 608973
rect 27521 608968 28060 608970
rect 27521 608912 27526 608968
rect 27582 608912 28060 608968
rect 27521 608910 28060 608912
rect 27521 608907 27587 608910
rect 284293 608834 284359 608837
rect 282686 608832 284359 608834
rect 282686 608776 284298 608832
rect 284354 608776 284359 608832
rect 282686 608774 284359 608776
rect 282686 608668 282746 608774
rect 284293 608771 284359 608774
rect 27613 608426 27679 608429
rect 27613 608424 28060 608426
rect 27613 608368 27618 608424
rect 27674 608368 28060 608424
rect 27613 608366 28060 608368
rect 27613 608363 27679 608366
rect 553025 608290 553091 608293
rect 551908 608288 553091 608290
rect 551908 608232 553030 608288
rect 553086 608232 553091 608288
rect 551908 608230 553091 608232
rect 553025 608227 553091 608230
rect 28582 607341 28642 607716
rect 28582 607336 28691 607341
rect 28582 607280 28630 607336
rect 28686 607280 28691 607336
rect 28582 607278 28691 607280
rect 28625 607275 28691 607278
rect 27153 607202 27219 607205
rect 27153 607200 28060 607202
rect 27153 607144 27158 607200
rect 27214 607144 28060 607200
rect 27153 607142 28060 607144
rect 27153 607139 27219 607142
rect 554497 607066 554563 607069
rect 551908 607064 554563 607066
rect 551908 607008 554502 607064
rect 554558 607008 554563 607064
rect 551908 607006 554563 607008
rect 554497 607003 554563 607006
rect 27429 606658 27495 606661
rect 27429 606656 28060 606658
rect 27429 606600 27434 606656
rect 27490 606600 28060 606656
rect 27429 606598 28060 606600
rect 27429 606595 27495 606598
rect 27245 605978 27311 605981
rect 27245 605976 28060 605978
rect 27245 605920 27250 605976
rect 27306 605920 28060 605976
rect 27245 605918 28060 605920
rect 27245 605915 27311 605918
rect 553117 605842 553183 605845
rect 551908 605840 553183 605842
rect 551908 605784 553122 605840
rect 553178 605784 553183 605840
rect 551908 605782 553183 605784
rect 553117 605779 553183 605782
rect 27797 605434 27863 605437
rect 27797 605432 28060 605434
rect 27797 605376 27802 605432
rect 27858 605376 28060 605432
rect 27797 605374 28060 605376
rect 27797 605371 27863 605374
rect 25998 604692 26004 604756
rect 26068 604754 26074 604756
rect 26068 604694 28060 604754
rect 26068 604692 26074 604694
rect 552657 604618 552723 604621
rect 551908 604616 552723 604618
rect 551908 604560 552662 604616
rect 552718 604560 552723 604616
rect 551908 604558 552723 604560
rect 552657 604555 552723 604558
rect 27337 604210 27403 604213
rect 578877 604210 578943 604213
rect 583520 604210 584960 604300
rect 27337 604208 28060 604210
rect 27337 604152 27342 604208
rect 27398 604152 28060 604208
rect 27337 604150 28060 604152
rect 578877 604208 584960 604210
rect 578877 604152 578882 604208
rect 578938 604152 584960 604208
rect 578877 604150 584960 604152
rect 27337 604147 27403 604150
rect 578877 604147 578943 604150
rect 583520 604060 584960 604150
rect 25814 603604 25820 603668
rect 25884 603666 25890 603668
rect 25884 603606 28060 603666
rect 25884 603604 25890 603606
rect 553209 603394 553275 603397
rect 551908 603392 553275 603394
rect 551908 603336 553214 603392
rect 553270 603336 553275 603392
rect 551908 603334 553275 603336
rect 553209 603331 553275 603334
rect 28582 602581 28642 602956
rect 28533 602576 28642 602581
rect 28533 602520 28538 602576
rect 28594 602520 28642 602576
rect 28533 602518 28642 602520
rect 28533 602515 28599 602518
rect 27889 602034 27955 602037
rect 28030 602034 28090 602412
rect 27889 602032 28090 602034
rect 27889 601976 27894 602032
rect 27950 601976 28090 602032
rect 27889 601974 28090 601976
rect 27889 601971 27955 601974
rect 28073 601898 28139 601901
rect 28030 601896 28139 601898
rect 28030 601840 28078 601896
rect 28134 601840 28139 601896
rect 28030 601835 28139 601840
rect 28030 601732 28090 601835
rect 551326 601629 551386 602140
rect 551326 601624 551435 601629
rect 551326 601568 551374 601624
rect 551430 601568 551435 601624
rect 551326 601566 551435 601568
rect 551369 601563 551435 601566
rect 27061 601218 27127 601221
rect 27061 601216 28060 601218
rect 27061 601160 27066 601216
rect 27122 601160 28060 601216
rect 27061 601158 28060 601160
rect 27061 601155 27127 601158
rect 551502 601156 551508 601220
rect 551572 601218 551578 601220
rect 551737 601218 551803 601221
rect 551572 601216 551803 601218
rect 551572 601160 551742 601216
rect 551798 601160 551803 601216
rect 551572 601158 551803 601160
rect 551572 601156 551578 601158
rect 551737 601155 551803 601158
rect 28582 600269 28642 600508
rect 551694 600405 551754 600916
rect 551694 600400 551803 600405
rect 551694 600344 551742 600400
rect 551798 600344 551803 600400
rect 551694 600342 551803 600344
rect 551737 600339 551803 600342
rect 28582 600264 28691 600269
rect 28582 600208 28630 600264
rect 28686 600208 28691 600264
rect 28582 600206 28691 600208
rect 28625 600203 28691 600206
rect 551369 599996 551435 599997
rect 25630 599932 25636 599996
rect 25700 599994 25706 599996
rect 25700 599934 28060 599994
rect 25700 599932 25706 599934
rect 551318 599932 551324 599996
rect 551388 599994 551435 599996
rect 551388 599992 551480 599994
rect 551430 599936 551480 599992
rect 551388 599934 551480 599936
rect 551388 599932 551435 599934
rect 551369 599931 551435 599932
rect 552749 599722 552815 599725
rect 551908 599720 552815 599722
rect 551908 599664 552754 599720
rect 552810 599664 552815 599720
rect 551908 599662 552815 599664
rect 552749 599659 552815 599662
rect 551318 599524 551324 599588
rect 551388 599586 551394 599588
rect 551686 599586 551692 599588
rect 551388 599526 551692 599586
rect 551388 599524 551394 599526
rect 551686 599524 551692 599526
rect 551756 599524 551762 599588
rect 28582 598909 28642 599420
rect 28533 598904 28642 598909
rect 28533 598848 28538 598904
rect 28594 598848 28642 598904
rect 28533 598846 28642 598848
rect 28533 598843 28599 598846
rect 26969 598770 27035 598773
rect 26969 598768 28060 598770
rect 26969 598712 26974 598768
rect 27030 598712 28060 598768
rect 26969 598710 28060 598712
rect 26969 598707 27035 598710
rect 28030 597685 28090 598196
rect 551878 597957 551938 598468
rect 551829 597952 551938 597957
rect 551829 597896 551834 597952
rect 551890 597896 551938 597952
rect 551829 597894 551938 597896
rect 551829 597891 551895 597894
rect 27981 597680 28090 597685
rect 27981 597624 27986 597680
rect 28042 597624 28090 597680
rect 27981 597622 28090 597624
rect 27981 597619 28047 597622
rect 28214 597141 28274 597516
rect 552841 597274 552907 597277
rect 551908 597272 552907 597274
rect 551908 597216 552846 597272
rect 552902 597216 552907 597272
rect 551908 597214 552907 597216
rect 552841 597211 552907 597214
rect 28165 597136 28274 597141
rect 28625 597138 28691 597141
rect 28165 597080 28170 597136
rect 28226 597080 28274 597136
rect 28165 597078 28274 597080
rect 28582 597136 28691 597138
rect 28582 597080 28630 597136
rect 28686 597080 28691 597136
rect 28165 597075 28231 597078
rect 28582 597075 28691 597080
rect 28582 596972 28642 597075
rect 26785 596458 26851 596461
rect 26785 596456 28060 596458
rect 26785 596400 26790 596456
rect 26846 596400 28060 596456
rect 26785 596398 28060 596400
rect 26785 596395 26851 596398
rect -960 596050 480 596140
rect 3509 596050 3575 596053
rect 553301 596050 553367 596053
rect -960 596048 3575 596050
rect -960 595992 3514 596048
rect 3570 595992 3575 596048
rect -960 595990 3575 595992
rect 551908 596048 553367 596050
rect 551908 595992 553306 596048
rect 553362 595992 553367 596048
rect 551908 595990 553367 595992
rect -960 595900 480 595990
rect 3509 595987 3575 595990
rect 553301 595987 553367 595990
rect 28398 595373 28458 595748
rect 28398 595368 28507 595373
rect 28398 595312 28446 595368
rect 28502 595312 28507 595368
rect 28398 595310 28507 595312
rect 28441 595307 28507 595310
rect 26877 595234 26943 595237
rect 551369 595234 551435 595237
rect 26877 595232 28060 595234
rect 26877 595176 26882 595232
rect 26938 595176 28060 595232
rect 26877 595174 28060 595176
rect 551369 595232 551754 595234
rect 551369 595176 551374 595232
rect 551430 595176 551754 595232
rect 551369 595174 551754 595176
rect 26877 595171 26943 595174
rect 551369 595171 551435 595174
rect 551369 595100 551435 595101
rect 551694 595100 551754 595174
rect 551318 595098 551324 595100
rect 551278 595038 551324 595098
rect 551388 595096 551435 595100
rect 551430 595040 551435 595096
rect 551318 595036 551324 595038
rect 551388 595036 551435 595040
rect 551686 595036 551692 595100
rect 551756 595036 551762 595100
rect 551369 595035 551435 595036
rect 139577 594826 139643 594829
rect 552933 594826 552999 594829
rect 139534 594824 139643 594826
rect 139534 594768 139582 594824
rect 139638 594768 139643 594824
rect 139534 594763 139643 594768
rect 551908 594824 552999 594826
rect 551908 594768 552938 594824
rect 552994 594768 552999 594824
rect 551908 594766 552999 594768
rect 552933 594763 552999 594766
rect 139534 594660 139594 594763
rect 28214 594149 28274 594524
rect 28214 594144 28323 594149
rect 28214 594088 28262 594144
rect 28318 594088 28323 594144
rect 28214 594086 28323 594088
rect 28257 594083 28323 594086
rect 24945 594010 25011 594013
rect 24945 594008 28060 594010
rect 24945 593952 24950 594008
rect 25006 593952 28060 594008
rect 24945 593950 28060 593952
rect 24945 593947 25011 593950
rect 554589 593738 554655 593741
rect 551908 593736 554655 593738
rect 551908 593680 554594 593736
rect 554650 593680 554655 593736
rect 551908 593678 554655 593680
rect 554589 593675 554655 593678
rect 28398 592925 28458 593300
rect 28349 592920 28458 592925
rect 28349 592864 28354 592920
rect 28410 592864 28458 592920
rect 28349 592862 28458 592864
rect 28349 592859 28415 592862
rect 26049 592786 26115 592789
rect 26049 592784 28060 592786
rect 26049 592728 26054 592784
rect 26110 592728 28060 592784
rect 26049 592726 28060 592728
rect 26049 592723 26115 592726
rect 554681 592514 554747 592517
rect 551908 592512 554747 592514
rect 551908 592456 554686 592512
rect 554742 592456 554747 592512
rect 551908 592454 554747 592456
rect 554681 592451 554747 592454
rect 580441 592514 580507 592517
rect 583520 592514 584960 592604
rect 580441 592512 584960 592514
rect 580441 592456 580446 592512
rect 580502 592456 584960 592512
rect 580441 592454 584960 592456
rect 580441 592451 580507 592454
rect 551369 592378 551435 592381
rect 551502 592378 551508 592380
rect 551369 592376 551508 592378
rect 551369 592320 551374 592376
rect 551430 592320 551508 592376
rect 551369 592318 551508 592320
rect 551369 592315 551435 592318
rect 551502 592316 551508 592318
rect 551572 592316 551578 592380
rect 583520 592364 584960 592454
rect 26693 592242 26759 592245
rect 551369 592244 551435 592245
rect 26693 592240 28060 592242
rect 26693 592184 26698 592240
rect 26754 592184 28060 592240
rect 26693 592182 28060 592184
rect 26693 592179 26759 592182
rect 551318 592180 551324 592244
rect 551388 592242 551435 592244
rect 551388 592240 551480 592242
rect 551430 592184 551480 592240
rect 551388 592182 551480 592184
rect 551388 592180 551435 592182
rect 551369 592179 551435 592180
rect 455413 591698 455479 591701
rect 454020 591696 455479 591698
rect 454020 591640 455418 591696
rect 455474 591640 455479 591696
rect 454020 591638 455479 591640
rect 455413 591635 455479 591638
rect 25865 591562 25931 591565
rect 25865 591560 28060 591562
rect 25865 591504 25870 591560
rect 25926 591504 28060 591560
rect 25865 591502 28060 591504
rect 25865 591499 25931 591502
rect 554773 591290 554839 591293
rect 551908 591288 554839 591290
rect 551908 591232 554778 591288
rect 554834 591232 554839 591288
rect 551908 591230 554839 591232
rect 554773 591227 554839 591230
rect 28582 590477 28642 590988
rect 28533 590472 28642 590477
rect 28533 590416 28538 590472
rect 28594 590416 28642 590472
rect 28533 590414 28642 590416
rect 28533 590411 28599 590414
rect 28582 590069 28642 590308
rect 28582 590064 28691 590069
rect 554589 590066 554655 590069
rect 28582 590008 28630 590064
rect 28686 590008 28691 590064
rect 28582 590006 28691 590008
rect 551908 590064 554655 590066
rect 551908 590008 554594 590064
rect 554650 590008 554655 590064
rect 551908 590006 554655 590008
rect 28625 590003 28691 590006
rect 554589 590003 554655 590006
rect 25957 589794 26023 589797
rect 25957 589792 28060 589794
rect 25957 589736 25962 589792
rect 26018 589736 28060 589792
rect 25957 589734 28060 589736
rect 25957 589731 26023 589734
rect 28398 588709 28458 589220
rect 554589 588842 554655 588845
rect 551908 588840 554655 588842
rect 551908 588784 554594 588840
rect 554650 588784 554655 588840
rect 551908 588782 554655 588784
rect 554589 588779 554655 588782
rect 28398 588704 28507 588709
rect 28398 588648 28446 588704
rect 28502 588648 28507 588704
rect 28398 588646 28507 588648
rect 28441 588643 28507 588646
rect 28214 588165 28274 588540
rect 28214 588160 28323 588165
rect 28214 588104 28262 588160
rect 28318 588104 28323 588160
rect 28214 588102 28323 588104
rect 28257 588099 28323 588102
rect 25773 588026 25839 588029
rect 25773 588024 28060 588026
rect 25773 587968 25778 588024
rect 25834 587968 28060 588024
rect 25773 587966 28060 587968
rect 25773 587963 25839 587966
rect 554589 587618 554655 587621
rect 551908 587616 554655 587618
rect 551908 587560 554594 587616
rect 554650 587560 554655 587616
rect 551908 587558 554655 587560
rect 554589 587555 554655 587558
rect 28398 586941 28458 587316
rect 551318 587148 551324 587212
rect 551388 587210 551394 587212
rect 552974 587210 552980 587212
rect 551388 587150 552980 587210
rect 551388 587148 551394 587150
rect 552974 587148 552980 587150
rect 553044 587148 553050 587212
rect 28349 586936 28458 586941
rect 28625 586938 28691 586941
rect 551369 586940 551435 586941
rect 551318 586938 551324 586940
rect 28349 586880 28354 586936
rect 28410 586880 28458 586936
rect 28349 586878 28458 586880
rect 28582 586936 28691 586938
rect 28582 586880 28630 586936
rect 28686 586880 28691 586936
rect 28349 586875 28415 586878
rect 28582 586875 28691 586880
rect 551278 586878 551324 586938
rect 551388 586936 551435 586940
rect 551430 586880 551435 586936
rect 551318 586876 551324 586878
rect 551388 586876 551435 586880
rect 551369 586875 551435 586876
rect 28582 586772 28642 586875
rect 554865 586394 554931 586397
rect 551908 586392 554931 586394
rect 551908 586336 554870 586392
rect 554926 586336 554931 586392
rect 551908 586334 554931 586336
rect 554865 586331 554931 586334
rect 551369 586260 551435 586261
rect 551318 586258 551324 586260
rect 551278 586198 551324 586258
rect 551388 586256 551435 586260
rect 551430 586200 551435 586256
rect 551318 586196 551324 586198
rect 551388 586196 551435 586200
rect 551369 586195 551435 586196
rect 282269 586122 282335 586125
rect 282269 586120 282378 586122
rect 28582 585717 28642 586092
rect 282269 586064 282274 586120
rect 282330 586064 282378 586120
rect 282269 586059 282378 586064
rect 28582 585712 28691 585717
rect 28582 585656 28630 585712
rect 28686 585656 28691 585712
rect 28582 585654 28691 585656
rect 28625 585651 28691 585654
rect 25681 585578 25747 585581
rect 25681 585576 28060 585578
rect 25681 585520 25686 585576
rect 25742 585520 28060 585576
rect 282318 585548 282378 586059
rect 25681 585518 28060 585520
rect 25681 585515 25747 585518
rect 554865 585170 554931 585173
rect 551908 585168 554931 585170
rect 551908 585112 554870 585168
rect 554926 585112 554931 585168
rect 551908 585110 554931 585112
rect 554865 585107 554931 585110
rect 26601 585034 26667 585037
rect 26601 585032 28060 585034
rect 26601 584976 26606 585032
rect 26662 584976 28060 585032
rect 26601 584974 28060 584976
rect 26601 584971 26667 584974
rect 25497 584354 25563 584357
rect 25497 584352 28060 584354
rect 25497 584296 25502 584352
rect 25558 584296 28060 584352
rect 25497 584294 28060 584296
rect 25497 584291 25563 584294
rect 25589 583810 25655 583813
rect 551878 583810 551938 583916
rect 554865 583810 554931 583813
rect 25589 583808 28060 583810
rect 25589 583752 25594 583808
rect 25650 583752 28060 583808
rect 25589 583750 28060 583752
rect 551878 583808 554931 583810
rect 551878 583752 554870 583808
rect 554926 583752 554931 583808
rect 551878 583750 554931 583752
rect 25589 583747 25655 583750
rect 554865 583747 554931 583750
rect 25313 583130 25379 583133
rect 25313 583128 28060 583130
rect 25313 583072 25318 583128
rect 25374 583072 28060 583128
rect 25313 583070 28060 583072
rect 25313 583067 25379 583070
rect 555417 582722 555483 582725
rect 551908 582720 555483 582722
rect 551908 582664 555422 582720
rect 555478 582664 555483 582720
rect 551908 582662 555483 582664
rect 555417 582659 555483 582662
rect 26509 582586 26575 582589
rect 26509 582584 28060 582586
rect 26509 582528 26514 582584
rect 26570 582528 28060 582584
rect 26509 582526 28060 582528
rect 26509 582523 26575 582526
rect 551502 582524 551508 582588
rect 551572 582586 551578 582588
rect 552974 582586 552980 582588
rect 551572 582526 552980 582586
rect 551572 582524 551578 582526
rect 552974 582524 552980 582526
rect 553044 582524 553050 582588
rect 551318 582116 551324 582180
rect 551388 582116 551394 582180
rect 551326 582045 551386 582116
rect 25221 582042 25287 582045
rect 25221 582040 28060 582042
rect 25221 581984 25226 582040
rect 25282 581984 28060 582040
rect 25221 581982 28060 581984
rect 551326 582040 551435 582045
rect 551326 581984 551374 582040
rect 551430 581984 551435 582040
rect 551326 581982 551435 581984
rect 25221 581979 25287 581982
rect 551369 581979 551435 581982
rect -960 581620 480 581860
rect 25405 581362 25471 581365
rect 25405 581360 28060 581362
rect 25405 581304 25410 581360
rect 25466 581304 28060 581360
rect 25405 581302 28060 581304
rect 25405 581299 25471 581302
rect 551878 581090 551938 581468
rect 554865 581090 554931 581093
rect 551878 581088 554931 581090
rect 551878 581032 554870 581088
rect 554926 581032 554931 581088
rect 551878 581030 554931 581032
rect 554865 581027 554931 581030
rect 25129 580818 25195 580821
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 25129 580816 28060 580818
rect 25129 580760 25134 580816
rect 25190 580760 28060 580816
rect 25129 580758 28060 580760
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 25129 580755 25195 580758
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 28582 579733 28642 580108
rect 28582 579728 28691 579733
rect 28582 579672 28630 579728
rect 28686 579672 28691 579728
rect 28582 579670 28691 579672
rect 551878 579730 551938 580244
rect 554865 579730 554931 579733
rect 551878 579728 554931 579730
rect 551878 579672 554870 579728
rect 554926 579672 554931 579728
rect 551878 579670 554931 579672
rect 28625 579667 28691 579670
rect 554865 579667 554931 579670
rect 25037 579594 25103 579597
rect 25037 579592 28060 579594
rect 25037 579536 25042 579592
rect 25098 579536 28060 579592
rect 25037 579534 28060 579536
rect 25037 579531 25103 579534
rect 26417 578914 26483 578917
rect 26417 578912 28060 578914
rect 26417 578856 26422 578912
rect 26478 578856 28060 578912
rect 26417 578854 28060 578856
rect 26417 578851 26483 578854
rect 551502 578444 551508 578508
rect 551572 578444 551578 578508
rect 551878 578506 551938 579020
rect 554865 578506 554931 578509
rect 551878 578504 554931 578506
rect 551878 578448 554870 578504
rect 554926 578448 554931 578504
rect 551878 578446 554931 578448
rect 26141 578370 26207 578373
rect 26141 578368 28060 578370
rect 26141 578312 26146 578368
rect 26202 578312 28060 578368
rect 26141 578310 28060 578312
rect 26141 578307 26207 578310
rect 283097 578234 283163 578237
rect 283281 578234 283347 578237
rect 283097 578232 283347 578234
rect 283097 578176 283102 578232
rect 283158 578176 283286 578232
rect 283342 578176 283347 578232
rect 283097 578174 283347 578176
rect 283097 578171 283163 578174
rect 283281 578171 283347 578174
rect 551318 578172 551324 578236
rect 551388 578234 551394 578236
rect 551510 578234 551570 578444
rect 554865 578443 554931 578446
rect 551388 578174 551570 578234
rect 551388 578172 551394 578174
rect 28582 577285 28642 577796
rect 551369 577556 551435 577557
rect 551318 577554 551324 577556
rect 551278 577494 551324 577554
rect 551388 577552 551435 577556
rect 551430 577496 551435 577552
rect 551318 577492 551324 577494
rect 551388 577492 551435 577496
rect 551369 577491 551435 577492
rect 28582 577280 28691 577285
rect 28582 577224 28630 577280
rect 28686 577224 28691 577280
rect 28582 577222 28691 577224
rect 551878 577282 551938 577796
rect 554865 577282 554931 577285
rect 551878 577280 554931 577282
rect 551878 577224 554870 577280
rect 554926 577224 554931 577280
rect 551878 577222 554931 577224
rect 28625 577219 28691 577222
rect 554865 577219 554931 577222
rect 28582 576741 28642 577116
rect 28582 576736 28691 576741
rect 28582 576680 28630 576736
rect 28686 576680 28691 576736
rect 28582 576678 28691 576680
rect 28625 576675 28691 576678
rect 28582 576061 28642 576572
rect 28582 576056 28691 576061
rect 28582 576000 28630 576056
rect 28686 576000 28691 576056
rect 28582 575998 28691 576000
rect 551878 576058 551938 576572
rect 553301 576058 553367 576061
rect 551878 576056 553367 576058
rect 551878 576000 553306 576056
rect 553362 576000 553367 576056
rect 551878 575998 553367 576000
rect 28625 575995 28691 575998
rect 553301 575995 553367 575998
rect 28582 575516 28642 575892
rect 28574 575452 28580 575516
rect 28644 575452 28650 575516
rect 28582 575109 28642 575348
rect 28582 575104 28691 575109
rect 28582 575048 28630 575104
rect 28686 575048 28691 575104
rect 28582 575046 28691 575048
rect 28625 575043 28691 575046
rect 28625 574970 28691 574973
rect 28582 574968 28691 574970
rect 28582 574912 28630 574968
rect 28686 574912 28691 574968
rect 28582 574907 28691 574912
rect 28582 574804 28642 574907
rect 551878 574834 551938 575348
rect 553301 574834 553367 574837
rect 551878 574832 553367 574834
rect 551878 574776 553306 574832
rect 553362 574776 553367 574832
rect 551878 574774 553367 574776
rect 553301 574771 553367 574774
rect 26233 574154 26299 574157
rect 553301 574154 553367 574157
rect 26233 574152 28060 574154
rect 26233 574096 26238 574152
rect 26294 574096 28060 574152
rect 26233 574094 28060 574096
rect 551908 574152 553367 574154
rect 551908 574096 553306 574152
rect 553362 574096 553367 574152
rect 551908 574094 553367 574096
rect 26233 574091 26299 574094
rect 553301 574091 553367 574094
rect 26325 573610 26391 573613
rect 26325 573608 28060 573610
rect 26325 573552 26330 573608
rect 26386 573552 28060 573608
rect 26325 573550 28060 573552
rect 26325 573547 26391 573550
rect 24853 572930 24919 572933
rect 553301 572930 553367 572933
rect 24853 572928 28060 572930
rect 24853 572872 24858 572928
rect 24914 572872 28060 572928
rect 24853 572870 28060 572872
rect 551908 572928 553367 572930
rect 551908 572872 553306 572928
rect 553362 572872 553367 572928
rect 551908 572870 553367 572872
rect 24853 572867 24919 572870
rect 553301 572867 553367 572870
rect 24761 572386 24827 572389
rect 24761 572384 28060 572386
rect 24761 572328 24766 572384
rect 24822 572328 28060 572384
rect 24761 572326 28060 572328
rect 24761 572323 24827 572326
rect 24669 571842 24735 571845
rect 24669 571840 28060 571842
rect 24669 571784 24674 571840
rect 24730 571784 28060 571840
rect 24669 571782 28060 571784
rect 24669 571779 24735 571782
rect 553301 571706 553367 571709
rect 551908 571704 553367 571706
rect 551908 571648 553306 571704
rect 553362 571648 553367 571704
rect 551908 571646 553367 571648
rect 553301 571643 553367 571646
rect 28574 571508 28580 571572
rect 28644 571570 28650 571572
rect 29177 571570 29243 571573
rect 28644 571568 29243 571570
rect 28644 571512 29182 571568
rect 29238 571512 29243 571568
rect 28644 571510 29243 571512
rect 28644 571508 28650 571510
rect 29177 571507 29243 571510
rect 551878 570074 551938 570588
rect 553301 570074 553367 570077
rect 551878 570072 553367 570074
rect 551878 570016 553306 570072
rect 553362 570016 553367 570072
rect 551878 570014 553367 570016
rect 553301 570011 553367 570014
rect 546350 569876 546356 569940
rect 546420 569938 546426 569940
rect 546420 569878 550650 569938
rect 546420 569876 546426 569878
rect 280286 569740 280292 569804
rect 280356 569802 280362 569804
rect 281390 569802 281396 569804
rect 280356 569742 281396 569802
rect 280356 569740 280362 569742
rect 281390 569740 281396 569742
rect 281460 569740 281466 569804
rect 550590 569802 550650 569878
rect 551502 569876 551508 569940
rect 551572 569876 551578 569940
rect 550817 569802 550883 569805
rect 550590 569800 550883 569802
rect 550590 569744 550822 569800
rect 550878 569744 550883 569800
rect 550590 569742 550883 569744
rect 550817 569739 550883 569742
rect 551001 569802 551067 569805
rect 551510 569802 551570 569876
rect 551001 569800 551570 569802
rect 551001 569744 551006 569800
rect 551062 569744 551570 569800
rect 551001 569742 551570 569744
rect 551001 569739 551067 569742
rect 551686 569740 551692 569804
rect 551756 569802 551762 569804
rect 551756 569742 551938 569802
rect 551756 569740 551762 569742
rect 550817 569530 550883 569533
rect 551878 569530 551938 569742
rect 550817 569528 551938 569530
rect 550817 569472 550822 569528
rect 550878 569472 551938 569528
rect 550817 569470 551938 569472
rect 550817 569467 550883 569470
rect 583520 568836 584960 569076
rect 326889 567898 326955 567901
rect 440509 567898 440575 567901
rect 326889 567896 440575 567898
rect 326889 567840 326894 567896
rect 326950 567840 440514 567896
rect 440570 567840 440575 567896
rect 326889 567838 440575 567840
rect 326889 567835 326955 567838
rect 440509 567835 440575 567838
rect -960 567354 480 567444
rect 3509 567354 3575 567357
rect -960 567352 3575 567354
rect -960 567296 3514 567352
rect 3570 567296 3575 567352
rect -960 567294 3575 567296
rect -960 567204 480 567294
rect 3509 567291 3575 567294
rect 280153 563818 280219 563821
rect 280286 563818 280292 563820
rect 280153 563816 280292 563818
rect 280153 563760 280158 563816
rect 280214 563760 280292 563816
rect 280153 563758 280292 563760
rect 280153 563755 280219 563758
rect 280286 563756 280292 563758
rect 280356 563756 280362 563820
rect 551001 563274 551067 563277
rect 551134 563274 551140 563276
rect 551001 563272 551140 563274
rect 551001 563216 551006 563272
rect 551062 563216 551140 563272
rect 551001 563214 551140 563216
rect 551001 563211 551067 563214
rect 551134 563212 551140 563214
rect 551204 563212 551210 563276
rect 550030 562260 550036 562324
rect 550100 562322 550106 562324
rect 551686 562322 551692 562324
rect 550100 562262 551692 562322
rect 550100 562260 550106 562262
rect 551686 562260 551692 562262
rect 551756 562260 551762 562324
rect 493961 560962 494027 560965
rect 548374 560962 548380 560964
rect 493961 560960 548380 560962
rect 493961 560904 493966 560960
rect 494022 560904 548380 560960
rect 493961 560902 548380 560904
rect 493961 560899 494027 560902
rect 548374 560900 548380 560902
rect 548444 560900 548450 560964
rect 551001 560284 551067 560285
rect 550766 560220 550772 560284
rect 550836 560220 550842 560284
rect 550950 560220 550956 560284
rect 551020 560282 551067 560284
rect 551020 560280 551112 560282
rect 551062 560224 551112 560280
rect 551020 560222 551112 560224
rect 551020 560220 551067 560222
rect 550774 560012 550834 560220
rect 551001 560219 551067 560220
rect 551134 560084 551140 560148
rect 551204 560146 551210 560148
rect 551502 560146 551508 560148
rect 551204 560086 551508 560146
rect 551204 560084 551210 560086
rect 551502 560084 551508 560086
rect 551572 560084 551578 560148
rect 550766 559948 550772 560012
rect 550836 559948 550842 560012
rect 29310 559540 29316 559604
rect 29380 559602 29386 559604
rect 100753 559602 100819 559605
rect 29380 559600 100819 559602
rect 29380 559544 100758 559600
rect 100814 559544 100819 559600
rect 29380 559542 100819 559544
rect 29380 559540 29386 559542
rect 100753 559539 100819 559542
rect 580165 557290 580231 557293
rect 583520 557290 584960 557380
rect 580165 557288 584960 557290
rect 580165 557232 580170 557288
rect 580226 557232 584960 557288
rect 580165 557230 584960 557232
rect 580165 557227 580231 557230
rect 583520 557140 584960 557230
rect 551001 555524 551067 555525
rect 550950 555522 550956 555524
rect 550910 555462 550956 555522
rect 551020 555520 551067 555524
rect 551062 555464 551067 555520
rect 550950 555460 550956 555462
rect 551020 555460 551067 555464
rect 551001 555459 551067 555460
rect 25446 554100 25452 554164
rect 25516 554162 25522 554164
rect 90541 554162 90607 554165
rect 25516 554160 90607 554162
rect 25516 554104 90546 554160
rect 90602 554104 90607 554160
rect 25516 554102 90607 554104
rect 25516 554100 25522 554102
rect 90541 554099 90607 554102
rect 25262 553964 25268 554028
rect 25332 554026 25338 554028
rect 90357 554026 90423 554029
rect 25332 554024 90423 554026
rect 25332 553968 90362 554024
rect 90418 553968 90423 554024
rect 25332 553966 90423 553968
rect 25332 553964 25338 553966
rect 90357 553963 90423 553966
rect 280153 553210 280219 553213
rect 280470 553210 280476 553212
rect 280153 553208 280476 553210
rect -960 553074 480 553164
rect 280153 553152 280158 553208
rect 280214 553152 280476 553208
rect 280153 553150 280476 553152
rect 280153 553147 280219 553150
rect 280470 553148 280476 553150
rect 280540 553148 280546 553212
rect 3141 553074 3207 553077
rect -960 553072 3207 553074
rect -960 553016 3146 553072
rect 3202 553016 3207 553072
rect -960 553014 3207 553016
rect -960 552924 480 553014
rect 3141 553011 3207 553014
rect 282913 550626 282979 550629
rect 283097 550626 283163 550629
rect 282913 550624 283163 550626
rect 282913 550568 282918 550624
rect 282974 550568 283102 550624
rect 283158 550568 283163 550624
rect 282913 550566 283163 550568
rect 282913 550563 282979 550566
rect 283097 550563 283163 550566
rect 550582 548524 550588 548588
rect 550652 548586 550658 548588
rect 551686 548586 551692 548588
rect 550652 548526 551692 548586
rect 550652 548524 550658 548526
rect 551686 548524 551692 548526
rect 551756 548524 551762 548588
rect 499481 545730 499547 545733
rect 552790 545730 552796 545732
rect 499481 545728 552796 545730
rect 499481 545672 499486 545728
rect 499542 545672 552796 545728
rect 499481 545670 552796 545672
rect 499481 545667 499547 545670
rect 552790 545668 552796 545670
rect 552860 545668 552866 545732
rect 580901 545594 580967 545597
rect 583520 545594 584960 545684
rect 580901 545592 584960 545594
rect 580901 545536 580906 545592
rect 580962 545536 584960 545592
rect 580901 545534 584960 545536
rect 580901 545531 580967 545534
rect 583520 545444 584960 545534
rect 551134 543764 551140 543828
rect 551204 543826 551210 543828
rect 551502 543826 551508 543828
rect 551204 543766 551508 543826
rect 551204 543764 551210 543766
rect 551502 543764 551508 543766
rect 551572 543764 551578 543828
rect 551134 543628 551140 543692
rect 551204 543690 551210 543692
rect 551686 543690 551692 543692
rect 551204 543630 551692 543690
rect 551204 543628 551210 543630
rect 551686 543628 551692 543630
rect 551756 543628 551762 543692
rect 280286 541180 280292 541244
rect 280356 541242 280362 541244
rect 280470 541242 280476 541244
rect 280356 541182 280476 541242
rect 280356 541180 280362 541182
rect 280470 541180 280476 541182
rect 280540 541180 280546 541244
rect 550582 538868 550588 538932
rect 550652 538930 550658 538932
rect 551502 538930 551508 538932
rect 550652 538870 551508 538930
rect 550652 538868 550658 538870
rect 551502 538868 551508 538870
rect 551572 538868 551578 538932
rect -960 538658 480 538748
rect 3509 538658 3575 538661
rect -960 538656 3575 538658
rect -960 538600 3514 538656
rect 3570 538600 3575 538656
rect -960 538598 3575 538600
rect -960 538508 480 538598
rect 3509 538595 3575 538598
rect 493777 534714 493843 534717
rect 549846 534714 549852 534716
rect 493777 534712 549852 534714
rect 493777 534656 493782 534712
rect 493838 534656 549852 534712
rect 493777 534654 549852 534656
rect 493777 534651 493843 534654
rect 549846 534652 549852 534654
rect 549916 534652 549922 534716
rect 280470 534306 280476 534308
rect 280294 534246 280476 534306
rect 280294 533900 280354 534246
rect 280470 534244 280476 534246
rect 280540 534244 280546 534308
rect 280286 533836 280292 533900
rect 280356 533836 280362 533900
rect 583520 533748 584960 533988
rect 25814 533564 25820 533628
rect 25884 533626 25890 533628
rect 80237 533626 80303 533629
rect 25884 533624 80303 533626
rect 25884 533568 80242 533624
rect 80298 533568 80303 533624
rect 25884 533566 80303 533568
rect 25884 533564 25890 533566
rect 80237 533563 80303 533566
rect 508221 533626 508287 533629
rect 552606 533626 552612 533628
rect 508221 533624 552612 533626
rect 508221 533568 508226 533624
rect 508282 533568 552612 533624
rect 508221 533566 552612 533568
rect 508221 533563 508287 533566
rect 552606 533564 552612 533566
rect 552676 533564 552682 533628
rect 25998 533428 26004 533492
rect 26068 533490 26074 533492
rect 82445 533490 82511 533493
rect 26068 533488 82511 533490
rect 26068 533432 82450 533488
rect 82506 533432 82511 533488
rect 26068 533430 82511 533432
rect 26068 533428 26074 533430
rect 82445 533427 82511 533430
rect 506105 533490 506171 533493
rect 552422 533490 552428 533492
rect 506105 533488 552428 533490
rect 506105 533432 506110 533488
rect 506166 533432 552428 533488
rect 506105 533430 552428 533432
rect 506105 533427 506171 533430
rect 552422 533428 552428 533430
rect 552492 533428 552498 533492
rect 28206 533292 28212 533356
rect 28276 533354 28282 533356
rect 97533 533354 97599 533357
rect 28276 533352 97599 533354
rect 28276 533296 97538 533352
rect 97594 533296 97599 533352
rect 28276 533294 97599 533296
rect 28276 533292 28282 533294
rect 97533 533291 97599 533294
rect 501781 533354 501847 533357
rect 552054 533354 552060 533356
rect 501781 533352 552060 533354
rect 501781 533296 501786 533352
rect 501842 533296 552060 533352
rect 501781 533294 552060 533296
rect 501781 533291 501847 533294
rect 552054 533292 552060 533294
rect 552124 533292 552130 533356
rect 175089 533218 175155 533221
rect 421373 533218 421439 533221
rect 175089 533216 421439 533218
rect 175089 533160 175094 533216
rect 175150 533160 421378 533216
rect 421434 533160 421439 533216
rect 175089 533158 421439 533160
rect 175089 533155 175155 533158
rect 421373 533155 421439 533158
rect 170765 533082 170831 533085
rect 425697 533082 425763 533085
rect 170765 533080 425763 533082
rect 170765 533024 170770 533080
rect 170826 533024 425702 533080
rect 425758 533024 425763 533080
rect 170765 533022 425763 533024
rect 170765 533019 170831 533022
rect 425697 533019 425763 533022
rect 166441 532946 166507 532949
rect 430021 532946 430087 532949
rect 166441 532944 430087 532946
rect 166441 532888 166446 532944
rect 166502 532888 430026 532944
rect 430082 532888 430087 532944
rect 166441 532886 430087 532888
rect 166441 532883 166507 532886
rect 430021 532883 430087 532886
rect 154665 532810 154731 532813
rect 441797 532810 441863 532813
rect 154665 532808 441863 532810
rect 154665 532752 154670 532808
rect 154726 532752 441802 532808
rect 441858 532752 441863 532808
rect 154665 532750 441863 532752
rect 154665 532747 154731 532750
rect 441797 532747 441863 532750
rect 25630 532612 25636 532676
rect 25700 532674 25706 532676
rect 73797 532674 73863 532677
rect 25700 532672 73863 532674
rect 25700 532616 73802 532672
rect 73858 532616 73863 532672
rect 25700 532614 73863 532616
rect 25700 532612 25706 532614
rect 73797 532611 73863 532614
rect 505001 532674 505067 532677
rect 552238 532674 552244 532676
rect 505001 532672 552244 532674
rect 505001 532616 505006 532672
rect 505062 532616 552244 532672
rect 505001 532614 552244 532616
rect 505001 532611 505067 532614
rect 552238 532612 552244 532614
rect 552308 532612 552314 532676
rect 28022 532476 28028 532540
rect 28092 532538 28098 532540
rect 96429 532538 96495 532541
rect 28092 532536 96495 532538
rect 28092 532480 96434 532536
rect 96490 532480 96495 532536
rect 28092 532478 96495 532480
rect 28092 532476 28098 532478
rect 96429 532475 96495 532478
rect 503621 532538 503687 532541
rect 550950 532538 550956 532540
rect 503621 532536 550956 532538
rect 503621 532480 503626 532536
rect 503682 532480 550956 532536
rect 503621 532478 550956 532480
rect 503621 532475 503687 532478
rect 550950 532476 550956 532478
rect 551020 532476 551026 532540
rect 27102 532340 27108 532404
rect 27172 532402 27178 532404
rect 98545 532402 98611 532405
rect 27172 532400 98611 532402
rect 27172 532344 98550 532400
rect 98606 532344 98611 532400
rect 27172 532342 98611 532344
rect 27172 532340 27178 532342
rect 98545 532339 98611 532342
rect 498561 532402 498627 532405
rect 553710 532402 553716 532404
rect 498561 532400 553716 532402
rect 498561 532344 498566 532400
rect 498622 532344 553716 532400
rect 498561 532342 553716 532344
rect 498561 532339 498627 532342
rect 553710 532340 553716 532342
rect 553780 532340 553786 532404
rect 27286 532204 27292 532268
rect 27356 532266 27362 532268
rect 100753 532266 100819 532269
rect 27356 532264 100819 532266
rect 27356 532208 100758 532264
rect 100814 532208 100819 532264
rect 27356 532206 100819 532208
rect 27356 532204 27362 532206
rect 100753 532203 100819 532206
rect 495341 532266 495407 532269
rect 551502 532266 551508 532268
rect 495341 532264 551508 532266
rect 495341 532208 495346 532264
rect 495402 532208 551508 532264
rect 495341 532206 551508 532208
rect 495341 532203 495407 532206
rect 551502 532204 551508 532206
rect 551572 532204 551578 532268
rect 27470 532068 27476 532132
rect 27540 532130 27546 532132
rect 102869 532130 102935 532133
rect 27540 532128 102935 532130
rect 27540 532072 102874 532128
rect 102930 532072 102935 532128
rect 27540 532070 102935 532072
rect 27540 532068 27546 532070
rect 102869 532067 102935 532070
rect 325049 532130 325115 532133
rect 441613 532130 441679 532133
rect 325049 532128 441679 532130
rect 325049 532072 325054 532128
rect 325110 532072 441618 532128
rect 441674 532072 441679 532128
rect 325049 532070 441679 532072
rect 325049 532067 325115 532070
rect 441613 532067 441679 532070
rect 497457 532130 497523 532133
rect 553526 532130 553532 532132
rect 497457 532128 553532 532130
rect 497457 532072 497462 532128
rect 497518 532072 553532 532128
rect 497457 532070 553532 532072
rect 497457 532067 497523 532070
rect 553526 532068 553532 532070
rect 553596 532068 553602 532132
rect 27654 531932 27660 531996
rect 27724 531994 27730 531996
rect 103973 531994 104039 531997
rect 27724 531992 104039 531994
rect 27724 531936 103978 531992
rect 104034 531936 104039 531992
rect 27724 531934 104039 531936
rect 27724 531932 27730 531934
rect 103973 531931 104039 531934
rect 188061 531994 188127 531997
rect 408585 531994 408651 531997
rect 188061 531992 408651 531994
rect 188061 531936 188066 531992
rect 188122 531936 408590 531992
rect 408646 531936 408651 531992
rect 188061 531934 408651 531936
rect 188061 531931 188127 531934
rect 408585 531931 408651 531934
rect 496353 531994 496419 531997
rect 553342 531994 553348 531996
rect 496353 531992 553348 531994
rect 496353 531936 496358 531992
rect 496414 531936 553348 531992
rect 496353 531934 553348 531936
rect 496353 531931 496419 531934
rect 553342 531932 553348 531934
rect 553412 531932 553418 531996
rect 162209 531858 162275 531861
rect 434253 531858 434319 531861
rect 162209 531856 434319 531858
rect 162209 531800 162214 531856
rect 162270 531800 434258 531856
rect 434314 531800 434319 531856
rect 162209 531798 434319 531800
rect 162209 531795 162275 531798
rect 434253 531795 434319 531798
rect 516869 531858 516935 531861
rect 551870 531858 551876 531860
rect 516869 531856 551876 531858
rect 516869 531800 516874 531856
rect 516930 531800 551876 531856
rect 516869 531798 551876 531800
rect 516869 531795 516935 531798
rect 551870 531796 551876 531798
rect 551940 531796 551946 531860
rect 155677 531722 155743 531725
rect 440785 531722 440851 531725
rect 155677 531720 440851 531722
rect 155677 531664 155682 531720
rect 155738 531664 440790 531720
rect 440846 531664 440851 531720
rect 155677 531662 440851 531664
rect 155677 531659 155743 531662
rect 440785 531659 440851 531662
rect 153561 531586 153627 531589
rect 442993 531586 443059 531589
rect 153561 531584 443059 531586
rect 153561 531528 153566 531584
rect 153622 531528 442998 531584
rect 443054 531528 443059 531584
rect 153561 531526 443059 531528
rect 153561 531523 153627 531526
rect 442993 531523 443059 531526
rect 141693 531450 141759 531453
rect 454769 531450 454835 531453
rect 141693 531448 454835 531450
rect 141693 531392 141698 531448
rect 141754 531392 454774 531448
rect 454830 531392 454835 531448
rect 141693 531390 454835 531392
rect 141693 531387 141759 531390
rect 454769 531387 454835 531390
rect 545941 531314 546007 531317
rect 546350 531314 546356 531316
rect 545941 531312 546356 531314
rect 545941 531256 545946 531312
rect 546002 531256 546356 531312
rect 545941 531254 546356 531256
rect 545941 531251 546007 531254
rect 546350 531252 546356 531254
rect 546420 531252 546426 531316
rect 492029 531178 492095 531181
rect 492438 531178 492444 531180
rect 492029 531176 492444 531178
rect 492029 531120 492034 531176
rect 492090 531120 492444 531176
rect 492029 531118 492444 531120
rect 492029 531115 492095 531118
rect 492438 531116 492444 531118
rect 492508 531116 492514 531180
rect 515765 531178 515831 531181
rect 551318 531178 551324 531180
rect 515765 531176 551324 531178
rect 515765 531120 515770 531176
rect 515826 531120 551324 531176
rect 515765 531118 551324 531120
rect 515765 531115 515831 531118
rect 551318 531116 551324 531118
rect 551388 531116 551394 531180
rect 507117 531042 507183 531045
rect 551686 531042 551692 531044
rect 507117 531040 551692 531042
rect 507117 530984 507122 531040
rect 507178 530984 551692 531040
rect 507117 530982 551692 530984
rect 507117 530979 507183 530982
rect 551686 530980 551692 530982
rect 551756 530980 551762 531044
rect 26734 530844 26740 530908
rect 26804 530906 26810 530908
rect 92105 530906 92171 530909
rect 26804 530904 92171 530906
rect 26804 530848 92110 530904
rect 92166 530848 92171 530904
rect 26804 530846 92171 530848
rect 26804 530844 26810 530846
rect 92105 530843 92171 530846
rect 509049 530906 509115 530909
rect 554078 530906 554084 530908
rect 509049 530904 554084 530906
rect 509049 530848 509054 530904
rect 509110 530848 554084 530904
rect 509049 530846 554084 530848
rect 509049 530843 509115 530846
rect 554078 530844 554084 530846
rect 554148 530844 554154 530908
rect 27838 530708 27844 530772
rect 27908 530770 27914 530772
rect 93209 530770 93275 530773
rect 27908 530768 93275 530770
rect 27908 530712 93214 530768
rect 93270 530712 93275 530768
rect 27908 530710 93275 530712
rect 27908 530708 27914 530710
rect 93209 530707 93275 530710
rect 500677 530770 500743 530773
rect 550766 530770 550772 530772
rect 500677 530768 550772 530770
rect 500677 530712 500682 530768
rect 500738 530712 550772 530768
rect 500677 530710 550772 530712
rect 500677 530707 500743 530710
rect 550766 530708 550772 530710
rect 550836 530708 550842 530772
rect 26918 530572 26924 530636
rect 26988 530634 26994 530636
rect 94221 530634 94287 530637
rect 26988 530632 94287 530634
rect 26988 530576 94226 530632
rect 94282 530576 94287 530632
rect 26988 530574 94287 530576
rect 26988 530572 26994 530574
rect 94221 530571 94287 530574
rect 502885 530634 502951 530637
rect 553894 530634 553900 530636
rect 502885 530632 553900 530634
rect 502885 530576 502890 530632
rect 502946 530576 553900 530632
rect 502885 530574 553900 530576
rect 502885 530571 502951 530574
rect 553894 530572 553900 530574
rect 553964 530572 553970 530636
rect 119061 530226 119127 530229
rect 477493 530226 477559 530229
rect 119061 530224 477559 530226
rect 119061 530168 119066 530224
rect 119122 530168 477498 530224
rect 477554 530168 477559 530224
rect 119061 530166 477559 530168
rect 119061 530163 119127 530166
rect 477493 530163 477559 530166
rect 115841 530090 115907 530093
rect 480621 530090 480687 530093
rect 115841 530088 480687 530090
rect 115841 530032 115846 530088
rect 115902 530032 480626 530088
rect 480682 530032 480687 530088
rect 115841 530030 480687 530032
rect 115841 530027 115907 530030
rect 480621 530027 480687 530030
rect 106089 529954 106155 529957
rect 490373 529954 490439 529957
rect 106089 529952 490439 529954
rect 106089 529896 106094 529952
rect 106150 529896 490378 529952
rect 490434 529896 490439 529952
rect 106089 529894 490439 529896
rect 106089 529891 106155 529894
rect 490373 529891 490439 529894
rect 107561 528594 107627 528597
rect 489269 528594 489335 528597
rect 107561 528592 489335 528594
rect 107561 528536 107566 528592
rect 107622 528536 489274 528592
rect 489330 528536 489335 528592
rect 107561 528534 489335 528536
rect 107561 528531 107627 528534
rect 489269 528531 489335 528534
rect 280286 528396 280292 528460
rect 280356 528458 280362 528460
rect 280521 528458 280587 528461
rect 280356 528456 280587 528458
rect 280356 528400 280526 528456
rect 280582 528400 280587 528456
rect 280356 528398 280587 528400
rect 280356 528396 280362 528398
rect 280521 528395 280587 528398
rect 115105 528322 115171 528325
rect 115933 528322 115999 528325
rect 471697 528322 471763 528325
rect 115105 528320 115999 528322
rect 115105 528264 115110 528320
rect 115166 528264 115938 528320
rect 115994 528264 115999 528320
rect 115105 528262 115999 528264
rect 115105 528259 115171 528262
rect 115933 528259 115999 528262
rect 471654 528320 471763 528322
rect 471654 528264 471702 528320
rect 471758 528264 471763 528320
rect 471654 528259 471763 528264
rect 125317 528220 125383 528223
rect 125317 528218 125426 528220
rect 125317 528162 125322 528218
rect 125378 528162 125426 528218
rect 125317 528157 125426 528162
rect 125366 527234 125426 528157
rect 260606 527854 267842 527914
rect 260606 527506 260666 527854
rect 267782 527642 267842 527854
rect 386462 527854 395906 527914
rect 267782 527582 269130 527642
rect 222334 527446 231594 527506
rect 144870 527310 147690 527370
rect 144870 527234 144930 527310
rect 125366 527174 144930 527234
rect 147630 527234 147690 527310
rect 154438 527310 157258 527370
rect 154438 527234 154498 527310
rect 147630 527174 154498 527234
rect 157198 527234 157258 527310
rect 186086 527310 191850 527370
rect 186086 527234 186146 527310
rect 157198 527174 186146 527234
rect 191790 527234 191850 527310
rect 210926 527310 215954 527370
rect 191790 527174 201602 527234
rect 201542 526962 201602 527174
rect 210926 526962 210986 527310
rect 215894 527234 215954 527310
rect 222334 527234 222394 527446
rect 215894 527174 222394 527234
rect 231534 527234 231594 527446
rect 239998 527446 241530 527506
rect 239998 527234 240058 527446
rect 231534 527174 240058 527234
rect 241470 527234 241530 527446
rect 251222 527446 260666 527506
rect 251222 527370 251282 527446
rect 251038 527310 251282 527370
rect 269070 527370 269130 527582
rect 296621 527506 296687 527509
rect 298093 527506 298159 527509
rect 296621 527504 298159 527506
rect 296621 527448 296626 527504
rect 296682 527448 298098 527504
rect 298154 527448 298159 527504
rect 296621 527446 298159 527448
rect 296621 527443 296687 527446
rect 298093 527443 298159 527446
rect 282821 527370 282887 527373
rect 269070 527368 282887 527370
rect 269070 527312 282826 527368
rect 282882 527312 282887 527368
rect 269070 527310 282887 527312
rect 251038 527234 251098 527310
rect 282821 527307 282887 527310
rect 326846 527310 331874 527370
rect 241470 527174 251098 527234
rect 283005 527234 283071 527237
rect 288525 527234 288591 527237
rect 283005 527232 288591 527234
rect 283005 527176 283010 527232
rect 283066 527176 288530 527232
rect 288586 527176 288591 527232
rect 283005 527174 288591 527176
rect 283005 527171 283071 527174
rect 288525 527171 288591 527174
rect 302969 527234 303035 527237
rect 317413 527234 317479 527237
rect 302969 527232 317479 527234
rect 302969 527176 302974 527232
rect 303030 527176 317418 527232
rect 317474 527176 317479 527232
rect 302969 527174 317479 527176
rect 302969 527171 303035 527174
rect 317413 527171 317479 527174
rect 201542 526902 210986 526962
rect 317413 526962 317479 526965
rect 326846 526962 326906 527310
rect 331814 527234 331874 527310
rect 340646 527310 350458 527370
rect 340646 527234 340706 527310
rect 331814 527174 340706 527234
rect 350398 527234 350458 527310
rect 362174 527310 365730 527370
rect 362174 527234 362234 527310
rect 350398 527174 362234 527234
rect 365670 527098 365730 527310
rect 375238 527310 381554 527370
rect 375238 527098 375298 527310
rect 381494 527234 381554 527310
rect 386462 527234 386522 527854
rect 381494 527174 386522 527234
rect 395846 527234 395906 527854
rect 423814 527718 427922 527778
rect 423814 527642 423874 527718
rect 408542 527582 414122 527642
rect 396214 527446 398850 527506
rect 396214 527234 396274 527446
rect 395846 527174 396274 527234
rect 398790 527234 398850 527446
rect 408542 527370 408602 527582
rect 404310 527310 408602 527370
rect 414062 527370 414122 527582
rect 418294 527582 423874 527642
rect 427862 527642 427922 527718
rect 442950 527718 452578 527778
rect 427862 527582 437306 527642
rect 418294 527370 418354 527582
rect 437246 527506 437306 527582
rect 442950 527506 443010 527718
rect 437246 527446 443010 527506
rect 452518 527506 452578 527718
rect 452518 527446 454234 527506
rect 414062 527310 418354 527370
rect 454174 527370 454234 527446
rect 454174 527310 454418 527370
rect 404310 527234 404370 527310
rect 398790 527174 404370 527234
rect 454358 527234 454418 527310
rect 471654 527234 471714 528259
rect 454358 527174 471714 527234
rect 365670 527038 375298 527098
rect 317413 526960 326906 526962
rect 317413 526904 317418 526960
rect 317474 526904 326906 526960
rect 317413 526902 326906 526904
rect 317413 526899 317479 526902
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 280521 518940 280587 518941
rect 280470 518876 280476 518940
rect 280540 518938 280587 518940
rect 282913 518938 282979 518941
rect 283189 518938 283255 518941
rect 280540 518936 280632 518938
rect 280582 518880 280632 518936
rect 280540 518878 280632 518880
rect 282913 518936 283255 518938
rect 282913 518880 282918 518936
rect 282974 518880 283194 518936
rect 283250 518880 283255 518936
rect 282913 518878 283255 518880
rect 280540 518876 280587 518878
rect 280521 518875 280587 518876
rect 282913 518875 282979 518878
rect 283189 518875 283255 518878
rect 281533 515946 281599 515949
rect 279036 515944 281599 515946
rect 279036 515888 281538 515944
rect 281594 515888 281599 515944
rect 279036 515886 281599 515888
rect 281533 515883 281599 515886
rect 314653 515810 314719 515813
rect 315941 515810 316007 515813
rect 314653 515808 317676 515810
rect 314653 515752 314658 515808
rect 314714 515752 315946 515808
rect 316002 515752 317676 515808
rect 314653 515750 317676 515752
rect 314653 515747 314719 515750
rect 315941 515747 316007 515750
rect 579613 510370 579679 510373
rect 583520 510370 584960 510460
rect 579613 510368 584960 510370
rect 579613 510312 579618 510368
rect 579674 510312 584960 510368
rect 579613 510310 584960 510312
rect 579613 510307 579679 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 2865 509962 2931 509965
rect -960 509960 2931 509962
rect -960 509904 2870 509960
rect 2926 509904 2931 509960
rect -960 509902 2931 509904
rect -960 509812 480 509902
rect 2865 509899 2931 509902
rect 280470 509282 280476 509284
rect 280294 509222 280476 509282
rect 280294 509146 280354 509222
rect 280470 509220 280476 509222
rect 280540 509220 280546 509284
rect 280470 509146 280476 509148
rect 280294 509086 280476 509146
rect 280470 509084 280476 509086
rect 280540 509084 280546 509148
rect 146894 500926 147322 500986
rect 118693 500852 118759 500853
rect 118693 500850 118740 500852
rect 118648 500848 118740 500850
rect 118648 500792 118698 500848
rect 118648 500790 118740 500792
rect 118693 500788 118740 500790
rect 118804 500788 118810 500852
rect 120073 500850 120139 500853
rect 132585 500850 132651 500853
rect 120073 500848 132651 500850
rect 120073 500792 120078 500848
rect 120134 500792 132590 500848
rect 132646 500792 132651 500848
rect 120073 500790 132651 500792
rect 118693 500787 118759 500788
rect 120073 500787 120139 500790
rect 132585 500787 132651 500790
rect 142061 500850 142127 500853
rect 144637 500850 144703 500853
rect 146894 500850 146954 500926
rect 142061 500848 144703 500850
rect 142061 500792 142066 500848
rect 142122 500792 144642 500848
rect 144698 500792 144703 500848
rect 142061 500790 144703 500792
rect 142061 500787 142127 500790
rect 144637 500787 144703 500790
rect 144870 500790 146954 500850
rect 147029 500852 147095 500853
rect 147029 500848 147076 500852
rect 147140 500850 147146 500852
rect 147262 500850 147322 500926
rect 148133 500852 148199 500853
rect 147806 500850 147812 500852
rect 147029 500792 147034 500848
rect 115933 500714 115999 500717
rect 144870 500714 144930 500790
rect 147029 500788 147076 500792
rect 147140 500790 147186 500850
rect 147262 500790 147812 500850
rect 147140 500788 147146 500790
rect 147806 500788 147812 500790
rect 147876 500788 147882 500852
rect 148133 500848 148180 500852
rect 148244 500850 148250 500852
rect 149237 500850 149303 500853
rect 149646 500850 149652 500852
rect 148133 500792 148138 500848
rect 148133 500788 148180 500792
rect 148244 500790 148290 500850
rect 149237 500848 149652 500850
rect 149237 500792 149242 500848
rect 149298 500792 149652 500848
rect 149237 500790 149652 500792
rect 148244 500788 148250 500790
rect 147029 500787 147095 500788
rect 148133 500787 148199 500788
rect 149237 500787 149303 500790
rect 149646 500788 149652 500790
rect 149716 500788 149722 500852
rect 149830 500788 149836 500852
rect 149900 500850 149906 500852
rect 150341 500850 150407 500853
rect 149900 500848 150407 500850
rect 149900 500792 150346 500848
rect 150402 500792 150407 500848
rect 149900 500790 150407 500792
rect 149900 500788 149906 500790
rect 150341 500787 150407 500790
rect 150934 500788 150940 500852
rect 151004 500850 151010 500852
rect 151353 500850 151419 500853
rect 152457 500852 152523 500853
rect 152406 500850 152412 500852
rect 151004 500848 151419 500850
rect 151004 500792 151358 500848
rect 151414 500792 151419 500848
rect 151004 500790 151419 500792
rect 151004 500788 151010 500790
rect 151353 500787 151419 500790
rect 151494 500790 152290 500850
rect 152366 500790 152412 500850
rect 152476 500848 152523 500852
rect 152518 500792 152523 500848
rect 115933 500712 144930 500714
rect 115933 500656 115938 500712
rect 115994 500656 144930 500712
rect 115933 500654 144930 500656
rect 146017 500714 146083 500717
rect 151494 500714 151554 500790
rect 146017 500712 151554 500714
rect 146017 500656 146022 500712
rect 146078 500656 151554 500712
rect 146017 500654 151554 500656
rect 115933 500651 115999 500654
rect 146017 500651 146083 500654
rect 114737 500578 114803 500581
rect 148358 500578 148364 500580
rect 114737 500576 148364 500578
rect 114737 500520 114742 500576
rect 114798 500520 148364 500576
rect 114737 500518 148364 500520
rect 114737 500515 114803 500518
rect 148358 500516 148364 500518
rect 148428 500516 148434 500580
rect 152230 500578 152290 500790
rect 152406 500788 152412 500790
rect 152476 500788 152523 500792
rect 153142 500788 153148 500852
rect 153212 500850 153218 500852
rect 153377 500850 153443 500853
rect 153212 500848 153443 500850
rect 153212 500792 153382 500848
rect 153438 500792 153443 500848
rect 153212 500790 153443 500792
rect 153212 500788 153218 500790
rect 152457 500787 152523 500788
rect 153377 500787 153443 500790
rect 189574 500788 189580 500852
rect 189644 500850 189650 500852
rect 190177 500850 190243 500853
rect 189644 500848 190243 500850
rect 189644 500792 190182 500848
rect 190238 500792 190243 500848
rect 189644 500790 190243 500792
rect 189644 500788 189650 500790
rect 190177 500787 190243 500790
rect 191046 500788 191052 500852
rect 191116 500850 191122 500852
rect 191281 500850 191347 500853
rect 191116 500848 191347 500850
rect 191116 500792 191286 500848
rect 191342 500792 191347 500848
rect 191116 500790 191347 500792
rect 191116 500788 191122 500790
rect 191281 500787 191347 500790
rect 189073 500714 189139 500717
rect 189758 500714 189764 500716
rect 189073 500712 189764 500714
rect 189073 500656 189078 500712
rect 189134 500656 189764 500712
rect 189073 500654 189764 500656
rect 189073 500651 189139 500654
rect 189758 500652 189764 500654
rect 189828 500652 189834 500716
rect 512545 500714 512611 500717
rect 548374 500714 548380 500716
rect 512545 500712 548380 500714
rect 512545 500656 512550 500712
rect 512606 500656 548380 500712
rect 512545 500654 548380 500656
rect 512545 500651 512611 500654
rect 548374 500652 548380 500654
rect 548444 500652 548450 500716
rect 153326 500578 153332 500580
rect 152230 500518 153332 500578
rect 153326 500516 153332 500518
rect 153396 500516 153402 500580
rect 153469 500578 153535 500581
rect 153878 500578 153884 500580
rect 153469 500576 153884 500578
rect 153469 500520 153474 500576
rect 153530 500520 153884 500576
rect 153469 500518 153884 500520
rect 153469 500515 153535 500518
rect 153878 500516 153884 500518
rect 153948 500516 153954 500580
rect 514661 500578 514727 500581
rect 549846 500578 549852 500580
rect 514661 500576 549852 500578
rect 514661 500520 514666 500576
rect 514722 500520 549852 500576
rect 514661 500518 549852 500520
rect 514661 500515 514727 500518
rect 549846 500516 549852 500518
rect 549916 500516 549922 500580
rect 113173 500442 113239 500445
rect 147990 500442 147996 500444
rect 113173 500440 147996 500442
rect 113173 500384 113178 500440
rect 113234 500384 147996 500440
rect 113173 500382 147996 500384
rect 113173 500379 113239 500382
rect 147990 500380 147996 500382
rect 148060 500380 148066 500444
rect 508221 500442 508287 500445
rect 546534 500442 546540 500444
rect 508221 500440 546540 500442
rect 508221 500384 508226 500440
rect 508282 500384 546540 500440
rect 508221 500382 546540 500384
rect 508221 500379 508287 500382
rect 546534 500380 546540 500382
rect 546604 500380 546610 500444
rect 112621 500306 112687 500309
rect 147254 500306 147260 500308
rect 112621 500304 147260 500306
rect 112621 500248 112626 500304
rect 112682 500248 147260 500304
rect 112621 500246 147260 500248
rect 112621 500243 112687 500246
rect 147254 500244 147260 500246
rect 147324 500244 147330 500308
rect 500677 500306 500743 500309
rect 550582 500306 550588 500308
rect 500677 500304 550588 500306
rect 500677 500248 500682 500304
rect 500738 500248 550588 500304
rect 500677 500246 550588 500248
rect 500677 500243 500743 500246
rect 550582 500244 550588 500246
rect 550652 500244 550658 500308
rect 114553 500170 114619 500173
rect 114686 500170 114692 500172
rect 114553 500168 114692 500170
rect 114553 500112 114558 500168
rect 114614 500112 114692 500168
rect 114553 500110 114692 500112
rect 114553 500107 114619 500110
rect 114686 500108 114692 500110
rect 114756 500108 114762 500172
rect 147622 500170 147628 500172
rect 114878 500110 147628 500170
rect 107193 500034 107259 500037
rect 114878 500034 114938 500110
rect 147622 500108 147628 500110
rect 147692 500108 147698 500172
rect 188838 500108 188844 500172
rect 188908 500170 188914 500172
rect 194501 500170 194567 500173
rect 188908 500168 194567 500170
rect 188908 500112 194506 500168
rect 194562 500112 194567 500168
rect 188908 500110 194567 500112
rect 188908 500108 188914 500110
rect 194501 500107 194567 500110
rect 497457 500170 497523 500173
rect 550766 500170 550772 500172
rect 497457 500168 550772 500170
rect 497457 500112 497462 500168
rect 497518 500112 550772 500168
rect 497457 500110 550772 500112
rect 497457 500107 497523 500110
rect 550766 500108 550772 500110
rect 550836 500108 550842 500172
rect 107193 500032 114938 500034
rect 107193 499976 107198 500032
rect 107254 499976 114938 500032
rect 107193 499974 114938 499976
rect 134149 500034 134215 500037
rect 150566 500034 150572 500036
rect 134149 500032 150572 500034
rect 134149 499976 134154 500032
rect 134210 499976 150572 500032
rect 134149 499974 150572 499976
rect 107193 499971 107259 499974
rect 134149 499971 134215 499974
rect 150566 499972 150572 499974
rect 150636 499972 150642 500036
rect 136265 499898 136331 499901
rect 150750 499898 150756 499900
rect 136265 499896 150756 499898
rect 136265 499840 136270 499896
rect 136326 499840 150756 499896
rect 136265 499838 150756 499840
rect 136265 499835 136331 499838
rect 150750 499836 150756 499838
rect 150820 499836 150826 499900
rect 138473 499762 138539 499765
rect 149278 499762 149284 499764
rect 138473 499760 149284 499762
rect 138473 499704 138478 499760
rect 138534 499704 149284 499760
rect 138473 499702 149284 499704
rect 138473 499699 138539 499702
rect 149278 499700 149284 499702
rect 149348 499700 149354 499764
rect 132585 499626 132651 499629
rect 142061 499626 142127 499629
rect 132585 499624 142127 499626
rect 132585 499568 132590 499624
rect 132646 499568 142066 499624
rect 142122 499568 142127 499624
rect 132585 499566 142127 499568
rect 132585 499563 132651 499566
rect 142061 499563 142127 499566
rect 144637 499626 144703 499629
rect 151118 499626 151124 499628
rect 144637 499624 151124 499626
rect 144637 499568 144642 499624
rect 144698 499568 151124 499624
rect 144637 499566 151124 499568
rect 144637 499563 144703 499566
rect 151118 499564 151124 499566
rect 151188 499564 151194 499628
rect 580901 498674 580967 498677
rect 583520 498674 584960 498764
rect 580901 498672 584960 498674
rect 580901 498616 580906 498672
rect 580962 498616 584960 498672
rect 580901 498614 584960 498616
rect 580901 498611 580967 498614
rect 583520 498524 584960 498614
rect 110413 497994 110479 497997
rect 150014 497994 150020 497996
rect 110413 497992 150020 497994
rect 110413 497936 110418 497992
rect 110474 497936 150020 497992
rect 110413 497934 150020 497936
rect 110413 497931 110479 497934
rect 150014 497932 150020 497934
rect 150084 497932 150090 497996
rect 110597 497858 110663 497861
rect 151302 497858 151308 497860
rect 110597 497856 151308 497858
rect 110597 497800 110602 497856
rect 110658 497800 151308 497856
rect 110597 497798 151308 497800
rect 110597 497795 110663 497798
rect 151302 497796 151308 497798
rect 151372 497796 151378 497860
rect 109033 497722 109099 497725
rect 150382 497722 150388 497724
rect 109033 497720 150388 497722
rect 109033 497664 109038 497720
rect 109094 497664 150388 497720
rect 109033 497662 150388 497664
rect 109033 497659 109099 497662
rect 150382 497660 150388 497662
rect 150452 497660 150458 497724
rect 107653 497586 107719 497589
rect 149094 497586 149100 497588
rect 107653 497584 149100 497586
rect 107653 497528 107658 497584
rect 107714 497528 149100 497584
rect 107653 497526 149100 497528
rect 107653 497523 107719 497526
rect 149094 497524 149100 497526
rect 149164 497524 149170 497588
rect 104893 497450 104959 497453
rect 147438 497450 147444 497452
rect 104893 497448 147444 497450
rect 104893 497392 104898 497448
rect 104954 497392 147444 497448
rect 104893 497390 147444 497392
rect 104893 497387 104959 497390
rect 147438 497388 147444 497390
rect 147508 497388 147514 497452
rect -960 495546 480 495636
rect 3509 495546 3575 495549
rect 280337 495548 280403 495549
rect 280286 495546 280292 495548
rect -960 495544 3575 495546
rect -960 495488 3514 495544
rect 3570 495488 3575 495544
rect -960 495486 3575 495488
rect 280246 495486 280292 495546
rect 280356 495544 280403 495548
rect 280398 495488 280403 495544
rect -960 495396 480 495486
rect 3509 495483 3575 495486
rect 280286 495484 280292 495486
rect 280356 495484 280403 495488
rect 280337 495483 280403 495484
rect 20478 492492 20484 492556
rect 20548 492554 20554 492556
rect 21357 492554 21423 492557
rect 20548 492552 21423 492554
rect 20548 492496 21362 492552
rect 21418 492496 21423 492552
rect 20548 492494 21423 492496
rect 20548 492492 20554 492494
rect 21357 492491 21423 492494
rect 280337 489970 280403 489973
rect 280654 489970 280660 489972
rect 280337 489968 280660 489970
rect 280337 489912 280342 489968
rect 280398 489912 280660 489968
rect 280337 489910 280660 489912
rect 280337 489907 280403 489910
rect 280654 489908 280660 489910
rect 280724 489908 280730 489972
rect 106181 489154 106247 489157
rect 153009 489154 153075 489157
rect 106181 489152 153075 489154
rect 106181 489096 106186 489152
rect 106242 489096 153014 489152
rect 153070 489096 153075 489152
rect 106181 489094 153075 489096
rect 106181 489091 106247 489094
rect 153009 489091 153075 489094
rect 583520 486692 584960 486932
rect 151905 486570 151971 486573
rect 152774 486570 152780 486572
rect 151905 486568 152780 486570
rect 151905 486512 151910 486568
rect 151966 486512 152780 486568
rect 151905 486510 152780 486512
rect 151905 486507 151971 486510
rect 152774 486508 152780 486510
rect 152844 486508 152850 486572
rect 151997 486436 152063 486437
rect 151997 486434 152044 486436
rect 151952 486432 152044 486434
rect 151952 486376 152002 486432
rect 151952 486374 152044 486376
rect 151997 486372 152044 486374
rect 152108 486372 152114 486436
rect 151997 486371 152063 486372
rect 20294 485012 20300 485076
rect 20364 485074 20370 485076
rect 21214 485074 21220 485076
rect 20364 485014 21220 485074
rect 20364 485012 20370 485014
rect 21214 485012 21220 485014
rect 21284 485012 21290 485076
rect 282913 483034 282979 483037
rect 283097 483034 283163 483037
rect 282913 483032 283163 483034
rect 282913 482976 282918 483032
rect 282974 482976 283102 483032
rect 283158 482976 283163 483032
rect 282913 482974 283163 482976
rect 282913 482971 282979 482974
rect 283097 482971 283163 482974
rect 320541 483034 320607 483037
rect 320725 483034 320791 483037
rect 320541 483032 320791 483034
rect 320541 482976 320546 483032
rect 320602 482976 320730 483032
rect 320786 482976 320791 483032
rect 320541 482974 320791 482976
rect 320541 482971 320607 482974
rect 320725 482971 320791 482974
rect -960 481130 480 481220
rect 3141 481130 3207 481133
rect -960 481128 3207 481130
rect -960 481072 3146 481128
rect 3202 481072 3207 481128
rect -960 481070 3207 481072
rect -960 480980 480 481070
rect 3141 481067 3207 481070
rect 280102 480252 280108 480316
rect 280172 480314 280178 480316
rect 280654 480314 280660 480316
rect 280172 480254 280660 480314
rect 280172 480252 280178 480254
rect 280654 480252 280660 480254
rect 280724 480252 280730 480316
rect 280153 480044 280219 480045
rect 280102 480042 280108 480044
rect 280062 479982 280108 480042
rect 280172 480040 280219 480044
rect 280214 479984 280219 480040
rect 280102 479980 280108 479982
rect 280172 479980 280219 479984
rect 280153 479979 280219 479980
rect 507761 475554 507827 475557
rect 553342 475554 553348 475556
rect 507761 475552 553348 475554
rect 507761 475496 507766 475552
rect 507822 475496 553348 475552
rect 507761 475494 553348 475496
rect 507761 475491 507827 475494
rect 553342 475492 553348 475494
rect 553412 475492 553418 475556
rect 493961 475418 494027 475421
rect 552054 475418 552060 475420
rect 493961 475416 552060 475418
rect 493961 475360 493966 475416
rect 494022 475360 552060 475416
rect 493961 475358 552060 475360
rect 493961 475355 494027 475358
rect 552054 475356 552060 475358
rect 552124 475356 552130 475420
rect 583520 474996 584960 475236
rect 551921 473922 551987 473925
rect 551921 473920 552122 473922
rect 551921 473864 551926 473920
rect 551982 473864 552122 473920
rect 551921 473862 552122 473864
rect 551921 473859 551987 473862
rect 546585 473516 546651 473517
rect 546534 473514 546540 473516
rect 546494 473454 546540 473514
rect 546604 473512 546651 473516
rect 546646 473456 546651 473512
rect 546534 473452 546540 473454
rect 546604 473452 546651 473456
rect 546585 473451 546651 473452
rect 552062 473348 552122 473862
rect 552105 473106 552171 473109
rect 552062 473104 552171 473106
rect 552062 473048 552110 473104
rect 552166 473048 552171 473104
rect 552062 473043 552171 473048
rect 552062 472804 552122 473043
rect 554773 472154 554839 472157
rect 552644 472152 554839 472154
rect 552644 472096 554778 472152
rect 554834 472096 554839 472152
rect 552644 472094 554839 472096
rect 554773 472091 554839 472094
rect 279601 471882 279667 471885
rect 279558 471880 279667 471882
rect 279558 471824 279606 471880
rect 279662 471824 279667 471880
rect 279558 471819 279667 471824
rect 552054 471820 552060 471884
rect 552124 471820 552130 471884
rect 279558 471308 279618 471819
rect 552062 471580 552122 471820
rect 552289 471338 552355 471341
rect 552565 471338 552631 471341
rect 552289 471336 552631 471338
rect 552289 471280 552294 471336
rect 552350 471280 552570 471336
rect 552626 471280 552631 471336
rect 552289 471278 552631 471280
rect 552289 471275 552355 471278
rect 552565 471275 552631 471278
rect 555693 471066 555759 471069
rect 552644 471064 555759 471066
rect 552644 471008 555698 471064
rect 555754 471008 555759 471064
rect 552644 471006 555759 471008
rect 555693 471003 555759 471006
rect 280153 470658 280219 470661
rect 280286 470658 280292 470660
rect 280153 470656 280292 470658
rect 280153 470600 280158 470656
rect 280214 470600 280292 470656
rect 280153 470598 280292 470600
rect 280153 470595 280219 470598
rect 280286 470596 280292 470598
rect 280356 470596 280362 470660
rect 555877 470386 555943 470389
rect 552644 470384 555943 470386
rect 552644 470328 555882 470384
rect 555938 470328 555943 470384
rect 552644 470326 555943 470328
rect 555877 470323 555943 470326
rect 552054 470052 552060 470116
rect 552124 470052 552130 470116
rect 552062 469812 552122 470052
rect 555969 469298 556035 469301
rect 552644 469296 556035 469298
rect 552644 469240 555974 469296
rect 556030 469240 556035 469296
rect 552644 469238 556035 469240
rect 555969 469235 556035 469238
rect 552933 468618 552999 468621
rect 552644 468616 552999 468618
rect 552644 468560 552938 468616
rect 552994 468560 552999 468616
rect 552644 468558 552999 468560
rect 552933 468555 552999 468558
rect 552054 468284 552060 468348
rect 552124 468284 552130 468348
rect 552062 468044 552122 468284
rect 554957 467530 555023 467533
rect 552644 467528 555023 467530
rect 552644 467472 554962 467528
rect 555018 467472 555023 467528
rect 552644 467470 555023 467472
rect 554957 467467 555023 467470
rect 552105 467258 552171 467261
rect 552062 467256 552171 467258
rect 552062 467200 552110 467256
rect 552166 467200 552171 467256
rect 552062 467195 552171 467200
rect -960 466700 480 466940
rect 552062 466820 552122 467195
rect 553209 466306 553275 466309
rect 552644 466304 553275 466306
rect 552644 466248 553214 466304
rect 553270 466248 553275 466304
rect 552644 466246 553275 466248
rect 553209 466243 553275 466246
rect 555233 465626 555299 465629
rect 552644 465624 555299 465626
rect 552644 465568 555238 465624
rect 555294 465568 555299 465624
rect 552644 465566 555299 465568
rect 555233 465563 555299 465566
rect 156045 465354 156111 465357
rect 153916 465352 156111 465354
rect 153916 465296 156050 465352
rect 156106 465296 156111 465352
rect 153916 465294 156111 465296
rect 156045 465291 156111 465294
rect 556061 465082 556127 465085
rect 552644 465080 556127 465082
rect 552644 465024 556066 465080
rect 556122 465024 556127 465080
rect 552644 465022 556127 465024
rect 556061 465019 556127 465022
rect 553342 464538 553348 464540
rect 552644 464478 553348 464538
rect 553342 464476 553348 464478
rect 553412 464476 553418 464540
rect 554773 463858 554839 463861
rect 552644 463856 554839 463858
rect 552644 463800 554778 463856
rect 554834 463800 554839 463856
rect 552644 463798 554839 463800
rect 554773 463795 554839 463798
rect 280286 463660 280292 463724
rect 280356 463722 280362 463724
rect 280654 463722 280660 463724
rect 280356 463662 280660 463722
rect 280356 463660 280362 463662
rect 280654 463660 280660 463662
rect 280724 463660 280730 463724
rect 553025 463586 553091 463589
rect 552614 463584 553091 463586
rect 552614 463528 553030 463584
rect 553086 463528 553091 463584
rect 552614 463526 553091 463528
rect 552614 463284 552674 463526
rect 553025 463523 553091 463526
rect 580165 463450 580231 463453
rect 583520 463450 584960 463540
rect 580165 463448 584960 463450
rect 580165 463392 580170 463448
rect 580226 463392 584960 463448
rect 580165 463390 584960 463392
rect 580165 463387 580231 463390
rect 583520 463300 584960 463390
rect 313273 462770 313339 462773
rect 553301 462770 553367 462773
rect 313273 462768 316020 462770
rect 313273 462712 313278 462768
rect 313334 462712 316020 462768
rect 313273 462710 316020 462712
rect 552644 462768 553367 462770
rect 552644 462712 553306 462768
rect 553362 462712 553367 462768
rect 552644 462710 553367 462712
rect 313273 462707 313339 462710
rect 553301 462707 553367 462710
rect 555141 462090 555207 462093
rect 552644 462088 555207 462090
rect 552644 462032 555146 462088
rect 555202 462032 555207 462088
rect 552644 462030 555207 462032
rect 555141 462027 555207 462030
rect 555182 461546 555188 461548
rect 552644 461486 555188 461546
rect 555182 461484 555188 461486
rect 555252 461484 555258 461548
rect 552841 461002 552907 461005
rect 552644 461000 552907 461002
rect 552644 460944 552846 461000
rect 552902 460944 552907 461000
rect 552644 460942 552907 460944
rect 552841 460939 552907 460942
rect 554814 460322 554820 460324
rect 552644 460262 554820 460322
rect 554814 460260 554820 460262
rect 554884 460260 554890 460324
rect 553025 459778 553091 459781
rect 552644 459776 553091 459778
rect 552644 459720 553030 459776
rect 553086 459720 553091 459776
rect 552644 459718 553091 459720
rect 553025 459715 553091 459718
rect 553117 459234 553183 459237
rect 552644 459232 553183 459234
rect 552644 459176 553122 459232
rect 553178 459176 553183 459232
rect 552644 459174 553183 459176
rect 553117 459171 553183 459174
rect 552105 458962 552171 458965
rect 552062 458960 552171 458962
rect 552062 458904 552110 458960
rect 552166 458904 552171 458960
rect 552062 458899 552171 458904
rect 552062 458524 552122 458899
rect 555417 458010 555483 458013
rect 552644 458008 555483 458010
rect 552644 457952 555422 458008
rect 555478 457952 555483 458008
rect 552644 457950 555483 457952
rect 555417 457947 555483 457950
rect 554589 457330 554655 457333
rect 552644 457328 554655 457330
rect 552644 457272 554594 457328
rect 554650 457272 554655 457328
rect 552644 457270 554655 457272
rect 554589 457267 554655 457270
rect 552841 456786 552907 456789
rect 552644 456784 552907 456786
rect 552644 456728 552846 456784
rect 552902 456728 552907 456784
rect 552644 456726 552907 456728
rect 552841 456723 552907 456726
rect 552105 456514 552171 456517
rect 552062 456512 552171 456514
rect 552062 456456 552110 456512
rect 552166 456456 552171 456512
rect 552062 456451 552171 456456
rect 552062 456212 552122 456451
rect 555325 455562 555391 455565
rect 552644 455560 555391 455562
rect 552644 455504 555330 455560
rect 555386 455504 555391 455560
rect 552644 455502 555391 455504
rect 555325 455499 555391 455502
rect 552105 455290 552171 455293
rect 552062 455288 552171 455290
rect 552062 455232 552110 455288
rect 552166 455232 552171 455288
rect 552062 455227 552171 455232
rect 552062 454988 552122 455227
rect 553209 454474 553275 454477
rect 552644 454472 553275 454474
rect 552644 454416 553214 454472
rect 553270 454416 553275 454472
rect 552644 454414 553275 454416
rect 553209 454411 553275 454414
rect 554497 453794 554563 453797
rect 552644 453792 554563 453794
rect 552644 453736 554502 453792
rect 554558 453736 554563 453792
rect 552644 453734 554563 453736
rect 554497 453731 554563 453734
rect 552381 453522 552447 453525
rect 552381 453520 552490 453522
rect 552381 453464 552386 453520
rect 552442 453464 552490 453520
rect 552381 453459 552490 453464
rect 552430 453220 552490 453459
rect 552749 452978 552815 452981
rect 552614 452976 552815 452978
rect 552614 452920 552754 452976
rect 552810 452920 552815 452976
rect 552614 452918 552815 452920
rect 552614 452676 552674 452918
rect 552749 452915 552815 452918
rect -960 452434 480 452524
rect 3417 452434 3483 452437
rect -960 452432 3483 452434
rect -960 452376 3422 452432
rect 3478 452376 3483 452432
rect -960 452374 3483 452376
rect -960 452284 480 452374
rect 3417 452371 3483 452374
rect 555785 452026 555851 452029
rect 552644 452024 555851 452026
rect 552644 451968 555790 452024
rect 555846 451968 555851 452024
rect 552644 451966 555851 451968
rect 555785 451963 555851 451966
rect 580901 451754 580967 451757
rect 583520 451754 584960 451844
rect 580901 451752 584960 451754
rect 580901 451696 580906 451752
rect 580962 451696 584960 451752
rect 580901 451694 584960 451696
rect 580901 451691 580967 451694
rect 583520 451604 584960 451694
rect 554405 451482 554471 451485
rect 552644 451480 554471 451482
rect 552644 451424 554410 451480
rect 554466 451424 554471 451480
rect 552644 451422 554471 451424
rect 554405 451419 554471 451422
rect 280245 451212 280311 451213
rect 280245 451210 280292 451212
rect 280200 451208 280292 451210
rect 280200 451152 280250 451208
rect 280200 451150 280292 451152
rect 280245 451148 280292 451150
rect 280356 451148 280362 451212
rect 552565 451210 552631 451213
rect 552565 451208 552674 451210
rect 552565 451152 552570 451208
rect 552626 451152 552674 451208
rect 280245 451147 280311 451148
rect 552565 451147 552674 451152
rect 185577 450938 185643 450941
rect 185577 450936 188140 450938
rect 185577 450880 185582 450936
rect 185638 450880 188140 450936
rect 552614 450908 552674 451147
rect 185577 450878 188140 450880
rect 185577 450875 185643 450878
rect 443637 450666 443703 450669
rect 552473 450666 552539 450669
rect 443637 450664 446108 450666
rect 443637 450608 443642 450664
rect 443698 450608 446108 450664
rect 443637 450606 446108 450608
rect 552430 450664 552539 450666
rect 552430 450608 552478 450664
rect 552534 450608 552539 450664
rect 443637 450603 443703 450606
rect 552430 450603 552539 450608
rect 552430 450228 552490 450603
rect 555693 449714 555759 449717
rect 552644 449712 555759 449714
rect 552644 449656 555698 449712
rect 555754 449656 555759 449712
rect 552644 449654 555759 449656
rect 555693 449651 555759 449654
rect 554313 449034 554379 449037
rect 552644 449032 554379 449034
rect 552644 448976 554318 449032
rect 554374 448976 554379 449032
rect 552644 448974 554379 448976
rect 554313 448971 554379 448974
rect 552289 448762 552355 448765
rect 552246 448760 552355 448762
rect 552246 448704 552294 448760
rect 552350 448704 552355 448760
rect 552246 448699 552355 448704
rect 552246 448460 552306 448699
rect 552197 448218 552263 448221
rect 552197 448216 552306 448218
rect 552197 448160 552202 448216
rect 552258 448160 552306 448216
rect 552197 448155 552306 448160
rect 552246 447916 552306 448155
rect 555049 447266 555115 447269
rect 552644 447264 555115 447266
rect 552644 447208 555054 447264
rect 555110 447208 555115 447264
rect 552644 447206 555115 447208
rect 555049 447203 555115 447206
rect 553945 446722 554011 446725
rect 552644 446720 554011 446722
rect 552644 446664 553950 446720
rect 554006 446664 554011 446720
rect 552644 446662 554011 446664
rect 553945 446659 554011 446662
rect 555601 446178 555667 446181
rect 552644 446176 555667 446178
rect 552644 446120 555606 446176
rect 555662 446120 555667 446176
rect 552644 446118 555667 446120
rect 555601 446115 555667 446118
rect 280245 445772 280311 445773
rect 280245 445768 280292 445772
rect 280356 445770 280362 445772
rect 280245 445712 280250 445768
rect 280245 445708 280292 445712
rect 280356 445710 280402 445770
rect 280356 445708 280362 445710
rect 280245 445707 280311 445708
rect 553669 445498 553735 445501
rect 552644 445496 553735 445498
rect 552644 445440 553674 445496
rect 553730 445440 553735 445496
rect 552644 445438 553735 445440
rect 553669 445435 553735 445438
rect 552013 445226 552079 445229
rect 552013 445224 552122 445226
rect 552013 445168 552018 445224
rect 552074 445168 552122 445224
rect 552013 445163 552122 445168
rect 552062 444924 552122 445163
rect 553853 444410 553919 444413
rect 552644 444408 553919 444410
rect 552644 444352 553858 444408
rect 553914 444352 553919 444408
rect 552644 444350 553919 444352
rect 553853 444347 553919 444350
rect 555969 443730 556035 443733
rect 552644 443728 556035 443730
rect 552644 443672 555974 443728
rect 556030 443672 556035 443728
rect 552644 443670 556035 443672
rect 555969 443667 556035 443670
rect 12525 443594 12591 443597
rect 12525 443592 16100 443594
rect 12525 443536 12530 443592
rect 12586 443536 16100 443592
rect 12525 443534 16100 443536
rect 12525 443531 12591 443534
rect 553577 443186 553643 443189
rect 552644 443184 553643 443186
rect 552644 443128 553582 443184
rect 553638 443128 553643 443184
rect 552644 443126 553643 443128
rect 553577 443123 553643 443126
rect 552933 442506 552999 442509
rect 552644 442504 552999 442506
rect 552644 442448 552938 442504
rect 552994 442448 552999 442504
rect 552644 442446 552999 442448
rect 552933 442443 552999 442446
rect 553761 441962 553827 441965
rect 552644 441960 553827 441962
rect 552644 441904 553766 441960
rect 553822 441904 553827 441960
rect 552644 441902 553827 441904
rect 553761 441899 553827 441902
rect 552013 441690 552079 441693
rect 552013 441688 552122 441690
rect 552013 441632 552018 441688
rect 552074 441632 552122 441688
rect 552013 441627 552122 441632
rect 552062 441388 552122 441627
rect 553393 440738 553459 440741
rect 552644 440736 553459 440738
rect 552644 440680 553398 440736
rect 553454 440680 553459 440736
rect 552644 440678 553459 440680
rect 553393 440675 553459 440678
rect 553485 440194 553551 440197
rect 552644 440192 553551 440194
rect 552644 440136 553490 440192
rect 553546 440136 553551 440192
rect 552644 440134 553551 440136
rect 553485 440131 553551 440134
rect 552197 439922 552263 439925
rect 552197 439920 552306 439922
rect 552197 439864 552202 439920
rect 552258 439864 552306 439920
rect 552197 439859 552306 439864
rect 314653 439650 314719 439653
rect 314653 439648 316020 439650
rect 314653 439592 314658 439648
rect 314714 439592 316020 439648
rect 552246 439620 552306 439859
rect 583520 439772 584960 440012
rect 314653 439590 316020 439592
rect 314653 439587 314719 439590
rect 280337 439516 280403 439517
rect 280286 439452 280292 439516
rect 280356 439514 280403 439516
rect 280356 439512 280448 439514
rect 280398 439456 280448 439512
rect 280356 439454 280448 439456
rect 280356 439452 280403 439454
rect 280337 439451 280403 439452
rect 554957 438970 555023 438973
rect 552644 438968 555023 438970
rect 552644 438912 554962 438968
rect 555018 438912 555023 438968
rect 552644 438910 555023 438912
rect 554957 438907 555023 438910
rect 555877 438426 555943 438429
rect 552644 438424 555943 438426
rect 552644 438368 555882 438424
rect 555938 438368 555943 438424
rect 552644 438366 555943 438368
rect 555877 438363 555943 438366
rect -960 438018 480 438108
rect 3417 438018 3483 438021
rect -960 438016 3483 438018
rect -960 437960 3422 438016
rect 3478 437960 3483 438016
rect -960 437958 3483 437960
rect -960 437868 480 437958
rect 3417 437955 3483 437958
rect 555509 437882 555575 437885
rect 552644 437880 555575 437882
rect 552644 437824 555514 437880
rect 555570 437824 555575 437880
rect 552644 437822 555575 437824
rect 555509 437819 555575 437822
rect 556061 437202 556127 437205
rect 552644 437200 556127 437202
rect 552644 437144 556066 437200
rect 556122 437144 556127 437200
rect 552644 437142 556127 437144
rect 556061 437139 556127 437142
rect 554773 436658 554839 436661
rect 552644 436656 554839 436658
rect 552644 436600 554778 436656
rect 554834 436600 554839 436656
rect 552644 436598 554839 436600
rect 554773 436595 554839 436598
rect 554957 436114 555023 436117
rect 552644 436112 555023 436114
rect 552644 436056 554962 436112
rect 555018 436056 555023 436112
rect 552644 436054 555023 436056
rect 554957 436051 555023 436054
rect 554773 435434 554839 435437
rect 552644 435432 554839 435434
rect 552644 435376 554778 435432
rect 554834 435376 554839 435432
rect 552644 435374 554839 435376
rect 554773 435371 554839 435374
rect 554865 434890 554931 434893
rect 552644 434888 554931 434890
rect 552644 434832 554870 434888
rect 554926 434832 554931 434888
rect 552644 434830 554931 434832
rect 554865 434827 554931 434830
rect 280337 434756 280403 434757
rect 280286 434754 280292 434756
rect 280246 434694 280292 434754
rect 280356 434752 280403 434756
rect 280398 434696 280403 434752
rect 280286 434692 280292 434694
rect 280356 434692 280403 434696
rect 280337 434691 280403 434692
rect 554773 434210 554839 434213
rect 552644 434208 554839 434210
rect 552644 434152 554778 434208
rect 554834 434152 554839 434208
rect 552644 434150 554839 434152
rect 554773 434147 554839 434150
rect 554865 433666 554931 433669
rect 552644 433664 554931 433666
rect 552644 433608 554870 433664
rect 554926 433608 554931 433664
rect 552644 433606 554931 433608
rect 554865 433603 554931 433606
rect 554773 433122 554839 433125
rect 552644 433120 554839 433122
rect 552644 433064 554778 433120
rect 554834 433064 554839 433120
rect 552644 433062 554839 433064
rect 554773 433059 554839 433062
rect 554865 432442 554931 432445
rect 552644 432440 554931 432442
rect 552644 432384 554870 432440
rect 554926 432384 554931 432440
rect 552644 432382 554931 432384
rect 554865 432379 554931 432382
rect 554773 431898 554839 431901
rect 552644 431896 554839 431898
rect 552644 431840 554778 431896
rect 554834 431840 554839 431896
rect 552644 431838 554839 431840
rect 554773 431835 554839 431838
rect 554865 431354 554931 431357
rect 552644 431352 554931 431354
rect 552644 431296 554870 431352
rect 554926 431296 554931 431352
rect 552644 431294 554931 431296
rect 554865 431291 554931 431294
rect 554957 430674 555023 430677
rect 552644 430672 555023 430674
rect 552644 430616 554962 430672
rect 555018 430616 555023 430672
rect 552644 430614 555023 430616
rect 554957 430611 555023 430614
rect 281533 430538 281599 430541
rect 282269 430538 282335 430541
rect 279956 430536 282335 430538
rect 279956 430480 281538 430536
rect 281594 430480 282274 430536
rect 282330 430480 282335 430536
rect 279956 430478 282335 430480
rect 281533 430475 281599 430478
rect 282269 430475 282335 430478
rect 554773 430130 554839 430133
rect 552644 430128 554839 430130
rect 552644 430072 554778 430128
rect 554834 430072 554839 430128
rect 552644 430070 554839 430072
rect 554773 430067 554839 430070
rect 554865 429586 554931 429589
rect 552644 429584 554931 429586
rect 552644 429528 554870 429584
rect 554926 429528 554931 429584
rect 552644 429526 554931 429528
rect 554865 429523 554931 429526
rect 554865 428906 554931 428909
rect 552644 428904 554931 428906
rect 552644 428848 554870 428904
rect 554926 428848 554931 428904
rect 552644 428846 554931 428848
rect 554865 428843 554931 428846
rect 317086 428708 317092 428772
rect 317156 428770 317162 428772
rect 338113 428770 338179 428773
rect 317156 428768 338179 428770
rect 317156 428712 338118 428768
rect 338174 428712 338179 428768
rect 317156 428710 338179 428712
rect 317156 428708 317162 428710
rect 338113 428707 338179 428710
rect 316902 428572 316908 428636
rect 316972 428634 316978 428636
rect 338389 428634 338455 428637
rect 316972 428632 338455 428634
rect 316972 428576 338394 428632
rect 338450 428576 338455 428632
rect 316972 428574 338455 428576
rect 316972 428572 316978 428574
rect 338389 428571 338455 428574
rect 280286 428436 280292 428500
rect 280356 428498 280362 428500
rect 281022 428498 281028 428500
rect 280356 428438 281028 428498
rect 280356 428436 280362 428438
rect 281022 428436 281028 428438
rect 281092 428436 281098 428500
rect 317270 428436 317276 428500
rect 317340 428498 317346 428500
rect 343633 428498 343699 428501
rect 317340 428496 343699 428498
rect 317340 428440 343638 428496
rect 343694 428440 343699 428496
rect 317340 428438 343699 428440
rect 317340 428436 317346 428438
rect 343633 428435 343699 428438
rect 554773 428362 554839 428365
rect 552644 428360 554839 428362
rect 552644 428304 554778 428360
rect 554834 428304 554839 428360
rect 552644 428302 554839 428304
rect 554773 428299 554839 428302
rect 583520 428076 584960 428316
rect 554773 427818 554839 427821
rect 552644 427816 554839 427818
rect 552644 427760 554778 427816
rect 554834 427760 554839 427816
rect 552644 427758 554839 427760
rect 554773 427755 554839 427758
rect -960 423738 480 423828
rect 3509 423738 3575 423741
rect -960 423736 3575 423738
rect -960 423680 3514 423736
rect 3570 423680 3575 423736
rect -960 423678 3575 423680
rect -960 423588 480 423678
rect 3509 423675 3575 423678
rect 280838 423540 280844 423604
rect 280908 423602 280914 423604
rect 281022 423602 281028 423604
rect 280908 423542 281028 423602
rect 280908 423540 280914 423542
rect 281022 423540 281028 423542
rect 281092 423540 281098 423604
rect 153886 421290 153946 421804
rect 281625 421292 281691 421293
rect 157190 421290 157196 421292
rect 153886 421230 157196 421290
rect 157190 421228 157196 421230
rect 157260 421228 157266 421292
rect 281574 421228 281580 421292
rect 281644 421290 281691 421292
rect 281644 421288 281736 421290
rect 281686 421232 281736 421288
rect 281644 421230 281736 421232
rect 281644 421228 281691 421230
rect 281625 421227 281691 421228
rect 580165 416530 580231 416533
rect 583520 416530 584960 416620
rect 580165 416528 584960 416530
rect 580165 416472 580170 416528
rect 580226 416472 584960 416528
rect 580165 416470 584960 416472
rect 580165 416467 580231 416470
rect 583520 416380 584960 416470
rect -960 409172 480 409412
rect 580901 404834 580967 404837
rect 583520 404834 584960 404924
rect 580901 404832 584960 404834
rect 580901 404776 580906 404832
rect 580962 404776 584960 404832
rect 580901 404774 584960 404776
rect 580901 404771 580967 404774
rect 583520 404684 584960 404774
rect 121361 401570 121427 401573
rect 151118 401570 151124 401572
rect 121361 401568 151124 401570
rect 121361 401512 121366 401568
rect 121422 401512 151124 401568
rect 121361 401510 151124 401512
rect 121361 401507 121427 401510
rect 151118 401508 151124 401510
rect 151188 401508 151194 401572
rect 115749 401434 115815 401437
rect 148358 401434 148364 401436
rect 115749 401432 148364 401434
rect 115749 401376 115754 401432
rect 115810 401376 148364 401432
rect 115749 401374 148364 401376
rect 115749 401371 115815 401374
rect 148358 401372 148364 401374
rect 148428 401372 148434 401436
rect 114461 401298 114527 401301
rect 147990 401298 147996 401300
rect 114461 401296 147996 401298
rect 114461 401240 114466 401296
rect 114522 401240 147996 401296
rect 114461 401238 147996 401240
rect 114461 401235 114527 401238
rect 147990 401236 147996 401238
rect 148060 401236 148066 401300
rect 115841 401162 115907 401165
rect 150198 401162 150204 401164
rect 115841 401160 150204 401162
rect 115841 401104 115846 401160
rect 115902 401104 150204 401160
rect 115841 401102 150204 401104
rect 115841 401099 115907 401102
rect 150198 401100 150204 401102
rect 150268 401100 150274 401164
rect 111701 401026 111767 401029
rect 150014 401026 150020 401028
rect 111701 401024 150020 401026
rect 111701 400968 111706 401024
rect 111762 400968 150020 401024
rect 111701 400966 150020 400968
rect 111701 400963 111767 400966
rect 150014 400964 150020 400966
rect 150084 400964 150090 401028
rect 111609 400890 111675 400893
rect 151302 400890 151308 400892
rect 111609 400888 151308 400890
rect 111609 400832 111614 400888
rect 111670 400832 151308 400888
rect 111609 400830 151308 400832
rect 111609 400827 111675 400830
rect 151302 400828 151308 400830
rect 151372 400828 151378 400892
rect 135161 400754 135227 400757
rect 150566 400754 150572 400756
rect 135161 400752 150572 400754
rect 135161 400696 135166 400752
rect 135222 400696 150572 400752
rect 135161 400694 150572 400696
rect 135161 400691 135227 400694
rect 150566 400692 150572 400694
rect 150636 400692 150642 400756
rect 136541 400618 136607 400621
rect 150750 400618 150756 400620
rect 136541 400616 150756 400618
rect 136541 400560 136546 400616
rect 136602 400560 150756 400616
rect 136541 400558 150756 400560
rect 136541 400555 136607 400558
rect 150750 400556 150756 400558
rect 150820 400556 150826 400620
rect 139301 400482 139367 400485
rect 149278 400482 149284 400484
rect 139301 400480 149284 400482
rect 139301 400424 139306 400480
rect 139362 400424 149284 400480
rect 139301 400422 149284 400424
rect 139301 400419 139367 400422
rect 149278 400420 149284 400422
rect 149348 400420 149354 400484
rect 146201 400346 146267 400349
rect 153326 400346 153332 400348
rect 146201 400344 153332 400346
rect 146201 400288 146206 400344
rect 146262 400288 153332 400344
rect 146201 400286 153332 400288
rect 146201 400283 146267 400286
rect 153326 400284 153332 400286
rect 153396 400284 153402 400348
rect -960 395042 480 395132
rect 4797 395042 4863 395045
rect -960 395040 4863 395042
rect -960 394984 4802 395040
rect 4858 394984 4863 395040
rect -960 394982 4863 394984
rect -960 394892 480 394982
rect 4797 394979 4863 394982
rect 583520 392852 584960 393092
rect 284293 392730 284359 392733
rect 282716 392728 284359 392730
rect 282716 392672 284298 392728
rect 284354 392672 284359 392728
rect 282716 392670 284359 392672
rect 284293 392667 284359 392670
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 2773 380626 2839 380629
rect -960 380624 2839 380626
rect -960 380568 2778 380624
rect 2834 380568 2839 380624
rect -960 380566 2839 380568
rect -960 380476 480 380566
rect 2773 380563 2839 380566
rect 75870 376818 75930 377332
rect 189942 376818 189948 376820
rect 75870 376758 189948 376818
rect 189942 376756 189948 376758
rect 190012 376756 190018 376820
rect 282453 369882 282519 369885
rect 282453 369880 282562 369882
rect 282453 369824 282458 369880
rect 282514 369824 282562 369880
rect 282453 369819 282562 369824
rect 282502 369580 282562 369819
rect 580165 369610 580231 369613
rect 583520 369610 584960 369700
rect 580165 369608 584960 369610
rect 580165 369552 580170 369608
rect 580226 369552 584960 369608
rect 580165 369550 584960 369552
rect 580165 369547 580231 369550
rect 583520 369460 584960 369550
rect -960 366210 480 366300
rect 2773 366210 2839 366213
rect -960 366208 2839 366210
rect -960 366152 2778 366208
rect 2834 366152 2839 366208
rect -960 366150 2839 366152
rect -960 366060 480 366150
rect 2773 366147 2839 366150
rect 77937 363762 78003 363765
rect 75900 363760 78003 363762
rect 75900 363704 77942 363760
rect 77998 363704 78003 363760
rect 75900 363702 78003 363704
rect 77937 363699 78003 363702
rect 189942 360028 189948 360092
rect 190012 360090 190018 360092
rect 282545 360090 282611 360093
rect 190012 360088 282611 360090
rect 190012 360032 282550 360088
rect 282606 360032 282611 360088
rect 190012 360030 282611 360032
rect 190012 360028 190018 360030
rect 282545 360027 282611 360030
rect 580901 357914 580967 357917
rect 583520 357914 584960 358004
rect 580901 357912 584960 357914
rect 580901 357856 580906 357912
rect 580962 357856 584960 357912
rect 580901 357854 584960 357856
rect 580901 357851 580967 357854
rect 583520 357764 584960 357854
rect 20294 357580 20300 357644
rect 20364 357642 20370 357644
rect 21357 357642 21423 357645
rect 20364 357640 21423 357642
rect 20364 357584 21362 357640
rect 21418 357584 21423 357640
rect 20364 357582 21423 357584
rect 20364 357580 20370 357582
rect 21357 357579 21423 357582
rect 280470 357580 280476 357644
rect 280540 357642 280546 357644
rect 281022 357642 281028 357644
rect 280540 357582 281028 357642
rect 280540 357580 280546 357582
rect 281022 357580 281028 357582
rect 281092 357580 281098 357644
rect 188838 357444 188844 357508
rect 188908 357506 188914 357508
rect 194133 357506 194199 357509
rect 188908 357504 194199 357506
rect 188908 357448 194138 357504
rect 194194 357448 194199 357504
rect 188908 357446 194199 357448
rect 188908 357444 188914 357446
rect 194133 357443 194199 357446
rect -960 351780 480 352020
rect 122238 351870 122850 351930
rect 119337 351794 119403 351797
rect 122238 351794 122298 351870
rect 119337 351792 122298 351794
rect 119337 351736 119342 351792
rect 119398 351736 122298 351792
rect 119337 351734 122298 351736
rect 122465 351794 122531 351797
rect 122598 351794 122604 351796
rect 122465 351792 122604 351794
rect 122465 351736 122470 351792
rect 122526 351736 122604 351792
rect 122465 351734 122604 351736
rect 119337 351731 119403 351734
rect 122465 351731 122531 351734
rect 122598 351732 122604 351734
rect 122668 351732 122674 351796
rect 122790 351794 122850 351870
rect 189441 351794 189507 351797
rect 189758 351794 189764 351796
rect 122790 351734 147506 351794
rect 112897 351658 112963 351661
rect 147254 351658 147260 351660
rect 112897 351656 147260 351658
rect 112897 351600 112902 351656
rect 112958 351600 147260 351656
rect 112897 351598 147260 351600
rect 112897 351595 112963 351598
rect 147254 351596 147260 351598
rect 147324 351596 147330 351660
rect 147446 351658 147506 351734
rect 189441 351792 189764 351794
rect 189441 351736 189446 351792
rect 189502 351736 189764 351792
rect 189441 351734 189764 351736
rect 189441 351731 189507 351734
rect 189758 351732 189764 351734
rect 189828 351732 189834 351796
rect 191046 351732 191052 351796
rect 191116 351794 191122 351796
rect 191189 351794 191255 351797
rect 191116 351792 191255 351794
rect 191116 351736 191194 351792
rect 191250 351736 191255 351792
rect 191116 351734 191255 351736
rect 191116 351732 191122 351734
rect 191189 351731 191255 351734
rect 151854 351658 151860 351660
rect 147446 351598 151860 351658
rect 151854 351596 151860 351598
rect 151924 351596 151930 351660
rect 189574 351596 189580 351660
rect 189644 351658 189650 351660
rect 189901 351658 189967 351661
rect 189644 351656 189967 351658
rect 189644 351600 189906 351656
rect 189962 351600 189967 351656
rect 189644 351598 189967 351600
rect 189644 351596 189650 351598
rect 189901 351595 189967 351598
rect 109585 351522 109651 351525
rect 146293 351522 146359 351525
rect 109585 351520 146359 351522
rect 109585 351464 109590 351520
rect 109646 351464 146298 351520
rect 146354 351464 146359 351520
rect 109585 351462 146359 351464
rect 109585 351459 109651 351462
rect 146293 351459 146359 351462
rect 146937 351522 147003 351525
rect 147070 351522 147076 351524
rect 146937 351520 147076 351522
rect 146937 351464 146942 351520
rect 146998 351464 147076 351520
rect 146937 351462 147076 351464
rect 146937 351459 147003 351462
rect 147070 351460 147076 351462
rect 147140 351460 147146 351524
rect 148041 351522 148107 351525
rect 148174 351522 148180 351524
rect 148041 351520 148180 351522
rect 148041 351464 148046 351520
rect 148102 351464 148180 351520
rect 148041 351462 148180 351464
rect 148041 351459 148107 351462
rect 148174 351460 148180 351462
rect 148244 351460 148250 351524
rect 149421 351522 149487 351525
rect 149646 351522 149652 351524
rect 149421 351520 149652 351522
rect 149421 351464 149426 351520
rect 149482 351464 149652 351520
rect 149421 351462 149652 351464
rect 149421 351459 149487 351462
rect 149646 351460 149652 351462
rect 149716 351460 149722 351524
rect 149830 351460 149836 351524
rect 149900 351522 149906 351524
rect 150065 351522 150131 351525
rect 149900 351520 150131 351522
rect 149900 351464 150070 351520
rect 150126 351464 150131 351520
rect 149900 351462 150131 351464
rect 149900 351460 149906 351462
rect 150065 351459 150131 351462
rect 150934 351460 150940 351524
rect 151004 351522 151010 351524
rect 151169 351522 151235 351525
rect 152365 351524 152431 351525
rect 152365 351522 152412 351524
rect 151004 351520 151235 351522
rect 151004 351464 151174 351520
rect 151230 351464 151235 351520
rect 151004 351462 151235 351464
rect 152320 351520 152412 351522
rect 152320 351464 152370 351520
rect 152320 351462 152412 351464
rect 151004 351460 151010 351462
rect 151169 351459 151235 351462
rect 152365 351460 152412 351462
rect 152476 351460 152482 351524
rect 152365 351459 152431 351460
rect 107561 351386 107627 351389
rect 147622 351386 147628 351388
rect 107561 351384 147628 351386
rect 107561 351328 107566 351384
rect 107622 351328 147628 351384
rect 107561 351326 147628 351328
rect 107561 351323 107627 351326
rect 147622 351324 147628 351326
rect 147692 351324 147698 351388
rect 108665 351250 108731 351253
rect 145557 351250 145623 351253
rect 108665 351248 145623 351250
rect 108665 351192 108670 351248
rect 108726 351192 145562 351248
rect 145618 351192 145623 351248
rect 108665 351190 145623 351192
rect 108665 351187 108731 351190
rect 145557 351187 145623 351190
rect 146293 351250 146359 351253
rect 150382 351250 150388 351252
rect 146293 351248 150388 351250
rect 146293 351192 146298 351248
rect 146354 351192 150388 351248
rect 146293 351190 150388 351192
rect 146293 351187 146359 351190
rect 150382 351188 150388 351190
rect 150452 351188 150458 351252
rect 75821 351114 75887 351117
rect 104893 351114 104959 351117
rect 75821 351112 104959 351114
rect 75821 351056 75826 351112
rect 75882 351056 104898 351112
rect 104954 351056 104959 351112
rect 75821 351054 104959 351056
rect 75821 351051 75887 351054
rect 104893 351051 104959 351054
rect 106181 351114 106247 351117
rect 147438 351114 147444 351116
rect 106181 351112 147444 351114
rect 106181 351056 106186 351112
rect 106242 351056 147444 351112
rect 106181 351054 147444 351056
rect 106181 351051 106247 351054
rect 147438 351052 147444 351054
rect 147508 351052 147514 351116
rect 117129 350978 117195 350981
rect 144913 350978 144979 350981
rect 117129 350976 144979 350978
rect 117129 350920 117134 350976
rect 117190 350920 144918 350976
rect 144974 350920 144979 350976
rect 117129 350918 144979 350920
rect 117129 350915 117195 350918
rect 144913 350915 144979 350918
rect 145557 350978 145623 350981
rect 149094 350978 149100 350980
rect 145557 350976 149100 350978
rect 145557 350920 145562 350976
rect 145618 350920 149100 350976
rect 145557 350918 149100 350920
rect 145557 350915 145623 350918
rect 149094 350916 149100 350918
rect 149164 350916 149170 350980
rect 129089 350842 129155 350845
rect 129590 350842 129596 350844
rect 129089 350840 129596 350842
rect 129089 350784 129094 350840
rect 129150 350784 129596 350840
rect 129089 350782 129596 350784
rect 129089 350779 129155 350782
rect 129590 350780 129596 350782
rect 129660 350780 129666 350844
rect 129733 350842 129799 350845
rect 152038 350842 152044 350844
rect 129733 350840 152044 350842
rect 129733 350784 129738 350840
rect 129794 350784 152044 350840
rect 129733 350782 152044 350784
rect 129733 350779 129799 350782
rect 152038 350780 152044 350782
rect 152108 350780 152114 350844
rect 126881 350706 126947 350709
rect 153142 350706 153148 350708
rect 126881 350704 153148 350706
rect 126881 350648 126886 350704
rect 126942 350648 153148 350704
rect 126881 350646 153148 350648
rect 126881 350643 126947 350646
rect 153142 350644 153148 350646
rect 153212 350644 153218 350708
rect 124673 350570 124739 350573
rect 129733 350570 129799 350573
rect 124673 350568 129799 350570
rect 124673 350512 124678 350568
rect 124734 350512 129738 350568
rect 129794 350512 129799 350568
rect 124673 350510 129799 350512
rect 124673 350507 124739 350510
rect 129733 350507 129799 350510
rect 144913 350570 144979 350573
rect 147806 350570 147812 350572
rect 144913 350568 147812 350570
rect 144913 350512 144918 350568
rect 144974 350512 147812 350568
rect 144913 350510 147812 350512
rect 144913 350507 144979 350510
rect 147806 350508 147812 350510
rect 147876 350508 147882 350572
rect 280286 350372 280292 350436
rect 280356 350434 280362 350436
rect 280838 350434 280844 350436
rect 280356 350374 280844 350434
rect 280356 350372 280362 350374
rect 280838 350372 280844 350374
rect 280908 350372 280914 350436
rect 280286 347652 280292 347716
rect 280356 347652 280362 347716
rect 280294 347581 280354 347652
rect 280294 347576 280403 347581
rect 280294 347520 280342 347576
rect 280398 347520 280403 347576
rect 280294 347518 280403 347520
rect 280337 347515 280403 347518
rect 583520 345932 584960 346172
rect 280337 338194 280403 338197
rect 280654 338194 280660 338196
rect 280337 338192 280660 338194
rect 280337 338136 280342 338192
rect 280398 338136 280660 338192
rect 280337 338134 280660 338136
rect 280337 338131 280403 338134
rect 280654 338132 280660 338134
rect 280724 338132 280730 338196
rect -960 337514 480 337604
rect 3141 337514 3207 337517
rect -960 337512 3207 337514
rect -960 337456 3146 337512
rect 3202 337456 3207 337512
rect -960 337454 3207 337456
rect -960 337364 480 337454
rect 3141 337451 3207 337454
rect 280654 336636 280660 336700
rect 280724 336636 280730 336700
rect 280286 336500 280292 336564
rect 280356 336562 280362 336564
rect 280662 336562 280722 336636
rect 280356 336502 280722 336562
rect 280356 336500 280362 336502
rect 282269 336018 282335 336021
rect 279006 336016 282335 336018
rect 279006 335960 282274 336016
rect 282330 335960 282335 336016
rect 279006 335958 282335 335960
rect 279006 335920 279066 335958
rect 282269 335955 282335 335958
rect 583520 334236 584960 334476
rect 304257 328266 304323 328269
rect 301668 328264 304323 328266
rect 301668 328208 304262 328264
rect 304318 328208 304323 328264
rect 301668 328206 304323 328208
rect 304257 328203 304323 328206
rect 280337 327044 280403 327045
rect 280286 326980 280292 327044
rect 280356 327042 280403 327044
rect 280356 327040 280448 327042
rect 280398 326984 280448 327040
rect 280356 326982 280448 326984
rect 280356 326980 280403 326982
rect 280337 326979 280403 326980
rect 303613 326362 303679 326365
rect 301668 326360 303679 326362
rect 301668 326304 303618 326360
rect 303674 326304 303679 326360
rect 301668 326302 303679 326304
rect 303613 326299 303679 326302
rect 289721 325274 289787 325277
rect 289721 325272 290812 325274
rect 289721 325216 289726 325272
rect 289782 325216 290812 325272
rect 289721 325214 290812 325216
rect 289721 325211 289787 325214
rect 303613 324458 303679 324461
rect 301668 324456 303679 324458
rect 301668 324400 303618 324456
rect 303674 324400 303679 324456
rect 301668 324398 303679 324400
rect 303613 324395 303679 324398
rect -960 323098 480 323188
rect 2773 323098 2839 323101
rect -960 323096 2839 323098
rect -960 323040 2778 323096
rect 2834 323040 2839 323096
rect -960 323038 2839 323040
rect -960 322948 480 323038
rect 2773 323035 2839 323038
rect 580165 322690 580231 322693
rect 583520 322690 584960 322780
rect 580165 322688 584960 322690
rect 580165 322632 580170 322688
rect 580226 322632 584960 322688
rect 580165 322630 584960 322632
rect 580165 322627 580231 322630
rect 304349 322554 304415 322557
rect 301668 322552 304415 322554
rect 301668 322496 304354 322552
rect 304410 322496 304415 322552
rect 583520 322540 584960 322630
rect 301668 322494 304415 322496
rect 304349 322491 304415 322494
rect 214414 322084 214420 322148
rect 214484 322146 214490 322148
rect 282177 322146 282243 322149
rect 214484 322144 282243 322146
rect 214484 322088 282182 322144
rect 282238 322088 282243 322144
rect 214484 322086 282243 322088
rect 214484 322084 214490 322086
rect 282177 322083 282243 322086
rect 20478 320724 20484 320788
rect 20548 320786 20554 320788
rect 51574 320786 51580 320788
rect 20548 320726 51580 320786
rect 20548 320724 20554 320726
rect 51574 320724 51580 320726
rect 51644 320724 51650 320788
rect 304441 320650 304507 320653
rect 301668 320648 304507 320650
rect 301668 320592 304446 320648
rect 304502 320592 304507 320648
rect 301668 320590 304507 320592
rect 304441 320587 304507 320590
rect 189073 320514 189139 320517
rect 195094 320514 195100 320516
rect 189073 320512 195100 320514
rect 189073 320456 189078 320512
rect 189134 320456 195100 320512
rect 189073 320454 195100 320456
rect 189073 320451 189139 320454
rect 195094 320452 195100 320454
rect 195164 320452 195170 320516
rect 192385 320378 192451 320381
rect 196566 320378 196572 320380
rect 192385 320376 196572 320378
rect 192385 320320 192390 320376
rect 192446 320320 196572 320376
rect 192385 320318 196572 320320
rect 192385 320315 192451 320318
rect 196566 320316 196572 320318
rect 196636 320316 196642 320380
rect 190177 320242 190243 320245
rect 190310 320242 190316 320244
rect 190177 320240 190316 320242
rect 190177 320184 190182 320240
rect 190238 320184 190316 320240
rect 190177 320182 190316 320184
rect 190177 320179 190243 320182
rect 190310 320180 190316 320182
rect 190380 320180 190386 320244
rect 191281 320242 191347 320245
rect 191598 320242 191604 320244
rect 191281 320240 191604 320242
rect 191281 320184 191286 320240
rect 191342 320184 191604 320240
rect 191281 320182 191604 320184
rect 191281 320179 191347 320182
rect 191598 320180 191604 320182
rect 191668 320180 191674 320244
rect 194358 320180 194364 320244
rect 194428 320242 194434 320244
rect 194501 320242 194567 320245
rect 194428 320240 194567 320242
rect 194428 320184 194506 320240
rect 194562 320184 194567 320240
rect 194428 320182 194567 320184
rect 194428 320180 194434 320182
rect 194501 320179 194567 320182
rect 193397 319426 193463 319429
rect 208342 319426 208348 319428
rect 193397 319424 208348 319426
rect 193397 319368 193402 319424
rect 193458 319368 208348 319424
rect 193397 319366 208348 319368
rect 193397 319363 193463 319366
rect 208342 319364 208348 319366
rect 208412 319364 208418 319428
rect 303613 318746 303679 318749
rect 301668 318744 303679 318746
rect 301668 318688 303618 318744
rect 303674 318688 303679 318744
rect 301668 318686 303679 318688
rect 303613 318683 303679 318686
rect 280337 317660 280403 317661
rect 280286 317658 280292 317660
rect 280246 317598 280292 317658
rect 280356 317656 280403 317660
rect 280398 317600 280403 317656
rect 280286 317596 280292 317598
rect 280356 317596 280403 317600
rect 280337 317595 280403 317596
rect 280337 317388 280403 317389
rect 280286 317324 280292 317388
rect 280356 317386 280403 317388
rect 280356 317384 280448 317386
rect 280398 317328 280448 317384
rect 280356 317326 280448 317328
rect 280356 317324 280403 317326
rect 280337 317323 280403 317324
rect 288893 317114 288959 317117
rect 288893 317112 290812 317114
rect 288893 317056 288898 317112
rect 288954 317056 290812 317112
rect 288893 317054 290812 317056
rect 288893 317051 288959 317054
rect 304349 316978 304415 316981
rect 301668 316976 304415 316978
rect 301668 316920 304354 316976
rect 304410 316920 304415 316976
rect 301668 316918 304415 316920
rect 304349 316915 304415 316918
rect 304257 315074 304323 315077
rect 301668 315072 304323 315074
rect 301668 315016 304262 315072
rect 304318 315016 304323 315072
rect 301668 315014 304323 315016
rect 304257 315011 304323 315014
rect 303613 313170 303679 313173
rect 301668 313168 303679 313170
rect 301668 313112 303618 313168
rect 303674 313112 303679 313168
rect 301668 313110 303679 313112
rect 303613 313107 303679 313110
rect 303613 311266 303679 311269
rect 301668 311264 303679 311266
rect 301668 311208 303618 311264
rect 303674 311208 303679 311264
rect 301668 311206 303679 311208
rect 303613 311203 303679 311206
rect 580349 310858 580415 310861
rect 580901 310858 580967 310861
rect 583520 310858 584960 310948
rect 580349 310856 584960 310858
rect 580349 310800 580354 310856
rect 580410 310800 580906 310856
rect 580962 310800 584960 310856
rect 580349 310798 584960 310800
rect 580349 310795 580415 310798
rect 580901 310795 580967 310798
rect 583520 310708 584960 310798
rect 280337 309636 280403 309637
rect 280286 309634 280292 309636
rect 280246 309574 280292 309634
rect 280356 309632 280403 309636
rect 280398 309576 280403 309632
rect 280286 309572 280292 309574
rect 280356 309572 280403 309576
rect 280337 309571 280403 309572
rect 303613 309362 303679 309365
rect 301668 309360 303679 309362
rect 301668 309304 303618 309360
rect 303674 309304 303679 309360
rect 301668 309302 303679 309304
rect 303613 309299 303679 309302
rect 2773 309090 2839 309093
rect 3509 309090 3575 309093
rect 2773 309088 3575 309090
rect 2773 309032 2778 309088
rect 2834 309032 3514 309088
rect 3570 309032 3575 309088
rect 2773 309030 3575 309032
rect 2773 309027 2839 309030
rect 3509 309027 3575 309030
rect 289629 308954 289695 308957
rect 289629 308952 290812 308954
rect -960 308818 480 308908
rect 289629 308896 289634 308952
rect 289690 308896 290812 308952
rect 289629 308894 290812 308896
rect 289629 308891 289695 308894
rect 2773 308818 2839 308821
rect -960 308816 2839 308818
rect -960 308760 2778 308816
rect 2834 308760 2839 308816
rect -960 308758 2839 308760
rect -960 308668 480 308758
rect 2773 308755 2839 308758
rect 303613 307458 303679 307461
rect 301668 307456 303679 307458
rect 301668 307400 303618 307456
rect 303674 307400 303679 307456
rect 301668 307398 303679 307400
rect 303613 307395 303679 307398
rect 280286 306308 280292 306372
rect 280356 306370 280362 306372
rect 280470 306370 280476 306372
rect 280356 306310 280476 306370
rect 280356 306308 280362 306310
rect 280470 306308 280476 306310
rect 280540 306308 280546 306372
rect 300902 305557 300962 305660
rect 300853 305552 300962 305557
rect 300853 305496 300858 305552
rect 300914 305496 300962 305552
rect 300853 305494 300962 305496
rect 300853 305491 300919 305494
rect 292573 302834 292639 302837
rect 332910 302834 332916 302836
rect 292573 302832 332916 302834
rect 292573 302776 292578 302832
rect 292634 302776 332916 302832
rect 292573 302774 332916 302776
rect 292573 302771 292639 302774
rect 332910 302772 332916 302774
rect 332980 302772 332986 302836
rect 583520 299012 584960 299252
rect 280654 296652 280660 296716
rect 280724 296714 280730 296716
rect 281022 296714 281028 296716
rect 280724 296654 281028 296714
rect 280724 296652 280730 296654
rect 281022 296652 281028 296654
rect 281092 296652 281098 296716
rect 279509 295898 279575 295901
rect 279509 295896 279618 295898
rect 279509 295840 279514 295896
rect 279570 295840 279618 295896
rect 279509 295835 279618 295840
rect 113357 295354 113423 295357
rect 111964 295352 113423 295354
rect 111964 295296 113362 295352
rect 113418 295296 113423 295352
rect 279558 295324 279618 295835
rect 111964 295294 113423 295296
rect 113357 295291 113423 295294
rect 281022 295156 281028 295220
rect 281092 295156 281098 295220
rect 280705 295082 280771 295085
rect 281030 295082 281090 295156
rect 280705 295080 281090 295082
rect 280705 295024 280710 295080
rect 280766 295024 281090 295080
rect 280705 295022 281090 295024
rect 280705 295019 280771 295022
rect -960 294402 480 294492
rect 3601 294402 3667 294405
rect -960 294400 3667 294402
rect -960 294344 3606 294400
rect 3662 294344 3667 294400
rect -960 294342 3667 294344
rect -960 294252 480 294342
rect 3601 294339 3667 294342
rect 583520 287316 584960 287556
rect -960 280122 480 280212
rect 2773 280122 2839 280125
rect -960 280120 2839 280122
rect -960 280064 2778 280120
rect 2834 280064 2839 280120
rect -960 280062 2839 280064
rect -960 279972 480 280062
rect 2773 280059 2839 280062
rect 280705 277674 280771 277677
rect 280478 277672 280771 277674
rect 280478 277616 280710 277672
rect 280766 277616 280771 277672
rect 280478 277614 280771 277616
rect 280478 277540 280538 277614
rect 280705 277611 280771 277614
rect 280470 277476 280476 277540
rect 280540 277476 280546 277540
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 17125 274954 17191 274957
rect 185577 274954 185643 274957
rect 17125 274952 20148 274954
rect 17125 274896 17130 274952
rect 17186 274896 20148 274952
rect 17125 274894 20148 274896
rect 185577 274952 188140 274954
rect 185577 274896 185582 274952
rect 185638 274896 188140 274952
rect 185577 274894 188140 274896
rect 17125 274891 17191 274894
rect 185577 274891 185643 274894
rect 280470 273458 280476 273460
rect 280294 273398 280476 273458
rect 280294 273188 280354 273398
rect 280470 273396 280476 273398
rect 280540 273396 280546 273460
rect 280286 273124 280292 273188
rect 280356 273124 280362 273188
rect -960 265706 480 265796
rect 2773 265706 2839 265709
rect -960 265704 2839 265706
rect -960 265648 2778 265704
rect 2834 265648 2839 265704
rect -960 265646 2839 265648
rect -960 265556 480 265646
rect 2773 265643 2839 265646
rect 580349 263938 580415 263941
rect 580901 263938 580967 263941
rect 583520 263938 584960 264028
rect 580349 263936 584960 263938
rect 580349 263880 580354 263936
rect 580410 263880 580906 263936
rect 580962 263880 584960 263936
rect 580349 263878 584960 263880
rect 580349 263875 580415 263878
rect 580901 263875 580967 263878
rect 583520 263788 584960 263878
rect 280286 259524 280292 259588
rect 280356 259586 280362 259588
rect 280470 259586 280476 259588
rect 280356 259526 280476 259586
rect 280356 259524 280362 259526
rect 280470 259524 280476 259526
rect 280540 259524 280546 259588
rect 282177 255098 282243 255101
rect 279926 255096 282243 255098
rect 279926 255040 282182 255096
rect 282238 255040 282243 255096
rect 279926 255038 282243 255040
rect 279926 254554 279986 255038
rect 282177 255035 282243 255038
rect 279404 254524 279986 254554
rect 111934 254010 111994 254524
rect 279374 254494 279956 254524
rect 146017 254146 146083 254149
rect 138062 254144 146083 254146
rect 138062 254088 146022 254144
rect 146078 254088 146083 254144
rect 138062 254086 146083 254088
rect 138062 254010 138122 254086
rect 146017 254083 146083 254086
rect 149513 254146 149579 254149
rect 149513 254144 154498 254146
rect 149513 254088 149518 254144
rect 149574 254088 154498 254144
rect 149513 254086 154498 254088
rect 149513 254083 149579 254086
rect 111934 253950 138122 254010
rect 154438 254010 154498 254086
rect 279374 254012 279434 254494
rect 181662 254010 181668 254012
rect 154438 253950 161490 254010
rect 161430 253874 161490 253950
rect 171182 253950 181668 254010
rect 161430 253814 167010 253874
rect 166950 253602 167010 253814
rect 171182 253602 171242 253950
rect 181662 253948 181668 253950
rect 181732 253948 181738 254012
rect 279366 253948 279372 254012
rect 279436 253948 279442 254012
rect 166950 253542 171242 253602
rect 583520 252092 584960 252332
rect -960 251140 480 251380
rect 280521 251156 280587 251157
rect 280470 251154 280476 251156
rect 280430 251094 280476 251154
rect 280540 251152 280587 251156
rect 280582 251096 280587 251152
rect 280470 251092 280476 251094
rect 280540 251092 280587 251096
rect 280521 251091 280587 251092
rect 280521 241634 280587 241637
rect 280654 241634 280660 241636
rect 280521 241632 280660 241634
rect 280521 241576 280526 241632
rect 280582 241576 280660 241632
rect 280521 241574 280660 241576
rect 280521 241571 280587 241574
rect 280654 241572 280660 241574
rect 280724 241572 280730 241636
rect 583520 240396 584960 240636
rect -960 237010 480 237100
rect 2773 237010 2839 237013
rect -960 237008 2839 237010
rect -960 236952 2778 237008
rect 2834 236952 2839 237008
rect -960 236950 2839 236952
rect -960 236860 480 236950
rect 2773 236947 2839 236950
rect 51574 235996 51580 236060
rect 51644 236058 51650 236060
rect 67173 236058 67239 236061
rect 51644 236056 67239 236058
rect 51644 236000 67178 236056
rect 67234 236000 67239 236056
rect 51644 235998 67239 236000
rect 51644 235996 51650 235998
rect 67173 235995 67239 235998
rect 194358 235180 194364 235244
rect 194428 235242 194434 235244
rect 209773 235242 209839 235245
rect 194428 235240 209839 235242
rect 194428 235184 209778 235240
rect 209834 235184 209839 235240
rect 194428 235182 209839 235184
rect 194428 235180 194434 235182
rect 209773 235179 209839 235182
rect 250437 235242 250503 235245
rect 280654 235242 280660 235244
rect 250437 235240 280660 235242
rect 250437 235184 250442 235240
rect 250498 235184 280660 235240
rect 250437 235182 280660 235184
rect 250437 235179 250503 235182
rect 280654 235180 280660 235182
rect 280724 235180 280730 235244
rect 191598 233820 191604 233884
rect 191668 233882 191674 233884
rect 205817 233882 205883 233885
rect 191668 233880 205883 233882
rect 191668 233824 205822 233880
rect 205878 233824 205883 233880
rect 191668 233822 205883 233824
rect 191668 233820 191674 233822
rect 205817 233819 205883 233822
rect 196566 232460 196572 232524
rect 196636 232522 196642 232524
rect 207013 232522 207079 232525
rect 196636 232520 207079 232522
rect 196636 232464 207018 232520
rect 207074 232464 207079 232520
rect 196636 232462 207079 232464
rect 196636 232460 196642 232462
rect 207013 232459 207079 232462
rect 190310 229740 190316 229804
rect 190380 229802 190386 229804
rect 205725 229802 205791 229805
rect 190380 229800 205791 229802
rect 190380 229744 205730 229800
rect 205786 229744 205791 229800
rect 190380 229742 205791 229744
rect 190380 229740 190386 229742
rect 205725 229739 205791 229742
rect 579981 228850 580047 228853
rect 583520 228850 584960 228940
rect 579981 228848 584960 228850
rect 579981 228792 579986 228848
rect 580042 228792 584960 228848
rect 579981 228790 584960 228792
rect 579981 228787 580047 228790
rect 583520 228700 584960 228790
rect 195094 228244 195100 228308
rect 195164 228306 195170 228308
rect 204529 228306 204595 228309
rect 195164 228304 204595 228306
rect 195164 228248 204534 228304
rect 204590 228248 204595 228304
rect 195164 228246 204595 228248
rect 195164 228244 195170 228246
rect 204529 228243 204595 228246
rect 208342 223620 208348 223684
rect 208412 223682 208418 223684
rect 208853 223682 208919 223685
rect 208412 223680 208919 223682
rect 208412 223624 208858 223680
rect 208914 223624 208919 223680
rect 208412 223622 208919 223624
rect 208412 223620 208418 223622
rect 208853 223619 208919 223622
rect -960 222594 480 222684
rect 2773 222594 2839 222597
rect -960 222592 2839 222594
rect -960 222536 2778 222592
rect 2834 222536 2839 222592
rect -960 222534 2839 222536
rect -960 222444 480 222534
rect 2773 222531 2839 222534
rect 213913 221370 213979 221373
rect 211508 221368 213979 221370
rect 211508 221312 213918 221368
rect 213974 221312 213979 221368
rect 211508 221310 213979 221312
rect 213913 221307 213979 221310
rect 229001 221370 229067 221373
rect 229001 221368 230092 221370
rect 229001 221312 229006 221368
rect 229062 221312 230092 221368
rect 229001 221310 230092 221312
rect 229001 221307 229067 221310
rect 116393 221234 116459 221237
rect 116393 221232 119692 221234
rect 116393 221176 116398 221232
rect 116454 221176 119692 221232
rect 116393 221174 119692 221176
rect 116393 221171 116459 221174
rect 226333 220826 226399 220829
rect 226333 220824 230092 220826
rect 226333 220768 226338 220824
rect 226394 220768 230092 220824
rect 226333 220766 230092 220768
rect 226333 220763 226399 220766
rect 214005 220554 214071 220557
rect 211508 220552 214071 220554
rect 211508 220496 214010 220552
rect 214066 220496 214071 220552
rect 211508 220494 214071 220496
rect 214005 220491 214071 220494
rect 226333 220146 226399 220149
rect 226333 220144 230092 220146
rect 226333 220088 226338 220144
rect 226394 220088 230092 220144
rect 226333 220086 230092 220088
rect 226333 220083 226399 220086
rect 116117 220010 116183 220013
rect 116117 220008 119692 220010
rect 116117 219952 116122 220008
rect 116178 219952 119692 220008
rect 116117 219950 119692 219952
rect 116117 219947 116183 219950
rect 213913 219738 213979 219741
rect 211508 219736 213979 219738
rect 211508 219680 213918 219736
rect 213974 219680 213979 219736
rect 211508 219678 213979 219680
rect 213913 219675 213979 219678
rect 226425 219602 226491 219605
rect 226425 219600 230092 219602
rect 226425 219544 226430 219600
rect 226486 219544 230092 219600
rect 226425 219542 230092 219544
rect 226425 219539 226491 219542
rect 104801 219330 104867 219333
rect 101078 219328 104867 219330
rect 101078 219272 104806 219328
rect 104862 219272 104867 219328
rect 101078 219270 104867 219272
rect 101078 219096 101138 219270
rect 104801 219267 104867 219270
rect 226333 219058 226399 219061
rect 226333 219056 230092 219058
rect 226333 219000 226338 219056
rect 226394 219000 230092 219056
rect 226333 218998 230092 219000
rect 226333 218995 226399 218998
rect 116393 218922 116459 218925
rect 213913 218922 213979 218925
rect 116393 218920 119692 218922
rect 116393 218864 116398 218920
rect 116454 218864 119692 218920
rect 116393 218862 119692 218864
rect 211508 218920 213979 218922
rect 211508 218864 213918 218920
rect 213974 218864 213979 218920
rect 211508 218862 213979 218864
rect 116393 218859 116459 218862
rect 213913 218859 213979 218862
rect 226425 218378 226491 218381
rect 226425 218376 230092 218378
rect 226425 218320 226430 218376
rect 226486 218320 230092 218376
rect 226425 218318 230092 218320
rect 226425 218315 226491 218318
rect 214005 218242 214071 218245
rect 211508 218240 214071 218242
rect 211508 218184 214010 218240
rect 214066 218184 214071 218240
rect 211508 218182 214071 218184
rect 214005 218179 214071 218182
rect 104801 217970 104867 217973
rect 101078 217968 104867 217970
rect 101078 217912 104806 217968
rect 104862 217912 104867 217968
rect 101078 217910 104867 217912
rect 101078 217872 101138 217910
rect 104801 217907 104867 217910
rect 226333 217834 226399 217837
rect 226333 217832 230092 217834
rect 226333 217776 226338 217832
rect 226394 217776 230092 217832
rect 226333 217774 230092 217776
rect 226333 217771 226399 217774
rect 116393 217698 116459 217701
rect 116393 217696 119692 217698
rect 116393 217640 116398 217696
rect 116454 217640 119692 217696
rect 116393 217638 119692 217640
rect 116393 217635 116459 217638
rect 213913 217426 213979 217429
rect 211508 217424 213979 217426
rect 211508 217368 213918 217424
rect 213974 217368 213979 217424
rect 211508 217366 213979 217368
rect 213913 217363 213979 217366
rect 226425 217290 226491 217293
rect 226425 217288 230092 217290
rect 226425 217232 226430 217288
rect 226486 217232 230092 217288
rect 226425 217230 230092 217232
rect 226425 217227 226491 217230
rect 580901 217018 580967 217021
rect 583520 217018 584960 217108
rect 580901 217016 584960 217018
rect 580901 216960 580906 217016
rect 580962 216960 584960 217016
rect 580901 216958 584960 216960
rect 580901 216955 580967 216958
rect 583520 216868 584960 216958
rect 101078 216610 101138 216648
rect 104801 216610 104867 216613
rect 101078 216608 104867 216610
rect 101078 216552 104806 216608
rect 104862 216552 104867 216608
rect 101078 216550 104867 216552
rect 104801 216547 104867 216550
rect 115933 216610 115999 216613
rect 213913 216610 213979 216613
rect 115933 216608 119692 216610
rect 115933 216552 115938 216608
rect 115994 216552 119692 216608
rect 115933 216550 119692 216552
rect 211508 216608 213979 216610
rect 211508 216552 213918 216608
rect 213974 216552 213979 216608
rect 211508 216550 213979 216552
rect 115933 216547 115999 216550
rect 213913 216547 213979 216550
rect 226333 216610 226399 216613
rect 226333 216608 230092 216610
rect 226333 216552 226338 216608
rect 226394 216552 230092 216608
rect 226333 216550 230092 216552
rect 226333 216547 226399 216550
rect 226425 216066 226491 216069
rect 226425 216064 230092 216066
rect 226425 216008 226430 216064
rect 226486 216008 230092 216064
rect 226425 216006 230092 216008
rect 226425 216003 226491 216006
rect 213913 215794 213979 215797
rect 211508 215792 213979 215794
rect 211508 215736 213918 215792
rect 213974 215736 213979 215792
rect 211508 215734 213979 215736
rect 213913 215731 213979 215734
rect 104801 215658 104867 215661
rect 101078 215656 104867 215658
rect 101078 215600 104806 215656
rect 104862 215600 104867 215656
rect 101078 215598 104867 215600
rect 101078 215424 101138 215598
rect 104801 215595 104867 215598
rect 226333 215522 226399 215525
rect 226333 215520 230092 215522
rect 226333 215464 226338 215520
rect 226394 215464 230092 215520
rect 226333 215462 230092 215464
rect 226333 215459 226399 215462
rect 116393 215386 116459 215389
rect 116393 215384 119692 215386
rect 116393 215328 116398 215384
rect 116454 215328 119692 215384
rect 116393 215326 119692 215328
rect 116393 215323 116459 215326
rect 213913 215114 213979 215117
rect 211508 215112 213979 215114
rect 211508 215056 213918 215112
rect 213974 215056 213979 215112
rect 211508 215054 213979 215056
rect 213913 215051 213979 215054
rect 226425 214842 226491 214845
rect 226425 214840 230092 214842
rect 226425 214784 226430 214840
rect 226486 214784 230092 214840
rect 226425 214782 230092 214784
rect 226425 214779 226491 214782
rect 104801 214706 104867 214709
rect 101078 214704 104867 214706
rect 101078 214648 104806 214704
rect 104862 214648 104867 214704
rect 101078 214646 104867 214648
rect 101078 214200 101138 214646
rect 104801 214643 104867 214646
rect 214005 214298 214071 214301
rect 211508 214296 214071 214298
rect 211508 214240 214010 214296
rect 214066 214240 214071 214296
rect 211508 214238 214071 214240
rect 214005 214235 214071 214238
rect 226333 214298 226399 214301
rect 226333 214296 230092 214298
rect 226333 214240 226338 214296
rect 226394 214240 230092 214296
rect 226333 214238 230092 214240
rect 226333 214235 226399 214238
rect 116393 214162 116459 214165
rect 116393 214160 119692 214162
rect 116393 214104 116398 214160
rect 116454 214104 119692 214160
rect 116393 214102 119692 214104
rect 116393 214099 116459 214102
rect 226425 213618 226491 213621
rect 226425 213616 230092 213618
rect 226425 213560 226430 213616
rect 226486 213560 230092 213616
rect 226425 213558 230092 213560
rect 226425 213555 226491 213558
rect 104801 213482 104867 213485
rect 213913 213482 213979 213485
rect 101078 213480 104867 213482
rect 101078 213424 104806 213480
rect 104862 213424 104867 213480
rect 101078 213422 104867 213424
rect 211508 213480 213979 213482
rect 211508 213424 213918 213480
rect 213974 213424 213979 213480
rect 211508 213422 213979 213424
rect 101078 212976 101138 213422
rect 104801 213419 104867 213422
rect 213913 213419 213979 213422
rect 115933 213074 115999 213077
rect 226333 213074 226399 213077
rect 115933 213072 119692 213074
rect 115933 213016 115938 213072
rect 115994 213016 119692 213072
rect 115933 213014 119692 213016
rect 226333 213072 230092 213074
rect 226333 213016 226338 213072
rect 226394 213016 230092 213072
rect 226333 213014 230092 213016
rect 115933 213011 115999 213014
rect 226333 213011 226399 213014
rect 214005 212666 214071 212669
rect 211508 212664 214071 212666
rect 211508 212608 214010 212664
rect 214066 212608 214071 212664
rect 211508 212606 214071 212608
rect 214005 212603 214071 212606
rect 226517 212530 226583 212533
rect 226517 212528 230092 212530
rect 226517 212472 226522 212528
rect 226578 212472 230092 212528
rect 226517 212470 230092 212472
rect 226517 212467 226583 212470
rect 104433 212122 104499 212125
rect 101078 212120 104499 212122
rect 101078 212064 104438 212120
rect 104494 212064 104499 212120
rect 101078 212062 104499 212064
rect 101078 211752 101138 212062
rect 104433 212059 104499 212062
rect 213913 211986 213979 211989
rect 211508 211984 213979 211986
rect 211508 211928 213918 211984
rect 213974 211928 213979 211984
rect 211508 211926 213979 211928
rect 213913 211923 213979 211926
rect 116301 211850 116367 211853
rect 226057 211850 226123 211853
rect 116301 211848 119692 211850
rect 116301 211792 116306 211848
rect 116362 211792 119692 211848
rect 116301 211790 119692 211792
rect 226057 211848 230092 211850
rect 226057 211792 226062 211848
rect 226118 211792 230092 211848
rect 226057 211790 230092 211792
rect 116301 211787 116367 211790
rect 226057 211787 226123 211790
rect 226241 211306 226307 211309
rect 226241 211304 230092 211306
rect 226241 211248 226246 211304
rect 226302 211248 230092 211304
rect 226241 211246 230092 211248
rect 226241 211243 226307 211246
rect 214005 211170 214071 211173
rect 211508 211168 214071 211170
rect 211508 211112 214010 211168
rect 214066 211112 214071 211168
rect 211508 211110 214071 211112
rect 214005 211107 214071 211110
rect 104801 210898 104867 210901
rect 101078 210896 104867 210898
rect 101078 210840 104806 210896
rect 104862 210840 104867 210896
rect 101078 210838 104867 210840
rect 101078 210528 101138 210838
rect 104801 210835 104867 210838
rect 116301 210762 116367 210765
rect 225965 210762 226031 210765
rect 116301 210760 119692 210762
rect 116301 210704 116306 210760
rect 116362 210704 119692 210760
rect 116301 210702 119692 210704
rect 225965 210760 230092 210762
rect 225965 210704 225970 210760
rect 226026 210704 230092 210760
rect 225965 210702 230092 210704
rect 116301 210699 116367 210702
rect 225965 210699 226031 210702
rect 213913 210354 213979 210357
rect 211508 210352 213979 210354
rect 211508 210296 213918 210352
rect 213974 210296 213979 210352
rect 211508 210294 213979 210296
rect 213913 210291 213979 210294
rect 226149 210082 226215 210085
rect 226149 210080 230092 210082
rect 226149 210024 226154 210080
rect 226210 210024 230092 210080
rect 226149 210022 230092 210024
rect 226149 210019 226215 210022
rect 104801 209538 104867 209541
rect 101078 209536 104867 209538
rect 101078 209480 104806 209536
rect 104862 209480 104867 209536
rect 101078 209478 104867 209480
rect 101078 209304 101138 209478
rect 104801 209475 104867 209478
rect 116025 209538 116091 209541
rect 213913 209538 213979 209541
rect 116025 209536 119692 209538
rect 116025 209480 116030 209536
rect 116086 209480 119692 209536
rect 116025 209478 119692 209480
rect 211508 209536 213979 209538
rect 211508 209480 213918 209536
rect 213974 209480 213979 209536
rect 211508 209478 213979 209480
rect 116025 209475 116091 209478
rect 213913 209475 213979 209478
rect 226057 209538 226123 209541
rect 226057 209536 230092 209538
rect 226057 209480 226062 209536
rect 226118 209480 230092 209536
rect 226057 209478 230092 209480
rect 226057 209475 226123 209478
rect 226241 208994 226307 208997
rect 226241 208992 230092 208994
rect 226241 208936 226246 208992
rect 226302 208936 230092 208992
rect 226241 208934 230092 208936
rect 226241 208931 226307 208934
rect 214005 208858 214071 208861
rect 211508 208856 214071 208858
rect 211508 208800 214010 208856
rect 214066 208800 214071 208856
rect 211508 208798 214071 208800
rect 214005 208795 214071 208798
rect 116393 208314 116459 208317
rect 116393 208312 119692 208314
rect -960 208028 480 208268
rect 116393 208256 116398 208312
rect 116454 208256 119692 208312
rect 116393 208254 119692 208256
rect 116393 208251 116459 208254
rect 104801 208178 104867 208181
rect 101078 208176 104867 208178
rect 101078 208120 104806 208176
rect 104862 208120 104867 208176
rect 101078 208118 104867 208120
rect 101078 208080 101138 208118
rect 104801 208115 104867 208118
rect 213913 208042 213979 208045
rect 211508 208040 213979 208042
rect 211508 207984 213918 208040
rect 213974 207984 213979 208040
rect 211508 207982 213979 207984
rect 213913 207979 213979 207982
rect 226149 208042 226215 208045
rect 230062 208042 230122 208284
rect 226149 208040 230122 208042
rect 226149 207984 226154 208040
rect 226210 207984 230122 208040
rect 226149 207982 230122 207984
rect 226149 207979 226215 207982
rect 225781 207770 225847 207773
rect 225781 207768 230092 207770
rect 225781 207712 225786 207768
rect 225842 207712 230092 207768
rect 225781 207710 230092 207712
rect 225781 207707 225847 207710
rect 116301 207226 116367 207229
rect 214005 207226 214071 207229
rect 116301 207224 119692 207226
rect 116301 207168 116306 207224
rect 116362 207168 119692 207224
rect 116301 207166 119692 207168
rect 211508 207224 214071 207226
rect 211508 207168 214010 207224
rect 214066 207168 214071 207224
rect 211508 207166 214071 207168
rect 116301 207163 116367 207166
rect 214005 207163 214071 207166
rect 225965 207226 226031 207229
rect 225965 207224 230092 207226
rect 225965 207168 225970 207224
rect 226026 207168 230092 207224
rect 225965 207166 230092 207168
rect 225965 207163 226031 207166
rect 104801 206954 104867 206957
rect 101078 206952 104867 206954
rect 101078 206896 104806 206952
rect 104862 206896 104867 206952
rect 101078 206894 104867 206896
rect 101078 206856 101138 206894
rect 104801 206891 104867 206894
rect 225873 206546 225939 206549
rect 225873 206544 230092 206546
rect 225873 206488 225878 206544
rect 225934 206488 230092 206544
rect 225873 206486 230092 206488
rect 225873 206483 225939 206486
rect 213913 206410 213979 206413
rect 211508 206408 213979 206410
rect 211508 206352 213918 206408
rect 213974 206352 213979 206408
rect 211508 206350 213979 206352
rect 213913 206347 213979 206350
rect 104709 206274 104775 206277
rect 101078 206272 104775 206274
rect 101078 206216 104714 206272
rect 104770 206216 104775 206272
rect 101078 206214 104775 206216
rect 101078 205632 101138 206214
rect 104709 206211 104775 206214
rect 115933 206002 115999 206005
rect 226241 206002 226307 206005
rect 115933 206000 119692 206002
rect 115933 205944 115938 206000
rect 115994 205944 119692 206000
rect 115933 205942 119692 205944
rect 226241 206000 230092 206002
rect 226241 205944 226246 206000
rect 226302 205944 230092 206000
rect 226241 205942 230092 205944
rect 115933 205939 115999 205942
rect 226241 205939 226307 205942
rect 214005 205730 214071 205733
rect 211508 205728 214071 205730
rect 211508 205672 214010 205728
rect 214066 205672 214071 205728
rect 211508 205670 214071 205672
rect 214005 205667 214071 205670
rect 225597 205322 225663 205325
rect 225597 205320 230092 205322
rect 225597 205264 225602 205320
rect 225658 205264 230092 205320
rect 225597 205262 230092 205264
rect 225597 205259 225663 205262
rect 583520 205172 584960 205412
rect 104801 205050 104867 205053
rect 101078 205048 104867 205050
rect 101078 204992 104806 205048
rect 104862 204992 104867 205048
rect 101078 204990 104867 204992
rect 101078 204408 101138 204990
rect 104801 204987 104867 204990
rect 116393 204914 116459 204917
rect 213913 204914 213979 204917
rect 116393 204912 119692 204914
rect 116393 204856 116398 204912
rect 116454 204856 119692 204912
rect 116393 204854 119692 204856
rect 211508 204912 213979 204914
rect 211508 204856 213918 204912
rect 213974 204856 213979 204912
rect 211508 204854 213979 204856
rect 116393 204851 116459 204854
rect 213913 204851 213979 204854
rect 225689 204778 225755 204781
rect 225689 204776 230092 204778
rect 225689 204720 225694 204776
rect 225750 204720 230092 204776
rect 225689 204718 230092 204720
rect 225689 204715 225755 204718
rect 226241 204234 226307 204237
rect 226241 204232 230092 204234
rect 226241 204176 226246 204232
rect 226302 204176 230092 204232
rect 226241 204174 230092 204176
rect 226241 204171 226307 204174
rect 213913 204098 213979 204101
rect 211508 204096 213979 204098
rect 211508 204040 213918 204096
rect 213974 204040 213979 204096
rect 211508 204038 213979 204040
rect 213913 204035 213979 204038
rect 104801 203690 104867 203693
rect 101078 203688 104867 203690
rect 101078 203632 104806 203688
rect 104862 203632 104867 203688
rect 101078 203630 104867 203632
rect 101078 203184 101138 203630
rect 104801 203627 104867 203630
rect 116301 203690 116367 203693
rect 116301 203688 119692 203690
rect 116301 203632 116306 203688
rect 116362 203632 119692 203688
rect 116301 203630 119692 203632
rect 116301 203627 116367 203630
rect 226057 203554 226123 203557
rect 226057 203552 230092 203554
rect 226057 203496 226062 203552
rect 226118 203496 230092 203552
rect 226057 203494 230092 203496
rect 226057 203491 226123 203494
rect 214005 203282 214071 203285
rect 211508 203280 214071 203282
rect 211508 203224 214010 203280
rect 214066 203224 214071 203280
rect 211508 203222 214071 203224
rect 214005 203219 214071 203222
rect 225965 203010 226031 203013
rect 225965 203008 230092 203010
rect 225965 202952 225970 203008
rect 226026 202952 230092 203008
rect 225965 202950 230092 202952
rect 225965 202947 226031 202950
rect 104801 202466 104867 202469
rect 101078 202464 104867 202466
rect 101078 202408 104806 202464
rect 104862 202408 104867 202464
rect 101078 202406 104867 202408
rect 101078 201960 101138 202406
rect 104801 202403 104867 202406
rect 116117 202466 116183 202469
rect 213913 202466 213979 202469
rect 116117 202464 119692 202466
rect 116117 202408 116122 202464
rect 116178 202408 119692 202464
rect 116117 202406 119692 202408
rect 211508 202464 213979 202466
rect 211508 202408 213918 202464
rect 213974 202408 213979 202464
rect 211508 202406 213979 202408
rect 116117 202403 116183 202406
rect 213913 202403 213979 202406
rect 225781 202466 225847 202469
rect 225781 202464 230092 202466
rect 225781 202408 225786 202464
rect 225842 202408 230092 202464
rect 225781 202406 230092 202408
rect 225781 202403 225847 202406
rect 214005 201786 214071 201789
rect 211508 201784 214071 201786
rect 211508 201728 214010 201784
rect 214066 201728 214071 201784
rect 211508 201726 214071 201728
rect 214005 201723 214071 201726
rect 226149 201786 226215 201789
rect 226149 201784 230092 201786
rect 226149 201728 226154 201784
rect 226210 201728 230092 201784
rect 226149 201726 230092 201728
rect 226149 201723 226215 201726
rect 116117 201378 116183 201381
rect 116117 201376 119692 201378
rect 116117 201320 116122 201376
rect 116178 201320 119692 201376
rect 116117 201318 119692 201320
rect 116117 201315 116183 201318
rect 226333 201242 226399 201245
rect 226333 201240 230092 201242
rect 226333 201184 226338 201240
rect 226394 201184 230092 201240
rect 226333 201182 230092 201184
rect 226333 201179 226399 201182
rect 104801 201106 104867 201109
rect 101078 201104 104867 201106
rect 101078 201048 104806 201104
rect 104862 201048 104867 201104
rect 101078 201046 104867 201048
rect 101078 200736 101138 201046
rect 104801 201043 104867 201046
rect 213913 200970 213979 200973
rect 211508 200968 213979 200970
rect 211508 200912 213918 200968
rect 213974 200912 213979 200968
rect 211508 200910 213979 200912
rect 213913 200907 213979 200910
rect 225873 200698 225939 200701
rect 225873 200696 230092 200698
rect 225873 200640 225878 200696
rect 225934 200640 230092 200696
rect 225873 200638 230092 200640
rect 225873 200635 225939 200638
rect 115933 200154 115999 200157
rect 214005 200154 214071 200157
rect 115933 200152 119692 200154
rect 115933 200096 115938 200152
rect 115994 200096 119692 200152
rect 115933 200094 119692 200096
rect 211508 200152 214071 200154
rect 211508 200096 214010 200152
rect 214066 200096 214071 200152
rect 211508 200094 214071 200096
rect 115933 200091 115999 200094
rect 214005 200091 214071 200094
rect 225689 200018 225755 200021
rect 225689 200016 230092 200018
rect 225689 199960 225694 200016
rect 225750 199960 230092 200016
rect 225689 199958 230092 199960
rect 225689 199955 225755 199958
rect 104801 199882 104867 199885
rect 101078 199880 104867 199882
rect 101078 199824 104806 199880
rect 104862 199824 104867 199880
rect 101078 199822 104867 199824
rect 101078 199512 101138 199822
rect 104801 199819 104867 199822
rect 226425 199474 226491 199477
rect 226425 199472 230092 199474
rect 226425 199416 226430 199472
rect 226486 199416 230092 199472
rect 226425 199414 230092 199416
rect 226425 199411 226491 199414
rect 213913 199338 213979 199341
rect 211508 199336 213979 199338
rect 211508 199280 213918 199336
rect 213974 199280 213979 199336
rect 211508 199278 213979 199280
rect 213913 199275 213979 199278
rect 115933 199066 115999 199069
rect 115933 199064 119692 199066
rect 115933 199008 115938 199064
rect 115994 199008 119692 199064
rect 115933 199006 119692 199008
rect 115933 199003 115999 199006
rect 226333 198930 226399 198933
rect 226333 198928 230092 198930
rect 226333 198872 226338 198928
rect 226394 198872 230092 198928
rect 226333 198870 230092 198872
rect 226333 198867 226399 198870
rect 213913 198658 213979 198661
rect 338113 198658 338179 198661
rect 211508 198656 213979 198658
rect 211508 198600 213918 198656
rect 213974 198600 213979 198656
rect 211508 198598 213979 198600
rect 336628 198656 338179 198658
rect 336628 198600 338118 198656
rect 338174 198600 338179 198656
rect 336628 198598 338179 198600
rect 213913 198595 213979 198598
rect 338113 198595 338179 198598
rect 104801 198522 104867 198525
rect 101078 198520 104867 198522
rect 101078 198464 104806 198520
rect 104862 198464 104867 198520
rect 101078 198462 104867 198464
rect 101078 198288 101138 198462
rect 104801 198459 104867 198462
rect 226425 198250 226491 198253
rect 226425 198248 230092 198250
rect 226425 198192 226430 198248
rect 226486 198192 230092 198248
rect 226425 198190 230092 198192
rect 226425 198187 226491 198190
rect 116117 197842 116183 197845
rect 214005 197842 214071 197845
rect 116117 197840 119692 197842
rect 116117 197784 116122 197840
rect 116178 197784 119692 197840
rect 116117 197782 119692 197784
rect 211508 197840 214071 197842
rect 211508 197784 214010 197840
rect 214066 197784 214071 197840
rect 211508 197782 214071 197784
rect 116117 197779 116183 197782
rect 214005 197779 214071 197782
rect 226333 197706 226399 197709
rect 226333 197704 230092 197706
rect 226333 197648 226338 197704
rect 226394 197648 230092 197704
rect 226333 197646 230092 197648
rect 226333 197643 226399 197646
rect 104801 197298 104867 197301
rect 101078 197296 104867 197298
rect 101078 197240 104806 197296
rect 104862 197240 104867 197296
rect 101078 197238 104867 197240
rect 101078 197200 101138 197238
rect 104801 197235 104867 197238
rect 213913 197026 213979 197029
rect 211508 197024 213979 197026
rect 211508 196968 213918 197024
rect 213974 196968 213979 197024
rect 211508 196966 213979 196968
rect 213913 196963 213979 196966
rect 226333 197026 226399 197029
rect 226333 197024 230092 197026
rect 226333 196968 226338 197024
rect 226394 196968 230092 197024
rect 226333 196966 230092 196968
rect 226333 196963 226399 196966
rect 116393 196754 116459 196757
rect 116393 196752 119692 196754
rect 116393 196696 116398 196752
rect 116454 196696 119692 196752
rect 116393 196694 119692 196696
rect 116393 196691 116459 196694
rect 104709 196618 104775 196621
rect 101078 196616 104775 196618
rect 101078 196560 104714 196616
rect 104770 196560 104775 196616
rect 101078 196558 104775 196560
rect 101078 195976 101138 196558
rect 104709 196555 104775 196558
rect 226701 196482 226767 196485
rect 226701 196480 230092 196482
rect 226701 196424 226706 196480
rect 226762 196424 230092 196480
rect 226701 196422 230092 196424
rect 226701 196419 226767 196422
rect 214005 196210 214071 196213
rect 211508 196208 214071 196210
rect 211508 196152 214010 196208
rect 214066 196152 214071 196208
rect 211508 196150 214071 196152
rect 214005 196147 214071 196150
rect 226517 195938 226583 195941
rect 226517 195936 230092 195938
rect 226517 195880 226522 195936
rect 226578 195880 230092 195936
rect 226517 195878 230092 195880
rect 226517 195875 226583 195878
rect 115933 195530 115999 195533
rect 213913 195530 213979 195533
rect 115933 195528 119692 195530
rect 115933 195472 115938 195528
rect 115994 195472 119692 195528
rect 115933 195470 119692 195472
rect 211508 195528 213979 195530
rect 211508 195472 213918 195528
rect 213974 195472 213979 195528
rect 211508 195470 213979 195472
rect 115933 195467 115999 195470
rect 213913 195467 213979 195470
rect 104801 195394 104867 195397
rect 101078 195392 104867 195394
rect 101078 195336 104806 195392
rect 104862 195336 104867 195392
rect 101078 195334 104867 195336
rect 101078 194752 101138 195334
rect 104801 195331 104867 195334
rect 226333 195258 226399 195261
rect 226333 195256 230092 195258
rect 226333 195200 226338 195256
rect 226394 195200 230092 195256
rect 226333 195198 230092 195200
rect 226333 195195 226399 195198
rect 214005 194714 214071 194717
rect 211508 194712 214071 194714
rect 211508 194656 214010 194712
rect 214066 194656 214071 194712
rect 211508 194654 214071 194656
rect 214005 194651 214071 194654
rect 226425 194714 226491 194717
rect 226425 194712 230092 194714
rect 226425 194656 226430 194712
rect 226486 194656 230092 194712
rect 226425 194654 230092 194656
rect 226425 194651 226491 194654
rect 116117 194306 116183 194309
rect 116117 194304 119692 194306
rect 116117 194248 116122 194304
rect 116178 194248 119692 194304
rect 116117 194246 119692 194248
rect 116117 194243 116183 194246
rect 226333 194170 226399 194173
rect 226333 194168 230092 194170
rect 226333 194112 226338 194168
rect 226394 194112 230092 194168
rect 226333 194110 230092 194112
rect 226333 194107 226399 194110
rect 104801 194034 104867 194037
rect 101078 194032 104867 194034
rect -960 193898 480 193988
rect 101078 193976 104806 194032
rect 104862 193976 104867 194032
rect 101078 193974 104867 193976
rect 2773 193898 2839 193901
rect -960 193896 2839 193898
rect -960 193840 2778 193896
rect 2834 193840 2839 193896
rect -960 193838 2839 193840
rect -960 193748 480 193838
rect 2773 193835 2839 193838
rect 101078 193528 101138 193974
rect 104801 193971 104867 193974
rect 213913 193898 213979 193901
rect 211508 193896 213979 193898
rect 211508 193840 213918 193896
rect 213974 193840 213979 193896
rect 211508 193838 213979 193840
rect 213913 193835 213979 193838
rect 226425 193490 226491 193493
rect 226425 193488 230092 193490
rect 226425 193432 226430 193488
rect 226486 193432 230092 193488
rect 583520 193476 584960 193716
rect 226425 193430 230092 193432
rect 226425 193427 226491 193430
rect 116393 193218 116459 193221
rect 116393 193216 119692 193218
rect 116393 193160 116398 193216
rect 116454 193160 119692 193216
rect 116393 193158 119692 193160
rect 116393 193155 116459 193158
rect 213913 193082 213979 193085
rect 211508 193080 213979 193082
rect 211508 193024 213918 193080
rect 213974 193024 213979 193080
rect 211508 193022 213979 193024
rect 213913 193019 213979 193022
rect 226425 192946 226491 192949
rect 226425 192944 230092 192946
rect 226425 192888 226430 192944
rect 226486 192888 230092 192944
rect 226425 192886 230092 192888
rect 226425 192883 226491 192886
rect 104433 192810 104499 192813
rect 101078 192808 104499 192810
rect 101078 192752 104438 192808
rect 104494 192752 104499 192808
rect 101078 192750 104499 192752
rect 101078 192304 101138 192750
rect 104433 192747 104499 192750
rect 214005 192402 214071 192405
rect 211508 192400 214071 192402
rect 211508 192344 214010 192400
rect 214066 192344 214071 192400
rect 211508 192342 214071 192344
rect 214005 192339 214071 192342
rect 226333 192402 226399 192405
rect 226333 192400 230092 192402
rect 226333 192344 226338 192400
rect 226394 192344 230092 192400
rect 226333 192342 230092 192344
rect 226333 192339 226399 192342
rect 116025 191994 116091 191997
rect 116025 191992 119692 191994
rect 116025 191936 116030 191992
rect 116086 191936 119692 191992
rect 116025 191934 119692 191936
rect 116025 191931 116091 191934
rect 226425 191722 226491 191725
rect 226425 191720 230092 191722
rect 226425 191664 226430 191720
rect 226486 191664 230092 191720
rect 226425 191662 230092 191664
rect 226425 191659 226491 191662
rect 213913 191586 213979 191589
rect 211508 191584 213979 191586
rect 211508 191528 213918 191584
rect 213974 191528 213979 191584
rect 211508 191526 213979 191528
rect 213913 191523 213979 191526
rect 104433 191450 104499 191453
rect 101078 191448 104499 191450
rect 101078 191392 104438 191448
rect 104494 191392 104499 191448
rect 101078 191390 104499 191392
rect 101078 191080 101138 191390
rect 104433 191387 104499 191390
rect 226517 191178 226583 191181
rect 226517 191176 230092 191178
rect 226517 191120 226522 191176
rect 226578 191120 230092 191176
rect 226517 191118 230092 191120
rect 226517 191115 226583 191118
rect 116485 190906 116551 190909
rect 116485 190904 119692 190906
rect 116485 190848 116490 190904
rect 116546 190848 119692 190904
rect 116485 190846 119692 190848
rect 116485 190843 116551 190846
rect 214005 190770 214071 190773
rect 211508 190768 214071 190770
rect 211508 190712 214010 190768
rect 214066 190712 214071 190768
rect 211508 190710 214071 190712
rect 214005 190707 214071 190710
rect 226333 190498 226399 190501
rect 226333 190496 230092 190498
rect 226333 190440 226338 190496
rect 226394 190440 230092 190496
rect 226333 190438 230092 190440
rect 226333 190435 226399 190438
rect 104709 190226 104775 190229
rect 101078 190224 104775 190226
rect 101078 190168 104714 190224
rect 104770 190168 104775 190224
rect 101078 190166 104775 190168
rect 101078 189856 101138 190166
rect 104709 190163 104775 190166
rect 213913 189954 213979 189957
rect 211508 189952 213979 189954
rect 211508 189896 213918 189952
rect 213974 189896 213979 189952
rect 211508 189894 213979 189896
rect 213913 189891 213979 189894
rect 226425 189954 226491 189957
rect 226425 189952 230092 189954
rect 226425 189896 226430 189952
rect 226486 189896 230092 189952
rect 226425 189894 230092 189896
rect 226425 189891 226491 189894
rect 116393 189682 116459 189685
rect 116393 189680 119692 189682
rect 116393 189624 116398 189680
rect 116454 189624 119692 189680
rect 116393 189622 119692 189624
rect 116393 189619 116459 189622
rect 226333 189410 226399 189413
rect 226333 189408 230092 189410
rect 226333 189352 226338 189408
rect 226394 189352 230092 189408
rect 226333 189350 230092 189352
rect 226333 189347 226399 189350
rect 214005 189274 214071 189277
rect 211508 189272 214071 189274
rect 211508 189216 214010 189272
rect 214066 189216 214071 189272
rect 211508 189214 214071 189216
rect 214005 189211 214071 189214
rect 104801 188866 104867 188869
rect 101078 188864 104867 188866
rect 101078 188808 104806 188864
rect 104862 188808 104867 188864
rect 101078 188806 104867 188808
rect 101078 188632 101138 188806
rect 104801 188803 104867 188806
rect 226333 188730 226399 188733
rect 226333 188728 230092 188730
rect 226333 188672 226338 188728
rect 226394 188672 230092 188728
rect 226333 188670 230092 188672
rect 226333 188667 226399 188670
rect 116393 188458 116459 188461
rect 213913 188458 213979 188461
rect 116393 188456 119692 188458
rect 116393 188400 116398 188456
rect 116454 188400 119692 188456
rect 116393 188398 119692 188400
rect 211508 188456 213979 188458
rect 211508 188400 213918 188456
rect 213974 188400 213979 188456
rect 211508 188398 213979 188400
rect 116393 188395 116459 188398
rect 213913 188395 213979 188398
rect 226425 188186 226491 188189
rect 226425 188184 230092 188186
rect 226425 188128 226430 188184
rect 226486 188128 230092 188184
rect 226425 188126 230092 188128
rect 226425 188123 226491 188126
rect 214189 187642 214255 187645
rect 211508 187640 214255 187642
rect 211508 187584 214194 187640
rect 214250 187584 214255 187640
rect 211508 187582 214255 187584
rect 214189 187579 214255 187582
rect 227069 187642 227135 187645
rect 227069 187640 230092 187642
rect 227069 187584 227074 187640
rect 227130 187584 230092 187640
rect 227069 187582 230092 187584
rect 227069 187579 227135 187582
rect 104801 187506 104867 187509
rect 101078 187504 104867 187506
rect 101078 187448 104806 187504
rect 104862 187448 104867 187504
rect 101078 187446 104867 187448
rect 101078 187408 101138 187446
rect 104801 187443 104867 187446
rect 115933 187370 115999 187373
rect 115933 187368 119692 187370
rect 115933 187312 115938 187368
rect 115994 187312 119692 187368
rect 115933 187310 119692 187312
rect 115933 187307 115999 187310
rect 226333 186962 226399 186965
rect 226333 186960 230092 186962
rect 226333 186904 226338 186960
rect 226394 186904 230092 186960
rect 226333 186902 230092 186904
rect 226333 186899 226399 186902
rect 213913 186826 213979 186829
rect 211508 186824 213979 186826
rect 211508 186768 213918 186824
rect 213974 186768 213979 186824
rect 211508 186766 213979 186768
rect 213913 186763 213979 186766
rect 226425 186418 226491 186421
rect 226425 186416 230092 186418
rect 226425 186360 226430 186416
rect 226486 186360 230092 186416
rect 226425 186358 230092 186360
rect 226425 186355 226491 186358
rect 104801 186282 104867 186285
rect 101078 186280 104867 186282
rect 101078 186224 104806 186280
rect 104862 186224 104867 186280
rect 101078 186222 104867 186224
rect 101078 186184 101138 186222
rect 104801 186219 104867 186222
rect 116025 186146 116091 186149
rect 116025 186144 119692 186146
rect 116025 186088 116030 186144
rect 116086 186088 119692 186144
rect 116025 186086 119692 186088
rect 116025 186083 116091 186086
rect 214465 186010 214531 186013
rect 211508 186008 214531 186010
rect 211508 185952 214470 186008
rect 214526 185952 214531 186008
rect 211508 185950 214531 185952
rect 214465 185947 214531 185950
rect 226333 185874 226399 185877
rect 226333 185872 230092 185874
rect 226333 185816 226338 185872
rect 226394 185816 230092 185872
rect 226333 185814 230092 185816
rect 226333 185811 226399 185814
rect 104709 185602 104775 185605
rect 101078 185600 104775 185602
rect 101078 185544 104714 185600
rect 104770 185544 104775 185600
rect 101078 185542 104775 185544
rect 101078 184960 101138 185542
rect 104709 185539 104775 185542
rect 213913 185330 213979 185333
rect 211508 185328 213979 185330
rect 211508 185272 213918 185328
rect 213974 185272 213979 185328
rect 211508 185270 213979 185272
rect 213913 185267 213979 185270
rect 226425 185194 226491 185197
rect 226425 185192 230092 185194
rect 226425 185136 226430 185192
rect 226486 185136 230092 185192
rect 226425 185134 230092 185136
rect 226425 185131 226491 185134
rect 116393 185058 116459 185061
rect 116393 185056 119692 185058
rect 116393 185000 116398 185056
rect 116454 185000 119692 185056
rect 116393 184998 119692 185000
rect 116393 184995 116459 184998
rect 226333 184650 226399 184653
rect 226333 184648 230092 184650
rect 226333 184592 226338 184648
rect 226394 184592 230092 184648
rect 226333 184590 230092 184592
rect 226333 184587 226399 184590
rect 214097 184514 214163 184517
rect 211508 184512 214163 184514
rect 211508 184456 214102 184512
rect 214158 184456 214163 184512
rect 211508 184454 214163 184456
rect 214097 184451 214163 184454
rect 104801 184378 104867 184381
rect 101078 184376 104867 184378
rect 101078 184320 104806 184376
rect 104862 184320 104867 184376
rect 101078 184318 104867 184320
rect 101078 183736 101138 184318
rect 104801 184315 104867 184318
rect 226977 184106 227043 184109
rect 226977 184104 230092 184106
rect 226977 184048 226982 184104
rect 227038 184048 230092 184104
rect 226977 184046 230092 184048
rect 226977 184043 227043 184046
rect 116393 183834 116459 183837
rect 116393 183832 119692 183834
rect 116393 183776 116398 183832
rect 116454 183776 119692 183832
rect 116393 183774 119692 183776
rect 116393 183771 116459 183774
rect 215201 183698 215267 183701
rect 211508 183696 215267 183698
rect 211508 183640 215206 183696
rect 215262 183640 215267 183696
rect 211508 183638 215267 183640
rect 215201 183635 215267 183638
rect 226425 183426 226491 183429
rect 226425 183424 230092 183426
rect 226425 183368 226430 183424
rect 226486 183368 230092 183424
rect 226425 183366 230092 183368
rect 226425 183363 226491 183366
rect 104801 183018 104867 183021
rect 101078 183016 104867 183018
rect 101078 182960 104806 183016
rect 104862 182960 104867 183016
rect 101078 182958 104867 182960
rect 101078 182512 101138 182958
rect 104801 182955 104867 182958
rect 215017 182882 215083 182885
rect 211508 182880 215083 182882
rect 211508 182824 215022 182880
rect 215078 182824 215083 182880
rect 211508 182822 215083 182824
rect 215017 182819 215083 182822
rect 225689 182882 225755 182885
rect 225689 182880 230092 182882
rect 225689 182824 225694 182880
rect 225750 182824 230092 182880
rect 225689 182822 230092 182824
rect 225689 182819 225755 182822
rect 115933 182610 115999 182613
rect 115933 182608 119692 182610
rect 115933 182552 115938 182608
rect 115994 182552 119692 182608
rect 115933 182550 119692 182552
rect 115933 182547 115999 182550
rect 215201 182202 215267 182205
rect 211508 182200 215267 182202
rect 211508 182144 215206 182200
rect 215262 182144 215267 182200
rect 211508 182142 215267 182144
rect 215201 182139 215267 182142
rect 226333 182202 226399 182205
rect 226333 182200 230092 182202
rect 226333 182144 226338 182200
rect 226394 182144 230092 182200
rect 226333 182142 230092 182144
rect 226333 182139 226399 182142
rect 214281 181930 214347 181933
rect 211478 181928 214347 181930
rect 211478 181872 214286 181928
rect 214342 181872 214347 181928
rect 211478 181870 214347 181872
rect 104801 181794 104867 181797
rect 101078 181792 104867 181794
rect 101078 181736 104806 181792
rect 104862 181736 104867 181792
rect 101078 181734 104867 181736
rect 101078 181288 101138 181734
rect 104801 181731 104867 181734
rect 115933 181522 115999 181525
rect 115933 181520 119692 181522
rect 115933 181464 115938 181520
rect 115994 181464 119692 181520
rect 115933 181462 119692 181464
rect 115933 181459 115999 181462
rect 211478 181356 211538 181870
rect 214281 181867 214347 181870
rect 579981 181930 580047 181933
rect 583520 181930 584960 182020
rect 579981 181928 584960 181930
rect 579981 181872 579986 181928
rect 580042 181872 584960 181928
rect 579981 181870 584960 181872
rect 579981 181867 580047 181870
rect 583520 181780 584960 181870
rect 226333 181658 226399 181661
rect 226333 181656 230092 181658
rect 226333 181600 226338 181656
rect 226394 181600 230092 181656
rect 226333 181598 230092 181600
rect 226333 181595 226399 181598
rect 226333 181114 226399 181117
rect 226333 181112 230092 181114
rect 226333 181056 226338 181112
rect 226394 181056 230092 181112
rect 226333 181054 230092 181056
rect 226333 181051 226399 181054
rect 213913 180570 213979 180573
rect 211508 180568 213979 180570
rect 211508 180512 213918 180568
rect 213974 180512 213979 180568
rect 211508 180510 213979 180512
rect 213913 180507 213979 180510
rect 104801 180434 104867 180437
rect 101078 180432 104867 180434
rect 101078 180376 104806 180432
rect 104862 180376 104867 180432
rect 101078 180374 104867 180376
rect 101078 180064 101138 180374
rect 104801 180371 104867 180374
rect 226425 180434 226491 180437
rect 226425 180432 230092 180434
rect 226425 180376 226430 180432
rect 226486 180376 230092 180432
rect 226425 180374 230092 180376
rect 226425 180371 226491 180374
rect 116393 180298 116459 180301
rect 116393 180296 119692 180298
rect 116393 180240 116398 180296
rect 116454 180240 119692 180296
rect 116393 180238 119692 180240
rect 116393 180235 116459 180238
rect 226333 179890 226399 179893
rect 226333 179888 230092 179890
rect 226333 179832 226338 179888
rect 226394 179832 230092 179888
rect 226333 179830 230092 179832
rect 226333 179827 226399 179830
rect 214373 179754 214439 179757
rect 211508 179752 214439 179754
rect 211508 179696 214378 179752
rect 214434 179696 214439 179752
rect 211508 179694 214439 179696
rect 214373 179691 214439 179694
rect -960 179482 480 179572
rect 2773 179482 2839 179485
rect -960 179480 2839 179482
rect -960 179424 2778 179480
rect 2834 179424 2839 179480
rect -960 179422 2839 179424
rect -960 179332 480 179422
rect 2773 179419 2839 179422
rect 226333 179346 226399 179349
rect 226333 179344 230092 179346
rect 226333 179288 226338 179344
rect 226394 179288 230092 179344
rect 226333 179286 230092 179288
rect 226333 179283 226399 179286
rect 115933 179210 115999 179213
rect 115933 179208 119692 179210
rect 115933 179152 115938 179208
rect 115994 179152 119692 179208
rect 115933 179150 119692 179152
rect 115933 179147 115999 179150
rect 104801 179074 104867 179077
rect 213913 179074 213979 179077
rect 101078 179072 104867 179074
rect 101078 179016 104806 179072
rect 104862 179016 104867 179072
rect 101078 179014 104867 179016
rect 211508 179072 213979 179074
rect 211508 179016 213918 179072
rect 213974 179016 213979 179072
rect 211508 179014 213979 179016
rect 101078 178840 101138 179014
rect 104801 179011 104867 179014
rect 213913 179011 213979 179014
rect 226425 178666 226491 178669
rect 226425 178664 230092 178666
rect 226425 178608 226430 178664
rect 226486 178608 230092 178664
rect 226425 178606 230092 178608
rect 226425 178603 226491 178606
rect 214005 178258 214071 178261
rect 211508 178256 214071 178258
rect 211508 178200 214010 178256
rect 214066 178200 214071 178256
rect 211508 178198 214071 178200
rect 214005 178195 214071 178198
rect 225597 178122 225663 178125
rect 225597 178120 230092 178122
rect 225597 178064 225602 178120
rect 225658 178064 230092 178120
rect 225597 178062 230092 178064
rect 225597 178059 225663 178062
rect 115933 177986 115999 177989
rect 115933 177984 119692 177986
rect 115933 177928 115938 177984
rect 115994 177928 119692 177984
rect 115933 177926 119692 177928
rect 115933 177923 115999 177926
rect 104157 177850 104223 177853
rect 101078 177848 104223 177850
rect 101078 177792 104162 177848
rect 104218 177792 104223 177848
rect 101078 177790 104223 177792
rect 101078 177616 101138 177790
rect 104157 177787 104223 177790
rect 226333 177578 226399 177581
rect 226333 177576 230092 177578
rect 226333 177520 226338 177576
rect 226394 177520 230092 177576
rect 226333 177518 230092 177520
rect 226333 177515 226399 177518
rect 213913 177442 213979 177445
rect 211508 177440 213979 177442
rect 211508 177384 213918 177440
rect 213974 177384 213979 177440
rect 211508 177382 213979 177384
rect 213913 177379 213979 177382
rect 116393 176898 116459 176901
rect 226425 176898 226491 176901
rect 116393 176896 119692 176898
rect 116393 176840 116398 176896
rect 116454 176840 119692 176896
rect 116393 176838 119692 176840
rect 226425 176896 230092 176898
rect 226425 176840 226430 176896
rect 226486 176840 230092 176896
rect 226425 176838 230092 176840
rect 116393 176835 116459 176838
rect 226425 176835 226491 176838
rect 214281 176626 214347 176629
rect 211508 176624 214347 176626
rect 211508 176568 214286 176624
rect 214342 176568 214347 176624
rect 211508 176566 214347 176568
rect 214281 176563 214347 176566
rect 104157 176490 104223 176493
rect 101078 176488 104223 176490
rect 101078 176432 104162 176488
rect 104218 176432 104223 176488
rect 101078 176430 104223 176432
rect 101078 176392 101138 176430
rect 104157 176427 104223 176430
rect 226885 176354 226951 176357
rect 226885 176352 230092 176354
rect 226885 176296 226890 176352
rect 226946 176296 230092 176352
rect 226885 176294 230092 176296
rect 226885 176291 226951 176294
rect 214005 175946 214071 175949
rect 211508 175944 214071 175946
rect 211508 175888 214010 175944
rect 214066 175888 214071 175944
rect 211508 175886 214071 175888
rect 214005 175883 214071 175886
rect 227437 175810 227503 175813
rect 227437 175808 230092 175810
rect 227437 175752 227442 175808
rect 227498 175752 230092 175808
rect 227437 175750 230092 175752
rect 227437 175747 227503 175750
rect 116393 175674 116459 175677
rect 116393 175672 119692 175674
rect 116393 175616 116398 175672
rect 116454 175616 119692 175672
rect 116393 175614 119692 175616
rect 116393 175611 116459 175614
rect 104801 175266 104867 175269
rect 101078 175264 104867 175266
rect 101078 175208 104806 175264
rect 104862 175208 104867 175264
rect 101078 175206 104867 175208
rect 101078 175168 101138 175206
rect 104801 175203 104867 175206
rect 214189 175130 214255 175133
rect 211508 175128 214255 175130
rect 211508 175072 214194 175128
rect 214250 175072 214255 175128
rect 211508 175070 214255 175072
rect 214189 175067 214255 175070
rect 104525 174586 104591 174589
rect 101078 174584 104591 174586
rect 101078 174528 104530 174584
rect 104586 174528 104591 174584
rect 101078 174526 104591 174528
rect 101078 174080 101138 174526
rect 104525 174523 104591 174526
rect 115933 174450 115999 174453
rect 115933 174448 119692 174450
rect 115933 174392 115938 174448
rect 115994 174392 119692 174448
rect 115933 174390 119692 174392
rect 115933 174387 115999 174390
rect 213913 174314 213979 174317
rect 211508 174312 213979 174314
rect 211508 174256 213918 174312
rect 213974 174256 213979 174312
rect 211508 174254 213979 174256
rect 213913 174251 213979 174254
rect 214189 173906 214255 173909
rect 214465 173906 214531 173909
rect 214189 173904 214531 173906
rect 214189 173848 214194 173904
rect 214250 173848 214470 173904
rect 214526 173848 214531 173904
rect 214189 173846 214531 173848
rect 214189 173843 214255 173846
rect 214465 173843 214531 173846
rect 283373 173906 283439 173909
rect 332910 173906 332916 173908
rect 283373 173904 332916 173906
rect 283373 173848 283378 173904
rect 283434 173848 332916 173904
rect 283373 173846 332916 173848
rect 283373 173843 283439 173846
rect 332910 173844 332916 173846
rect 332980 173844 332986 173908
rect 4797 173770 4863 173773
rect 4797 173768 9322 173770
rect 4797 173712 4802 173768
rect 4858 173712 9322 173768
rect 4797 173710 9322 173712
rect 4797 173707 4863 173710
rect 9262 173536 9322 173710
rect 214005 173498 214071 173501
rect 211508 173496 214071 173498
rect 211508 173440 214010 173496
rect 214066 173440 214071 173496
rect 211508 173438 214071 173440
rect 214005 173435 214071 173438
rect 104801 173362 104867 173365
rect 101078 173360 104867 173362
rect 101078 173304 104806 173360
rect 104862 173304 104867 173360
rect 101078 173302 104867 173304
rect 101078 172856 101138 173302
rect 104801 173299 104867 173302
rect 116393 173362 116459 173365
rect 116393 173360 119692 173362
rect 116393 173304 116398 173360
rect 116454 173304 119692 173360
rect 116393 173302 119692 173304
rect 116393 173299 116459 173302
rect 232221 173226 232287 173229
rect 283373 173226 283439 173229
rect 232221 173224 283439 173226
rect 232221 173168 232226 173224
rect 232282 173168 283378 173224
rect 283434 173168 283439 173224
rect 232221 173166 283439 173168
rect 232221 173163 232287 173166
rect 283373 173163 283439 173166
rect 213913 172818 213979 172821
rect 211508 172816 213979 172818
rect 211508 172760 213918 172816
rect 213974 172760 213979 172816
rect 211508 172758 213979 172760
rect 213913 172755 213979 172758
rect 104433 172138 104499 172141
rect 101078 172136 104499 172138
rect 101078 172080 104438 172136
rect 104494 172080 104499 172136
rect 101078 172078 104499 172080
rect 101078 171632 101138 172078
rect 104433 172075 104499 172078
rect 116117 172138 116183 172141
rect 116117 172136 119692 172138
rect 116117 172080 116122 172136
rect 116178 172080 119692 172136
rect 116117 172078 119692 172080
rect 116117 172075 116183 172078
rect 214373 172002 214439 172005
rect 211508 172000 214439 172002
rect 211508 171944 214378 172000
rect 214434 171944 214439 172000
rect 211508 171942 214439 171944
rect 214373 171939 214439 171942
rect 213913 171186 213979 171189
rect 211508 171184 213979 171186
rect 211508 171128 213918 171184
rect 213974 171128 213979 171184
rect 211508 171126 213979 171128
rect 213913 171123 213979 171126
rect 116301 171050 116367 171053
rect 116301 171048 119692 171050
rect 116301 170992 116306 171048
rect 116362 170992 119692 171048
rect 116301 170990 119692 170992
rect 116301 170987 116367 170990
rect 104801 170778 104867 170781
rect 101078 170776 104867 170778
rect 101078 170720 104806 170776
rect 104862 170720 104867 170776
rect 101078 170718 104867 170720
rect 101078 170408 101138 170718
rect 104801 170715 104867 170718
rect 215017 170370 215083 170373
rect 211508 170368 215083 170370
rect 211508 170312 215022 170368
rect 215078 170312 215083 170368
rect 211508 170310 215083 170312
rect 215017 170307 215083 170310
rect 580901 170098 580967 170101
rect 583520 170098 584960 170188
rect 580901 170096 584960 170098
rect 580901 170040 580906 170096
rect 580962 170040 584960 170096
rect 580901 170038 584960 170040
rect 580901 170035 580967 170038
rect 583520 169948 584960 170038
rect 116393 169826 116459 169829
rect 116393 169824 119692 169826
rect 116393 169768 116398 169824
rect 116454 169768 119692 169824
rect 116393 169766 119692 169768
rect 116393 169763 116459 169766
rect 213913 169554 213979 169557
rect 211508 169552 213979 169554
rect 211508 169496 213918 169552
rect 213974 169496 213979 169552
rect 211508 169494 213979 169496
rect 213913 169491 213979 169494
rect 104801 169418 104867 169421
rect 101078 169416 104867 169418
rect 101078 169360 104806 169416
rect 104862 169360 104867 169416
rect 101078 169358 104867 169360
rect 101078 169184 101138 169358
rect 104801 169355 104867 169358
rect 215109 168874 215175 168877
rect 211508 168872 215175 168874
rect 211508 168816 215114 168872
rect 215170 168816 215175 168872
rect 211508 168814 215175 168816
rect 215109 168811 215175 168814
rect 116393 168602 116459 168605
rect 116393 168600 119692 168602
rect 116393 168544 116398 168600
rect 116454 168544 119692 168600
rect 116393 168542 119692 168544
rect 116393 168539 116459 168542
rect 104157 168194 104223 168197
rect 101078 168192 104223 168194
rect 101078 168136 104162 168192
rect 104218 168136 104223 168192
rect 101078 168134 104223 168136
rect 101078 167960 101138 168134
rect 104157 168131 104223 168134
rect 213913 168058 213979 168061
rect 211508 168056 213979 168058
rect 211508 168000 213918 168056
rect 213974 168000 213979 168056
rect 211508 167998 213979 168000
rect 213913 167995 213979 167998
rect 115933 167514 115999 167517
rect 115933 167512 119692 167514
rect 115933 167456 115938 167512
rect 115994 167456 119692 167512
rect 115933 167454 119692 167456
rect 115933 167451 115999 167454
rect 214833 167242 214899 167245
rect 211508 167240 214899 167242
rect 211508 167184 214838 167240
rect 214894 167184 214899 167240
rect 211508 167182 214899 167184
rect 214833 167179 214899 167182
rect 104249 166970 104315 166973
rect 101078 166968 104315 166970
rect 101078 166912 104254 166968
rect 104310 166912 104315 166968
rect 101078 166910 104315 166912
rect 101078 166736 101138 166910
rect 104249 166907 104315 166910
rect 213913 166426 213979 166429
rect 211508 166424 213979 166426
rect 211508 166368 213918 166424
rect 213974 166368 213979 166424
rect 211508 166366 213979 166368
rect 213913 166363 213979 166366
rect 115933 166290 115999 166293
rect 115933 166288 119692 166290
rect 115933 166232 115938 166288
rect 115994 166232 119692 166288
rect 115933 166230 119692 166232
rect 115933 166227 115999 166230
rect 214005 165746 214071 165749
rect 211508 165744 214071 165746
rect 211508 165688 214010 165744
rect 214066 165688 214071 165744
rect 211508 165686 214071 165688
rect 214005 165683 214071 165686
rect 104801 165610 104867 165613
rect 101078 165608 104867 165610
rect 101078 165552 104806 165608
rect 104862 165552 104867 165608
rect 101078 165550 104867 165552
rect 101078 165512 101138 165550
rect 104801 165547 104867 165550
rect 116117 165202 116183 165205
rect 116117 165200 119692 165202
rect -960 164916 480 165156
rect 116117 165144 116122 165200
rect 116178 165144 119692 165200
rect 116117 165142 119692 165144
rect 116117 165139 116183 165142
rect 104617 164930 104683 164933
rect 213913 164930 213979 164933
rect 101078 164928 104683 164930
rect 101078 164872 104622 164928
rect 104678 164872 104683 164928
rect 101078 164870 104683 164872
rect 211508 164928 213979 164930
rect 211508 164872 213918 164928
rect 213974 164872 213979 164928
rect 211508 164870 213979 164872
rect 101078 164288 101138 164870
rect 104617 164867 104683 164870
rect 213913 164867 213979 164870
rect 213913 164114 213979 164117
rect 211508 164112 213979 164114
rect 211508 164056 213918 164112
rect 213974 164056 213979 164112
rect 211508 164054 213979 164056
rect 213913 164051 213979 164054
rect 116393 163978 116459 163981
rect 116393 163976 119692 163978
rect 116393 163920 116398 163976
rect 116454 163920 119692 163976
rect 116393 163918 119692 163920
rect 116393 163915 116459 163918
rect 104801 163706 104867 163709
rect 101078 163704 104867 163706
rect 101078 163648 104806 163704
rect 104862 163648 104867 163704
rect 101078 163646 104867 163648
rect 101078 163064 101138 163646
rect 104801 163643 104867 163646
rect 213913 163298 213979 163301
rect 211508 163296 213979 163298
rect 211508 163240 213918 163296
rect 213974 163240 213979 163296
rect 211508 163238 213979 163240
rect 213913 163235 213979 163238
rect 116209 162754 116275 162757
rect 116209 162752 119692 162754
rect 116209 162696 116214 162752
rect 116270 162696 119692 162752
rect 116209 162694 119692 162696
rect 116209 162691 116275 162694
rect 213913 162618 213979 162621
rect 211508 162616 213979 162618
rect 211508 162560 213918 162616
rect 213974 162560 213979 162616
rect 211508 162558 213979 162560
rect 213913 162555 213979 162558
rect 104801 162346 104867 162349
rect 101078 162344 104867 162346
rect 101078 162288 104806 162344
rect 104862 162288 104867 162344
rect 101078 162286 104867 162288
rect 101078 161840 101138 162286
rect 104801 162283 104867 162286
rect 213913 161802 213979 161805
rect 211508 161800 213979 161802
rect 211508 161744 213918 161800
rect 213974 161744 213979 161800
rect 211508 161742 213979 161744
rect 213913 161739 213979 161742
rect 116393 161666 116459 161669
rect 116393 161664 119692 161666
rect 116393 161608 116398 161664
rect 116454 161608 119692 161664
rect 116393 161606 119692 161608
rect 116393 161603 116459 161606
rect 104801 160986 104867 160989
rect 213913 160986 213979 160989
rect 101078 160984 104867 160986
rect 101078 160928 104806 160984
rect 104862 160928 104867 160984
rect 101078 160926 104867 160928
rect 211508 160984 213979 160986
rect 211508 160928 213918 160984
rect 213974 160928 213979 160984
rect 211508 160926 213979 160928
rect 101078 160616 101138 160926
rect 104801 160923 104867 160926
rect 213913 160923 213979 160926
rect 116393 160442 116459 160445
rect 116393 160440 119692 160442
rect 116393 160384 116398 160440
rect 116454 160384 119692 160440
rect 116393 160382 119692 160384
rect 116393 160379 116459 160382
rect 213913 160170 213979 160173
rect 211508 160168 213979 160170
rect 211508 160112 213918 160168
rect 213974 160112 213979 160168
rect 211508 160110 213979 160112
rect 213913 160107 213979 160110
rect 104801 159762 104867 159765
rect 101078 159760 104867 159762
rect 101078 159704 104806 159760
rect 104862 159704 104867 159760
rect 101078 159702 104867 159704
rect 101078 159392 101138 159702
rect 104801 159699 104867 159702
rect 214414 159490 214420 159492
rect 211508 159430 214420 159490
rect 214414 159428 214420 159430
rect 214484 159428 214490 159492
rect 116393 159354 116459 159357
rect 116393 159352 119692 159354
rect 116393 159296 116398 159352
rect 116454 159296 119692 159352
rect 116393 159294 119692 159296
rect 116393 159291 116459 159294
rect 103697 158674 103763 158677
rect 214741 158674 214807 158677
rect 101078 158672 103763 158674
rect 101078 158616 103702 158672
rect 103758 158616 103763 158672
rect 101078 158614 103763 158616
rect 211508 158672 214807 158674
rect 211508 158616 214746 158672
rect 214802 158616 214807 158672
rect 211508 158614 214807 158616
rect 101078 158168 101138 158614
rect 103697 158611 103763 158614
rect 214741 158611 214807 158614
rect 583520 158252 584960 158492
rect 116393 158130 116459 158133
rect 116393 158128 119692 158130
rect 116393 158072 116398 158128
rect 116454 158072 119692 158128
rect 116393 158070 119692 158072
rect 116393 158067 116459 158070
rect 214925 157858 214991 157861
rect 211508 157856 214991 157858
rect 211508 157800 214930 157856
rect 214986 157800 214991 157856
rect 211508 157798 214991 157800
rect 214925 157795 214991 157798
rect 104249 157314 104315 157317
rect 101078 157312 104315 157314
rect 101078 157256 104254 157312
rect 104310 157256 104315 157312
rect 101078 157254 104315 157256
rect 101078 156944 101138 157254
rect 104249 157251 104315 157254
rect 116025 157042 116091 157045
rect 213913 157042 213979 157045
rect 116025 157040 119692 157042
rect 116025 156984 116030 157040
rect 116086 156984 119692 157040
rect 116025 156982 119692 156984
rect 211508 157040 213979 157042
rect 211508 156984 213918 157040
rect 213974 156984 213979 157040
rect 211508 156982 213979 156984
rect 116025 156979 116091 156982
rect 213913 156979 213979 156982
rect 214097 156362 214163 156365
rect 211508 156360 214163 156362
rect 211508 156304 214102 156360
rect 214158 156304 214163 156360
rect 211508 156302 214163 156304
rect 214097 156299 214163 156302
rect 104801 155954 104867 155957
rect 101078 155952 104867 155954
rect 101078 155896 104806 155952
rect 104862 155896 104867 155952
rect 101078 155894 104867 155896
rect 101078 155720 101138 155894
rect 104801 155891 104867 155894
rect 116025 155818 116091 155821
rect 116025 155816 119692 155818
rect 116025 155760 116030 155816
rect 116086 155760 119692 155816
rect 116025 155758 119692 155760
rect 116025 155755 116091 155758
rect 213913 155546 213979 155549
rect 211508 155544 213979 155546
rect 211508 155488 213918 155544
rect 213974 155488 213979 155544
rect 211508 155486 213979 155488
rect 213913 155483 213979 155486
rect 214925 154730 214991 154733
rect 211508 154728 214991 154730
rect 211508 154672 214930 154728
rect 214986 154672 214991 154728
rect 211508 154670 214991 154672
rect 214925 154667 214991 154670
rect 116393 154594 116459 154597
rect 232313 154594 232379 154597
rect 232497 154594 232563 154597
rect 116393 154592 119692 154594
rect 116393 154536 116398 154592
rect 116454 154536 119692 154592
rect 116393 154534 119692 154536
rect 232313 154592 232563 154594
rect 232313 154536 232318 154592
rect 232374 154536 232502 154592
rect 232558 154536 232563 154592
rect 232313 154534 232563 154536
rect 116393 154531 116459 154534
rect 232313 154531 232379 154534
rect 232497 154531 232563 154534
rect 101078 154458 101138 154496
rect 104341 154458 104407 154461
rect 101078 154456 104407 154458
rect 101078 154400 104346 154456
rect 104402 154400 104407 154456
rect 101078 154398 104407 154400
rect 104341 154395 104407 154398
rect 104617 153914 104683 153917
rect 214005 153914 214071 153917
rect 101078 153912 104683 153914
rect 101078 153856 104622 153912
rect 104678 153856 104683 153912
rect 101078 153854 104683 153856
rect 211508 153912 214071 153914
rect 211508 153856 214010 153912
rect 214066 153856 214071 153912
rect 211508 153854 214071 153856
rect 101078 153272 101138 153854
rect 104617 153851 104683 153854
rect 214005 153851 214071 153854
rect 115933 153506 115999 153509
rect 115933 153504 119692 153506
rect 115933 153448 115938 153504
rect 115994 153448 119692 153504
rect 115933 153446 119692 153448
rect 115933 153443 115999 153446
rect 213913 153234 213979 153237
rect 211508 153232 213979 153234
rect 211508 153176 213918 153232
rect 213974 153176 213979 153232
rect 211508 153174 213979 153176
rect 213913 153171 213979 153174
rect 104801 152690 104867 152693
rect 101078 152688 104867 152690
rect 101078 152632 104806 152688
rect 104862 152632 104867 152688
rect 101078 152630 104867 152632
rect 101078 152048 101138 152630
rect 104801 152627 104867 152630
rect 213913 152418 213979 152421
rect 211508 152416 213979 152418
rect 211508 152360 213918 152416
rect 213974 152360 213979 152416
rect 211508 152358 213979 152360
rect 213913 152355 213979 152358
rect 116393 152282 116459 152285
rect 116393 152280 119692 152282
rect 116393 152224 116398 152280
rect 116454 152224 119692 152280
rect 116393 152222 119692 152224
rect 116393 152219 116459 152222
rect 104249 151602 104315 151605
rect 213913 151602 213979 151605
rect 101078 151600 104315 151602
rect 101078 151544 104254 151600
rect 104310 151544 104315 151600
rect 101078 151542 104315 151544
rect 211508 151600 213979 151602
rect 211508 151544 213918 151600
rect 213974 151544 213979 151600
rect 211508 151542 213979 151544
rect 101078 150960 101138 151542
rect 104249 151539 104315 151542
rect 213913 151539 213979 151542
rect 116393 151194 116459 151197
rect 116393 151192 119692 151194
rect 116393 151136 116398 151192
rect 116454 151136 119692 151192
rect 116393 151134 119692 151136
rect 116393 151131 116459 151134
rect -960 150786 480 150876
rect 2773 150786 2839 150789
rect 213913 150786 213979 150789
rect -960 150784 2839 150786
rect -960 150728 2778 150784
rect 2834 150728 2839 150784
rect -960 150726 2839 150728
rect 211508 150784 213979 150786
rect 211508 150728 213918 150784
rect 213974 150728 213979 150784
rect 211508 150726 213979 150728
rect -960 150636 480 150726
rect 2773 150723 2839 150726
rect 213913 150723 213979 150726
rect 103789 150378 103855 150381
rect 101078 150376 103855 150378
rect 101078 150320 103794 150376
rect 103850 150320 103855 150376
rect 101078 150318 103855 150320
rect 101078 149736 101138 150318
rect 103789 150315 103855 150318
rect 116393 149970 116459 149973
rect 213913 149970 213979 149973
rect 116393 149968 119692 149970
rect 116393 149912 116398 149968
rect 116454 149912 119692 149968
rect 116393 149910 119692 149912
rect 211508 149968 213979 149970
rect 211508 149912 213918 149968
rect 213974 149912 213979 149968
rect 211508 149910 213979 149912
rect 116393 149907 116459 149910
rect 213913 149907 213979 149910
rect 227437 149426 227503 149429
rect 227437 149424 230092 149426
rect 227437 149368 227442 149424
rect 227498 149368 230092 149424
rect 227437 149366 230092 149368
rect 227437 149363 227503 149366
rect 213913 149290 213979 149293
rect 211508 149288 213979 149290
rect 211508 149232 213918 149288
rect 213974 149232 213979 149288
rect 211508 149230 213979 149232
rect 213913 149227 213979 149230
rect 103697 149018 103763 149021
rect 101078 149016 103763 149018
rect 101078 148960 103702 149016
rect 103758 148960 103763 149016
rect 101078 148958 103763 148960
rect 101078 148512 101138 148958
rect 103697 148955 103763 148958
rect 227437 148882 227503 148885
rect 227437 148880 230092 148882
rect 227437 148824 227442 148880
rect 227498 148824 230092 148880
rect 227437 148822 230092 148824
rect 227437 148819 227503 148822
rect 116393 148746 116459 148749
rect 116393 148744 119692 148746
rect 116393 148688 116398 148744
rect 116454 148688 119692 148744
rect 116393 148686 119692 148688
rect 116393 148683 116459 148686
rect 213913 148474 213979 148477
rect 211508 148472 213979 148474
rect 211508 148416 213918 148472
rect 213974 148416 213979 148472
rect 211508 148414 213979 148416
rect 213913 148411 213979 148414
rect 227529 148202 227595 148205
rect 227529 148200 230092 148202
rect 227529 148144 227534 148200
rect 227590 148144 230092 148200
rect 227529 148142 230092 148144
rect 227529 148139 227595 148142
rect 104341 147658 104407 147661
rect 101078 147656 104407 147658
rect 101078 147600 104346 147656
rect 104402 147600 104407 147656
rect 101078 147598 104407 147600
rect 101078 147288 101138 147598
rect 104341 147595 104407 147598
rect 115933 147658 115999 147661
rect 214005 147658 214071 147661
rect 115933 147656 119692 147658
rect 115933 147600 115938 147656
rect 115994 147600 119692 147656
rect 115933 147598 119692 147600
rect 211508 147656 214071 147658
rect 211508 147600 214010 147656
rect 214066 147600 214071 147656
rect 211508 147598 214071 147600
rect 115933 147595 115999 147598
rect 214005 147595 214071 147598
rect 227437 147658 227503 147661
rect 227437 147656 230092 147658
rect 227437 147600 227442 147656
rect 227498 147600 230092 147656
rect 227437 147598 230092 147600
rect 227437 147595 227503 147598
rect 226977 146978 227043 146981
rect 226977 146976 230092 146978
rect 226977 146920 226982 146976
rect 227038 146920 230092 146976
rect 226977 146918 230092 146920
rect 226977 146915 227043 146918
rect 213913 146842 213979 146845
rect 211508 146840 213979 146842
rect 211508 146784 213918 146840
rect 213974 146784 213979 146840
rect 211508 146782 213979 146784
rect 213913 146779 213979 146782
rect 583520 146556 584960 146796
rect 116393 146434 116459 146437
rect 227529 146434 227595 146437
rect 116393 146432 119692 146434
rect 116393 146376 116398 146432
rect 116454 146376 119692 146432
rect 116393 146374 119692 146376
rect 227529 146432 230092 146434
rect 227529 146376 227534 146432
rect 227590 146376 230092 146432
rect 227529 146374 230092 146376
rect 116393 146371 116459 146374
rect 227529 146371 227595 146374
rect 104801 146298 104867 146301
rect 101078 146296 104867 146298
rect 101078 146240 104806 146296
rect 104862 146240 104867 146296
rect 101078 146238 104867 146240
rect 101078 146064 101138 146238
rect 104801 146235 104867 146238
rect 214005 146162 214071 146165
rect 211508 146160 214071 146162
rect 211508 146104 214010 146160
rect 214066 146104 214071 146160
rect 211508 146102 214071 146104
rect 214005 146099 214071 146102
rect 227437 145890 227503 145893
rect 227437 145888 230092 145890
rect 227437 145832 227442 145888
rect 227498 145832 230092 145888
rect 227437 145830 230092 145832
rect 227437 145827 227503 145830
rect 116025 145346 116091 145349
rect 213913 145346 213979 145349
rect 116025 145344 119692 145346
rect 116025 145288 116030 145344
rect 116086 145288 119692 145344
rect 116025 145286 119692 145288
rect 211508 145344 213979 145346
rect 211508 145288 213918 145344
rect 213974 145288 213979 145344
rect 211508 145286 213979 145288
rect 116025 145283 116091 145286
rect 213913 145283 213979 145286
rect 226701 145210 226767 145213
rect 226701 145208 230092 145210
rect 226701 145152 226706 145208
rect 226762 145152 230092 145208
rect 226701 145150 230092 145152
rect 226701 145147 226767 145150
rect 101078 144802 101138 144840
rect 104709 144802 104775 144805
rect 101078 144800 104775 144802
rect 101078 144744 104714 144800
rect 104770 144744 104775 144800
rect 101078 144742 104775 144744
rect 104709 144739 104775 144742
rect 227437 144666 227503 144669
rect 227437 144664 230092 144666
rect 227437 144608 227442 144664
rect 227498 144608 230092 144664
rect 227437 144606 230092 144608
rect 227437 144603 227503 144606
rect 214005 144530 214071 144533
rect 211508 144528 214071 144530
rect 211508 144472 214010 144528
rect 214066 144472 214071 144528
rect 211508 144470 214071 144472
rect 214005 144467 214071 144470
rect 104617 144258 104683 144261
rect 101078 144256 104683 144258
rect 101078 144200 104622 144256
rect 104678 144200 104683 144256
rect 101078 144198 104683 144200
rect 101078 143616 101138 144198
rect 104617 144195 104683 144198
rect 116393 144122 116459 144125
rect 116393 144120 119692 144122
rect 116393 144064 116398 144120
rect 116454 144064 119692 144120
rect 116393 144062 119692 144064
rect 116393 144059 116459 144062
rect 226517 143986 226583 143989
rect 226517 143984 230092 143986
rect 226517 143928 226522 143984
rect 226578 143928 230092 143984
rect 226517 143926 230092 143928
rect 226517 143923 226583 143926
rect 213913 143714 213979 143717
rect 211508 143712 213979 143714
rect 211508 143656 213918 143712
rect 213974 143656 213979 143712
rect 211508 143654 213979 143656
rect 213913 143651 213979 143654
rect 214557 143578 214623 143581
rect 214741 143578 214807 143581
rect 214557 143576 214807 143578
rect 214557 143520 214562 143576
rect 214618 143520 214746 143576
rect 214802 143520 214807 143576
rect 214557 143518 214807 143520
rect 214557 143515 214623 143518
rect 214741 143515 214807 143518
rect 227437 143442 227503 143445
rect 227437 143440 230092 143442
rect 227437 143384 227442 143440
rect 227498 143384 230092 143440
rect 227437 143382 230092 143384
rect 227437 143379 227503 143382
rect 104525 143034 104591 143037
rect 214005 143034 214071 143037
rect 101078 143032 104591 143034
rect 101078 142976 104530 143032
rect 104586 142976 104591 143032
rect 101078 142974 104591 142976
rect 211508 143032 214071 143034
rect 211508 142976 214010 143032
rect 214066 142976 214071 143032
rect 211508 142974 214071 142976
rect 101078 142392 101138 142974
rect 104525 142971 104591 142974
rect 214005 142971 214071 142974
rect 116393 142898 116459 142901
rect 226885 142898 226951 142901
rect 116393 142896 119692 142898
rect 116393 142840 116398 142896
rect 116454 142840 119692 142896
rect 116393 142838 119692 142840
rect 226885 142896 230092 142898
rect 226885 142840 226890 142896
rect 226946 142840 230092 142896
rect 226885 142838 230092 142840
rect 116393 142835 116459 142838
rect 226885 142835 226951 142838
rect 213913 142218 213979 142221
rect 211508 142216 213979 142218
rect 211508 142160 213918 142216
rect 213974 142160 213979 142216
rect 211508 142158 213979 142160
rect 213913 142155 213979 142158
rect 227621 142218 227687 142221
rect 227621 142216 230092 142218
rect 227621 142160 227626 142216
rect 227682 142160 230092 142216
rect 227621 142158 230092 142160
rect 227621 142155 227687 142158
rect 104157 141810 104223 141813
rect 101078 141808 104223 141810
rect 101078 141752 104162 141808
rect 104218 141752 104223 141808
rect 101078 141750 104223 141752
rect 101078 141168 101138 141750
rect 104157 141747 104223 141750
rect 116393 141810 116459 141813
rect 116393 141808 119692 141810
rect 116393 141752 116398 141808
rect 116454 141752 119692 141808
rect 116393 141750 119692 141752
rect 116393 141747 116459 141750
rect 226701 141674 226767 141677
rect 226701 141672 230092 141674
rect 226701 141616 226706 141672
rect 226762 141616 230092 141672
rect 226701 141614 230092 141616
rect 226701 141611 226767 141614
rect 213913 141402 213979 141405
rect 211508 141400 213979 141402
rect 211508 141344 213918 141400
rect 213974 141344 213979 141400
rect 211508 141342 213979 141344
rect 213913 141339 213979 141342
rect 227253 140994 227319 140997
rect 227253 140992 230092 140994
rect 227253 140936 227258 140992
rect 227314 140936 230092 140992
rect 227253 140934 230092 140936
rect 227253 140931 227319 140934
rect 103513 140586 103579 140589
rect 101078 140584 103579 140586
rect 101078 140528 103518 140584
rect 103574 140528 103579 140584
rect 101078 140526 103579 140528
rect 101078 139944 101138 140526
rect 103513 140523 103579 140526
rect 116393 140586 116459 140589
rect 214005 140586 214071 140589
rect 116393 140584 119692 140586
rect 116393 140528 116398 140584
rect 116454 140528 119692 140584
rect 116393 140526 119692 140528
rect 211508 140584 214071 140586
rect 211508 140528 214010 140584
rect 214066 140528 214071 140584
rect 211508 140526 214071 140528
rect 116393 140523 116459 140526
rect 214005 140523 214071 140526
rect 227069 140450 227135 140453
rect 227069 140448 230092 140450
rect 227069 140392 227074 140448
rect 227130 140392 230092 140448
rect 227069 140390 230092 140392
rect 227069 140387 227135 140390
rect 213913 139906 213979 139909
rect 211508 139904 213979 139906
rect 211508 139848 213918 139904
rect 213974 139848 213979 139904
rect 211508 139846 213979 139848
rect 213913 139843 213979 139846
rect 227529 139770 227595 139773
rect 227529 139768 230092 139770
rect 227529 139712 227534 139768
rect 227590 139712 230092 139768
rect 227529 139710 230092 139712
rect 227529 139707 227595 139710
rect 116301 139498 116367 139501
rect 116301 139496 119692 139498
rect 116301 139440 116306 139496
rect 116362 139440 119692 139496
rect 116301 139438 119692 139440
rect 116301 139435 116367 139438
rect 103697 139362 103763 139365
rect 101078 139360 103763 139362
rect 101078 139304 103702 139360
rect 103758 139304 103763 139360
rect 101078 139302 103763 139304
rect 101078 138720 101138 139302
rect 103697 139299 103763 139302
rect 227437 139226 227503 139229
rect 227437 139224 230092 139226
rect 227437 139168 227442 139224
rect 227498 139168 230092 139224
rect 227437 139166 230092 139168
rect 227437 139163 227503 139166
rect 214005 139090 214071 139093
rect 211508 139088 214071 139090
rect 211508 139032 214010 139088
rect 214066 139032 214071 139088
rect 211508 139030 214071 139032
rect 214005 139027 214071 139030
rect 227345 138682 227411 138685
rect 227345 138680 230092 138682
rect 227345 138624 227350 138680
rect 227406 138624 230092 138680
rect 227345 138622 230092 138624
rect 227345 138619 227411 138622
rect 115841 138274 115907 138277
rect 213913 138274 213979 138277
rect 115841 138272 119692 138274
rect 115841 138216 115846 138272
rect 115902 138216 119692 138272
rect 115841 138214 119692 138216
rect 211508 138272 213979 138274
rect 211508 138216 213918 138272
rect 213974 138216 213979 138272
rect 211508 138214 213979 138216
rect 115841 138211 115907 138214
rect 213913 138211 213979 138214
rect 104341 138002 104407 138005
rect 101078 138000 104407 138002
rect 101078 137944 104346 138000
rect 104402 137944 104407 138000
rect 101078 137942 104407 137944
rect 101078 137496 101138 137942
rect 104341 137939 104407 137942
rect 227437 138002 227503 138005
rect 227437 138000 230092 138002
rect 227437 137944 227442 138000
rect 227498 137944 230092 138000
rect 227437 137942 230092 137944
rect 227437 137939 227503 137942
rect 214005 137458 214071 137461
rect 211508 137456 214071 137458
rect 211508 137400 214010 137456
rect 214066 137400 214071 137456
rect 211508 137398 214071 137400
rect 214005 137395 214071 137398
rect 226701 137458 226767 137461
rect 226701 137456 230092 137458
rect 226701 137400 226706 137456
rect 226762 137400 230092 137456
rect 226701 137398 230092 137400
rect 226701 137395 226767 137398
rect 116393 137186 116459 137189
rect 116393 137184 119692 137186
rect 116393 137128 116398 137184
rect 116454 137128 119692 137184
rect 116393 137126 119692 137128
rect 116393 137123 116459 137126
rect 213913 136778 213979 136781
rect 211508 136776 213979 136778
rect 211508 136720 213918 136776
rect 213974 136720 213979 136776
rect 211508 136718 213979 136720
rect 213913 136715 213979 136718
rect 226517 136778 226583 136781
rect 226517 136776 230092 136778
rect 226517 136720 226522 136776
rect 226578 136720 230092 136776
rect 226517 136718 230092 136720
rect 226517 136715 226583 136718
rect 104801 136642 104867 136645
rect 101078 136640 104867 136642
rect 101078 136584 104806 136640
rect 104862 136584 104867 136640
rect 101078 136582 104867 136584
rect -960 136370 480 136460
rect 2773 136370 2839 136373
rect -960 136368 2839 136370
rect -960 136312 2778 136368
rect 2834 136312 2839 136368
rect -960 136310 2839 136312
rect -960 136220 480 136310
rect 2773 136307 2839 136310
rect 101078 136272 101138 136582
rect 104801 136579 104867 136582
rect 226609 136234 226675 136237
rect 226609 136232 230092 136234
rect 226609 136176 226614 136232
rect 226670 136176 230092 136232
rect 226609 136174 230092 136176
rect 226609 136171 226675 136174
rect 115933 135962 115999 135965
rect 213913 135962 213979 135965
rect 115933 135960 119692 135962
rect 115933 135904 115938 135960
rect 115994 135904 119692 135960
rect 115933 135902 119692 135904
rect 211508 135960 213979 135962
rect 211508 135904 213918 135960
rect 213974 135904 213979 135960
rect 211508 135902 213979 135904
rect 115933 135899 115999 135902
rect 213913 135899 213979 135902
rect 226425 135690 226491 135693
rect 226425 135688 230092 135690
rect 226425 135632 226430 135688
rect 226486 135632 230092 135688
rect 226425 135630 230092 135632
rect 226425 135627 226491 135630
rect 104801 135146 104867 135149
rect 214005 135146 214071 135149
rect 101078 135144 104867 135146
rect 101078 135088 104806 135144
rect 104862 135088 104867 135144
rect 101078 135086 104867 135088
rect 211508 135144 214071 135146
rect 211508 135088 214010 135144
rect 214066 135088 214071 135144
rect 211508 135086 214071 135088
rect 101078 135048 101138 135086
rect 104801 135083 104867 135086
rect 214005 135083 214071 135086
rect 226793 135010 226859 135013
rect 226793 135008 230092 135010
rect 226793 134952 226798 135008
rect 226854 134952 230092 135008
rect 226793 134950 230092 134952
rect 226793 134947 226859 134950
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 116393 134738 116459 134741
rect 116393 134736 119692 134738
rect 116393 134680 116398 134736
rect 116454 134680 119692 134736
rect 583520 134724 584960 134814
rect 116393 134678 119692 134680
rect 116393 134675 116459 134678
rect 227437 134466 227503 134469
rect 227437 134464 230092 134466
rect 227437 134408 227442 134464
rect 227498 134408 230092 134464
rect 227437 134406 230092 134408
rect 227437 134403 227503 134406
rect 213913 134330 213979 134333
rect 211508 134328 213979 134330
rect 211508 134272 213918 134328
rect 213974 134272 213979 134328
rect 211508 134270 213979 134272
rect 213913 134267 213979 134270
rect 101078 133786 101138 133824
rect 104801 133786 104867 133789
rect 101078 133784 104867 133786
rect 101078 133728 104806 133784
rect 104862 133728 104867 133784
rect 101078 133726 104867 133728
rect 104801 133723 104867 133726
rect 227069 133786 227135 133789
rect 227069 133784 230092 133786
rect 227069 133728 227074 133784
rect 227130 133728 230092 133784
rect 227069 133726 230092 133728
rect 227069 133723 227135 133726
rect 117129 133650 117195 133653
rect 117129 133648 119692 133650
rect 117129 133592 117134 133648
rect 117190 133592 119692 133648
rect 117129 133590 119692 133592
rect 117129 133587 117195 133590
rect 214005 133514 214071 133517
rect 211508 133512 214071 133514
rect 211508 133456 214010 133512
rect 214066 133456 214071 133512
rect 211508 133454 214071 133456
rect 214005 133451 214071 133454
rect 104709 133242 104775 133245
rect 101078 133240 104775 133242
rect 101078 133184 104714 133240
rect 104770 133184 104775 133240
rect 101078 133182 104775 133184
rect 101078 132600 101138 133182
rect 104709 133179 104775 133182
rect 227621 133242 227687 133245
rect 227621 133240 230092 133242
rect 227621 133184 227626 133240
rect 227682 133184 230092 133240
rect 227621 133182 230092 133184
rect 227621 133179 227687 133182
rect 213913 132834 213979 132837
rect 211508 132832 213979 132834
rect 211508 132776 213918 132832
rect 213974 132776 213979 132832
rect 211508 132774 213979 132776
rect 213913 132771 213979 132774
rect 227529 132562 227595 132565
rect 227529 132560 230092 132562
rect 227529 132504 227534 132560
rect 227590 132504 230092 132560
rect 227529 132502 230092 132504
rect 227529 132499 227595 132502
rect 116393 132426 116459 132429
rect 116393 132424 119692 132426
rect 116393 132368 116398 132424
rect 116454 132368 119692 132424
rect 116393 132366 119692 132368
rect 116393 132363 116459 132366
rect 104341 132018 104407 132021
rect 214005 132018 214071 132021
rect 101078 132016 104407 132018
rect 101078 131960 104346 132016
rect 104402 131960 104407 132016
rect 101078 131958 104407 131960
rect 211508 132016 214071 132018
rect 211508 131960 214010 132016
rect 214066 131960 214071 132016
rect 211508 131958 214071 131960
rect 101078 131376 101138 131958
rect 104341 131955 104407 131958
rect 214005 131955 214071 131958
rect 227345 132018 227411 132021
rect 227345 132016 230092 132018
rect 227345 131960 227350 132016
rect 227406 131960 230092 132016
rect 227345 131958 230092 131960
rect 227345 131955 227411 131958
rect 227437 131474 227503 131477
rect 227437 131472 230092 131474
rect 227437 131416 227442 131472
rect 227498 131416 230092 131472
rect 227437 131414 230092 131416
rect 227437 131411 227503 131414
rect 115933 131338 115999 131341
rect 115933 131336 119692 131338
rect 115933 131280 115938 131336
rect 115994 131280 119692 131336
rect 115933 131278 119692 131280
rect 115933 131275 115999 131278
rect 213913 131202 213979 131205
rect 211508 131200 213979 131202
rect 211508 131144 213918 131200
rect 213974 131144 213979 131200
rect 211508 131142 213979 131144
rect 213913 131139 213979 131142
rect 226701 130794 226767 130797
rect 226701 130792 230092 130794
rect 226701 130736 226706 130792
rect 226762 130736 230092 130792
rect 226701 130734 230092 130736
rect 226701 130731 226767 130734
rect 103973 130658 104039 130661
rect 101078 130656 104039 130658
rect 101078 130600 103978 130656
rect 104034 130600 104039 130656
rect 101078 130598 104039 130600
rect 101078 130152 101138 130598
rect 103973 130595 104039 130598
rect 213913 130386 213979 130389
rect 211508 130384 213979 130386
rect 211508 130328 213918 130384
rect 213974 130328 213979 130384
rect 211508 130326 213979 130328
rect 213913 130323 213979 130326
rect 227069 130250 227135 130253
rect 227069 130248 230092 130250
rect 227069 130192 227074 130248
rect 227130 130192 230092 130248
rect 227069 130190 230092 130192
rect 227069 130187 227135 130190
rect 116669 130114 116735 130117
rect 116669 130112 119692 130114
rect 116669 130056 116674 130112
rect 116730 130056 119692 130112
rect 116669 130054 119692 130056
rect 116669 130051 116735 130054
rect 213913 129706 213979 129709
rect 211508 129704 213979 129706
rect 211508 129648 213918 129704
rect 213974 129648 213979 129704
rect 211508 129646 213979 129648
rect 213913 129643 213979 129646
rect 226517 129570 226583 129573
rect 226517 129568 230092 129570
rect 226517 129512 226522 129568
rect 226578 129512 230092 129568
rect 226517 129510 230092 129512
rect 226517 129507 226583 129510
rect 104801 129298 104867 129301
rect 101078 129296 104867 129298
rect 101078 129240 104806 129296
rect 104862 129240 104867 129296
rect 101078 129238 104867 129240
rect 101078 128928 101138 129238
rect 104801 129235 104867 129238
rect 227529 129026 227595 129029
rect 227529 129024 230092 129026
rect 227529 128968 227534 129024
rect 227590 128968 230092 129024
rect 227529 128966 230092 128968
rect 227529 128963 227595 128966
rect 116393 128890 116459 128893
rect 213913 128890 213979 128893
rect 116393 128888 119692 128890
rect 116393 128832 116398 128888
rect 116454 128832 119692 128888
rect 116393 128830 119692 128832
rect 211508 128888 213979 128890
rect 211508 128832 213918 128888
rect 213974 128832 213979 128888
rect 211508 128830 213979 128832
rect 116393 128827 116459 128830
rect 213913 128827 213979 128830
rect 227437 128482 227503 128485
rect 227437 128480 230092 128482
rect 227437 128424 227442 128480
rect 227498 128424 230092 128480
rect 227437 128422 230092 128424
rect 227437 128419 227503 128422
rect 104801 128074 104867 128077
rect 213913 128074 213979 128077
rect 101078 128072 104867 128074
rect 101078 128016 104806 128072
rect 104862 128016 104867 128072
rect 101078 128014 104867 128016
rect 211508 128072 213979 128074
rect 211508 128016 213918 128072
rect 213974 128016 213979 128072
rect 211508 128014 213979 128016
rect 101078 127840 101138 128014
rect 104801 128011 104867 128014
rect 213913 128011 213979 128014
rect 116393 127802 116459 127805
rect 226333 127802 226399 127805
rect 116393 127800 119692 127802
rect 116393 127744 116398 127800
rect 116454 127744 119692 127800
rect 116393 127742 119692 127744
rect 226333 127800 230092 127802
rect 226333 127744 226338 127800
rect 226394 127744 230092 127800
rect 226333 127742 230092 127744
rect 116393 127739 116459 127742
rect 226333 127739 226399 127742
rect 213913 127258 213979 127261
rect 211508 127256 213979 127258
rect 211508 127200 213918 127256
rect 213974 127200 213979 127256
rect 211508 127198 213979 127200
rect 213913 127195 213979 127198
rect 227437 127258 227503 127261
rect 227437 127256 230092 127258
rect 227437 127200 227442 127256
rect 227498 127200 230092 127256
rect 227437 127198 230092 127200
rect 227437 127195 227503 127198
rect 343633 126714 343699 126717
rect 342148 126712 343699 126714
rect 342148 126656 343638 126712
rect 343694 126656 343699 126712
rect 342148 126654 343699 126656
rect 343633 126651 343699 126654
rect 116393 126578 116459 126581
rect 213913 126578 213979 126581
rect 116393 126576 119692 126578
rect 116393 126520 116398 126576
rect 116454 126520 119692 126576
rect 116393 126518 119692 126520
rect 211508 126576 213979 126578
rect 211508 126520 213918 126576
rect 213974 126520 213979 126576
rect 211508 126518 213979 126520
rect 116393 126515 116459 126518
rect 213913 126515 213979 126518
rect 227437 126578 227503 126581
rect 227437 126576 230092 126578
rect 227437 126520 227442 126576
rect 227498 126520 230092 126576
rect 227437 126518 230092 126520
rect 227437 126515 227503 126518
rect 227437 126034 227503 126037
rect 227437 126032 230092 126034
rect 227437 125976 227442 126032
rect 227498 125976 230092 126032
rect 227437 125974 230092 125976
rect 227437 125971 227503 125974
rect 213913 125762 213979 125765
rect 211508 125760 213979 125762
rect 211508 125704 213918 125760
rect 213974 125704 213979 125760
rect 211508 125702 213979 125704
rect 213913 125699 213979 125702
rect 116393 125490 116459 125493
rect 116393 125488 119692 125490
rect 116393 125432 116398 125488
rect 116454 125432 119692 125488
rect 116393 125430 119692 125432
rect 116393 125427 116459 125430
rect 227437 125354 227503 125357
rect 227437 125352 230092 125354
rect 227437 125296 227442 125352
rect 227498 125296 230092 125352
rect 227437 125294 230092 125296
rect 227437 125291 227503 125294
rect 32213 125084 32279 125085
rect 32213 125080 32260 125084
rect 32324 125082 32330 125084
rect 32213 125024 32218 125080
rect 32213 125020 32260 125024
rect 32324 125022 32370 125082
rect 32324 125020 32330 125022
rect 32213 125019 32279 125020
rect 213913 124946 213979 124949
rect 211508 124944 213979 124946
rect 211508 124888 213918 124944
rect 213974 124888 213979 124944
rect 211508 124886 213979 124888
rect 213913 124883 213979 124886
rect 227253 124810 227319 124813
rect 227253 124808 230092 124810
rect 227253 124752 227258 124808
rect 227314 124752 230092 124808
rect 227253 124750 230092 124752
rect 227253 124747 227319 124750
rect 116301 124266 116367 124269
rect 227253 124266 227319 124269
rect 116301 124264 119692 124266
rect 116301 124208 116306 124264
rect 116362 124208 119692 124264
rect 116301 124206 119692 124208
rect 227253 124264 230092 124266
rect 227253 124208 227258 124264
rect 227314 124208 230092 124264
rect 227253 124206 230092 124208
rect 116301 124203 116367 124206
rect 227253 124203 227319 124206
rect 213913 124130 213979 124133
rect 211508 124128 213979 124130
rect 211508 124072 213918 124128
rect 213974 124072 213979 124128
rect 211508 124070 213979 124072
rect 213913 124067 213979 124070
rect 227253 123586 227319 123589
rect 227253 123584 230092 123586
rect 227253 123528 227258 123584
rect 227314 123528 230092 123584
rect 227253 123526 230092 123528
rect 227253 123523 227319 123526
rect 213913 123450 213979 123453
rect 211508 123448 213979 123450
rect 211508 123392 213918 123448
rect 213974 123392 213979 123448
rect 211508 123390 213979 123392
rect 213913 123387 213979 123390
rect 580901 123178 580967 123181
rect 583520 123178 584960 123268
rect 580901 123176 584960 123178
rect 580901 123120 580906 123176
rect 580962 123120 584960 123176
rect 580901 123118 584960 123120
rect 580901 123115 580967 123118
rect 116577 123042 116643 123045
rect 227437 123042 227503 123045
rect 116577 123040 119692 123042
rect 116577 122984 116582 123040
rect 116638 122984 119692 123040
rect 116577 122982 119692 122984
rect 227437 123040 230092 123042
rect 227437 122984 227442 123040
rect 227498 122984 230092 123040
rect 583520 123028 584960 123118
rect 227437 122982 230092 122984
rect 116577 122979 116643 122982
rect 227437 122979 227503 122982
rect 213913 122634 213979 122637
rect 211508 122632 213979 122634
rect 211508 122576 213918 122632
rect 213974 122576 213979 122632
rect 211508 122574 213979 122576
rect 213913 122571 213979 122574
rect 227437 122362 227503 122365
rect 227437 122360 230092 122362
rect 227437 122304 227442 122360
rect 227498 122304 230092 122360
rect 227437 122302 230092 122304
rect 227437 122299 227503 122302
rect -960 121940 480 122180
rect 116393 121954 116459 121957
rect 116393 121952 119692 121954
rect 116393 121896 116398 121952
rect 116454 121896 119692 121952
rect 116393 121894 119692 121896
rect 116393 121891 116459 121894
rect 213913 121818 213979 121821
rect 211508 121816 213979 121818
rect 211508 121760 213918 121816
rect 213974 121760 213979 121816
rect 211508 121758 213979 121760
rect 213913 121755 213979 121758
rect 227437 121818 227503 121821
rect 227437 121816 230092 121818
rect 227437 121760 227442 121816
rect 227498 121760 230092 121816
rect 227437 121758 230092 121760
rect 227437 121755 227503 121758
rect 227437 121274 227503 121277
rect 227437 121272 230092 121274
rect 227437 121216 227442 121272
rect 227498 121216 230092 121272
rect 227437 121214 230092 121216
rect 227437 121211 227503 121214
rect 213913 121002 213979 121005
rect 211508 121000 213979 121002
rect 211508 120944 213918 121000
rect 213974 120944 213979 121000
rect 211508 120942 213979 120944
rect 213913 120939 213979 120942
rect 116393 120730 116459 120733
rect 116393 120728 119692 120730
rect 116393 120672 116398 120728
rect 116454 120672 119692 120728
rect 116393 120670 119692 120672
rect 116393 120667 116459 120670
rect 227437 120594 227503 120597
rect 227437 120592 230092 120594
rect 227437 120536 227442 120592
rect 227498 120536 230092 120592
rect 227437 120534 230092 120536
rect 227437 120531 227503 120534
rect 213913 120322 213979 120325
rect 211508 120320 213979 120322
rect 211508 120264 213918 120320
rect 213974 120264 213979 120320
rect 211508 120262 213979 120264
rect 213913 120259 213979 120262
rect 226425 120050 226491 120053
rect 226425 120048 230092 120050
rect 226425 119992 226430 120048
rect 226486 119992 230092 120048
rect 226425 119990 230092 119992
rect 226425 119987 226491 119990
rect 116393 119642 116459 119645
rect 116393 119640 119692 119642
rect 116393 119584 116398 119640
rect 116454 119584 119692 119640
rect 116393 119582 119692 119584
rect 116393 119579 116459 119582
rect 213913 119506 213979 119509
rect 211508 119504 213979 119506
rect 211508 119448 213918 119504
rect 213974 119448 213979 119504
rect 211508 119446 213979 119448
rect 213913 119443 213979 119446
rect 226333 119370 226399 119373
rect 226333 119368 230092 119370
rect 226333 119312 226338 119368
rect 226394 119312 230092 119368
rect 226333 119310 230092 119312
rect 226333 119307 226399 119310
rect 226241 118826 226307 118829
rect 226241 118824 230092 118826
rect 226241 118768 226246 118824
rect 226302 118768 230092 118824
rect 226241 118766 230092 118768
rect 226241 118763 226307 118766
rect 213913 118690 213979 118693
rect 211508 118688 213979 118690
rect 211508 118632 213918 118688
rect 213974 118632 213979 118688
rect 211508 118630 213979 118632
rect 213913 118627 213979 118630
rect 116393 118418 116459 118421
rect 116393 118416 119692 118418
rect 116393 118360 116398 118416
rect 116454 118360 119692 118416
rect 116393 118358 119692 118360
rect 116393 118355 116459 118358
rect 227437 118146 227503 118149
rect 227437 118144 230092 118146
rect 227437 118088 227442 118144
rect 227498 118088 230092 118144
rect 227437 118086 230092 118088
rect 227437 118083 227503 118086
rect 214005 117874 214071 117877
rect 211508 117872 214071 117874
rect 211508 117816 214010 117872
rect 214066 117816 214071 117872
rect 211508 117814 214071 117816
rect 214005 117811 214071 117814
rect 226149 117602 226215 117605
rect 226149 117600 230092 117602
rect 226149 117544 226154 117600
rect 226210 117544 230092 117600
rect 226149 117542 230092 117544
rect 226149 117539 226215 117542
rect 116393 117194 116459 117197
rect 116393 117192 119692 117194
rect 116393 117136 116398 117192
rect 116454 117136 119692 117192
rect 116393 117134 119692 117136
rect 116393 117131 116459 117134
rect 213913 117058 213979 117061
rect 211508 117056 213979 117058
rect 211508 117000 213918 117056
rect 213974 117000 213979 117056
rect 211508 116998 213979 117000
rect 213913 116995 213979 116998
rect 227437 117058 227503 117061
rect 227437 117056 230092 117058
rect 227437 117000 227442 117056
rect 227498 117000 230092 117056
rect 227437 116998 230092 117000
rect 227437 116995 227503 116998
rect 214005 116378 214071 116381
rect 211508 116376 214071 116378
rect 211508 116320 214010 116376
rect 214066 116320 214071 116376
rect 211508 116318 214071 116320
rect 214005 116315 214071 116318
rect 226241 116378 226307 116381
rect 226241 116376 230092 116378
rect 226241 116320 226246 116376
rect 226302 116320 230092 116376
rect 226241 116318 230092 116320
rect 226241 116315 226307 116318
rect 116117 116106 116183 116109
rect 116117 116104 119692 116106
rect 116117 116048 116122 116104
rect 116178 116048 119692 116104
rect 116117 116046 119692 116048
rect 116117 116043 116183 116046
rect 227069 115834 227135 115837
rect 227069 115832 230092 115834
rect 227069 115776 227074 115832
rect 227130 115776 230092 115832
rect 227069 115774 230092 115776
rect 227069 115771 227135 115774
rect 213913 115562 213979 115565
rect 211508 115560 213979 115562
rect 211508 115504 213918 115560
rect 213974 115504 213979 115560
rect 211508 115502 213979 115504
rect 213913 115499 213979 115502
rect 226149 115154 226215 115157
rect 226149 115152 230092 115154
rect 226149 115096 226154 115152
rect 226210 115096 230092 115152
rect 226149 115094 230092 115096
rect 226149 115091 226215 115094
rect 116393 114882 116459 114885
rect 116393 114880 119692 114882
rect 116393 114824 116398 114880
rect 116454 114824 119692 114880
rect 116393 114822 119692 114824
rect 116393 114819 116459 114822
rect 214005 114746 214071 114749
rect 211508 114744 214071 114746
rect 211508 114688 214010 114744
rect 214066 114688 214071 114744
rect 211508 114686 214071 114688
rect 214005 114683 214071 114686
rect 226057 114610 226123 114613
rect 226057 114608 230092 114610
rect 226057 114552 226062 114608
rect 226118 114552 230092 114608
rect 226057 114550 230092 114552
rect 226057 114547 226123 114550
rect 226241 114066 226307 114069
rect 226241 114064 230092 114066
rect 226241 114008 226246 114064
rect 226302 114008 230092 114064
rect 226241 114006 230092 114008
rect 226241 114003 226307 114006
rect 213913 113930 213979 113933
rect 211508 113928 213979 113930
rect 211508 113872 213918 113928
rect 213974 113872 213979 113928
rect 211508 113870 213979 113872
rect 213913 113867 213979 113870
rect 116393 113794 116459 113797
rect 116393 113792 119692 113794
rect 116393 113736 116398 113792
rect 116454 113736 119692 113792
rect 116393 113734 119692 113736
rect 116393 113731 116459 113734
rect 225965 113386 226031 113389
rect 225965 113384 230092 113386
rect 225965 113328 225970 113384
rect 226026 113328 230092 113384
rect 225965 113326 230092 113328
rect 225965 113323 226031 113326
rect 214005 113250 214071 113253
rect 211508 113248 214071 113250
rect 211508 113192 214010 113248
rect 214066 113192 214071 113248
rect 211508 113190 214071 113192
rect 214005 113187 214071 113190
rect 226149 112842 226215 112845
rect 226149 112840 230092 112842
rect 226149 112784 226154 112840
rect 226210 112784 230092 112840
rect 226149 112782 230092 112784
rect 226149 112779 226215 112782
rect 116393 112570 116459 112573
rect 116393 112568 119692 112570
rect 116393 112512 116398 112568
rect 116454 112512 119692 112568
rect 116393 112510 119692 112512
rect 116393 112507 116459 112510
rect 213913 112434 213979 112437
rect 211508 112432 213979 112434
rect 211508 112376 213918 112432
rect 213974 112376 213979 112432
rect 211508 112374 213979 112376
rect 213913 112371 213979 112374
rect 225873 112162 225939 112165
rect 225873 112160 230092 112162
rect 225873 112104 225878 112160
rect 225934 112104 230092 112160
rect 225873 112102 230092 112104
rect 225873 112099 225939 112102
rect 213913 111618 213979 111621
rect 211508 111616 213979 111618
rect 211508 111560 213918 111616
rect 213974 111560 213979 111616
rect 211508 111558 213979 111560
rect 213913 111555 213979 111558
rect 226241 111618 226307 111621
rect 226241 111616 230092 111618
rect 226241 111560 226246 111616
rect 226302 111560 230092 111616
rect 226241 111558 230092 111560
rect 226241 111555 226307 111558
rect 116393 111482 116459 111485
rect 116393 111480 119692 111482
rect 116393 111424 116398 111480
rect 116454 111424 119692 111480
rect 116393 111422 119692 111424
rect 116393 111419 116459 111422
rect 583520 111332 584960 111572
rect 226057 110938 226123 110941
rect 226057 110936 230092 110938
rect 226057 110880 226062 110936
rect 226118 110880 230092 110936
rect 226057 110878 230092 110880
rect 226057 110875 226123 110878
rect 214005 110802 214071 110805
rect 211508 110800 214071 110802
rect 211508 110744 214010 110800
rect 214066 110744 214071 110800
rect 211508 110742 214071 110744
rect 214005 110739 214071 110742
rect 225781 110394 225847 110397
rect 225781 110392 230092 110394
rect 225781 110336 225786 110392
rect 225842 110336 230092 110392
rect 225781 110334 230092 110336
rect 225781 110331 225847 110334
rect 116393 110258 116459 110261
rect 116393 110256 119692 110258
rect 116393 110200 116398 110256
rect 116454 110200 119692 110256
rect 116393 110198 119692 110200
rect 116393 110195 116459 110198
rect 213913 110122 213979 110125
rect 211508 110120 213979 110122
rect 211508 110064 213918 110120
rect 213974 110064 213979 110120
rect 211508 110062 213979 110064
rect 213913 110059 213979 110062
rect 226333 109850 226399 109853
rect 226333 109848 230092 109850
rect 226333 109792 226338 109848
rect 226394 109792 230092 109848
rect 226333 109790 230092 109792
rect 226333 109787 226399 109790
rect 214005 109306 214071 109309
rect 211508 109304 214071 109306
rect 211508 109248 214010 109304
rect 214066 109248 214071 109304
rect 211508 109246 214071 109248
rect 214005 109243 214071 109246
rect 225597 109170 225663 109173
rect 225597 109168 230092 109170
rect 225597 109112 225602 109168
rect 225658 109112 230092 109168
rect 225597 109110 230092 109112
rect 225597 109107 225663 109110
rect 116301 109034 116367 109037
rect 214465 109034 214531 109037
rect 214741 109034 214807 109037
rect 116301 109032 119692 109034
rect 116301 108976 116306 109032
rect 116362 108976 119692 109032
rect 116301 108974 119692 108976
rect 214465 109032 214807 109034
rect 214465 108976 214470 109032
rect 214526 108976 214746 109032
rect 214802 108976 214807 109032
rect 214465 108974 214807 108976
rect 116301 108971 116367 108974
rect 214465 108971 214531 108974
rect 214741 108971 214807 108974
rect 226149 108626 226215 108629
rect 226149 108624 230092 108626
rect 226149 108568 226154 108624
rect 226210 108568 230092 108624
rect 226149 108566 230092 108568
rect 226149 108563 226215 108566
rect 213913 108490 213979 108493
rect 211508 108488 213979 108490
rect 211508 108432 213918 108488
rect 213974 108432 213979 108488
rect 211508 108430 213979 108432
rect 213913 108427 213979 108430
rect 116393 107946 116459 107949
rect 225689 107946 225755 107949
rect 116393 107944 119692 107946
rect 116393 107888 116398 107944
rect 116454 107888 119692 107944
rect 116393 107886 119692 107888
rect 225689 107944 230092 107946
rect 225689 107888 225694 107944
rect 225750 107888 230092 107944
rect 225689 107886 230092 107888
rect 116393 107883 116459 107886
rect 225689 107883 225755 107886
rect -960 107674 480 107764
rect 2773 107674 2839 107677
rect 214005 107674 214071 107677
rect -960 107672 2839 107674
rect -960 107616 2778 107672
rect 2834 107616 2839 107672
rect -960 107614 2839 107616
rect 211508 107672 214071 107674
rect 211508 107616 214010 107672
rect 214066 107616 214071 107672
rect 211508 107614 214071 107616
rect -960 107524 480 107614
rect 2773 107611 2839 107614
rect 214005 107611 214071 107614
rect 225965 107402 226031 107405
rect 225965 107400 230092 107402
rect 225965 107344 225970 107400
rect 226026 107344 230092 107400
rect 225965 107342 230092 107344
rect 225965 107339 226031 107342
rect 213913 106994 213979 106997
rect 211508 106992 213979 106994
rect 211508 106936 213918 106992
rect 213974 106936 213979 106992
rect 211508 106934 213979 106936
rect 213913 106931 213979 106934
rect 225873 106858 225939 106861
rect 225873 106856 230092 106858
rect 225873 106800 225878 106856
rect 225934 106800 230092 106856
rect 225873 106798 230092 106800
rect 225873 106795 225939 106798
rect 116393 106722 116459 106725
rect 116393 106720 119692 106722
rect 116393 106664 116398 106720
rect 116454 106664 119692 106720
rect 116393 106662 119692 106664
rect 116393 106659 116459 106662
rect 213913 106178 213979 106181
rect 211508 106176 213979 106178
rect 211508 106120 213918 106176
rect 213974 106120 213979 106176
rect 211508 106118 213979 106120
rect 213913 106115 213979 106118
rect 226241 105770 226307 105773
rect 230062 105770 230122 106148
rect 226241 105768 230122 105770
rect 226241 105712 226246 105768
rect 226302 105712 230122 105768
rect 226241 105710 230122 105712
rect 226241 105707 226307 105710
rect 116393 105634 116459 105637
rect 226057 105634 226123 105637
rect 116393 105632 119692 105634
rect 116393 105576 116398 105632
rect 116454 105576 119692 105632
rect 116393 105574 119692 105576
rect 226057 105632 230092 105634
rect 226057 105576 226062 105632
rect 226118 105576 230092 105632
rect 226057 105574 230092 105576
rect 116393 105571 116459 105574
rect 226057 105571 226123 105574
rect 214005 105362 214071 105365
rect 211508 105360 214071 105362
rect 211508 105304 214010 105360
rect 214066 105304 214071 105360
rect 211508 105302 214071 105304
rect 214005 105299 214071 105302
rect 227437 104954 227503 104957
rect 227437 104952 230092 104954
rect 227437 104896 227442 104952
rect 227498 104896 230092 104952
rect 227437 104894 230092 104896
rect 227437 104891 227503 104894
rect 213913 104546 213979 104549
rect 211508 104544 213979 104546
rect 211508 104488 213918 104544
rect 213974 104488 213979 104544
rect 211508 104486 213979 104488
rect 213913 104483 213979 104486
rect 116393 104410 116459 104413
rect 226241 104410 226307 104413
rect 116393 104408 119692 104410
rect 116393 104352 116398 104408
rect 116454 104352 119692 104408
rect 116393 104350 119692 104352
rect 226241 104408 230092 104410
rect 226241 104352 226246 104408
rect 226302 104352 230092 104408
rect 226241 104350 230092 104352
rect 116393 104347 116459 104350
rect 226241 104347 226307 104350
rect 214005 103866 214071 103869
rect 211508 103864 214071 103866
rect 211508 103808 214010 103864
rect 214066 103808 214071 103864
rect 211508 103806 214071 103808
rect 214005 103803 214071 103806
rect 227437 103866 227503 103869
rect 227437 103864 230092 103866
rect 227437 103808 227442 103864
rect 227498 103808 230092 103864
rect 227437 103806 230092 103808
rect 227437 103803 227503 103806
rect 116301 103186 116367 103189
rect 116301 103184 119692 103186
rect 116301 103128 116306 103184
rect 116362 103128 119692 103184
rect 116301 103126 119692 103128
rect 116301 103123 116367 103126
rect 213913 103050 213979 103053
rect 211508 103048 213979 103050
rect 211508 102992 213918 103048
rect 213974 102992 213979 103048
rect 211508 102990 213979 102992
rect 213913 102987 213979 102990
rect 214005 102234 214071 102237
rect 211508 102232 214071 102234
rect 211508 102176 214010 102232
rect 214066 102176 214071 102232
rect 211508 102174 214071 102176
rect 214005 102171 214071 102174
rect 116301 102098 116367 102101
rect 116301 102096 119692 102098
rect 116301 102040 116306 102096
rect 116362 102040 119692 102096
rect 116301 102038 119692 102040
rect 116301 102035 116367 102038
rect 213913 101418 213979 101421
rect 211508 101416 213979 101418
rect 211508 101360 213918 101416
rect 213974 101360 213979 101416
rect 211508 101358 213979 101360
rect 213913 101355 213979 101358
rect 116393 100874 116459 100877
rect 116393 100872 119692 100874
rect 116393 100816 116398 100872
rect 116454 100816 119692 100872
rect 116393 100814 119692 100816
rect 116393 100811 116459 100814
rect 213913 100602 213979 100605
rect 211508 100600 213979 100602
rect 211508 100544 213918 100600
rect 213974 100544 213979 100600
rect 211508 100542 213979 100544
rect 213913 100539 213979 100542
rect 214005 99922 214071 99925
rect 211508 99920 214071 99922
rect 211508 99864 214010 99920
rect 214066 99864 214071 99920
rect 211508 99862 214071 99864
rect 214005 99859 214071 99862
rect 116393 99786 116459 99789
rect 116393 99784 119692 99786
rect 116393 99728 116398 99784
rect 116454 99728 119692 99784
rect 116393 99726 119692 99728
rect 116393 99723 116459 99726
rect 583520 99636 584960 99876
rect 215109 99106 215175 99109
rect 211508 99104 215175 99106
rect 211508 99048 215114 99104
rect 215170 99048 215175 99104
rect 211508 99046 215175 99048
rect 215109 99043 215175 99046
rect 94497 98970 94563 98973
rect 91908 98968 94563 98970
rect 91908 98912 94502 98968
rect 94558 98912 94563 98968
rect 91908 98910 94563 98912
rect 94497 98907 94563 98910
rect 116393 98562 116459 98565
rect 116393 98560 119692 98562
rect 116393 98504 116398 98560
rect 116454 98504 119692 98560
rect 116393 98502 119692 98504
rect 116393 98499 116459 98502
rect 214649 98290 214715 98293
rect 211508 98288 214715 98290
rect 211508 98232 214654 98288
rect 214710 98232 214715 98288
rect 211508 98230 214715 98232
rect 214649 98227 214715 98230
rect 94681 98018 94747 98021
rect 91908 98016 94747 98018
rect 91908 97960 94686 98016
rect 94742 97960 94747 98016
rect 91908 97958 94747 97960
rect 94681 97955 94747 97958
rect 214097 97474 214163 97477
rect 211508 97472 214163 97474
rect 211508 97416 214102 97472
rect 214158 97416 214163 97472
rect 211508 97414 214163 97416
rect 214097 97411 214163 97414
rect 116393 97338 116459 97341
rect 116393 97336 119692 97338
rect 116393 97280 116398 97336
rect 116454 97280 119692 97336
rect 116393 97278 119692 97280
rect 116393 97275 116459 97278
rect 94589 97202 94655 97205
rect 91908 97200 94655 97202
rect 91908 97144 94594 97200
rect 94650 97144 94655 97200
rect 91908 97142 94655 97144
rect 94589 97139 94655 97142
rect 213913 96794 213979 96797
rect 211508 96792 213979 96794
rect 211508 96736 213918 96792
rect 213974 96736 213979 96792
rect 211508 96734 213979 96736
rect 213913 96731 213979 96734
rect 94773 96250 94839 96253
rect 91908 96248 94839 96250
rect 91908 96192 94778 96248
rect 94834 96192 94839 96248
rect 91908 96190 94839 96192
rect 94773 96187 94839 96190
rect 116301 96250 116367 96253
rect 116301 96248 119692 96250
rect 116301 96192 116306 96248
rect 116362 96192 119692 96248
rect 116301 96190 119692 96192
rect 116301 96187 116367 96190
rect 214557 95978 214623 95981
rect 211508 95976 214623 95978
rect 211508 95920 214562 95976
rect 214618 95920 214623 95976
rect 211508 95918 214623 95920
rect 214557 95915 214623 95918
rect 94957 95434 95023 95437
rect 91908 95432 95023 95434
rect 91908 95376 94962 95432
rect 95018 95376 95023 95432
rect 91908 95374 95023 95376
rect 94957 95371 95023 95374
rect 214741 95162 214807 95165
rect 211508 95160 214807 95162
rect 211508 95104 214746 95160
rect 214802 95104 214807 95160
rect 211508 95102 214807 95104
rect 214741 95099 214807 95102
rect 116485 95026 116551 95029
rect 116485 95024 119692 95026
rect 116485 94968 116490 95024
rect 116546 94968 119692 95024
rect 116485 94966 119692 94968
rect 116485 94963 116551 94966
rect 94865 94482 94931 94485
rect 91908 94480 94931 94482
rect 91908 94424 94870 94480
rect 94926 94424 94931 94480
rect 91908 94422 94931 94424
rect 94865 94419 94931 94422
rect 215109 94346 215175 94349
rect 211508 94344 215175 94346
rect 211508 94288 215114 94344
rect 215170 94288 215175 94344
rect 211508 94286 215175 94288
rect 215109 94283 215175 94286
rect 116393 93938 116459 93941
rect 116393 93936 119692 93938
rect 116393 93880 116398 93936
rect 116454 93880 119692 93936
rect 116393 93878 119692 93880
rect 116393 93875 116459 93878
rect 215109 93666 215175 93669
rect 211508 93664 215175 93666
rect 211508 93608 215114 93664
rect 215170 93608 215175 93664
rect 211508 93606 215175 93608
rect 215109 93603 215175 93606
rect 95141 93530 95207 93533
rect 91908 93528 95207 93530
rect 91908 93472 95146 93528
rect 95202 93472 95207 93528
rect 91908 93470 95207 93472
rect 95141 93467 95207 93470
rect -960 93258 480 93348
rect 2773 93258 2839 93261
rect -960 93256 2839 93258
rect -960 93200 2778 93256
rect 2834 93200 2839 93256
rect -960 93198 2839 93200
rect -960 93108 480 93198
rect 2773 93195 2839 93198
rect 215201 92850 215267 92853
rect 211508 92848 215267 92850
rect 211508 92792 215206 92848
rect 215262 92792 215267 92848
rect 211508 92790 215267 92792
rect 215201 92787 215267 92790
rect 94405 92714 94471 92717
rect 91908 92712 94471 92714
rect 91908 92656 94410 92712
rect 94466 92656 94471 92712
rect 91908 92654 94471 92656
rect 94405 92651 94471 92654
rect 116393 92714 116459 92717
rect 116393 92712 119692 92714
rect 116393 92656 116398 92712
rect 116454 92656 119692 92712
rect 116393 92654 119692 92656
rect 116393 92651 116459 92654
rect 214833 92034 214899 92037
rect 211508 92032 214899 92034
rect 211508 91976 214838 92032
rect 214894 91976 214899 92032
rect 211508 91974 214899 91976
rect 214833 91971 214899 91974
rect 94589 91762 94655 91765
rect 91908 91760 94655 91762
rect 91908 91704 94594 91760
rect 94650 91704 94655 91760
rect 91908 91702 94655 91704
rect 94589 91699 94655 91702
rect 116393 91626 116459 91629
rect 116393 91624 119692 91626
rect 116393 91568 116398 91624
rect 116454 91568 119692 91624
rect 116393 91566 119692 91568
rect 116393 91563 116459 91566
rect 215017 91218 215083 91221
rect 211508 91216 215083 91218
rect 211508 91160 215022 91216
rect 215078 91160 215083 91216
rect 211508 91158 215083 91160
rect 215017 91155 215083 91158
rect 95049 90946 95115 90949
rect 91908 90944 95115 90946
rect 91908 90888 95054 90944
rect 95110 90888 95115 90944
rect 91908 90886 95115 90888
rect 95049 90883 95115 90886
rect 214557 90538 214623 90541
rect 211508 90536 214623 90538
rect 211508 90480 214562 90536
rect 214618 90480 214623 90536
rect 211508 90478 214623 90480
rect 214557 90475 214623 90478
rect 116393 90402 116459 90405
rect 116393 90400 119692 90402
rect 116393 90344 116398 90400
rect 116454 90344 119692 90400
rect 116393 90342 119692 90344
rect 116393 90339 116459 90342
rect 94773 89994 94839 89997
rect 91908 89992 94839 89994
rect 91908 89936 94778 89992
rect 94834 89936 94839 89992
rect 91908 89934 94839 89936
rect 94773 89931 94839 89934
rect 214281 89722 214347 89725
rect 211508 89720 214347 89722
rect 211508 89664 214286 89720
rect 214342 89664 214347 89720
rect 211508 89662 214347 89664
rect 214281 89659 214347 89662
rect 94957 89178 95023 89181
rect 91908 89176 95023 89178
rect 91908 89120 94962 89176
rect 95018 89120 95023 89176
rect 91908 89118 95023 89120
rect 94957 89115 95023 89118
rect 115933 89178 115999 89181
rect 115933 89176 119692 89178
rect 115933 89120 115938 89176
rect 115994 89120 119692 89176
rect 115933 89118 119692 89120
rect 115933 89115 115999 89118
rect 214741 88906 214807 88909
rect 211508 88904 214807 88906
rect 211508 88848 214746 88904
rect 214802 88848 214807 88904
rect 211508 88846 214807 88848
rect 214741 88843 214807 88846
rect 95141 88226 95207 88229
rect 91908 88224 95207 88226
rect 91908 88168 95146 88224
rect 95202 88168 95207 88224
rect 91908 88166 95207 88168
rect 95141 88163 95207 88166
rect 116393 88090 116459 88093
rect 214189 88090 214255 88093
rect 116393 88088 119692 88090
rect 116393 88032 116398 88088
rect 116454 88032 119692 88088
rect 116393 88030 119692 88032
rect 211508 88088 214255 88090
rect 211508 88032 214194 88088
rect 214250 88032 214255 88088
rect 211508 88030 214255 88032
rect 116393 88027 116459 88030
rect 214189 88027 214255 88030
rect 580165 87954 580231 87957
rect 583520 87954 584960 88044
rect 580165 87952 584960 87954
rect 580165 87896 580170 87952
rect 580226 87896 584960 87952
rect 580165 87894 584960 87896
rect 580165 87891 580231 87894
rect 583520 87804 584960 87894
rect 214649 87410 214715 87413
rect 211508 87408 214715 87410
rect 211508 87352 214654 87408
rect 214710 87352 214715 87408
rect 211508 87350 214715 87352
rect 214649 87347 214715 87350
rect 94313 87274 94379 87277
rect 91908 87272 94379 87274
rect 91908 87216 94318 87272
rect 94374 87216 94379 87272
rect 91908 87214 94379 87216
rect 94313 87211 94379 87214
rect 116301 86866 116367 86869
rect 116301 86864 119692 86866
rect 116301 86808 116306 86864
rect 116362 86808 119692 86864
rect 116301 86806 119692 86808
rect 116301 86803 116367 86806
rect 214465 86594 214531 86597
rect 211508 86592 214531 86594
rect 211508 86536 214470 86592
rect 214526 86536 214531 86592
rect 211508 86534 214531 86536
rect 214465 86531 214531 86534
rect 94405 86458 94471 86461
rect 91908 86456 94471 86458
rect 91908 86400 94410 86456
rect 94466 86400 94471 86456
rect 91908 86398 94471 86400
rect 94405 86395 94471 86398
rect 116393 85778 116459 85781
rect 215109 85778 215175 85781
rect 116393 85776 119692 85778
rect 116393 85720 116398 85776
rect 116454 85720 119692 85776
rect 116393 85718 119692 85720
rect 211508 85776 215175 85778
rect 211508 85720 215114 85776
rect 215170 85720 215175 85776
rect 211508 85718 215175 85720
rect 116393 85715 116459 85718
rect 215109 85715 215175 85718
rect 94221 85506 94287 85509
rect 91908 85504 94287 85506
rect 91908 85448 94226 85504
rect 94282 85448 94287 85504
rect 91908 85446 94287 85448
rect 94221 85443 94287 85446
rect 214373 84962 214439 84965
rect 211508 84960 214439 84962
rect 211508 84904 214378 84960
rect 214434 84904 214439 84960
rect 211508 84902 214439 84904
rect 214373 84899 214439 84902
rect 95141 84690 95207 84693
rect 91908 84688 95207 84690
rect 91908 84632 95146 84688
rect 95202 84632 95207 84688
rect 91908 84630 95207 84632
rect 95141 84627 95207 84630
rect 116393 84554 116459 84557
rect 116393 84552 119692 84554
rect 116393 84496 116398 84552
rect 116454 84496 119692 84552
rect 116393 84494 119692 84496
rect 116393 84491 116459 84494
rect 215109 84282 215175 84285
rect 211508 84280 215175 84282
rect 211508 84224 215114 84280
rect 215170 84224 215175 84280
rect 211508 84222 215175 84224
rect 215109 84219 215175 84222
rect 95141 83738 95207 83741
rect 91908 83736 95207 83738
rect 91908 83680 95146 83736
rect 95202 83680 95207 83736
rect 91908 83678 95207 83680
rect 95141 83675 95207 83678
rect 214373 83466 214439 83469
rect 211508 83464 214439 83466
rect 211508 83408 214378 83464
rect 214434 83408 214439 83464
rect 211508 83406 214439 83408
rect 214373 83403 214439 83406
rect 116393 83330 116459 83333
rect 116393 83328 119692 83330
rect 116393 83272 116398 83328
rect 116454 83272 119692 83328
rect 116393 83270 119692 83272
rect 116393 83267 116459 83270
rect 94221 82922 94287 82925
rect 91908 82920 94287 82922
rect 91908 82864 94226 82920
rect 94282 82864 94287 82920
rect 91908 82862 94287 82864
rect 94221 82859 94287 82862
rect 214189 82650 214255 82653
rect 211508 82648 214255 82650
rect 211508 82592 214194 82648
rect 214250 82592 214255 82648
rect 211508 82590 214255 82592
rect 214189 82587 214255 82590
rect 115933 82242 115999 82245
rect 115933 82240 119692 82242
rect 115933 82184 115938 82240
rect 115994 82184 119692 82240
rect 115933 82182 119692 82184
rect 115933 82179 115999 82182
rect 94129 81970 94195 81973
rect 91908 81968 94195 81970
rect 91908 81912 94134 81968
rect 94190 81912 94195 81968
rect 91908 81910 94195 81912
rect 94129 81907 94195 81910
rect 215201 81834 215267 81837
rect 211508 81832 215267 81834
rect 211508 81776 215206 81832
rect 215262 81776 215267 81832
rect 211508 81774 215267 81776
rect 215201 81771 215267 81774
rect 227437 81154 227503 81157
rect 227437 81152 230092 81154
rect 227437 81096 227442 81152
rect 227498 81096 230092 81152
rect 227437 81094 230092 81096
rect 227437 81091 227503 81094
rect 94405 81018 94471 81021
rect 91908 81016 94471 81018
rect 91908 80960 94410 81016
rect 94466 80960 94471 81016
rect 91908 80958 94471 80960
rect 94405 80955 94471 80958
rect 116393 81018 116459 81021
rect 215109 81018 215175 81021
rect 116393 81016 119692 81018
rect 116393 80960 116398 81016
rect 116454 80960 119692 81016
rect 116393 80958 119692 80960
rect 211508 81016 215175 81018
rect 211508 80960 215114 81016
rect 215170 80960 215175 81016
rect 211508 80958 215175 80960
rect 116393 80955 116459 80958
rect 215109 80955 215175 80958
rect 227345 80474 227411 80477
rect 227345 80472 230092 80474
rect 227345 80416 227350 80472
rect 227406 80416 230092 80472
rect 227345 80414 230092 80416
rect 227345 80411 227411 80414
rect 214925 80338 214991 80341
rect 211508 80336 214991 80338
rect 211508 80280 214930 80336
rect 214986 80280 214991 80336
rect 211508 80278 214991 80280
rect 214925 80275 214991 80278
rect 94681 80202 94747 80205
rect 91908 80200 94747 80202
rect 91908 80144 94686 80200
rect 94742 80144 94747 80200
rect 91908 80142 94747 80144
rect 94681 80139 94747 80142
rect 116209 79930 116275 79933
rect 116209 79928 119692 79930
rect 116209 79872 116214 79928
rect 116270 79872 119692 79928
rect 116209 79870 119692 79872
rect 116209 79867 116275 79870
rect 227437 79794 227503 79797
rect 227437 79792 230092 79794
rect 227437 79736 227442 79792
rect 227498 79736 230092 79792
rect 227437 79734 230092 79736
rect 227437 79731 227503 79734
rect 213913 79522 213979 79525
rect 211508 79520 213979 79522
rect 211508 79464 213918 79520
rect 213974 79464 213979 79520
rect 211508 79462 213979 79464
rect 213913 79459 213979 79462
rect 94405 79250 94471 79253
rect 91908 79248 94471 79250
rect 91908 79192 94410 79248
rect 94466 79192 94471 79248
rect 91908 79190 94471 79192
rect 94405 79187 94471 79190
rect 227529 79114 227595 79117
rect 227529 79112 230092 79114
rect -960 78828 480 79068
rect 227529 79056 227534 79112
rect 227590 79056 230092 79112
rect 227529 79054 230092 79056
rect 227529 79051 227595 79054
rect 116393 78706 116459 78709
rect 214833 78706 214899 78709
rect 116393 78704 119692 78706
rect 116393 78648 116398 78704
rect 116454 78648 119692 78704
rect 116393 78646 119692 78648
rect 211508 78704 214899 78706
rect 211508 78648 214838 78704
rect 214894 78648 214899 78704
rect 211508 78646 214899 78648
rect 116393 78643 116459 78646
rect 214833 78643 214899 78646
rect 227437 78570 227503 78573
rect 227437 78568 230092 78570
rect 227437 78512 227442 78568
rect 227498 78512 230092 78568
rect 227437 78510 230092 78512
rect 227437 78507 227503 78510
rect 94497 78434 94563 78437
rect 91908 78432 94563 78434
rect 91908 78376 94502 78432
rect 94558 78376 94563 78432
rect 91908 78374 94563 78376
rect 94497 78371 94563 78374
rect 213913 77890 213979 77893
rect 211508 77888 213979 77890
rect 211508 77832 213918 77888
rect 213974 77832 213979 77888
rect 211508 77830 213979 77832
rect 213913 77827 213979 77830
rect 227529 77890 227595 77893
rect 227529 77888 230092 77890
rect 227529 77832 227534 77888
rect 227590 77832 230092 77888
rect 227529 77830 230092 77832
rect 227529 77827 227595 77830
rect 94221 77482 94287 77485
rect 91908 77480 94287 77482
rect 91908 77424 94226 77480
rect 94282 77424 94287 77480
rect 91908 77422 94287 77424
rect 94221 77419 94287 77422
rect 116393 77482 116459 77485
rect 116393 77480 119692 77482
rect 116393 77424 116398 77480
rect 116454 77424 119692 77480
rect 116393 77422 119692 77424
rect 116393 77419 116459 77422
rect 215017 77210 215083 77213
rect 211508 77208 215083 77210
rect 211508 77152 215022 77208
rect 215078 77152 215083 77208
rect 211508 77150 215083 77152
rect 215017 77147 215083 77150
rect 227437 77210 227503 77213
rect 227437 77208 230092 77210
rect 227437 77152 227442 77208
rect 227498 77152 230092 77208
rect 227437 77150 230092 77152
rect 227437 77147 227503 77150
rect 94589 76530 94655 76533
rect 91908 76528 94655 76530
rect 91908 76472 94594 76528
rect 94650 76472 94655 76528
rect 91908 76470 94655 76472
rect 94589 76467 94655 76470
rect 227529 76530 227595 76533
rect 227529 76528 230092 76530
rect 227529 76472 227534 76528
rect 227590 76472 230092 76528
rect 227529 76470 230092 76472
rect 227529 76467 227595 76470
rect 116393 76394 116459 76397
rect 213913 76394 213979 76397
rect 116393 76392 119692 76394
rect 116393 76336 116398 76392
rect 116454 76336 119692 76392
rect 116393 76334 119692 76336
rect 211508 76392 213979 76394
rect 211508 76336 213918 76392
rect 213974 76336 213979 76392
rect 211508 76334 213979 76336
rect 116393 76331 116459 76334
rect 213913 76331 213979 76334
rect 580901 76258 580967 76261
rect 583520 76258 584960 76348
rect 580901 76256 584960 76258
rect 580901 76200 580906 76256
rect 580962 76200 584960 76256
rect 580901 76198 584960 76200
rect 580901 76195 580967 76198
rect 583520 76108 584960 76198
rect 227437 75850 227503 75853
rect 227437 75848 230092 75850
rect 227437 75792 227442 75848
rect 227498 75792 230092 75848
rect 227437 75790 230092 75792
rect 227437 75787 227503 75790
rect 94589 75714 94655 75717
rect 91908 75712 94655 75714
rect 91908 75656 94594 75712
rect 94650 75656 94655 75712
rect 91908 75654 94655 75656
rect 94589 75651 94655 75654
rect 214741 75578 214807 75581
rect 211508 75576 214807 75578
rect 211508 75520 214746 75576
rect 214802 75520 214807 75576
rect 211508 75518 214807 75520
rect 214741 75515 214807 75518
rect 227437 75306 227503 75309
rect 227437 75304 230092 75306
rect 227437 75248 227442 75304
rect 227498 75248 230092 75304
rect 227437 75246 230092 75248
rect 227437 75243 227503 75246
rect 116393 75170 116459 75173
rect 116393 75168 119692 75170
rect 116393 75112 116398 75168
rect 116454 75112 119692 75168
rect 116393 75110 119692 75112
rect 116393 75107 116459 75110
rect 94957 74762 95023 74765
rect 213913 74762 213979 74765
rect 91908 74760 95023 74762
rect 91908 74704 94962 74760
rect 95018 74704 95023 74760
rect 91908 74702 95023 74704
rect 211508 74760 213979 74762
rect 211508 74704 213918 74760
rect 213974 74704 213979 74760
rect 211508 74702 213979 74704
rect 94957 74699 95023 74702
rect 213913 74699 213979 74702
rect 225597 74626 225663 74629
rect 225597 74624 230092 74626
rect 225597 74568 225602 74624
rect 225658 74568 230092 74624
rect 225597 74566 230092 74568
rect 225597 74563 225663 74566
rect 116393 74082 116459 74085
rect 214097 74082 214163 74085
rect 116393 74080 119692 74082
rect 116393 74024 116398 74080
rect 116454 74024 119692 74080
rect 116393 74022 119692 74024
rect 211508 74080 214163 74082
rect 211508 74024 214102 74080
rect 214158 74024 214163 74080
rect 211508 74022 214163 74024
rect 116393 74019 116459 74022
rect 214097 74019 214163 74022
rect 94589 73946 94655 73949
rect 91908 73944 94655 73946
rect 91908 73888 94594 73944
rect 94650 73888 94655 73944
rect 91908 73886 94655 73888
rect 94589 73883 94655 73886
rect 227437 73946 227503 73949
rect 227437 73944 230092 73946
rect 227437 73888 227442 73944
rect 227498 73888 230092 73944
rect 227437 73886 230092 73888
rect 227437 73883 227503 73886
rect 213913 73266 213979 73269
rect 211508 73264 213979 73266
rect 211508 73208 213918 73264
rect 213974 73208 213979 73264
rect 211508 73206 213979 73208
rect 213913 73203 213979 73206
rect 226977 73266 227043 73269
rect 226977 73264 230092 73266
rect 226977 73208 226982 73264
rect 227038 73208 230092 73264
rect 226977 73206 230092 73208
rect 226977 73203 227043 73206
rect 94773 72994 94839 72997
rect 91908 72992 94839 72994
rect 91908 72936 94778 72992
rect 94834 72936 94839 72992
rect 91908 72934 94839 72936
rect 94773 72931 94839 72934
rect 116393 72858 116459 72861
rect 116393 72856 119692 72858
rect 116393 72800 116398 72856
rect 116454 72800 119692 72856
rect 116393 72798 119692 72800
rect 116393 72795 116459 72798
rect 227437 72722 227503 72725
rect 227437 72720 230092 72722
rect 227437 72664 227442 72720
rect 227498 72664 230092 72720
rect 227437 72662 230092 72664
rect 227437 72659 227503 72662
rect 214557 72450 214623 72453
rect 211508 72448 214623 72450
rect 211508 72392 214562 72448
rect 214618 72392 214623 72448
rect 211508 72390 214623 72392
rect 214557 72387 214623 72390
rect 94405 72178 94471 72181
rect 91908 72176 94471 72178
rect 91908 72120 94410 72176
rect 94466 72120 94471 72176
rect 91908 72118 94471 72120
rect 94405 72115 94471 72118
rect 227529 72042 227595 72045
rect 227529 72040 230092 72042
rect 227529 71984 227534 72040
rect 227590 71984 230092 72040
rect 227529 71982 230092 71984
rect 227529 71979 227595 71982
rect 116577 71770 116643 71773
rect 116577 71768 119692 71770
rect 116577 71712 116582 71768
rect 116638 71712 119692 71768
rect 116577 71710 119692 71712
rect 116577 71707 116643 71710
rect 214005 71634 214071 71637
rect 211508 71632 214071 71634
rect 211508 71576 214010 71632
rect 214066 71576 214071 71632
rect 211508 71574 214071 71576
rect 214005 71571 214071 71574
rect 227437 71362 227503 71365
rect 227437 71360 230092 71362
rect 227437 71304 227442 71360
rect 227498 71304 230092 71360
rect 227437 71302 230092 71304
rect 227437 71299 227503 71302
rect 94865 71226 94931 71229
rect 91908 71224 94931 71226
rect 91908 71168 94870 71224
rect 94926 71168 94931 71224
rect 91908 71166 94931 71168
rect 94865 71163 94931 71166
rect 213913 70954 213979 70957
rect 211508 70952 213979 70954
rect 211508 70896 213918 70952
rect 213974 70896 213979 70952
rect 211508 70894 213979 70896
rect 213913 70891 213979 70894
rect 227529 70682 227595 70685
rect 227529 70680 230092 70682
rect 227529 70624 227534 70680
rect 227590 70624 230092 70680
rect 227529 70622 230092 70624
rect 227529 70619 227595 70622
rect 116393 70546 116459 70549
rect 116393 70544 119692 70546
rect 116393 70488 116398 70544
rect 116454 70488 119692 70544
rect 116393 70486 119692 70488
rect 116393 70483 116459 70486
rect 94865 70274 94931 70277
rect 91908 70272 94931 70274
rect 91908 70216 94870 70272
rect 94926 70216 94931 70272
rect 91908 70214 94931 70216
rect 94865 70211 94931 70214
rect 214649 70138 214715 70141
rect 211508 70136 214715 70138
rect 211508 70080 214654 70136
rect 214710 70080 214715 70136
rect 211508 70078 214715 70080
rect 214649 70075 214715 70078
rect 227437 70002 227503 70005
rect 227437 70000 230092 70002
rect 227437 69944 227442 70000
rect 227498 69944 230092 70000
rect 227437 69942 230092 69944
rect 227437 69939 227503 69942
rect 95049 69458 95115 69461
rect 91908 69456 95115 69458
rect 91908 69400 95054 69456
rect 95110 69400 95115 69456
rect 91908 69398 95115 69400
rect 95049 69395 95115 69398
rect 226517 69458 226583 69461
rect 226517 69456 230092 69458
rect 226517 69400 226522 69456
rect 226578 69400 230092 69456
rect 226517 69398 230092 69400
rect 226517 69395 226583 69398
rect 116393 69322 116459 69325
rect 215109 69322 215175 69325
rect 116393 69320 119692 69322
rect 116393 69264 116398 69320
rect 116454 69264 119692 69320
rect 116393 69262 119692 69264
rect 211508 69320 215175 69322
rect 211508 69264 215114 69320
rect 215170 69264 215175 69320
rect 211508 69262 215175 69264
rect 116393 69259 116459 69262
rect 215109 69259 215175 69262
rect 227437 68778 227503 68781
rect 227437 68776 230092 68778
rect 227437 68720 227442 68776
rect 227498 68720 230092 68776
rect 227437 68718 230092 68720
rect 227437 68715 227503 68718
rect 93853 68506 93919 68509
rect 214465 68506 214531 68509
rect 91908 68504 93919 68506
rect 91908 68448 93858 68504
rect 93914 68448 93919 68504
rect 91908 68446 93919 68448
rect 211508 68504 214531 68506
rect 211508 68448 214470 68504
rect 214526 68448 214531 68504
rect 211508 68446 214531 68448
rect 93853 68443 93919 68446
rect 214465 68443 214531 68446
rect 116393 68234 116459 68237
rect 116393 68232 119692 68234
rect 116393 68176 116398 68232
rect 116454 68176 119692 68232
rect 116393 68174 119692 68176
rect 116393 68171 116459 68174
rect 227529 68098 227595 68101
rect 227529 68096 230092 68098
rect 227529 68040 227534 68096
rect 227590 68040 230092 68096
rect 227529 68038 230092 68040
rect 227529 68035 227595 68038
rect 215109 67826 215175 67829
rect 211508 67824 215175 67826
rect 211508 67768 215114 67824
rect 215170 67768 215175 67824
rect 211508 67766 215175 67768
rect 215109 67763 215175 67766
rect 95141 67690 95207 67693
rect 91908 67688 95207 67690
rect 91908 67632 95146 67688
rect 95202 67632 95207 67688
rect 91908 67630 95207 67632
rect 95141 67627 95207 67630
rect 227437 67418 227503 67421
rect 227437 67416 230092 67418
rect 227437 67360 227442 67416
rect 227498 67360 230092 67416
rect 227437 67358 230092 67360
rect 227437 67355 227503 67358
rect 116393 67010 116459 67013
rect 215109 67010 215175 67013
rect 116393 67008 119692 67010
rect 116393 66952 116398 67008
rect 116454 66952 119692 67008
rect 116393 66950 119692 66952
rect 211508 67008 215175 67010
rect 211508 66952 215114 67008
rect 215170 66952 215175 67008
rect 211508 66950 215175 66952
rect 116393 66947 116459 66950
rect 215109 66947 215175 66950
rect 227529 66874 227595 66877
rect 227529 66872 230092 66874
rect 227529 66816 227534 66872
rect 227590 66816 230092 66872
rect 227529 66814 230092 66816
rect 227529 66811 227595 66814
rect 95141 66738 95207 66741
rect 91908 66736 95207 66738
rect 91908 66680 95146 66736
rect 95202 66680 95207 66736
rect 91908 66678 95207 66680
rect 95141 66675 95207 66678
rect 214373 66194 214439 66197
rect 211508 66192 214439 66194
rect 211508 66136 214378 66192
rect 214434 66136 214439 66192
rect 211508 66134 214439 66136
rect 214373 66131 214439 66134
rect 227437 66194 227503 66197
rect 227437 66192 230092 66194
rect 227437 66136 227442 66192
rect 227498 66136 230092 66192
rect 227437 66134 230092 66136
rect 227437 66131 227503 66134
rect 94681 65922 94747 65925
rect 91908 65920 94747 65922
rect 91908 65864 94686 65920
rect 94742 65864 94747 65920
rect 91908 65862 94747 65864
rect 94681 65859 94747 65862
rect 116393 65922 116459 65925
rect 116393 65920 119692 65922
rect 116393 65864 116398 65920
rect 116454 65864 119692 65920
rect 116393 65862 119692 65864
rect 116393 65859 116459 65862
rect 6177 65514 6243 65517
rect 227529 65514 227595 65517
rect 6177 65512 9292 65514
rect 6177 65456 6182 65512
rect 6238 65456 9292 65512
rect 6177 65454 9292 65456
rect 227529 65512 230092 65514
rect 227529 65456 227534 65512
rect 227590 65456 230092 65512
rect 227529 65454 230092 65456
rect 6177 65451 6243 65454
rect 227529 65451 227595 65454
rect 214005 65378 214071 65381
rect 211508 65376 214071 65378
rect 211508 65320 214010 65376
rect 214066 65320 214071 65376
rect 211508 65318 214071 65320
rect 214005 65315 214071 65318
rect 94681 64970 94747 64973
rect 91908 64968 94747 64970
rect 91908 64912 94686 64968
rect 94742 64912 94747 64968
rect 91908 64910 94747 64912
rect 94681 64907 94747 64910
rect 227437 64834 227503 64837
rect 227437 64832 230092 64834
rect 227437 64776 227442 64832
rect 227498 64776 230092 64832
rect 227437 64774 230092 64776
rect 227437 64771 227503 64774
rect 115933 64698 115999 64701
rect 115933 64696 119692 64698
rect -960 64562 480 64652
rect 115933 64640 115938 64696
rect 115994 64640 119692 64696
rect 115933 64638 119692 64640
rect 115933 64635 115999 64638
rect 2773 64562 2839 64565
rect 214557 64562 214623 64565
rect -960 64560 2839 64562
rect -960 64504 2778 64560
rect 2834 64504 2839 64560
rect -960 64502 2839 64504
rect 211508 64560 214623 64562
rect 211508 64504 214562 64560
rect 214618 64504 214623 64560
rect 211508 64502 214623 64504
rect -960 64412 480 64502
rect 2773 64499 2839 64502
rect 214557 64499 214623 64502
rect 583520 64412 584960 64652
rect 227437 64154 227503 64157
rect 227437 64152 230092 64154
rect 227437 64096 227442 64152
rect 227498 64096 230092 64152
rect 227437 64094 230092 64096
rect 227437 64091 227503 64094
rect 94497 64018 94563 64021
rect 91908 64016 94563 64018
rect 91908 63960 94502 64016
rect 94558 63960 94563 64016
rect 91908 63958 94563 63960
rect 94497 63955 94563 63958
rect 215109 63882 215175 63885
rect 211508 63880 215175 63882
rect 211508 63824 215114 63880
rect 215170 63824 215175 63880
rect 211508 63822 215175 63824
rect 215109 63819 215175 63822
rect 227529 63610 227595 63613
rect 227529 63608 230092 63610
rect 227529 63552 227534 63608
rect 227590 63552 230092 63608
rect 227529 63550 230092 63552
rect 227529 63547 227595 63550
rect 116209 63474 116275 63477
rect 116209 63472 119692 63474
rect 116209 63416 116214 63472
rect 116270 63416 119692 63472
rect 116209 63414 119692 63416
rect 116209 63411 116275 63414
rect 94865 63202 94931 63205
rect 91908 63200 94931 63202
rect 91908 63144 94870 63200
rect 94926 63144 94931 63200
rect 91908 63142 94931 63144
rect 94865 63139 94931 63142
rect 214649 63066 214715 63069
rect 211508 63064 214715 63066
rect 211508 63008 214654 63064
rect 214710 63008 214715 63064
rect 211508 63006 214715 63008
rect 214649 63003 214715 63006
rect 227437 62930 227503 62933
rect 227437 62928 230092 62930
rect 227437 62872 227442 62928
rect 227498 62872 230092 62928
rect 227437 62870 230092 62872
rect 227437 62867 227503 62870
rect 116393 62386 116459 62389
rect 116393 62384 119692 62386
rect 116393 62328 116398 62384
rect 116454 62328 119692 62384
rect 116393 62326 119692 62328
rect 116393 62323 116459 62326
rect 94957 62250 95023 62253
rect 215109 62250 215175 62253
rect 91908 62248 95023 62250
rect 91908 62192 94962 62248
rect 95018 62192 95023 62248
rect 91908 62190 95023 62192
rect 211508 62248 215175 62250
rect 211508 62192 215114 62248
rect 215170 62192 215175 62248
rect 211508 62190 215175 62192
rect 94957 62187 95023 62190
rect 215109 62187 215175 62190
rect 227529 62250 227595 62253
rect 227529 62248 230092 62250
rect 227529 62192 227534 62248
rect 227590 62192 230092 62248
rect 227529 62190 230092 62192
rect 227529 62187 227595 62190
rect 227529 61570 227595 61573
rect 227529 61568 230092 61570
rect 227529 61512 227534 61568
rect 227590 61512 230092 61568
rect 227529 61510 230092 61512
rect 227529 61507 227595 61510
rect 93945 61434 94011 61437
rect 214557 61434 214623 61437
rect 91908 61432 94011 61434
rect 91908 61376 93950 61432
rect 94006 61376 94011 61432
rect 91908 61374 94011 61376
rect 211508 61432 214623 61434
rect 211508 61376 214562 61432
rect 214618 61376 214623 61432
rect 211508 61374 214623 61376
rect 93945 61371 94011 61374
rect 214557 61371 214623 61374
rect 116393 61162 116459 61165
rect 116393 61160 119692 61162
rect 116393 61104 116398 61160
rect 116454 61104 119692 61160
rect 116393 61102 119692 61104
rect 116393 61099 116459 61102
rect 226701 61026 226767 61029
rect 226701 61024 230092 61026
rect 226701 60968 226706 61024
rect 226762 60968 230092 61024
rect 226701 60966 230092 60968
rect 226701 60963 226767 60966
rect 215109 60754 215175 60757
rect 211508 60752 215175 60754
rect 211508 60696 215114 60752
rect 215170 60696 215175 60752
rect 211508 60694 215175 60696
rect 215109 60691 215175 60694
rect 94589 60482 94655 60485
rect 91908 60480 94655 60482
rect 91908 60424 94594 60480
rect 94650 60424 94655 60480
rect 91908 60422 94655 60424
rect 94589 60419 94655 60422
rect 227069 60346 227135 60349
rect 227069 60344 230092 60346
rect 227069 60288 227074 60344
rect 227130 60288 230092 60344
rect 227069 60286 230092 60288
rect 227069 60283 227135 60286
rect 116393 60074 116459 60077
rect 116393 60072 119692 60074
rect 116393 60016 116398 60072
rect 116454 60016 119692 60072
rect 116393 60014 119692 60016
rect 116393 60011 116459 60014
rect 214557 59938 214623 59941
rect 211508 59936 214623 59938
rect 211508 59880 214562 59936
rect 214618 59880 214623 59936
rect 211508 59878 214623 59880
rect 214557 59875 214623 59878
rect 227437 59666 227503 59669
rect 227437 59664 230092 59666
rect 227437 59608 227442 59664
rect 227498 59608 230092 59664
rect 227437 59606 230092 59608
rect 227437 59603 227503 59606
rect 94405 59530 94471 59533
rect 91908 59528 94471 59530
rect 91908 59472 94410 59528
rect 94466 59472 94471 59528
rect 91908 59470 94471 59472
rect 94405 59467 94471 59470
rect 214097 59122 214163 59125
rect 211508 59120 214163 59122
rect 211508 59064 214102 59120
rect 214158 59064 214163 59120
rect 211508 59062 214163 59064
rect 214097 59059 214163 59062
rect 227437 58986 227503 58989
rect 227437 58984 230092 58986
rect 227437 58928 227442 58984
rect 227498 58928 230092 58984
rect 227437 58926 230092 58928
rect 227437 58923 227503 58926
rect 116393 58850 116459 58853
rect 116393 58848 119692 58850
rect 116393 58792 116398 58848
rect 116454 58792 119692 58848
rect 116393 58790 119692 58792
rect 116393 58787 116459 58790
rect 94773 58714 94839 58717
rect 91908 58712 94839 58714
rect 91908 58656 94778 58712
rect 94834 58656 94839 58712
rect 91908 58654 94839 58656
rect 94773 58651 94839 58654
rect 214189 58306 214255 58309
rect 211508 58304 214255 58306
rect 211508 58248 214194 58304
rect 214250 58248 214255 58304
rect 211508 58246 214255 58248
rect 214189 58243 214255 58246
rect 227529 58306 227595 58309
rect 227529 58304 230092 58306
rect 227529 58248 227534 58304
rect 227590 58248 230092 58304
rect 227529 58246 230092 58248
rect 227529 58243 227595 58246
rect 94221 57762 94287 57765
rect 91908 57760 94287 57762
rect 91908 57704 94226 57760
rect 94282 57704 94287 57760
rect 91908 57702 94287 57704
rect 94221 57699 94287 57702
rect 227253 57762 227319 57765
rect 227253 57760 230092 57762
rect 227253 57704 227258 57760
rect 227314 57704 230092 57760
rect 227253 57702 230092 57704
rect 227253 57699 227319 57702
rect 116301 57626 116367 57629
rect 213913 57626 213979 57629
rect 116301 57624 119692 57626
rect 116301 57568 116306 57624
rect 116362 57568 119692 57624
rect 116301 57566 119692 57568
rect 211508 57624 213979 57626
rect 211508 57568 213918 57624
rect 213974 57568 213979 57624
rect 211508 57566 213979 57568
rect 116301 57563 116367 57566
rect 213913 57563 213979 57566
rect 227437 57082 227503 57085
rect 227437 57080 230092 57082
rect 227437 57024 227442 57080
rect 227498 57024 230092 57080
rect 227437 57022 230092 57024
rect 227437 57019 227503 57022
rect 94313 56946 94379 56949
rect 91908 56944 94379 56946
rect 91908 56888 94318 56944
rect 94374 56888 94379 56944
rect 91908 56886 94379 56888
rect 94313 56883 94379 56886
rect 214005 56810 214071 56813
rect 211508 56808 214071 56810
rect 211508 56752 214010 56808
rect 214066 56752 214071 56808
rect 211508 56750 214071 56752
rect 214005 56747 214071 56750
rect 116301 56538 116367 56541
rect 116301 56536 119692 56538
rect 116301 56480 116306 56536
rect 116362 56480 119692 56536
rect 116301 56478 119692 56480
rect 116301 56475 116367 56478
rect 227253 56402 227319 56405
rect 227253 56400 230092 56402
rect 227253 56344 227258 56400
rect 227314 56344 230092 56400
rect 227253 56342 230092 56344
rect 227253 56339 227319 56342
rect 95141 55994 95207 55997
rect 215109 55994 215175 55997
rect 91908 55992 95207 55994
rect 91908 55936 95146 55992
rect 95202 55936 95207 55992
rect 91908 55934 95207 55936
rect 211508 55992 215175 55994
rect 211508 55936 215114 55992
rect 215170 55936 215175 55992
rect 211508 55934 215175 55936
rect 95141 55931 95207 55934
rect 215109 55931 215175 55934
rect 227437 55722 227503 55725
rect 227437 55720 230092 55722
rect 227437 55664 227442 55720
rect 227498 55664 230092 55720
rect 227437 55662 230092 55664
rect 227437 55659 227503 55662
rect 116393 55314 116459 55317
rect 116393 55312 119692 55314
rect 116393 55256 116398 55312
rect 116454 55256 119692 55312
rect 116393 55254 119692 55256
rect 116393 55251 116459 55254
rect 94681 55178 94747 55181
rect 214741 55178 214807 55181
rect 91908 55176 94747 55178
rect 91908 55120 94686 55176
rect 94742 55120 94747 55176
rect 91908 55118 94747 55120
rect 211508 55176 214807 55178
rect 211508 55120 214746 55176
rect 214802 55120 214807 55176
rect 211508 55118 214807 55120
rect 94681 55115 94747 55118
rect 214741 55115 214807 55118
rect 227437 55178 227503 55181
rect 227437 55176 230092 55178
rect 227437 55120 227442 55176
rect 227498 55120 230092 55176
rect 227437 55118 230092 55120
rect 227437 55115 227503 55118
rect 215109 54498 215175 54501
rect 211508 54496 215175 54498
rect 211508 54440 215114 54496
rect 215170 54440 215175 54496
rect 211508 54438 215175 54440
rect 215109 54435 215175 54438
rect 226517 54498 226583 54501
rect 226517 54496 230092 54498
rect 226517 54440 226522 54496
rect 226578 54440 230092 54496
rect 226517 54438 230092 54440
rect 226517 54435 226583 54438
rect 94497 54226 94563 54229
rect 91908 54224 94563 54226
rect 91908 54168 94502 54224
rect 94558 54168 94563 54224
rect 91908 54166 94563 54168
rect 94497 54163 94563 54166
rect 116393 54226 116459 54229
rect 116393 54224 119692 54226
rect 116393 54168 116398 54224
rect 116454 54168 119692 54224
rect 116393 54166 119692 54168
rect 116393 54163 116459 54166
rect 227437 53818 227503 53821
rect 227437 53816 230092 53818
rect 227437 53760 227442 53816
rect 227498 53760 230092 53816
rect 227437 53758 230092 53760
rect 227437 53755 227503 53758
rect 214741 53682 214807 53685
rect 211508 53680 214807 53682
rect 211508 53624 214746 53680
rect 214802 53624 214807 53680
rect 211508 53622 214807 53624
rect 214741 53619 214807 53622
rect 94957 53274 95023 53277
rect 91908 53272 95023 53274
rect 91908 53216 94962 53272
rect 95018 53216 95023 53272
rect 91908 53214 95023 53216
rect 94957 53211 95023 53214
rect 226517 53138 226583 53141
rect 226517 53136 230092 53138
rect 226517 53080 226522 53136
rect 226578 53080 230092 53136
rect 226517 53078 230092 53080
rect 226517 53075 226583 53078
rect 116393 53002 116459 53005
rect 116393 53000 119692 53002
rect 116393 52944 116398 53000
rect 116454 52944 119692 53000
rect 116393 52942 119692 52944
rect 116393 52939 116459 52942
rect 215109 52866 215175 52869
rect 211508 52864 215175 52866
rect 211508 52808 215114 52864
rect 215170 52808 215175 52864
rect 211508 52806 215175 52808
rect 215109 52803 215175 52806
rect 583520 52716 584960 52956
rect 95049 52458 95115 52461
rect 91908 52456 95115 52458
rect 91908 52400 95054 52456
rect 95110 52400 95115 52456
rect 91908 52398 95115 52400
rect 95049 52395 95115 52398
rect 227253 52458 227319 52461
rect 227253 52456 230092 52458
rect 227253 52400 227258 52456
rect 227314 52400 230092 52456
rect 227253 52398 230092 52400
rect 227253 52395 227319 52398
rect 215109 52050 215175 52053
rect 211508 52048 215175 52050
rect 211508 51992 215114 52048
rect 215170 51992 215175 52048
rect 211508 51990 215175 51992
rect 215109 51987 215175 51990
rect 115933 51914 115999 51917
rect 227437 51914 227503 51917
rect 115933 51912 119692 51914
rect 115933 51856 115938 51912
rect 115994 51856 119692 51912
rect 115933 51854 119692 51856
rect 227437 51912 230092 51914
rect 227437 51856 227442 51912
rect 227498 51856 230092 51912
rect 227437 51854 230092 51856
rect 115933 51851 115999 51854
rect 227437 51851 227503 51854
rect 94405 51506 94471 51509
rect 91908 51504 94471 51506
rect 91908 51448 94410 51504
rect 94466 51448 94471 51504
rect 91908 51446 94471 51448
rect 94405 51443 94471 51446
rect 214097 51370 214163 51373
rect 211508 51368 214163 51370
rect 211508 51312 214102 51368
rect 214158 51312 214163 51368
rect 211508 51310 214163 51312
rect 214097 51307 214163 51310
rect 227529 51234 227595 51237
rect 227529 51232 230092 51234
rect 227529 51176 227534 51232
rect 227590 51176 230092 51232
rect 227529 51174 230092 51176
rect 227529 51171 227595 51174
rect 93853 50690 93919 50693
rect 91908 50688 93919 50690
rect 91908 50632 93858 50688
rect 93914 50632 93919 50688
rect 91908 50630 93919 50632
rect 93853 50627 93919 50630
rect 116393 50690 116459 50693
rect 116393 50688 119692 50690
rect 116393 50632 116398 50688
rect 116454 50632 119692 50688
rect 116393 50630 119692 50632
rect 116393 50627 116459 50630
rect 215201 50554 215267 50557
rect 211508 50552 215267 50554
rect 211508 50496 215206 50552
rect 215262 50496 215267 50552
rect 211508 50494 215267 50496
rect 215201 50491 215267 50494
rect 226609 50554 226675 50557
rect 226609 50552 230092 50554
rect 226609 50496 226614 50552
rect 226670 50496 230092 50552
rect 226609 50494 230092 50496
rect 226609 50491 226675 50494
rect -960 50146 480 50236
rect 2773 50146 2839 50149
rect -960 50144 2839 50146
rect -960 50088 2778 50144
rect 2834 50088 2839 50144
rect -960 50086 2839 50088
rect -960 49996 480 50086
rect 2773 50083 2839 50086
rect 226977 49874 227043 49877
rect 411897 49874 411963 49877
rect 226977 49872 230092 49874
rect 226977 49816 226982 49872
rect 227038 49816 230092 49872
rect 226977 49814 230092 49816
rect 411897 49872 414092 49874
rect 411897 49816 411902 49872
rect 411958 49816 414092 49872
rect 411897 49814 414092 49816
rect 226977 49811 227043 49814
rect 411897 49811 411963 49814
rect 93945 49738 94011 49741
rect 215109 49738 215175 49741
rect 91908 49736 94011 49738
rect 91908 49680 93950 49736
rect 94006 49680 94011 49736
rect 91908 49678 94011 49680
rect 211508 49736 215175 49738
rect 211508 49680 215114 49736
rect 215170 49680 215175 49736
rect 211508 49678 215175 49680
rect 93945 49675 94011 49678
rect 215109 49675 215175 49678
rect 116393 49466 116459 49469
rect 116393 49464 119692 49466
rect 116393 49408 116398 49464
rect 116454 49408 119692 49464
rect 116393 49406 119692 49408
rect 116393 49403 116459 49406
rect 226701 49330 226767 49333
rect 226701 49328 230092 49330
rect 226701 49272 226706 49328
rect 226762 49272 230092 49328
rect 226701 49270 230092 49272
rect 226701 49267 226767 49270
rect 94037 48922 94103 48925
rect 215109 48922 215175 48925
rect 91908 48920 94103 48922
rect 91908 48864 94042 48920
rect 94098 48864 94103 48920
rect 91908 48862 94103 48864
rect 211508 48920 215175 48922
rect 211508 48864 215114 48920
rect 215170 48864 215175 48920
rect 211508 48862 215175 48864
rect 94037 48859 94103 48862
rect 215109 48859 215175 48862
rect 226793 48650 226859 48653
rect 226793 48648 230092 48650
rect 226793 48592 226798 48648
rect 226854 48592 230092 48648
rect 226793 48590 230092 48592
rect 226793 48587 226859 48590
rect 116117 48378 116183 48381
rect 116117 48376 119692 48378
rect 116117 48320 116122 48376
rect 116178 48320 119692 48376
rect 116117 48318 119692 48320
rect 116117 48315 116183 48318
rect 214741 48106 214807 48109
rect 211508 48104 214807 48106
rect 211508 48048 214746 48104
rect 214802 48048 214807 48104
rect 211508 48046 214807 48048
rect 214741 48043 214807 48046
rect 94773 47970 94839 47973
rect 91908 47968 94839 47970
rect 91908 47912 94778 47968
rect 94834 47912 94839 47968
rect 91908 47910 94839 47912
rect 94773 47907 94839 47910
rect 226333 47970 226399 47973
rect 226333 47968 230092 47970
rect 226333 47912 226338 47968
rect 226394 47912 230092 47968
rect 226333 47910 230092 47912
rect 226333 47907 226399 47910
rect 214005 47426 214071 47429
rect 211508 47424 214071 47426
rect 211508 47368 214010 47424
rect 214066 47368 214071 47424
rect 211508 47366 214071 47368
rect 214005 47363 214071 47366
rect 226517 47290 226583 47293
rect 226517 47288 230092 47290
rect 226517 47232 226522 47288
rect 226578 47232 230092 47288
rect 226517 47230 230092 47232
rect 226517 47227 226583 47230
rect 116393 47154 116459 47157
rect 116393 47152 119692 47154
rect 116393 47096 116398 47152
rect 116454 47096 119692 47152
rect 116393 47094 119692 47096
rect 116393 47091 116459 47094
rect 95141 47018 95207 47021
rect 91908 47016 95207 47018
rect 91908 46960 95146 47016
rect 95202 46960 95207 47016
rect 91908 46958 95207 46960
rect 95141 46955 95207 46958
rect 215201 46610 215267 46613
rect 211508 46608 215267 46610
rect 211508 46552 215206 46608
rect 215262 46552 215267 46608
rect 211508 46550 215267 46552
rect 215201 46547 215267 46550
rect 227529 46610 227595 46613
rect 227529 46608 230092 46610
rect 227529 46552 227534 46608
rect 227590 46552 230092 46608
rect 227529 46550 230092 46552
rect 227529 46547 227595 46550
rect 94221 46202 94287 46205
rect 91908 46200 94287 46202
rect 91908 46144 94226 46200
rect 94282 46144 94287 46200
rect 91908 46142 94287 46144
rect 94221 46139 94287 46142
rect 116393 46066 116459 46069
rect 227621 46066 227687 46069
rect 116393 46064 119692 46066
rect 116393 46008 116398 46064
rect 116454 46008 119692 46064
rect 116393 46006 119692 46008
rect 227621 46064 230092 46066
rect 227621 46008 227626 46064
rect 227682 46008 230092 46064
rect 227621 46006 230092 46008
rect 116393 46003 116459 46006
rect 227621 46003 227687 46006
rect 215109 45794 215175 45797
rect 211508 45792 215175 45794
rect 211508 45736 215114 45792
rect 215170 45736 215175 45792
rect 211508 45734 215175 45736
rect 215109 45731 215175 45734
rect 227345 45386 227411 45389
rect 227345 45384 230092 45386
rect 227345 45328 227350 45384
rect 227406 45328 230092 45384
rect 227345 45326 230092 45328
rect 227345 45323 227411 45326
rect 95049 45250 95115 45253
rect 91908 45248 95115 45250
rect 91908 45192 95054 45248
rect 95110 45192 95115 45248
rect 91908 45190 95115 45192
rect 95049 45187 95115 45190
rect 215201 44978 215267 44981
rect 211508 44976 215267 44978
rect 211508 44920 215206 44976
rect 215262 44920 215267 44976
rect 211508 44918 215267 44920
rect 215201 44915 215267 44918
rect 116393 44842 116459 44845
rect 116393 44840 119692 44842
rect 116393 44784 116398 44840
rect 116454 44784 119692 44840
rect 116393 44782 119692 44784
rect 116393 44779 116459 44782
rect 227437 44706 227503 44709
rect 227437 44704 230092 44706
rect 227437 44648 227442 44704
rect 227498 44648 230092 44704
rect 227437 44646 230092 44648
rect 227437 44643 227503 44646
rect 94405 44434 94471 44437
rect 91908 44432 94471 44434
rect 91908 44376 94410 44432
rect 94466 44376 94471 44432
rect 91908 44374 94471 44376
rect 94405 44371 94471 44374
rect 215109 44298 215175 44301
rect 211508 44296 215175 44298
rect 211508 44240 215114 44296
rect 215170 44240 215175 44296
rect 211508 44238 215175 44240
rect 215109 44235 215175 44238
rect 226701 44026 226767 44029
rect 226701 44024 230092 44026
rect 226701 43968 226706 44024
rect 226762 43968 230092 44024
rect 226701 43966 230092 43968
rect 226701 43963 226767 43966
rect 115933 43618 115999 43621
rect 115933 43616 119692 43618
rect 115933 43560 115938 43616
rect 115994 43560 119692 43616
rect 115933 43558 119692 43560
rect 115933 43555 115999 43558
rect 94497 43482 94563 43485
rect 214373 43482 214439 43485
rect 91908 43480 94563 43482
rect 91908 43424 94502 43480
rect 94558 43424 94563 43480
rect 91908 43422 94563 43424
rect 211508 43480 214439 43482
rect 211508 43424 214378 43480
rect 214434 43424 214439 43480
rect 211508 43422 214439 43424
rect 94497 43419 94563 43422
rect 214373 43419 214439 43422
rect 227069 43482 227135 43485
rect 227069 43480 230092 43482
rect 227069 43424 227074 43480
rect 227130 43424 230092 43480
rect 227069 43422 230092 43424
rect 227069 43419 227135 43422
rect 227253 42802 227319 42805
rect 227253 42800 230092 42802
rect 227253 42744 227258 42800
rect 227314 42744 230092 42800
rect 227253 42742 230092 42744
rect 227253 42739 227319 42742
rect 214097 42666 214163 42669
rect 211508 42664 214163 42666
rect 211508 42608 214102 42664
rect 214158 42608 214163 42664
rect 211508 42606 214163 42608
rect 214097 42603 214163 42606
rect 94129 42530 94195 42533
rect 91908 42528 94195 42530
rect 91908 42472 94134 42528
rect 94190 42472 94195 42528
rect 91908 42470 94195 42472
rect 94129 42467 94195 42470
rect 116393 42530 116459 42533
rect 116393 42528 119692 42530
rect 116393 42472 116398 42528
rect 116454 42472 119692 42528
rect 116393 42470 119692 42472
rect 116393 42467 116459 42470
rect 227437 42122 227503 42125
rect 227437 42120 230092 42122
rect 227437 42064 227442 42120
rect 227498 42064 230092 42120
rect 227437 42062 230092 42064
rect 227437 42059 227503 42062
rect 215109 41850 215175 41853
rect 211508 41848 215175 41850
rect 211508 41792 215114 41848
rect 215170 41792 215175 41848
rect 211508 41790 215175 41792
rect 215109 41787 215175 41790
rect 93945 41714 94011 41717
rect 91908 41712 94011 41714
rect 91908 41656 93950 41712
rect 94006 41656 94011 41712
rect 91908 41654 94011 41656
rect 93945 41651 94011 41654
rect 227529 41442 227595 41445
rect 227529 41440 230092 41442
rect 227529 41384 227534 41440
rect 227590 41384 230092 41440
rect 227529 41382 230092 41384
rect 227529 41379 227595 41382
rect 116301 41306 116367 41309
rect 116301 41304 119692 41306
rect 116301 41248 116306 41304
rect 116362 41248 119692 41304
rect 116301 41246 119692 41248
rect 116301 41243 116367 41246
rect 214649 41170 214715 41173
rect 211508 41168 214715 41170
rect 211508 41112 214654 41168
rect 214710 41112 214715 41168
rect 211508 41110 214715 41112
rect 214649 41107 214715 41110
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect 94773 40762 94839 40765
rect 91908 40760 94839 40762
rect 91908 40704 94778 40760
rect 94834 40704 94839 40760
rect 91908 40702 94839 40704
rect 94773 40699 94839 40702
rect 226425 40762 226491 40765
rect 226425 40760 230092 40762
rect 226425 40704 226430 40760
rect 226486 40704 230092 40760
rect 226425 40702 230092 40704
rect 226425 40699 226491 40702
rect 215109 40354 215175 40357
rect 211508 40352 215175 40354
rect 211508 40296 215114 40352
rect 215170 40296 215175 40352
rect 211508 40294 215175 40296
rect 215109 40291 215175 40294
rect 116393 40218 116459 40221
rect 226333 40218 226399 40221
rect 116393 40216 119692 40218
rect 116393 40160 116398 40216
rect 116454 40160 119692 40216
rect 116393 40158 119692 40160
rect 226333 40216 230092 40218
rect 226333 40160 226338 40216
rect 226394 40160 230092 40216
rect 226333 40158 230092 40160
rect 116393 40155 116459 40158
rect 226333 40155 226399 40158
rect 94589 39946 94655 39949
rect 91908 39944 94655 39946
rect 91908 39888 94594 39944
rect 94650 39888 94655 39944
rect 91908 39886 94655 39888
rect 94589 39883 94655 39886
rect 214557 39538 214623 39541
rect 211508 39536 214623 39538
rect 211508 39480 214562 39536
rect 214618 39480 214623 39536
rect 211508 39478 214623 39480
rect 214557 39475 214623 39478
rect 226609 39538 226675 39541
rect 226609 39536 230092 39538
rect 226609 39480 226614 39536
rect 226670 39480 230092 39536
rect 226609 39478 230092 39480
rect 226609 39475 226675 39478
rect 95141 38994 95207 38997
rect 91908 38992 95207 38994
rect 91908 38936 95146 38992
rect 95202 38936 95207 38992
rect 91908 38934 95207 38936
rect 95141 38931 95207 38934
rect 116393 38994 116459 38997
rect 116393 38992 119692 38994
rect 116393 38936 116398 38992
rect 116454 38936 119692 38992
rect 116393 38934 119692 38936
rect 116393 38931 116459 38934
rect 227069 38858 227135 38861
rect 227069 38856 230092 38858
rect 227069 38800 227074 38856
rect 227130 38800 230092 38856
rect 227069 38798 230092 38800
rect 227069 38795 227135 38798
rect 215109 38722 215175 38725
rect 563697 38722 563763 38725
rect 211508 38720 215175 38722
rect 211508 38664 215114 38720
rect 215170 38664 215175 38720
rect 211508 38662 215175 38664
rect 561108 38720 563763 38722
rect 561108 38664 563702 38720
rect 563758 38664 563763 38720
rect 561108 38662 563763 38664
rect 215109 38659 215175 38662
rect 563697 38659 563763 38662
rect 94497 38178 94563 38181
rect 91908 38176 94563 38178
rect 91908 38120 94502 38176
rect 94558 38120 94563 38176
rect 91908 38118 94563 38120
rect 94497 38115 94563 38118
rect 227437 38178 227503 38181
rect 227437 38176 230092 38178
rect 227437 38120 227442 38176
rect 227498 38120 230092 38176
rect 227437 38118 230092 38120
rect 227437 38115 227503 38118
rect 215109 38042 215175 38045
rect 211508 38040 215175 38042
rect 211508 37984 215114 38040
rect 215170 37984 215175 38040
rect 211508 37982 215175 37984
rect 215109 37979 215175 37982
rect 116393 37770 116459 37773
rect 116393 37768 119692 37770
rect 116393 37712 116398 37768
rect 116454 37712 119692 37768
rect 116393 37710 119692 37712
rect 116393 37707 116459 37710
rect 226701 37634 226767 37637
rect 226701 37632 230092 37634
rect 226701 37576 226706 37632
rect 226762 37576 230092 37632
rect 226701 37574 230092 37576
rect 226701 37571 226767 37574
rect 95049 37226 95115 37229
rect 214097 37226 214163 37229
rect 91908 37224 95115 37226
rect 91908 37168 95054 37224
rect 95110 37168 95115 37224
rect 91908 37166 95115 37168
rect 211508 37224 214163 37226
rect 211508 37168 214102 37224
rect 214158 37168 214163 37224
rect 211508 37166 214163 37168
rect 95049 37163 95115 37166
rect 214097 37163 214163 37166
rect 227529 36954 227595 36957
rect 227529 36952 230092 36954
rect 227529 36896 227534 36952
rect 227590 36896 230092 36952
rect 227529 36894 230092 36896
rect 227529 36891 227595 36894
rect 116393 36682 116459 36685
rect 116393 36680 119692 36682
rect 116393 36624 116398 36680
rect 116454 36624 119692 36680
rect 116393 36622 119692 36624
rect 116393 36619 116459 36622
rect 215109 36410 215175 36413
rect 211508 36408 215175 36410
rect 211508 36352 215114 36408
rect 215170 36352 215175 36408
rect 211508 36350 215175 36352
rect 215109 36347 215175 36350
rect 94589 36274 94655 36277
rect 91908 36272 94655 36274
rect 91908 36216 94594 36272
rect 94650 36216 94655 36272
rect 91908 36214 94655 36216
rect 94589 36211 94655 36214
rect 227437 36274 227503 36277
rect 227437 36272 230092 36274
rect 227437 36216 227442 36272
rect 227498 36216 230092 36272
rect 227437 36214 230092 36216
rect 227437 36211 227503 36214
rect -960 35866 480 35956
rect 3509 35866 3575 35869
rect -960 35864 3575 35866
rect -960 35808 3514 35864
rect 3570 35808 3575 35864
rect -960 35806 3575 35808
rect -960 35716 480 35806
rect 3509 35803 3575 35806
rect 214649 35594 214715 35597
rect 211508 35592 214715 35594
rect 211508 35536 214654 35592
rect 214710 35536 214715 35592
rect 211508 35534 214715 35536
rect 214649 35531 214715 35534
rect 226701 35594 226767 35597
rect 226701 35592 230092 35594
rect 226701 35536 226706 35592
rect 226762 35536 230092 35592
rect 226701 35534 230092 35536
rect 226701 35531 226767 35534
rect 93853 35458 93919 35461
rect 91908 35456 93919 35458
rect 91908 35400 93858 35456
rect 93914 35400 93919 35456
rect 91908 35398 93919 35400
rect 93853 35395 93919 35398
rect 116393 35458 116459 35461
rect 116393 35456 119692 35458
rect 116393 35400 116398 35456
rect 116454 35400 119692 35456
rect 116393 35398 119692 35400
rect 116393 35395 116459 35398
rect 215109 34914 215175 34917
rect 211508 34912 215175 34914
rect 211508 34856 215114 34912
rect 215170 34856 215175 34912
rect 211508 34854 215175 34856
rect 215109 34851 215175 34854
rect 227437 34914 227503 34917
rect 227437 34912 230092 34914
rect 227437 34856 227442 34912
rect 227498 34856 230092 34912
rect 227437 34854 230092 34856
rect 227437 34851 227503 34854
rect 93945 34506 94011 34509
rect 91908 34504 94011 34506
rect 91908 34448 93950 34504
rect 94006 34448 94011 34504
rect 91908 34446 94011 34448
rect 93945 34443 94011 34446
rect 116301 34370 116367 34373
rect 227437 34370 227503 34373
rect 116301 34368 119692 34370
rect 116301 34312 116306 34368
rect 116362 34312 119692 34368
rect 116301 34310 119692 34312
rect 227437 34368 230092 34370
rect 227437 34312 227442 34368
rect 227498 34312 230092 34368
rect 227437 34310 230092 34312
rect 116301 34307 116367 34310
rect 227437 34307 227503 34310
rect 214557 34098 214623 34101
rect 211508 34096 214623 34098
rect 211508 34040 214562 34096
rect 214618 34040 214623 34096
rect 211508 34038 214623 34040
rect 214557 34035 214623 34038
rect 95141 33690 95207 33693
rect 91908 33688 95207 33690
rect 91908 33632 95146 33688
rect 95202 33632 95207 33688
rect 91908 33630 95207 33632
rect 95141 33627 95207 33630
rect 227345 33690 227411 33693
rect 227345 33688 230092 33690
rect 227345 33632 227350 33688
rect 227406 33632 230092 33688
rect 227345 33630 230092 33632
rect 227345 33627 227411 33630
rect 215109 33282 215175 33285
rect 211508 33280 215175 33282
rect 211508 33224 215114 33280
rect 215170 33224 215175 33280
rect 211508 33222 215175 33224
rect 215109 33219 215175 33222
rect 116393 33146 116459 33149
rect 116393 33144 119692 33146
rect 116393 33088 116398 33144
rect 116454 33088 119692 33144
rect 116393 33086 119692 33088
rect 116393 33083 116459 33086
rect 227437 33010 227503 33013
rect 227437 33008 230092 33010
rect 227437 32952 227442 33008
rect 227498 32952 230092 33008
rect 227437 32950 230092 32952
rect 227437 32947 227503 32950
rect 95141 32738 95207 32741
rect 91908 32736 95207 32738
rect 91908 32680 95146 32736
rect 95202 32680 95207 32736
rect 91908 32678 95207 32680
rect 95141 32675 95207 32678
rect 215109 32466 215175 32469
rect 211508 32464 215175 32466
rect 211508 32408 215114 32464
rect 215170 32408 215175 32464
rect 211508 32406 215175 32408
rect 215109 32403 215175 32406
rect 227529 32330 227595 32333
rect 227529 32328 230092 32330
rect 227529 32272 227534 32328
rect 227590 32272 230092 32328
rect 227529 32270 230092 32272
rect 227529 32267 227595 32270
rect 116393 32058 116459 32061
rect 116393 32056 119692 32058
rect 116393 32000 116398 32056
rect 116454 32000 119692 32056
rect 116393 31998 119692 32000
rect 116393 31995 116459 31998
rect 95141 31922 95207 31925
rect 91908 31920 95207 31922
rect 91908 31864 95146 31920
rect 95202 31864 95207 31920
rect 91908 31862 95207 31864
rect 95141 31859 95207 31862
rect 32305 31788 32371 31789
rect 32254 31786 32260 31788
rect 32214 31726 32260 31786
rect 32324 31784 32371 31788
rect 213913 31786 213979 31789
rect 32366 31728 32371 31784
rect 32254 31724 32260 31726
rect 32324 31724 32371 31728
rect 211508 31784 213979 31786
rect 211508 31728 213918 31784
rect 213974 31728 213979 31784
rect 211508 31726 213979 31728
rect 32305 31723 32371 31724
rect 213913 31723 213979 31726
rect 227437 31786 227503 31789
rect 227437 31784 230092 31786
rect 227437 31728 227442 31784
rect 227498 31728 230092 31784
rect 227437 31726 230092 31728
rect 227437 31723 227503 31726
rect 119981 30290 120047 30293
rect 231945 30290 232011 30293
rect 284569 30290 284635 30293
rect 119981 30288 284635 30290
rect 119981 30232 119986 30288
rect 120042 30232 231950 30288
rect 232006 30232 284574 30288
rect 284630 30232 284635 30288
rect 119981 30230 284635 30232
rect 119981 30227 120047 30230
rect 231945 30227 232011 30230
rect 284569 30227 284635 30230
rect 580901 29338 580967 29341
rect 583520 29338 584960 29428
rect 580901 29336 584960 29338
rect 580901 29280 580906 29336
rect 580962 29280 584960 29336
rect 580901 29278 584960 29280
rect 580901 29275 580967 29278
rect 583520 29188 584960 29278
rect 411253 27570 411319 27573
rect 411253 27568 414092 27570
rect 411253 27512 411258 27568
rect 411314 27512 414092 27568
rect 411253 27510 414092 27512
rect 411253 27507 411319 27510
rect -960 21450 480 21540
rect 2773 21450 2839 21453
rect -960 21448 2839 21450
rect -960 21392 2778 21448
rect 2834 21392 2839 21448
rect -960 21390 2839 21392
rect -960 21300 480 21390
rect 2773 21387 2839 21390
rect 583520 17492 584960 17732
rect 144177 14650 144243 14653
rect 419533 14650 419599 14653
rect 144177 14648 419599 14650
rect 144177 14592 144182 14648
rect 144238 14592 419538 14648
rect 419594 14592 419599 14648
rect 144177 14590 419599 14592
rect 144177 14587 144243 14590
rect 419533 14587 419599 14590
rect 140681 14514 140747 14517
rect 418337 14514 418403 14517
rect 140681 14512 418403 14514
rect 140681 14456 140686 14512
rect 140742 14456 418342 14512
rect 418398 14456 418403 14512
rect 140681 14454 418403 14456
rect 140681 14451 140747 14454
rect 418337 14451 418403 14454
rect 422293 13834 422359 13837
rect 425421 13834 425487 13837
rect 422293 13832 425487 13834
rect 422293 13776 422298 13832
rect 422354 13776 425426 13832
rect 425482 13776 425487 13832
rect 422293 13774 425487 13776
rect 422293 13771 422359 13774
rect 425421 13771 425487 13774
rect 250437 13426 250503 13429
rect 430297 13426 430363 13429
rect 250437 13424 430363 13426
rect 250437 13368 250442 13424
rect 250498 13368 430302 13424
rect 430358 13368 430363 13424
rect 250437 13366 430363 13368
rect 250437 13363 250503 13366
rect 430297 13363 430363 13366
rect 243537 13290 243603 13293
rect 427997 13290 428063 13293
rect 243537 13288 428063 13290
rect 243537 13232 243542 13288
rect 243598 13232 428002 13288
rect 428058 13232 428063 13288
rect 243537 13230 428063 13232
rect 243537 13227 243603 13230
rect 427997 13227 428063 13230
rect 239397 13154 239463 13157
rect 425697 13154 425763 13157
rect 239397 13152 425763 13154
rect 239397 13096 239402 13152
rect 239458 13096 425702 13152
rect 425758 13096 425763 13152
rect 239397 13094 425763 13096
rect 239397 13091 239463 13094
rect 425697 13091 425763 13094
rect 232497 13018 232563 13021
rect 426801 13018 426867 13021
rect 232497 13016 426867 13018
rect 232497 12960 232502 13016
rect 232558 12960 426806 13016
rect 426862 12960 426867 13016
rect 232497 12958 426867 12960
rect 232497 12955 232563 12958
rect 426801 12955 426867 12958
rect 410425 12882 410491 12885
rect 412541 12882 412607 12885
rect 410425 12880 412607 12882
rect 410425 12824 410430 12880
rect 410486 12824 412546 12880
rect 412602 12824 412607 12880
rect 410425 12822 412607 12824
rect 410425 12819 410491 12822
rect 412541 12819 412607 12822
rect 422293 12882 422359 12885
rect 431861 12882 431927 12885
rect 422293 12880 431927 12882
rect 422293 12824 422298 12880
rect 422354 12824 431866 12880
rect 431922 12824 431927 12880
rect 422293 12822 431927 12824
rect 422293 12819 422359 12822
rect 431861 12819 431927 12822
rect 246297 12202 246363 12205
rect 422569 12202 422635 12205
rect 246297 12200 422635 12202
rect 246297 12144 246302 12200
rect 246358 12144 422574 12200
rect 422630 12144 422635 12200
rect 246297 12142 422635 12144
rect 246297 12139 246363 12142
rect 422569 12139 422635 12142
rect 171777 12066 171843 12069
rect 428733 12066 428799 12069
rect 171777 12064 428799 12066
rect 171777 12008 171782 12064
rect 171838 12008 428738 12064
rect 428794 12008 428799 12064
rect 171777 12006 428799 12008
rect 171777 12003 171843 12006
rect 428733 12003 428799 12006
rect 164693 11930 164759 11933
rect 426433 11930 426499 11933
rect 164693 11928 426499 11930
rect 164693 11872 164698 11928
rect 164754 11872 426438 11928
rect 426494 11872 426499 11928
rect 164693 11870 426499 11872
rect 164693 11867 164759 11870
rect 426433 11867 426499 11870
rect 156321 11794 156387 11797
rect 423765 11794 423831 11797
rect 156321 11792 423831 11794
rect 156321 11736 156326 11792
rect 156382 11736 423770 11792
rect 423826 11736 423831 11792
rect 156321 11734 423831 11736
rect 156321 11731 156387 11734
rect 423765 11731 423831 11734
rect 128997 11658 129063 11661
rect 414933 11658 414999 11661
rect 128997 11656 414999 11658
rect 128997 11600 129002 11656
rect 129058 11600 414938 11656
rect 414994 11600 414999 11656
rect 128997 11598 414999 11600
rect 128997 11595 129063 11598
rect 414933 11595 414999 11598
rect 145649 10570 145715 10573
rect 420269 10570 420335 10573
rect 145649 10568 420335 10570
rect 145649 10512 145654 10568
rect 145710 10512 420274 10568
rect 420330 10512 420335 10568
rect 145649 10510 420335 10512
rect 145649 10507 145715 10510
rect 420269 10507 420335 10510
rect 142061 10434 142127 10437
rect 419165 10434 419231 10437
rect 142061 10432 419231 10434
rect 142061 10376 142066 10432
rect 142122 10376 419170 10432
rect 419226 10376 419231 10432
rect 142061 10374 419231 10376
rect 142061 10371 142127 10374
rect 419165 10371 419231 10374
rect 136081 10298 136147 10301
rect 417233 10298 417299 10301
rect 136081 10296 417299 10298
rect 136081 10240 136086 10296
rect 136142 10240 417238 10296
rect 417294 10240 417299 10296
rect 136081 10238 417299 10240
rect 136081 10235 136147 10238
rect 417233 10235 417299 10238
rect 435449 9890 435515 9893
rect 434670 9888 435515 9890
rect 434670 9832 435454 9888
rect 435510 9832 435515 9888
rect 434670 9830 435515 9832
rect 184565 9754 184631 9757
rect 184749 9754 184815 9757
rect 184565 9752 184815 9754
rect 184565 9696 184570 9752
rect 184626 9696 184754 9752
rect 184810 9696 184815 9752
rect 184565 9694 184815 9696
rect 434670 9754 434730 9830
rect 435449 9827 435515 9830
rect 446949 9890 447015 9893
rect 446949 9888 447426 9890
rect 446949 9832 446954 9888
rect 447010 9832 447426 9888
rect 446949 9830 447426 9832
rect 446949 9827 447015 9830
rect 434805 9754 434871 9757
rect 434670 9752 434871 9754
rect 434670 9696 434810 9752
rect 434866 9696 434871 9752
rect 434670 9694 434871 9696
rect 184565 9691 184631 9694
rect 184749 9691 184815 9694
rect 434805 9691 434871 9694
rect 447225 9754 447291 9757
rect 447366 9754 447426 9830
rect 447225 9752 447426 9754
rect 447225 9696 447230 9752
rect 447286 9696 447426 9752
rect 447225 9694 447426 9696
rect 447225 9691 447291 9694
rect 206277 9210 206343 9213
rect 439865 9210 439931 9213
rect 206277 9208 439931 9210
rect 206277 9152 206282 9208
rect 206338 9152 439870 9208
rect 439926 9152 439931 9208
rect 206277 9150 439931 9152
rect 206277 9147 206343 9150
rect 439865 9147 439931 9150
rect 138473 9074 138539 9077
rect 417693 9074 417759 9077
rect 138473 9072 417759 9074
rect 138473 9016 138478 9072
rect 138534 9016 417698 9072
rect 417754 9016 417759 9072
rect 138473 9014 417759 9016
rect 138473 9011 138539 9014
rect 417693 9011 417759 9014
rect 134885 8938 134951 8941
rect 416865 8938 416931 8941
rect 134885 8936 416931 8938
rect 134885 8880 134890 8936
rect 134946 8880 416870 8936
rect 416926 8880 416931 8936
rect 134885 8878 416931 8880
rect 134885 8875 134951 8878
rect 416865 8875 416931 8878
rect 158713 8258 158779 8261
rect 424501 8258 424567 8261
rect 158713 8256 424567 8258
rect 158713 8200 158718 8256
rect 158774 8200 424506 8256
rect 424562 8200 424567 8256
rect 158713 8198 424567 8200
rect 158713 8195 158779 8198
rect 424501 8195 424567 8198
rect 155125 8122 155191 8125
rect 423397 8122 423463 8125
rect 155125 8120 423463 8122
rect 155125 8064 155130 8120
rect 155186 8064 423402 8120
rect 423458 8064 423463 8120
rect 155125 8062 423463 8064
rect 155125 8059 155191 8062
rect 423397 8059 423463 8062
rect 151537 7986 151603 7989
rect 422201 7986 422267 7989
rect 151537 7984 422267 7986
rect 151537 7928 151542 7984
rect 151598 7928 422206 7984
rect 422262 7928 422267 7984
rect 151537 7926 422267 7928
rect 151537 7923 151603 7926
rect 422201 7923 422267 7926
rect 148041 7850 148107 7853
rect 421097 7850 421163 7853
rect 148041 7848 421163 7850
rect 148041 7792 148046 7848
rect 148102 7792 421102 7848
rect 421158 7792 421163 7848
rect 148041 7790 421163 7792
rect 148041 7787 148107 7790
rect 421097 7787 421163 7790
rect 131389 7714 131455 7717
rect 415669 7714 415735 7717
rect 131389 7712 415735 7714
rect 131389 7656 131394 7712
rect 131450 7656 415674 7712
rect 415730 7656 415735 7712
rect 131389 7654 415735 7656
rect 131389 7651 131455 7654
rect 415669 7651 415735 7654
rect 127801 7578 127867 7581
rect 414565 7578 414631 7581
rect 127801 7576 414631 7578
rect 127801 7520 127806 7576
rect 127862 7520 414570 7576
rect 414626 7520 414631 7576
rect 127801 7518 414631 7520
rect 127801 7515 127867 7518
rect 414565 7515 414631 7518
rect -960 7170 480 7260
rect 2773 7170 2839 7173
rect -960 7168 2839 7170
rect -960 7112 2778 7168
rect 2834 7112 2839 7168
rect -960 7110 2839 7112
rect -960 7020 480 7110
rect 2773 7107 2839 7110
rect 283649 6354 283715 6357
rect 463785 6354 463851 6357
rect 283649 6352 463851 6354
rect 283649 6296 283654 6352
rect 283710 6296 463790 6352
rect 463846 6296 463851 6352
rect 283649 6294 463851 6296
rect 283649 6291 283715 6294
rect 463785 6291 463851 6294
rect 140957 6218 141023 6221
rect 418521 6218 418587 6221
rect 140957 6216 418587 6218
rect 140957 6160 140962 6216
rect 141018 6160 418526 6216
rect 418582 6160 418587 6216
rect 140957 6158 418587 6160
rect 140957 6155 141023 6158
rect 418521 6155 418587 6158
rect 583520 5796 584960 6036
rect 212257 5130 212323 5133
rect 441797 5130 441863 5133
rect 212257 5128 441863 5130
rect 212257 5072 212262 5128
rect 212318 5072 441802 5128
rect 441858 5072 441863 5128
rect 212257 5070 441863 5072
rect 212257 5067 212323 5070
rect 441797 5067 441863 5070
rect 205081 4994 205147 4997
rect 438853 4994 438919 4997
rect 205081 4992 438919 4994
rect 205081 4936 205086 4992
rect 205142 4936 438858 4992
rect 438914 4936 438919 4992
rect 205081 4934 438919 4936
rect 205081 4931 205147 4934
rect 438853 4931 438919 4934
rect 12433 4858 12499 4861
rect 128353 4858 128419 4861
rect 12433 4856 128419 4858
rect 12433 4800 12438 4856
rect 12494 4800 128358 4856
rect 128414 4800 128419 4856
rect 12433 4798 128419 4800
rect 12433 4795 12499 4798
rect 128353 4795 128419 4798
rect 201493 4858 201559 4861
rect 437473 4858 437539 4861
rect 201493 4856 437539 4858
rect 201493 4800 201498 4856
rect 201554 4800 437478 4856
rect 437534 4800 437539 4856
rect 201493 4798 437539 4800
rect 201493 4795 201559 4798
rect 437473 4795 437539 4798
rect 122925 4314 122991 4317
rect 125685 4314 125751 4317
rect 122925 4312 125751 4314
rect 122925 4256 122930 4312
rect 122986 4256 125690 4312
rect 125746 4256 125751 4312
rect 122925 4254 125751 4256
rect 122925 4251 122991 4254
rect 125685 4251 125751 4254
rect 113173 3906 113239 3909
rect 118693 3906 118759 3909
rect 113173 3904 118759 3906
rect 113173 3848 113178 3904
rect 113234 3848 118698 3904
rect 118754 3848 118759 3904
rect 113173 3846 118759 3848
rect 113173 3843 113239 3846
rect 118693 3843 118759 3846
rect 421373 3770 421439 3773
rect 426525 3770 426591 3773
rect 421373 3768 426591 3770
rect 421373 3712 421378 3768
rect 421434 3712 426530 3768
rect 426586 3712 426591 3768
rect 421373 3710 426591 3712
rect 421373 3707 421439 3710
rect 426525 3707 426591 3710
rect 113449 3634 113515 3637
rect 116025 3634 116091 3637
rect 113449 3632 116091 3634
rect 113449 3576 113454 3632
rect 113510 3576 116030 3632
rect 116086 3576 116091 3632
rect 113449 3574 116091 3576
rect 113449 3571 113515 3574
rect 116025 3571 116091 3574
rect 129825 3634 129891 3637
rect 133229 3634 133295 3637
rect 129825 3632 133295 3634
rect 129825 3576 129830 3632
rect 129886 3576 133234 3632
rect 133290 3576 133295 3632
rect 129825 3574 133295 3576
rect 129825 3571 129891 3574
rect 133229 3571 133295 3574
rect 182173 3634 182239 3637
rect 182633 3634 182699 3637
rect 182173 3632 182699 3634
rect 182173 3576 182178 3632
rect 182234 3576 182638 3632
rect 182694 3576 182699 3632
rect 182173 3574 182699 3576
rect 182173 3571 182239 3574
rect 182633 3571 182699 3574
rect 293125 3634 293191 3637
rect 431677 3634 431743 3637
rect 293125 3632 431743 3634
rect 293125 3576 293130 3632
rect 293186 3576 431682 3632
rect 431738 3576 431743 3632
rect 293125 3574 431743 3576
rect 293125 3571 293191 3574
rect 431677 3571 431743 3574
rect 285949 3498 286015 3501
rect 430481 3498 430547 3501
rect 285949 3496 430547 3498
rect 285949 3440 285954 3496
rect 286010 3440 430486 3496
rect 430542 3440 430547 3496
rect 285949 3438 430547 3440
rect 285949 3435 286015 3438
rect 430481 3435 430547 3438
rect 25497 3362 25563 3365
rect 138197 3362 138263 3365
rect 25497 3360 138263 3362
rect 25497 3304 25502 3360
rect 25558 3304 138202 3360
rect 138258 3304 138263 3360
rect 25497 3302 138263 3304
rect 25497 3299 25563 3302
rect 138197 3299 138263 3302
rect 278865 3362 278931 3365
rect 429101 3362 429167 3365
rect 278865 3360 429167 3362
rect 278865 3304 278870 3360
rect 278926 3304 429106 3360
rect 429162 3304 429167 3360
rect 278865 3302 429167 3304
rect 278865 3299 278931 3302
rect 429101 3299 429167 3302
rect 342897 2410 342963 2413
rect 347681 2410 347747 2413
rect 342897 2408 347747 2410
rect 342897 2352 342902 2408
rect 342958 2352 347686 2408
rect 347742 2352 347747 2408
rect 342897 2350 347747 2352
rect 342897 2347 342963 2350
rect 347681 2347 347747 2350
rect 415393 2410 415459 2413
rect 424961 2410 425027 2413
rect 415393 2408 425027 2410
rect 415393 2352 415398 2408
rect 415454 2352 424966 2408
rect 425022 2352 425027 2408
rect 415393 2350 425027 2352
rect 415393 2347 415459 2350
rect 424961 2347 425027 2350
rect 434713 2410 434779 2413
rect 442073 2410 442139 2413
rect 434713 2408 442139 2410
rect 434713 2352 434718 2408
rect 434774 2352 442078 2408
rect 442134 2352 442139 2408
rect 434713 2350 442139 2352
rect 434713 2347 434779 2350
rect 442073 2347 442139 2350
rect 381537 2138 381603 2141
rect 386321 2138 386387 2141
rect 381537 2136 386387 2138
rect 381537 2080 381542 2136
rect 381598 2080 386326 2136
rect 386382 2080 386387 2136
rect 381537 2078 386387 2080
rect 381537 2075 381603 2078
rect 386321 2075 386387 2078
<< via3 >>
rect 317092 700572 317156 700636
rect 317276 700436 317340 700500
rect 316908 700300 316972 700364
rect 492444 663852 492508 663916
rect 548380 662084 548444 662148
rect 551324 660044 551388 660108
rect 551508 658820 551572 658884
rect 553348 658140 553412 658204
rect 553532 656916 553596 656980
rect 553716 655692 553780 655756
rect 552796 654468 552860 654532
rect 551324 653108 551388 653172
rect 552060 651476 552124 651540
rect 553900 650796 553964 650860
rect 551324 649028 551388 649092
rect 552244 648348 552308 648412
rect 552428 647124 552492 647188
rect 551324 645764 551388 645828
rect 552612 644676 552676 644740
rect 554084 643452 554148 643516
rect 551324 639644 551388 639708
rect 551508 639508 551572 639572
rect 551324 639372 551388 639436
rect 551324 635972 551388 636036
rect 551876 634884 551940 634948
rect 551324 628008 551388 628012
rect 551324 627952 551374 628008
rect 551374 627952 551388 628008
rect 551324 627948 551388 627952
rect 551692 628008 551756 628012
rect 551692 627952 551706 628008
rect 551706 627952 551756 628008
rect 551692 627948 551756 627952
rect 113404 622372 113468 622436
rect 551324 618624 551388 618628
rect 551324 618568 551374 618624
rect 551374 618568 551388 618624
rect 551324 618564 551388 618568
rect 280660 618292 280724 618356
rect 551324 618292 551388 618356
rect 551692 618292 551756 618356
rect 106228 617612 106292 617676
rect 113404 617612 113468 617676
rect 551324 617536 551388 617540
rect 551324 617480 551374 617536
rect 551374 617480 551388 617536
rect 551324 617476 551388 617480
rect 25452 617340 25516 617404
rect 27660 616796 27724 616860
rect 551324 616388 551388 616452
rect 27476 616116 27540 616180
rect 21220 615708 21284 615772
rect 22140 615708 22204 615772
rect 28580 615708 28644 615772
rect 27292 614892 27356 614956
rect 25268 614348 25332 614412
rect 27108 613804 27172 613868
rect 551324 613804 551388 613868
rect 551324 613668 551388 613732
rect 28212 612716 28276 612780
rect 551508 612308 551572 612372
rect 551692 612308 551756 612372
rect 551324 612172 551388 612236
rect 28028 612036 28092 612100
rect 26924 611356 26988 611420
rect 27844 610812 27908 610876
rect 26740 610132 26804 610196
rect 26004 604692 26068 604756
rect 25820 603604 25884 603668
rect 551508 601156 551572 601220
rect 25636 599932 25700 599996
rect 551324 599992 551388 599996
rect 551324 599936 551374 599992
rect 551374 599936 551388 599992
rect 551324 599932 551388 599936
rect 551324 599524 551388 599588
rect 551692 599524 551756 599588
rect 551324 595096 551388 595100
rect 551324 595040 551374 595096
rect 551374 595040 551388 595096
rect 551324 595036 551388 595040
rect 551692 595036 551756 595100
rect 551508 592316 551572 592380
rect 551324 592240 551388 592244
rect 551324 592184 551374 592240
rect 551374 592184 551388 592240
rect 551324 592180 551388 592184
rect 551324 587148 551388 587212
rect 552980 587148 553044 587212
rect 551324 586936 551388 586940
rect 551324 586880 551374 586936
rect 551374 586880 551388 586936
rect 551324 586876 551388 586880
rect 551324 586256 551388 586260
rect 551324 586200 551374 586256
rect 551374 586200 551388 586256
rect 551324 586196 551388 586200
rect 551508 582524 551572 582588
rect 552980 582524 553044 582588
rect 551324 582116 551388 582180
rect 551508 578444 551572 578508
rect 551324 578172 551388 578236
rect 551324 577552 551388 577556
rect 551324 577496 551374 577552
rect 551374 577496 551388 577552
rect 551324 577492 551388 577496
rect 28580 575452 28644 575516
rect 28580 571508 28644 571572
rect 546356 569876 546420 569940
rect 280292 569740 280356 569804
rect 281396 569740 281460 569804
rect 551508 569876 551572 569940
rect 551692 569740 551756 569804
rect 280292 563756 280356 563820
rect 551140 563212 551204 563276
rect 550036 562260 550100 562324
rect 551692 562260 551756 562324
rect 548380 560900 548444 560964
rect 550772 560220 550836 560284
rect 550956 560280 551020 560284
rect 550956 560224 551006 560280
rect 551006 560224 551020 560280
rect 550956 560220 551020 560224
rect 551140 560084 551204 560148
rect 551508 560084 551572 560148
rect 550772 559948 550836 560012
rect 29316 559540 29380 559604
rect 550956 555520 551020 555524
rect 550956 555464 551006 555520
rect 551006 555464 551020 555520
rect 550956 555460 551020 555464
rect 25452 554100 25516 554164
rect 25268 553964 25332 554028
rect 280476 553148 280540 553212
rect 550588 548524 550652 548588
rect 551692 548524 551756 548588
rect 552796 545668 552860 545732
rect 551140 543764 551204 543828
rect 551508 543764 551572 543828
rect 551140 543628 551204 543692
rect 551692 543628 551756 543692
rect 280292 541180 280356 541244
rect 280476 541180 280540 541244
rect 550588 538868 550652 538932
rect 551508 538868 551572 538932
rect 549852 534652 549916 534716
rect 280476 534244 280540 534308
rect 280292 533836 280356 533900
rect 25820 533564 25884 533628
rect 552612 533564 552676 533628
rect 26004 533428 26068 533492
rect 552428 533428 552492 533492
rect 28212 533292 28276 533356
rect 552060 533292 552124 533356
rect 25636 532612 25700 532676
rect 552244 532612 552308 532676
rect 28028 532476 28092 532540
rect 550956 532476 551020 532540
rect 27108 532340 27172 532404
rect 553716 532340 553780 532404
rect 27292 532204 27356 532268
rect 551508 532204 551572 532268
rect 27476 532068 27540 532132
rect 553532 532068 553596 532132
rect 27660 531932 27724 531996
rect 553348 531932 553412 531996
rect 551876 531796 551940 531860
rect 546356 531252 546420 531316
rect 492444 531116 492508 531180
rect 551324 531116 551388 531180
rect 551692 530980 551756 531044
rect 26740 530844 26804 530908
rect 554084 530844 554148 530908
rect 27844 530708 27908 530772
rect 550772 530708 550836 530772
rect 26924 530572 26988 530636
rect 553900 530572 553964 530636
rect 280292 528396 280356 528460
rect 280476 518936 280540 518940
rect 280476 518880 280526 518936
rect 280526 518880 280540 518936
rect 280476 518876 280540 518880
rect 280476 509220 280540 509284
rect 280476 509084 280540 509148
rect 118740 500848 118804 500852
rect 118740 500792 118754 500848
rect 118754 500792 118804 500848
rect 118740 500788 118804 500792
rect 147076 500848 147140 500852
rect 147076 500792 147090 500848
rect 147090 500792 147140 500848
rect 147076 500788 147140 500792
rect 147812 500788 147876 500852
rect 148180 500848 148244 500852
rect 148180 500792 148194 500848
rect 148194 500792 148244 500848
rect 148180 500788 148244 500792
rect 149652 500788 149716 500852
rect 149836 500788 149900 500852
rect 150940 500788 151004 500852
rect 152412 500848 152476 500852
rect 152412 500792 152462 500848
rect 152462 500792 152476 500848
rect 148364 500516 148428 500580
rect 152412 500788 152476 500792
rect 153148 500788 153212 500852
rect 189580 500788 189644 500852
rect 191052 500788 191116 500852
rect 189764 500652 189828 500716
rect 548380 500652 548444 500716
rect 153332 500516 153396 500580
rect 153884 500516 153948 500580
rect 549852 500516 549916 500580
rect 147996 500380 148060 500444
rect 546540 500380 546604 500444
rect 147260 500244 147324 500308
rect 550588 500244 550652 500308
rect 114692 500108 114756 500172
rect 147628 500108 147692 500172
rect 188844 500108 188908 500172
rect 550772 500108 550836 500172
rect 150572 499972 150636 500036
rect 150756 499836 150820 499900
rect 149284 499700 149348 499764
rect 151124 499564 151188 499628
rect 150020 497932 150084 497996
rect 151308 497796 151372 497860
rect 150388 497660 150452 497724
rect 149100 497524 149164 497588
rect 147444 497388 147508 497452
rect 280292 495544 280356 495548
rect 280292 495488 280342 495544
rect 280342 495488 280356 495544
rect 280292 495484 280356 495488
rect 20484 492492 20548 492556
rect 280660 489908 280724 489972
rect 152780 486508 152844 486572
rect 152044 486432 152108 486436
rect 152044 486376 152058 486432
rect 152058 486376 152108 486432
rect 152044 486372 152108 486376
rect 20300 485012 20364 485076
rect 21220 485012 21284 485076
rect 280108 480252 280172 480316
rect 280660 480252 280724 480316
rect 280108 480040 280172 480044
rect 280108 479984 280158 480040
rect 280158 479984 280172 480040
rect 280108 479980 280172 479984
rect 553348 475492 553412 475556
rect 552060 475356 552124 475420
rect 546540 473512 546604 473516
rect 546540 473456 546590 473512
rect 546590 473456 546604 473512
rect 546540 473452 546604 473456
rect 552060 471820 552124 471884
rect 280292 470596 280356 470660
rect 552060 470052 552124 470116
rect 552060 468284 552124 468348
rect 553348 464476 553412 464540
rect 280292 463660 280356 463724
rect 280660 463660 280724 463724
rect 555188 461484 555252 461548
rect 554820 460260 554884 460324
rect 280292 451208 280356 451212
rect 280292 451152 280306 451208
rect 280306 451152 280356 451208
rect 280292 451148 280356 451152
rect 280292 445768 280356 445772
rect 280292 445712 280306 445768
rect 280306 445712 280356 445768
rect 280292 445708 280356 445712
rect 280292 439512 280356 439516
rect 280292 439456 280342 439512
rect 280342 439456 280356 439512
rect 280292 439452 280356 439456
rect 280292 434752 280356 434756
rect 280292 434696 280342 434752
rect 280342 434696 280356 434752
rect 280292 434692 280356 434696
rect 317092 428708 317156 428772
rect 316908 428572 316972 428636
rect 280292 428436 280356 428500
rect 281028 428436 281092 428500
rect 317276 428436 317340 428500
rect 280844 423540 280908 423604
rect 281028 423540 281092 423604
rect 157196 421228 157260 421292
rect 281580 421288 281644 421292
rect 281580 421232 281630 421288
rect 281630 421232 281644 421288
rect 281580 421228 281644 421232
rect 151124 401508 151188 401572
rect 148364 401372 148428 401436
rect 147996 401236 148060 401300
rect 150204 401100 150268 401164
rect 150020 400964 150084 401028
rect 151308 400828 151372 400892
rect 150572 400692 150636 400756
rect 150756 400556 150820 400620
rect 149284 400420 149348 400484
rect 153332 400284 153396 400348
rect 189948 376756 190012 376820
rect 189948 360028 190012 360092
rect 20300 357580 20364 357644
rect 280476 357580 280540 357644
rect 281028 357580 281092 357644
rect 188844 357444 188908 357508
rect 122604 351732 122668 351796
rect 147260 351596 147324 351660
rect 189764 351732 189828 351796
rect 191052 351732 191116 351796
rect 151860 351596 151924 351660
rect 189580 351596 189644 351660
rect 147076 351460 147140 351524
rect 148180 351460 148244 351524
rect 149652 351460 149716 351524
rect 149836 351460 149900 351524
rect 150940 351460 151004 351524
rect 152412 351520 152476 351524
rect 152412 351464 152426 351520
rect 152426 351464 152476 351520
rect 152412 351460 152476 351464
rect 147628 351324 147692 351388
rect 150388 351188 150452 351252
rect 147444 351052 147508 351116
rect 149100 350916 149164 350980
rect 129596 350780 129660 350844
rect 152044 350780 152108 350844
rect 153148 350644 153212 350708
rect 147812 350508 147876 350572
rect 280292 350372 280356 350436
rect 280844 350372 280908 350436
rect 280292 347652 280356 347716
rect 280660 338132 280724 338196
rect 280660 336636 280724 336700
rect 280292 336500 280356 336564
rect 280292 327040 280356 327044
rect 280292 326984 280342 327040
rect 280342 326984 280356 327040
rect 280292 326980 280356 326984
rect 214420 322084 214484 322148
rect 20484 320724 20548 320788
rect 51580 320724 51644 320788
rect 195100 320452 195164 320516
rect 196572 320316 196636 320380
rect 190316 320180 190380 320244
rect 191604 320180 191668 320244
rect 194364 320180 194428 320244
rect 208348 319364 208412 319428
rect 280292 317656 280356 317660
rect 280292 317600 280342 317656
rect 280342 317600 280356 317656
rect 280292 317596 280356 317600
rect 280292 317384 280356 317388
rect 280292 317328 280342 317384
rect 280342 317328 280356 317384
rect 280292 317324 280356 317328
rect 280292 309632 280356 309636
rect 280292 309576 280342 309632
rect 280342 309576 280356 309632
rect 280292 309572 280356 309576
rect 280292 306308 280356 306372
rect 280476 306308 280540 306372
rect 332916 302772 332980 302836
rect 280660 296652 280724 296716
rect 281028 296652 281092 296716
rect 281028 295156 281092 295220
rect 280476 277476 280540 277540
rect 280476 273396 280540 273460
rect 280292 273124 280356 273188
rect 280292 259524 280356 259588
rect 280476 259524 280540 259588
rect 181668 253948 181732 254012
rect 279372 253948 279436 254012
rect 280476 251152 280540 251156
rect 280476 251096 280526 251152
rect 280526 251096 280540 251152
rect 280476 251092 280540 251096
rect 280660 241572 280724 241636
rect 51580 235996 51644 236060
rect 194364 235180 194428 235244
rect 280660 235180 280724 235244
rect 191604 233820 191668 233884
rect 196572 232460 196636 232524
rect 190316 229740 190380 229804
rect 195100 228244 195164 228308
rect 208348 223620 208412 223684
rect 332916 173844 332980 173908
rect 214420 159428 214484 159492
rect 32260 125080 32324 125084
rect 32260 125024 32274 125080
rect 32274 125024 32324 125080
rect 32260 125020 32324 125024
rect 32260 31784 32324 31788
rect 32260 31728 32310 31784
rect 32310 31728 32324 31784
rect 32260 31724 32324 31728
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 -6926 -7976 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 -5986 -7036 709922
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 -5046 -6096 708982
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 -4106 -5156 708042
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 -3166 -4216 707102
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 -2226 -3276 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 617680 37404 649898
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 617680 55404 631898
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 617680 73404 649898
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 617680 91404 631898
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 617680 109404 649898
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 113403 622436 113469 622437
rect 113403 622372 113404 622436
rect 113468 622372 113469 622436
rect 113403 622371 113469 622372
rect 113406 617677 113466 622371
rect 126804 617680 127404 631898
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 106227 617676 106293 617677
rect 106227 617612 106228 617676
rect 106292 617612 106293 617676
rect 106227 617611 106293 617612
rect 113403 617676 113469 617677
rect 113403 617612 113404 617676
rect 113468 617612 113469 617676
rect 113403 617611 113469 617612
rect 25451 617404 25517 617405
rect 25451 617340 25452 617404
rect 25516 617340 25517 617404
rect 25451 617339 25517 617340
rect 21219 615772 21285 615773
rect 21219 615708 21220 615772
rect 21284 615708 21285 615772
rect 21219 615707 21285 615708
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 20483 492556 20549 492557
rect 20483 492492 20484 492556
rect 20548 492492 20549 492556
rect 20483 492491 20549 492492
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 487040 19404 487898
rect 20299 485076 20365 485077
rect 20299 485012 20300 485076
rect 20364 485012 20365 485076
rect 20299 485011 20365 485012
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 18804 380454 19404 400000
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 20302 357645 20362 485011
rect 20299 357644 20365 357645
rect 20299 357580 20300 357644
rect 20364 357580 20365 357644
rect 20299 357579 20365 357580
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 20486 320789 20546 492491
rect 21222 485077 21282 615707
rect 25267 614412 25333 614413
rect 25267 614348 25268 614412
rect 25332 614348 25333 614412
rect 25267 614347 25333 614348
rect 25270 554029 25330 614347
rect 25454 554165 25514 617339
rect 106230 617218 106290 617611
rect 27659 616860 27725 616861
rect 27659 616796 27660 616860
rect 27724 616796 27725 616860
rect 27659 616795 27725 616796
rect 27475 616180 27541 616181
rect 27475 616116 27476 616180
rect 27540 616116 27541 616180
rect 27475 616115 27541 616116
rect 27291 614956 27357 614957
rect 27291 614892 27292 614956
rect 27356 614892 27357 614956
rect 27291 614891 27357 614892
rect 27107 613868 27173 613869
rect 27107 613804 27108 613868
rect 27172 613804 27173 613868
rect 27107 613803 27173 613804
rect 26923 611420 26989 611421
rect 26923 611356 26924 611420
rect 26988 611356 26989 611420
rect 26923 611355 26989 611356
rect 26739 610196 26805 610197
rect 26739 610132 26740 610196
rect 26804 610132 26805 610196
rect 26739 610131 26805 610132
rect 26003 604756 26069 604757
rect 26003 604692 26004 604756
rect 26068 604692 26069 604756
rect 26003 604691 26069 604692
rect 25819 603668 25885 603669
rect 25819 603604 25820 603668
rect 25884 603604 25885 603668
rect 25819 603603 25885 603604
rect 25635 599996 25701 599997
rect 25635 599932 25636 599996
rect 25700 599932 25701 599996
rect 25635 599931 25701 599932
rect 25451 554164 25517 554165
rect 25451 554100 25452 554164
rect 25516 554100 25517 554164
rect 25451 554099 25517 554100
rect 25267 554028 25333 554029
rect 25267 553964 25268 554028
rect 25332 553964 25333 554028
rect 25267 553963 25333 553964
rect 25638 532677 25698 599931
rect 25822 533629 25882 603603
rect 25819 533628 25885 533629
rect 25819 533564 25820 533628
rect 25884 533564 25885 533628
rect 25819 533563 25885 533564
rect 26006 533493 26066 604691
rect 26003 533492 26069 533493
rect 26003 533428 26004 533492
rect 26068 533428 26069 533492
rect 26003 533427 26069 533428
rect 25635 532676 25701 532677
rect 25635 532612 25636 532676
rect 25700 532612 25701 532676
rect 25635 532611 25701 532612
rect 26742 530909 26802 610131
rect 26739 530908 26805 530909
rect 26739 530844 26740 530908
rect 26804 530844 26805 530908
rect 26739 530843 26805 530844
rect 26926 530637 26986 611355
rect 27110 532405 27170 613803
rect 27107 532404 27173 532405
rect 27107 532340 27108 532404
rect 27172 532340 27173 532404
rect 27107 532339 27173 532340
rect 27294 532269 27354 614891
rect 27291 532268 27357 532269
rect 27291 532204 27292 532268
rect 27356 532204 27357 532268
rect 27291 532203 27357 532204
rect 27478 532133 27538 616115
rect 27475 532132 27541 532133
rect 27475 532068 27476 532132
rect 27540 532068 27541 532132
rect 27475 532067 27541 532068
rect 27662 531997 27722 616795
rect 28579 615772 28645 615773
rect 28579 615708 28580 615772
rect 28644 615770 28645 615772
rect 28644 615710 29010 615770
rect 28644 615708 28645 615710
rect 28579 615707 28645 615708
rect 28950 615178 29010 615710
rect 28211 612780 28277 612781
rect 28211 612716 28212 612780
rect 28276 612716 28277 612780
rect 28211 612715 28277 612716
rect 28027 612100 28093 612101
rect 28027 612036 28028 612100
rect 28092 612036 28093 612100
rect 28027 612035 28093 612036
rect 27843 610876 27909 610877
rect 27843 610812 27844 610876
rect 27908 610812 27909 610876
rect 27843 610811 27909 610812
rect 27659 531996 27725 531997
rect 27659 531932 27660 531996
rect 27724 531932 27725 531996
rect 27659 531931 27725 531932
rect 27846 530773 27906 610811
rect 28030 532541 28090 612035
rect 28214 533357 28274 612715
rect 29502 581770 29562 614942
rect 29318 581710 29562 581770
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 28579 575516 28645 575517
rect 28579 575452 28580 575516
rect 28644 575452 28645 575516
rect 28579 575451 28645 575452
rect 28582 571573 28642 575451
rect 28579 571572 28645 571573
rect 28579 571508 28580 571572
rect 28644 571508 28645 571572
rect 28579 571507 28645 571508
rect 29318 559605 29378 581710
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 29315 559604 29381 559605
rect 29315 559540 29316 559604
rect 29380 559540 29381 559604
rect 29315 559539 29381 559540
rect 36804 542454 37404 571440
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 28211 533356 28277 533357
rect 28211 533292 28212 533356
rect 28276 533292 28277 533356
rect 28211 533291 28277 533292
rect 28027 532540 28093 532541
rect 28027 532476 28028 532540
rect 28092 532476 28093 532540
rect 28027 532475 28093 532476
rect 27843 530772 27909 530773
rect 27843 530708 27844 530772
rect 27908 530708 27909 530772
rect 27843 530707 27909 530708
rect 26923 530636 26989 530637
rect 26923 530572 26924 530636
rect 26988 530572 26989 530636
rect 26923 530571 26989 530572
rect 36804 528912 37404 541898
rect 54804 560454 55404 571440
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 528912 55404 559898
rect 72804 542454 73404 571440
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 528912 73404 541898
rect 90804 560454 91404 571440
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 528912 91404 559898
rect 108804 542454 109404 571440
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 528912 109404 541898
rect 126804 560454 127404 571440
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 528912 127404 559898
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 528912 145404 541898
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 528912 163404 559898
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 618224 199404 631898
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 618224 217404 649898
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 618224 235404 631898
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 618224 253404 649898
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 618224 271404 631898
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 280659 618356 280725 618357
rect 280659 618292 280660 618356
rect 280724 618292 280725 618356
rect 280659 618291 280725 618292
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 280662 611690 280722 618291
rect 280478 611630 280722 611690
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 280478 605570 280538 611630
rect 280478 605510 280722 605570
rect 280662 597410 280722 605510
rect 280662 597350 281458 597410
rect 281398 589250 281458 597350
rect 280110 589190 281458 589250
rect 280110 585850 280170 589190
rect 280110 585790 280538 585850
rect 280478 585170 280538 585790
rect 280478 585110 281090 585170
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 281030 577010 281090 585110
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 281030 576950 281458 577010
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 528912 181404 541898
rect 198804 560454 199404 574112
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 528912 199404 559898
rect 216804 542454 217404 574112
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 528912 217404 541898
rect 234804 560454 235404 574112
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 528912 235404 559898
rect 252804 542454 253404 574112
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 528912 253404 541898
rect 270804 560454 271404 574112
rect 281398 569805 281458 576950
rect 280291 569804 280357 569805
rect 280291 569740 280292 569804
rect 280356 569740 280357 569804
rect 280291 569739 280357 569740
rect 281395 569804 281461 569805
rect 281395 569740 281396 569804
rect 281460 569740 281461 569804
rect 281395 569739 281461 569740
rect 280294 563821 280354 569739
rect 280291 563820 280357 563821
rect 280291 563756 280292 563820
rect 280356 563756 280357 563820
rect 280291 563755 280357 563756
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 528912 271404 559898
rect 280475 553212 280541 553213
rect 280475 553148 280476 553212
rect 280540 553148 280541 553212
rect 280475 553147 280541 553148
rect 280478 550490 280538 553147
rect 280294 550430 280538 550490
rect 280294 541245 280354 550430
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 280291 541244 280357 541245
rect 280291 541180 280292 541244
rect 280356 541180 280357 541244
rect 280291 541179 280357 541180
rect 280475 541244 280541 541245
rect 280475 541180 280476 541244
rect 280540 541180 280541 541244
rect 280475 541179 280541 541180
rect 280478 534309 280538 541179
rect 280475 534308 280541 534309
rect 280475 534244 280476 534308
rect 280540 534244 280541 534308
rect 280475 534243 280541 534244
rect 280291 533900 280357 533901
rect 280291 533836 280292 533900
rect 280356 533836 280357 533900
rect 280291 533835 280357 533836
rect 280294 528461 280354 533835
rect 280291 528460 280357 528461
rect 280291 528396 280292 528460
rect 280356 528396 280357 528460
rect 280291 528395 280357 528396
rect 107675 524454 107995 524476
rect 107675 524218 107717 524454
rect 107953 524218 107995 524454
rect 107675 524134 107995 524218
rect 107675 523898 107717 524134
rect 107953 523898 107995 524134
rect 107675 523876 107995 523898
rect 192805 524454 193125 524476
rect 192805 524218 192847 524454
rect 193083 524218 193125 524454
rect 192805 524134 193125 524218
rect 192805 523898 192847 524134
rect 193083 523898 193125 524134
rect 192805 523876 193125 523898
rect 280475 518940 280541 518941
rect 280475 518876 280476 518940
rect 280540 518876 280541 518940
rect 280475 518875 280541 518876
rect 280478 509285 280538 518875
rect 280475 509284 280541 509285
rect 280475 509220 280476 509284
rect 280540 509220 280541 509284
rect 280475 509219 280541 509220
rect 280475 509148 280541 509149
rect 280475 509084 280476 509148
rect 280540 509084 280541 509148
rect 280475 509083 280541 509084
rect 65109 506454 65429 506476
rect 65109 506218 65151 506454
rect 65387 506218 65429 506454
rect 65109 506134 65429 506218
rect 65109 505898 65151 506134
rect 65387 505898 65429 506134
rect 65109 505876 65429 505898
rect 150240 506454 150560 506476
rect 150240 506218 150282 506454
rect 150518 506218 150560 506454
rect 150240 506134 150560 506218
rect 150240 505898 150282 506134
rect 150518 505898 150560 506134
rect 150240 505876 150560 505898
rect 235370 506454 235690 506476
rect 235370 506218 235412 506454
rect 235648 506218 235690 506454
rect 235370 506134 235690 506218
rect 235370 505898 235412 506134
rect 235648 505898 235690 506134
rect 235370 505876 235690 505898
rect 280478 504930 280538 509083
rect 280294 504870 280538 504930
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 36804 487040 37404 502800
rect 54804 488454 55404 502800
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 487040 55404 487898
rect 72804 487040 73404 502800
rect 90804 488454 91404 502800
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 487040 91404 487898
rect 108804 487040 109404 502800
rect 126804 488454 127404 502800
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 487040 127404 487898
rect 144804 487040 145404 502800
rect 147075 500852 147141 500853
rect 147075 500788 147076 500852
rect 147140 500788 147141 500852
rect 147075 500787 147141 500788
rect 147811 500852 147877 500853
rect 147811 500788 147812 500852
rect 147876 500788 147877 500852
rect 147811 500787 147877 500788
rect 148179 500852 148245 500853
rect 148179 500788 148180 500852
rect 148244 500788 148245 500852
rect 148179 500787 148245 500788
rect 149651 500852 149717 500853
rect 149651 500788 149652 500852
rect 149716 500788 149717 500852
rect 149651 500787 149717 500788
rect 149835 500852 149901 500853
rect 149835 500788 149836 500852
rect 149900 500788 149901 500852
rect 149835 500787 149901 500788
rect 150939 500852 151005 500853
rect 150939 500788 150940 500852
rect 151004 500788 151005 500852
rect 150939 500787 151005 500788
rect 21219 485076 21285 485077
rect 21219 485012 21220 485076
rect 21284 485012 21285 485076
rect 21219 485011 21285 485012
rect 23684 470454 24004 470476
rect 23684 470218 23726 470454
rect 23962 470218 24004 470454
rect 23684 470134 24004 470218
rect 23684 469898 23726 470134
rect 23962 469898 24004 470134
rect 23684 469876 24004 469898
rect 54404 470454 54724 470476
rect 54404 470218 54446 470454
rect 54682 470218 54724 470454
rect 54404 470134 54724 470218
rect 54404 469898 54446 470134
rect 54682 469898 54724 470134
rect 54404 469876 54724 469898
rect 85124 470454 85444 470476
rect 85124 470218 85166 470454
rect 85402 470218 85444 470454
rect 85124 470134 85444 470218
rect 85124 469898 85166 470134
rect 85402 469898 85444 470134
rect 85124 469876 85444 469898
rect 115844 470454 116164 470476
rect 115844 470218 115886 470454
rect 116122 470218 116164 470454
rect 115844 470134 116164 470218
rect 115844 469898 115886 470134
rect 116122 469898 116164 470134
rect 115844 469876 116164 469898
rect 146564 470454 146884 470476
rect 146564 470218 146606 470454
rect 146842 470218 146884 470454
rect 146564 470134 146884 470218
rect 146564 469898 146606 470134
rect 146842 469898 146884 470134
rect 146564 469876 146884 469898
rect 39044 452454 39364 452476
rect 39044 452218 39086 452454
rect 39322 452218 39364 452454
rect 39044 452134 39364 452218
rect 39044 451898 39086 452134
rect 39322 451898 39364 452134
rect 39044 451876 39364 451898
rect 69764 452454 70084 452476
rect 69764 452218 69806 452454
rect 70042 452218 70084 452454
rect 69764 452134 70084 452218
rect 69764 451898 69806 452134
rect 70042 451898 70084 452134
rect 69764 451876 70084 451898
rect 100484 452454 100804 452476
rect 100484 452218 100526 452454
rect 100762 452218 100804 452454
rect 100484 452134 100804 452218
rect 100484 451898 100526 452134
rect 100762 451898 100804 452134
rect 100484 451876 100804 451898
rect 131204 452454 131524 452476
rect 131204 452218 131246 452454
rect 131482 452218 131524 452454
rect 131204 452134 131524 452218
rect 131204 451898 131246 452134
rect 131482 451898 131524 452134
rect 131204 451876 131524 451898
rect 23684 434454 24004 434476
rect 23684 434218 23726 434454
rect 23962 434218 24004 434454
rect 23684 434134 24004 434218
rect 23684 433898 23726 434134
rect 23962 433898 24004 434134
rect 23684 433876 24004 433898
rect 54404 434454 54724 434476
rect 54404 434218 54446 434454
rect 54682 434218 54724 434454
rect 54404 434134 54724 434218
rect 54404 433898 54446 434134
rect 54682 433898 54724 434134
rect 54404 433876 54724 433898
rect 85124 434454 85444 434476
rect 85124 434218 85166 434454
rect 85402 434218 85444 434454
rect 85124 434134 85444 434218
rect 85124 433898 85166 434134
rect 85402 433898 85444 434134
rect 85124 433876 85444 433898
rect 115844 434454 116164 434476
rect 115844 434218 115886 434454
rect 116122 434218 116164 434454
rect 115844 434134 116164 434218
rect 115844 433898 115886 434134
rect 116122 433898 116164 434134
rect 115844 433876 116164 433898
rect 146564 434454 146884 434476
rect 146564 434218 146606 434454
rect 146842 434218 146884 434454
rect 146564 434134 146884 434218
rect 146564 433898 146606 434134
rect 146842 433898 146884 434134
rect 146564 433876 146884 433898
rect 39044 416454 39364 416476
rect 39044 416218 39086 416454
rect 39322 416218 39364 416454
rect 39044 416134 39364 416218
rect 39044 415898 39086 416134
rect 39322 415898 39364 416134
rect 39044 415876 39364 415898
rect 69764 416454 70084 416476
rect 69764 416218 69806 416454
rect 70042 416218 70084 416454
rect 69764 416134 70084 416218
rect 69764 415898 69806 416134
rect 70042 415898 70084 416134
rect 69764 415876 70084 415898
rect 100484 416454 100804 416476
rect 100484 416218 100526 416454
rect 100762 416218 100804 416454
rect 100484 416134 100804 416218
rect 100484 415898 100526 416134
rect 100762 415898 100804 416134
rect 100484 415876 100804 415898
rect 131204 416454 131524 416476
rect 131204 416218 131246 416454
rect 131482 416218 131524 416454
rect 131204 416134 131524 416218
rect 131204 415898 131246 416134
rect 131482 415898 131524 416134
rect 131204 415876 131524 415898
rect 36804 398454 37404 400000
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 384200 37404 397898
rect 54804 384200 55404 400000
rect 72804 398454 73404 400000
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 384200 73404 397898
rect 38875 380454 39195 380476
rect 38875 380218 38917 380454
rect 39153 380218 39195 380454
rect 38875 380134 39195 380218
rect 38875 379898 38917 380134
rect 39153 379898 39195 380134
rect 38875 379876 39195 379898
rect 56805 380454 57125 380476
rect 56805 380218 56847 380454
rect 57083 380218 57125 380454
rect 56805 380134 57125 380218
rect 56805 379898 56847 380134
rect 57083 379898 57125 380134
rect 56805 379876 57125 379898
rect 90804 380454 91404 400000
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 29909 362454 30229 362476
rect 29909 362218 29951 362454
rect 30187 362218 30229 362454
rect 29909 362134 30229 362218
rect 29909 361898 29951 362134
rect 30187 361898 30229 362134
rect 29909 361876 30229 361898
rect 47840 362454 48160 362476
rect 47840 362218 47882 362454
rect 48118 362218 48160 362454
rect 47840 362134 48160 362218
rect 47840 361898 47882 362134
rect 48118 361898 48160 362134
rect 47840 361876 48160 361898
rect 65770 362454 66090 362476
rect 65770 362218 65812 362454
rect 66048 362218 66090 362454
rect 65770 362134 66090 362218
rect 65770 361898 65812 362134
rect 66048 361898 66090 362134
rect 65770 361876 66090 361898
rect 36804 348912 37404 357000
rect 54804 348912 55404 357000
rect 72804 348912 73404 357000
rect 90804 348912 91404 379898
rect 108804 398454 109404 400000
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 348912 109404 361898
rect 122606 351797 122666 400742
rect 126804 380454 127404 400000
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 122603 351796 122669 351797
rect 122603 351732 122604 351796
rect 122668 351732 122669 351796
rect 122603 351731 122669 351732
rect 126804 348912 127404 379898
rect 129598 350845 129658 401422
rect 144804 398454 145404 400000
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 129595 350844 129661 350845
rect 129595 350780 129596 350844
rect 129660 350780 129661 350844
rect 129595 350779 129661 350780
rect 144804 348912 145404 361898
rect 147078 351525 147138 500787
rect 147259 500308 147325 500309
rect 147259 500244 147260 500308
rect 147324 500244 147325 500308
rect 147259 500243 147325 500244
rect 147262 351661 147322 500243
rect 147627 500172 147693 500173
rect 147627 500108 147628 500172
rect 147692 500108 147693 500172
rect 147627 500107 147693 500108
rect 147443 497452 147509 497453
rect 147443 497388 147444 497452
rect 147508 497388 147509 497452
rect 147443 497387 147509 497388
rect 147259 351660 147325 351661
rect 147259 351596 147260 351660
rect 147324 351596 147325 351660
rect 147259 351595 147325 351596
rect 147075 351524 147141 351525
rect 147075 351460 147076 351524
rect 147140 351460 147141 351524
rect 147075 351459 147141 351460
rect 147446 351117 147506 497387
rect 147630 351389 147690 500107
rect 147627 351388 147693 351389
rect 147627 351324 147628 351388
rect 147692 351324 147693 351388
rect 147627 351323 147693 351324
rect 147443 351116 147509 351117
rect 147443 351052 147444 351116
rect 147508 351052 147509 351116
rect 147443 351051 147509 351052
rect 147814 350573 147874 500787
rect 147995 500444 148061 500445
rect 147995 500380 147996 500444
rect 148060 500380 148061 500444
rect 147995 500379 148061 500380
rect 147998 401301 148058 500379
rect 147995 401300 148061 401301
rect 147995 401236 147996 401300
rect 148060 401236 148061 401300
rect 147995 401235 148061 401236
rect 148182 351525 148242 500787
rect 148363 500580 148429 500581
rect 148363 500516 148364 500580
rect 148428 500516 148429 500580
rect 148363 500515 148429 500516
rect 148366 401437 148426 500515
rect 149283 499764 149349 499765
rect 149283 499700 149284 499764
rect 149348 499700 149349 499764
rect 149283 499699 149349 499700
rect 149099 497588 149165 497589
rect 149099 497524 149100 497588
rect 149164 497524 149165 497588
rect 149099 497523 149165 497524
rect 148363 401436 148429 401437
rect 148363 401372 148364 401436
rect 148428 401372 148429 401436
rect 148363 401371 148429 401372
rect 148179 351524 148245 351525
rect 148179 351460 148180 351524
rect 148244 351460 148245 351524
rect 148179 351459 148245 351460
rect 149102 350981 149162 497523
rect 149286 400485 149346 499699
rect 149283 400484 149349 400485
rect 149283 400420 149284 400484
rect 149348 400420 149349 400484
rect 149283 400419 149349 400420
rect 149654 351525 149714 500787
rect 149838 351525 149898 500787
rect 150571 500036 150637 500037
rect 150019 497996 150085 497997
rect 150019 497932 150020 497996
rect 150084 497932 150085 497996
rect 150019 497931 150085 497932
rect 150022 401029 150082 497931
rect 150206 401165 150266 500022
rect 150571 499972 150572 500036
rect 150636 499972 150637 500036
rect 150571 499971 150637 499972
rect 150387 497724 150453 497725
rect 150387 497660 150388 497724
rect 150452 497660 150453 497724
rect 150387 497659 150453 497660
rect 150203 401164 150269 401165
rect 150203 401100 150204 401164
rect 150268 401100 150269 401164
rect 150203 401099 150269 401100
rect 150019 401028 150085 401029
rect 150019 400964 150020 401028
rect 150084 400964 150085 401028
rect 150019 400963 150085 400964
rect 149651 351524 149717 351525
rect 149651 351460 149652 351524
rect 149716 351460 149717 351524
rect 149651 351459 149717 351460
rect 149835 351524 149901 351525
rect 149835 351460 149836 351524
rect 149900 351460 149901 351524
rect 149835 351459 149901 351460
rect 150390 351253 150450 497659
rect 150574 400757 150634 499971
rect 150755 499900 150821 499901
rect 150755 499836 150756 499900
rect 150820 499836 150821 499900
rect 150755 499835 150821 499836
rect 150571 400756 150637 400757
rect 150571 400692 150572 400756
rect 150636 400692 150637 400756
rect 150571 400691 150637 400692
rect 150758 400621 150818 499835
rect 150755 400620 150821 400621
rect 150755 400556 150756 400620
rect 150820 400556 150821 400620
rect 150755 400555 150821 400556
rect 150942 351525 151002 500787
rect 152411 500852 152477 500853
rect 152411 500788 152412 500852
rect 152476 500788 152477 500852
rect 152411 500787 152477 500788
rect 153147 500852 153213 500853
rect 153147 500788 153148 500852
rect 153212 500788 153213 500852
rect 153147 500787 153213 500788
rect 151123 499628 151189 499629
rect 151123 499564 151124 499628
rect 151188 499564 151189 499628
rect 151123 499563 151189 499564
rect 151126 401573 151186 499563
rect 151307 497860 151373 497861
rect 151307 497796 151308 497860
rect 151372 497796 151373 497860
rect 151307 497795 151373 497796
rect 151123 401572 151189 401573
rect 151123 401508 151124 401572
rect 151188 401508 151189 401572
rect 151123 401507 151189 401508
rect 151310 400893 151370 497795
rect 151307 400892 151373 400893
rect 151307 400828 151308 400892
rect 151372 400828 151373 400892
rect 151307 400827 151373 400828
rect 151862 351661 151922 500702
rect 152043 486436 152109 486437
rect 152043 486372 152044 486436
rect 152108 486372 152109 486436
rect 152043 486371 152109 486372
rect 151859 351660 151925 351661
rect 151859 351596 151860 351660
rect 151924 351596 151925 351660
rect 151859 351595 151925 351596
rect 150939 351524 151005 351525
rect 150939 351460 150940 351524
rect 151004 351460 151005 351524
rect 150939 351459 151005 351460
rect 150387 351252 150453 351253
rect 150387 351188 150388 351252
rect 150452 351188 150453 351252
rect 150387 351187 150453 351188
rect 149099 350980 149165 350981
rect 149099 350916 149100 350980
rect 149164 350916 149165 350980
rect 149099 350915 149165 350916
rect 152046 350845 152106 486371
rect 152414 351525 152474 500787
rect 152779 486572 152845 486573
rect 152779 486508 152780 486572
rect 152844 486508 152845 486572
rect 152779 486507 152845 486508
rect 152782 401658 152842 486507
rect 152411 351524 152477 351525
rect 152411 351460 152412 351524
rect 152476 351460 152477 351524
rect 152411 351459 152477 351460
rect 152043 350844 152109 350845
rect 152043 350780 152044 350844
rect 152108 350780 152109 350844
rect 152043 350779 152109 350780
rect 153150 350709 153210 500787
rect 153331 500580 153397 500581
rect 153331 500516 153332 500580
rect 153396 500516 153397 500580
rect 153331 500515 153397 500516
rect 153883 500580 153949 500581
rect 153883 500516 153884 500580
rect 153948 500516 153949 500580
rect 153883 500515 153949 500516
rect 153334 400349 153394 500515
rect 153886 400978 153946 500515
rect 162804 488454 163404 502800
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 153331 400348 153397 400349
rect 153331 400284 153332 400348
rect 153396 400284 153397 400348
rect 153331 400283 153397 400284
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 153147 350708 153213 350709
rect 153147 350644 153148 350708
rect 153212 350644 153213 350708
rect 153147 350643 153213 350644
rect 147811 350572 147877 350573
rect 147811 350508 147812 350572
rect 147876 350508 147877 350572
rect 147811 350507 147877 350508
rect 162804 348912 163404 379898
rect 180804 470454 181404 502800
rect 189579 500852 189645 500853
rect 189579 500788 189580 500852
rect 189644 500788 189645 500852
rect 189579 500787 189645 500788
rect 191051 500852 191117 500853
rect 191051 500788 191052 500852
rect 191116 500788 191117 500852
rect 191051 500787 191117 500788
rect 188843 500172 188909 500173
rect 188843 500108 188844 500172
rect 188908 500108 188909 500172
rect 188843 500107 188909 500108
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 348912 181404 361898
rect 188846 357509 188906 500107
rect 188843 357508 188909 357509
rect 188843 357444 188844 357508
rect 188908 357444 188909 357508
rect 188843 357443 188909 357444
rect 189582 351661 189642 500787
rect 189763 500716 189829 500717
rect 189763 500652 189764 500716
rect 189828 500652 189829 500716
rect 189763 500651 189829 500652
rect 189766 351797 189826 500651
rect 189947 376820 190013 376821
rect 189947 376756 189948 376820
rect 190012 376756 190013 376820
rect 189947 376755 190013 376756
rect 189950 360093 190010 376755
rect 189947 360092 190013 360093
rect 189947 360028 189948 360092
rect 190012 360028 190013 360092
rect 189947 360027 190013 360028
rect 191054 351797 191114 500787
rect 198804 491600 199404 502800
rect 216804 491600 217404 502800
rect 234804 491600 235404 502800
rect 252804 491600 253404 502800
rect 270804 491600 271404 502800
rect 280294 495549 280354 504870
rect 280291 495548 280357 495549
rect 280291 495484 280292 495548
rect 280356 495484 280357 495548
rect 280291 495483 280357 495484
rect 280659 489972 280725 489973
rect 280659 489908 280660 489972
rect 280724 489908 280725 489972
rect 280659 489907 280725 489908
rect 207614 488454 207934 488476
rect 207614 488218 207656 488454
rect 207892 488218 207934 488454
rect 207614 488134 207934 488218
rect 207614 487898 207656 488134
rect 207892 487898 207934 488134
rect 207614 487876 207934 487898
rect 238334 488454 238654 488476
rect 238334 488218 238376 488454
rect 238612 488218 238654 488454
rect 238334 488134 238654 488218
rect 238334 487898 238376 488134
rect 238612 487898 238654 488134
rect 238334 487876 238654 487898
rect 269054 488454 269374 488476
rect 269054 488218 269096 488454
rect 269332 488218 269374 488454
rect 269054 488134 269374 488218
rect 269054 487898 269096 488134
rect 269332 487898 269374 488134
rect 269054 487876 269374 487898
rect 280662 480317 280722 489907
rect 280107 480316 280173 480317
rect 280107 480252 280108 480316
rect 280172 480252 280173 480316
rect 280107 480251 280173 480252
rect 280659 480316 280725 480317
rect 280659 480252 280660 480316
rect 280724 480252 280725 480316
rect 280659 480251 280725 480252
rect 280110 480045 280170 480251
rect 280107 480044 280173 480045
rect 280107 479980 280108 480044
rect 280172 479980 280173 480044
rect 280107 479979 280173 479980
rect 280291 470660 280357 470661
rect 280291 470596 280292 470660
rect 280356 470596 280357 470660
rect 280291 470595 280357 470596
rect 192254 470454 192574 470476
rect 192254 470218 192296 470454
rect 192532 470218 192574 470454
rect 192254 470134 192574 470218
rect 192254 469898 192296 470134
rect 192532 469898 192574 470134
rect 192254 469876 192574 469898
rect 222974 470454 223294 470476
rect 222974 470218 223016 470454
rect 223252 470218 223294 470454
rect 222974 470134 223294 470218
rect 222974 469898 223016 470134
rect 223252 469898 223294 470134
rect 222974 469876 223294 469898
rect 253694 470454 254014 470476
rect 253694 470218 253736 470454
rect 253972 470218 254014 470454
rect 253694 470134 254014 470218
rect 253694 469898 253736 470134
rect 253972 469898 254014 470134
rect 253694 469876 254014 469898
rect 280294 463725 280354 470595
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 280291 463724 280357 463725
rect 280291 463660 280292 463724
rect 280356 463660 280357 463724
rect 280291 463659 280357 463660
rect 280659 463724 280725 463725
rect 280659 463660 280660 463724
rect 280724 463660 280725 463724
rect 280659 463659 280725 463660
rect 280662 456650 280722 463659
rect 280294 456590 280722 456650
rect 207614 452454 207934 452476
rect 207614 452218 207656 452454
rect 207892 452218 207934 452454
rect 207614 452134 207934 452218
rect 207614 451898 207656 452134
rect 207892 451898 207934 452134
rect 207614 451876 207934 451898
rect 238334 452454 238654 452476
rect 238334 452218 238376 452454
rect 238612 452218 238654 452454
rect 238334 452134 238654 452218
rect 238334 451898 238376 452134
rect 238612 451898 238654 452134
rect 238334 451876 238654 451898
rect 269054 452454 269374 452476
rect 269054 452218 269096 452454
rect 269332 452218 269374 452454
rect 269054 452134 269374 452218
rect 269054 451898 269096 452134
rect 269332 451898 269374 452134
rect 269054 451876 269374 451898
rect 280294 451213 280354 456590
rect 280291 451212 280357 451213
rect 280291 451148 280292 451212
rect 280356 451148 280357 451212
rect 280291 451147 280357 451148
rect 280291 445772 280357 445773
rect 280291 445708 280292 445772
rect 280356 445708 280357 445772
rect 280291 445707 280357 445708
rect 280294 439517 280354 445707
rect 280291 439516 280357 439517
rect 280291 439452 280292 439516
rect 280356 439452 280357 439516
rect 280291 439451 280357 439452
rect 280291 434756 280357 434757
rect 280291 434692 280292 434756
rect 280356 434692 280357 434756
rect 280291 434691 280357 434692
rect 192254 434454 192574 434476
rect 192254 434218 192296 434454
rect 192532 434218 192574 434454
rect 192254 434134 192574 434218
rect 192254 433898 192296 434134
rect 192532 433898 192574 434134
rect 192254 433876 192574 433898
rect 222974 434454 223294 434476
rect 222974 434218 223016 434454
rect 223252 434218 223294 434454
rect 222974 434134 223294 434218
rect 222974 433898 223016 434134
rect 223252 433898 223294 434134
rect 222974 433876 223294 433898
rect 253694 434454 254014 434476
rect 253694 434218 253736 434454
rect 253972 434218 254014 434454
rect 253694 434134 254014 434218
rect 253694 433898 253736 434134
rect 253972 433898 254014 434134
rect 253694 433876 254014 433898
rect 280294 428501 280354 434691
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 280291 428500 280357 428501
rect 280291 428436 280292 428500
rect 280356 428436 280357 428500
rect 280291 428435 280357 428436
rect 281027 428500 281093 428501
rect 281027 428436 281028 428500
rect 281092 428436 281093 428500
rect 281027 428435 281093 428436
rect 281030 423605 281090 428435
rect 280843 423604 280909 423605
rect 280843 423540 280844 423604
rect 280908 423540 280909 423604
rect 280843 423539 280909 423540
rect 281027 423604 281093 423605
rect 281027 423540 281028 423604
rect 281092 423540 281093 423604
rect 281027 423539 281093 423540
rect 280846 417890 280906 423539
rect 280662 417830 280906 417890
rect 207614 416454 207934 416476
rect 207614 416218 207656 416454
rect 207892 416218 207934 416454
rect 207614 416134 207934 416218
rect 207614 415898 207656 416134
rect 207892 415898 207934 416134
rect 207614 415876 207934 415898
rect 238334 416454 238654 416476
rect 238334 416218 238376 416454
rect 238612 416218 238654 416454
rect 238334 416134 238654 416218
rect 238334 415898 238376 416134
rect 238612 415898 238654 416134
rect 238334 415876 238654 415898
rect 269054 416454 269374 416476
rect 269054 416218 269096 416454
rect 269332 416218 269374 416454
rect 269054 416134 269374 416218
rect 269054 415898 269096 416134
rect 269332 415898 269374 416134
rect 269054 415876 269374 415898
rect 198804 402224 199404 410000
rect 216804 402224 217404 410000
rect 234804 402224 235404 410000
rect 252804 402224 253404 410000
rect 270804 402224 271404 410000
rect 280662 407010 280722 417830
rect 280294 406950 280722 407010
rect 280294 396130 280354 406950
rect 280110 396070 280354 396130
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 280110 389330 280170 396070
rect 280110 389270 280354 389330
rect 280294 379130 280354 389270
rect 280294 379070 280722 379130
rect 280662 369610 280722 379070
rect 280478 369550 280722 369610
rect 280478 366890 280538 369550
rect 280478 366830 281090 366890
rect 189763 351796 189829 351797
rect 189763 351732 189764 351796
rect 189828 351732 189829 351796
rect 189763 351731 189829 351732
rect 191051 351796 191117 351797
rect 191051 351732 191052 351796
rect 191116 351732 191117 351796
rect 191051 351731 191117 351732
rect 189579 351660 189645 351661
rect 189579 351596 189580 351660
rect 189644 351596 189645 351660
rect 189579 351595 189645 351596
rect 198804 348912 199404 358112
rect 216804 348912 217404 358112
rect 234804 348912 235404 358112
rect 252804 348912 253404 358112
rect 270804 348912 271404 358112
rect 281030 357645 281090 366830
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 280475 357644 280541 357645
rect 280475 357580 280476 357644
rect 280540 357580 280541 357644
rect 280475 357579 280541 357580
rect 281027 357644 281093 357645
rect 281027 357580 281028 357644
rect 281092 357580 281093 357644
rect 281027 357579 281093 357580
rect 280478 357370 280538 357579
rect 280478 357310 280906 357370
rect 280846 350437 280906 357310
rect 280291 350436 280357 350437
rect 280291 350372 280292 350436
rect 280356 350372 280357 350436
rect 280291 350371 280357 350372
rect 280843 350436 280909 350437
rect 280843 350372 280844 350436
rect 280908 350372 280909 350436
rect 280843 350371 280909 350372
rect 280294 347717 280354 350371
rect 280291 347716 280357 347717
rect 280291 347652 280292 347716
rect 280356 347652 280357 347716
rect 280291 347651 280357 347652
rect 107675 344454 107995 344476
rect 107675 344218 107717 344454
rect 107953 344218 107995 344454
rect 107675 344134 107995 344218
rect 107675 343898 107717 344134
rect 107953 343898 107995 344134
rect 107675 343876 107995 343898
rect 192805 344454 193125 344476
rect 192805 344218 192847 344454
rect 193083 344218 193125 344454
rect 192805 344134 193125 344218
rect 192805 343898 192847 344134
rect 193083 343898 193125 344134
rect 192805 343876 193125 343898
rect 280659 338196 280725 338197
rect 280659 338132 280660 338196
rect 280724 338132 280725 338196
rect 280659 338131 280725 338132
rect 280662 336701 280722 338131
rect 280659 336700 280725 336701
rect 280659 336636 280660 336700
rect 280724 336636 280725 336700
rect 280659 336635 280725 336636
rect 280291 336564 280357 336565
rect 280291 336500 280292 336564
rect 280356 336500 280357 336564
rect 280291 336499 280357 336500
rect 280294 327045 280354 336499
rect 280291 327044 280357 327045
rect 280291 326980 280292 327044
rect 280356 326980 280357 327044
rect 280291 326979 280357 326980
rect 65109 326454 65429 326476
rect 65109 326218 65151 326454
rect 65387 326218 65429 326454
rect 65109 326134 65429 326218
rect 65109 325898 65151 326134
rect 65387 325898 65429 326134
rect 65109 325876 65429 325898
rect 150240 326454 150560 326476
rect 150240 326218 150282 326454
rect 150518 326218 150560 326454
rect 150240 326134 150560 326218
rect 150240 325898 150282 326134
rect 150518 325898 150560 326134
rect 150240 325876 150560 325898
rect 235370 326454 235690 326476
rect 235370 326218 235412 326454
rect 235648 326218 235690 326454
rect 235370 326134 235690 326218
rect 235370 325898 235412 326134
rect 235648 325898 235690 326134
rect 235370 325876 235690 325898
rect 288804 326454 289404 361898
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 317091 700636 317157 700637
rect 317091 700572 317092 700636
rect 317156 700572 317157 700636
rect 317091 700571 317157 700572
rect 316907 700364 316973 700365
rect 316907 700300 316908 700364
rect 316972 700300 316973 700364
rect 316907 700299 316973 700300
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 316910 428637 316970 700299
rect 317094 428773 317154 700571
rect 317275 700500 317341 700501
rect 317275 700436 317276 700500
rect 317340 700436 317341 700500
rect 317275 700435 317341 700436
rect 317091 428772 317157 428773
rect 317091 428708 317092 428772
rect 317156 428708 317157 428772
rect 317091 428707 317157 428708
rect 316907 428636 316973 428637
rect 316907 428572 316908 428636
rect 316972 428572 316973 428636
rect 316907 428571 316973 428572
rect 317278 428501 317338 700435
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 657040 325404 685898
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 657040 343404 667898
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 657040 361404 685898
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 657040 379404 667898
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 657040 397404 685898
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 657040 415404 667898
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 657040 433404 685898
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 657040 451404 667898
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 662480 469404 685898
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 662480 487404 667898
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 492443 663916 492509 663917
rect 492443 663852 492444 663916
rect 492508 663852 492509 663916
rect 492443 663851 492509 663852
rect 323730 650454 324050 650476
rect 323730 650218 323772 650454
rect 324008 650218 324050 650454
rect 323730 650134 324050 650218
rect 323730 649898 323772 650134
rect 324008 649898 324050 650134
rect 323730 649876 324050 649898
rect 354450 650454 354770 650476
rect 354450 650218 354492 650454
rect 354728 650218 354770 650454
rect 354450 650134 354770 650218
rect 354450 649898 354492 650134
rect 354728 649898 354770 650134
rect 354450 649876 354770 649898
rect 385170 650454 385490 650476
rect 385170 650218 385212 650454
rect 385448 650218 385490 650454
rect 385170 650134 385490 650218
rect 385170 649898 385212 650134
rect 385448 649898 385490 650134
rect 385170 649876 385490 649898
rect 415890 650454 416210 650476
rect 415890 650218 415932 650454
rect 416168 650218 416210 650454
rect 415890 650134 416210 650218
rect 415890 649898 415932 650134
rect 416168 649898 416210 650134
rect 415890 649876 416210 649898
rect 446610 650454 446930 650476
rect 446610 650218 446652 650454
rect 446888 650218 446930 650454
rect 446610 650134 446930 650218
rect 446610 649898 446652 650134
rect 446888 649898 446930 650134
rect 446610 649876 446930 649898
rect 464208 650454 464528 650476
rect 464208 650218 464250 650454
rect 464486 650218 464528 650454
rect 464208 650134 464528 650218
rect 464208 649898 464250 650134
rect 464486 649898 464528 650134
rect 464208 649876 464528 649898
rect 339090 632454 339410 632476
rect 339090 632218 339132 632454
rect 339368 632218 339410 632454
rect 339090 632134 339410 632218
rect 339090 631898 339132 632134
rect 339368 631898 339410 632134
rect 339090 631876 339410 631898
rect 369810 632454 370130 632476
rect 369810 632218 369852 632454
rect 370088 632218 370130 632454
rect 369810 632134 370130 632218
rect 369810 631898 369852 632134
rect 370088 631898 370130 632134
rect 369810 631876 370130 631898
rect 400530 632454 400850 632476
rect 400530 632218 400572 632454
rect 400808 632218 400850 632454
rect 400530 632134 400850 632218
rect 400530 631898 400572 632134
rect 400808 631898 400850 632134
rect 400530 631876 400850 631898
rect 431250 632454 431570 632476
rect 431250 632218 431292 632454
rect 431528 632218 431570 632454
rect 431250 632134 431570 632218
rect 431250 631898 431292 632134
rect 431528 631898 431570 632134
rect 431250 631876 431570 631898
rect 479568 632454 479888 632476
rect 479568 632218 479610 632454
rect 479846 632218 479888 632454
rect 479568 632134 479888 632218
rect 479568 631898 479610 632134
rect 479846 631898 479888 632134
rect 479568 631876 479888 631898
rect 323730 614454 324050 614476
rect 323730 614218 323772 614454
rect 324008 614218 324050 614454
rect 323730 614134 324050 614218
rect 323730 613898 323772 614134
rect 324008 613898 324050 614134
rect 323730 613876 324050 613898
rect 354450 614454 354770 614476
rect 354450 614218 354492 614454
rect 354728 614218 354770 614454
rect 354450 614134 354770 614218
rect 354450 613898 354492 614134
rect 354728 613898 354770 614134
rect 354450 613876 354770 613898
rect 385170 614454 385490 614476
rect 385170 614218 385212 614454
rect 385448 614218 385490 614454
rect 385170 614134 385490 614218
rect 385170 613898 385212 614134
rect 385448 613898 385490 614134
rect 385170 613876 385490 613898
rect 415890 614454 416210 614476
rect 415890 614218 415932 614454
rect 416168 614218 416210 614454
rect 415890 614134 416210 614218
rect 415890 613898 415932 614134
rect 416168 613898 416210 614134
rect 415890 613876 416210 613898
rect 446610 614454 446930 614476
rect 446610 614218 446652 614454
rect 446888 614218 446930 614454
rect 446610 614134 446930 614218
rect 446610 613898 446652 614134
rect 446888 613898 446930 614134
rect 446610 613876 446930 613898
rect 464208 614454 464528 614476
rect 464208 614218 464250 614454
rect 464486 614218 464528 614454
rect 464208 614134 464528 614218
rect 464208 613898 464250 614134
rect 464486 613898 464528 614134
rect 464208 613876 464528 613898
rect 339090 596454 339410 596476
rect 339090 596218 339132 596454
rect 339368 596218 339410 596454
rect 339090 596134 339410 596218
rect 339090 595898 339132 596134
rect 339368 595898 339410 596134
rect 339090 595876 339410 595898
rect 369810 596454 370130 596476
rect 369810 596218 369852 596454
rect 370088 596218 370130 596454
rect 369810 596134 370130 596218
rect 369810 595898 369852 596134
rect 370088 595898 370130 596134
rect 369810 595876 370130 595898
rect 400530 596454 400850 596476
rect 400530 596218 400572 596454
rect 400808 596218 400850 596454
rect 400530 596134 400850 596218
rect 400530 595898 400572 596134
rect 400808 595898 400850 596134
rect 400530 595876 400850 595898
rect 431250 596454 431570 596476
rect 431250 596218 431292 596454
rect 431528 596218 431570 596454
rect 431250 596134 431570 596218
rect 431250 595898 431292 596134
rect 431528 595898 431570 596134
rect 431250 595876 431570 595898
rect 479568 596454 479888 596476
rect 479568 596218 479610 596454
rect 479846 596218 479888 596454
rect 479568 596134 479888 596218
rect 479568 595898 479610 596134
rect 479846 595898 479888 596134
rect 479568 595876 479888 595898
rect 323730 578454 324050 578476
rect 323730 578218 323772 578454
rect 324008 578218 324050 578454
rect 323730 578134 324050 578218
rect 323730 577898 323772 578134
rect 324008 577898 324050 578134
rect 323730 577876 324050 577898
rect 354450 578454 354770 578476
rect 354450 578218 354492 578454
rect 354728 578218 354770 578454
rect 354450 578134 354770 578218
rect 354450 577898 354492 578134
rect 354728 577898 354770 578134
rect 354450 577876 354770 577898
rect 385170 578454 385490 578476
rect 385170 578218 385212 578454
rect 385448 578218 385490 578454
rect 385170 578134 385490 578218
rect 385170 577898 385212 578134
rect 385448 577898 385490 578134
rect 385170 577876 385490 577898
rect 415890 578454 416210 578476
rect 415890 578218 415932 578454
rect 416168 578218 416210 578454
rect 415890 578134 416210 578218
rect 415890 577898 415932 578134
rect 416168 577898 416210 578134
rect 415890 577876 416210 577898
rect 446610 578454 446930 578476
rect 446610 578218 446652 578454
rect 446888 578218 446930 578454
rect 446610 578134 446930 578218
rect 446610 577898 446652 578134
rect 446888 577898 446930 578134
rect 446610 577876 446930 577898
rect 464208 578454 464528 578476
rect 464208 578218 464250 578454
rect 464486 578218 464528 578454
rect 464208 578134 464528 578218
rect 464208 577898 464250 578134
rect 464486 577898 464528 578134
rect 464208 577876 464528 577898
rect 324804 542454 325404 570000
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 528912 325404 541898
rect 342804 560454 343404 570000
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 528912 343404 559898
rect 360804 542454 361404 570000
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 528912 361404 541898
rect 378804 560454 379404 570000
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 528912 379404 559898
rect 396804 542454 397404 570000
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 528912 397404 541898
rect 414804 560454 415404 570000
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 528912 415404 559898
rect 432804 542454 433404 570000
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 528912 433404 541898
rect 450804 560454 451404 570000
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 528912 451404 559898
rect 468804 542454 469404 570000
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 528912 469404 541898
rect 486804 560454 487404 570000
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 528912 487404 559898
rect 492446 531181 492506 663851
rect 504804 662480 505404 685898
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 662480 523404 667898
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 662480 541404 685898
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 548379 662148 548445 662149
rect 548379 662084 548380 662148
rect 548444 662084 548445 662148
rect 548379 662083 548445 662084
rect 494928 650454 495248 650476
rect 494928 650218 494970 650454
rect 495206 650218 495248 650454
rect 494928 650134 495248 650218
rect 494928 649898 494970 650134
rect 495206 649898 495248 650134
rect 494928 649876 495248 649898
rect 525648 650454 525968 650476
rect 525648 650218 525690 650454
rect 525926 650218 525968 650454
rect 525648 650134 525968 650218
rect 525648 649898 525690 650134
rect 525926 649898 525968 650134
rect 525648 649876 525968 649898
rect 510288 632454 510608 632476
rect 510288 632218 510330 632454
rect 510566 632218 510608 632454
rect 510288 632134 510608 632218
rect 510288 631898 510330 632134
rect 510566 631898 510608 632134
rect 510288 631876 510608 631898
rect 541008 632454 541328 632476
rect 541008 632218 541050 632454
rect 541286 632218 541328 632454
rect 541008 632134 541328 632218
rect 541008 631898 541050 632134
rect 541286 631898 541328 632134
rect 541008 631876 541328 631898
rect 494928 614454 495248 614476
rect 494928 614218 494970 614454
rect 495206 614218 495248 614454
rect 494928 614134 495248 614218
rect 494928 613898 494970 614134
rect 495206 613898 495248 614134
rect 494928 613876 495248 613898
rect 525648 614454 525968 614476
rect 525648 614218 525690 614454
rect 525926 614218 525968 614454
rect 525648 614134 525968 614218
rect 525648 613898 525690 614134
rect 525926 613898 525968 614134
rect 525648 613876 525968 613898
rect 510288 596454 510608 596476
rect 510288 596218 510330 596454
rect 510566 596218 510608 596454
rect 510288 596134 510608 596218
rect 510288 595898 510330 596134
rect 510566 595898 510608 596134
rect 510288 595876 510608 595898
rect 541008 596454 541328 596476
rect 541008 596218 541050 596454
rect 541286 596218 541328 596454
rect 541008 596134 541328 596218
rect 541008 595898 541050 596134
rect 541286 595898 541328 596134
rect 541008 595876 541328 595898
rect 494928 578454 495248 578476
rect 494928 578218 494970 578454
rect 495206 578218 495248 578454
rect 494928 578134 495248 578218
rect 494928 577898 494970 578134
rect 495206 577898 495248 578134
rect 494928 577876 495248 577898
rect 525648 578454 525968 578476
rect 525648 578218 525690 578454
rect 525926 578218 525968 578454
rect 525648 578134 525968 578218
rect 525648 577898 525690 578134
rect 525926 577898 525968 578134
rect 525648 577876 525968 577898
rect 504804 542454 505404 570000
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 492443 531180 492509 531181
rect 492443 531116 492444 531180
rect 492508 531116 492509 531180
rect 492443 531115 492509 531116
rect 504804 528912 505404 541898
rect 522804 560454 523404 570000
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 528912 523404 559898
rect 540804 542454 541404 570000
rect 546355 569940 546421 569941
rect 546355 569876 546356 569940
rect 546420 569876 546421 569940
rect 546355 569875 546421 569876
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 528912 541404 541898
rect 546358 531317 546418 569875
rect 548382 560965 548442 662083
rect 551323 660108 551389 660109
rect 551323 660044 551324 660108
rect 551388 660044 551389 660108
rect 551323 660043 551389 660044
rect 551326 659970 551386 660043
rect 549854 659910 551386 659970
rect 549486 598858 549546 610862
rect 548379 560964 548445 560965
rect 548379 560900 548380 560964
rect 548444 560900 548445 560964
rect 548379 560899 548445 560900
rect 549854 534717 549914 659910
rect 551507 658884 551573 658885
rect 551507 658820 551508 658884
rect 551572 658820 551573 658884
rect 551507 658819 551573 658820
rect 551323 653172 551389 653173
rect 551323 653170 551324 653172
rect 550590 653110 551324 653170
rect 550590 649090 550650 653110
rect 551323 653108 551324 653110
rect 551388 653108 551389 653172
rect 551323 653107 551389 653108
rect 551510 649770 551570 658819
rect 553347 658204 553413 658205
rect 553347 658140 553348 658204
rect 553412 658140 553413 658204
rect 553347 658139 553413 658140
rect 552795 654532 552861 654533
rect 552795 654468 552796 654532
rect 552860 654468 552861 654532
rect 552795 654467 552861 654468
rect 552059 651540 552125 651541
rect 552059 651476 552060 651540
rect 552124 651476 552125 651540
rect 552059 651475 552125 651476
rect 550958 649710 551570 649770
rect 550590 649030 550834 649090
rect 550774 641610 550834 649030
rect 550590 641550 550834 641610
rect 550590 632770 550650 641550
rect 550958 636170 551018 649710
rect 551323 649092 551389 649093
rect 551323 649090 551324 649092
rect 551142 649030 551324 649090
rect 551142 639570 551202 649030
rect 551323 649028 551324 649030
rect 551388 649028 551389 649092
rect 551323 649027 551389 649028
rect 551323 645828 551389 645829
rect 551323 645764 551324 645828
rect 551388 645764 551389 645828
rect 551323 645763 551389 645764
rect 551326 639709 551386 645763
rect 551323 639708 551389 639709
rect 551323 639644 551324 639708
rect 551388 639644 551389 639708
rect 551323 639643 551389 639644
rect 551507 639572 551573 639573
rect 551507 639570 551508 639572
rect 551142 639510 551508 639570
rect 551507 639508 551508 639510
rect 551572 639508 551573 639572
rect 551507 639507 551573 639508
rect 551323 639436 551389 639437
rect 551323 639372 551324 639436
rect 551388 639372 551389 639436
rect 551323 639371 551389 639372
rect 551326 638890 551386 639371
rect 550038 632710 550650 632770
rect 550774 636110 551018 636170
rect 551142 638830 551386 638890
rect 550038 629370 550098 632710
rect 550774 629458 550834 636110
rect 550038 629310 550282 629370
rect 550222 628690 550282 629310
rect 550222 628630 550834 628690
rect 550222 610330 550282 627862
rect 550774 611098 550834 628630
rect 551142 624610 551202 638830
rect 551323 636036 551389 636037
rect 551323 635972 551324 636036
rect 551388 635972 551389 636036
rect 551323 635971 551389 635972
rect 551326 628013 551386 635971
rect 551875 634948 551941 634949
rect 551875 634884 551876 634948
rect 551940 634884 551941 634948
rect 551875 634883 551941 634884
rect 551323 628012 551389 628013
rect 551323 627948 551324 628012
rect 551388 627948 551389 628012
rect 551323 627947 551389 627948
rect 551691 628012 551757 628013
rect 551691 627948 551692 628012
rect 551756 627948 551757 628012
rect 551691 627947 551757 627948
rect 551142 624550 551386 624610
rect 551326 618629 551386 624550
rect 551323 618628 551389 618629
rect 551323 618564 551324 618628
rect 551388 618564 551389 618628
rect 551323 618563 551389 618564
rect 551694 618357 551754 627947
rect 551323 618356 551389 618357
rect 551323 618292 551324 618356
rect 551388 618292 551389 618356
rect 551323 618291 551389 618292
rect 551691 618356 551757 618357
rect 551691 618292 551692 618356
rect 551756 618292 551757 618356
rect 551691 618291 551757 618292
rect 551326 617810 551386 618291
rect 550958 617750 551386 617810
rect 550958 612370 551018 617750
rect 551323 617540 551389 617541
rect 551323 617476 551324 617540
rect 551388 617476 551389 617540
rect 551323 617475 551389 617476
rect 551326 617130 551386 617475
rect 551142 617070 551386 617130
rect 551142 613730 551202 617070
rect 551323 616452 551389 616453
rect 551323 616388 551324 616452
rect 551388 616388 551389 616452
rect 551323 616387 551389 616388
rect 551326 613869 551386 616387
rect 551323 613868 551389 613869
rect 551323 613804 551324 613868
rect 551388 613804 551389 613868
rect 551323 613803 551389 613804
rect 551323 613732 551389 613733
rect 551323 613730 551324 613732
rect 551142 613670 551324 613730
rect 551323 613668 551324 613670
rect 551388 613668 551389 613732
rect 551323 613667 551389 613668
rect 551507 612372 551573 612373
rect 551507 612370 551508 612372
rect 550958 612310 551508 612370
rect 551507 612308 551508 612310
rect 551572 612308 551573 612372
rect 551507 612307 551573 612308
rect 551691 612372 551757 612373
rect 551691 612308 551692 612372
rect 551756 612308 551757 612372
rect 551691 612307 551757 612308
rect 551323 612236 551389 612237
rect 551323 612172 551324 612236
rect 551388 612172 551389 612236
rect 551323 612171 551389 612172
rect 550222 610270 551018 610330
rect 550958 602986 551018 610270
rect 550406 602926 551018 602986
rect 550406 587210 550466 602926
rect 551326 599997 551386 612171
rect 551507 601220 551573 601221
rect 551507 601156 551508 601220
rect 551572 601156 551573 601220
rect 551507 601155 551573 601156
rect 551323 599996 551389 599997
rect 551323 599932 551324 599996
rect 551388 599932 551389 599996
rect 551323 599931 551389 599932
rect 551323 599588 551389 599589
rect 551323 599524 551324 599588
rect 551388 599524 551389 599588
rect 551323 599523 551389 599524
rect 550038 587150 550466 587210
rect 550038 585850 550098 587150
rect 550038 585790 550282 585850
rect 550222 575650 550282 585790
rect 550774 581770 550834 598622
rect 551326 596730 551386 599523
rect 551142 596670 551386 596730
rect 551142 588570 551202 596670
rect 551323 595100 551389 595101
rect 551323 595036 551324 595100
rect 551388 595036 551389 595100
rect 551323 595035 551389 595036
rect 551326 592245 551386 595035
rect 551510 592381 551570 601155
rect 551694 599589 551754 612307
rect 551691 599588 551757 599589
rect 551691 599524 551692 599588
rect 551756 599524 551757 599588
rect 551691 599523 551757 599524
rect 551691 595100 551757 595101
rect 551691 595036 551692 595100
rect 551756 595036 551757 595100
rect 551691 595035 551757 595036
rect 551507 592380 551573 592381
rect 551507 592316 551508 592380
rect 551572 592316 551573 592380
rect 551507 592315 551573 592316
rect 551323 592244 551389 592245
rect 551323 592180 551324 592244
rect 551388 592180 551389 592244
rect 551323 592179 551389 592180
rect 551142 588510 551386 588570
rect 551326 587213 551386 588510
rect 551323 587212 551389 587213
rect 551323 587148 551324 587212
rect 551388 587148 551389 587212
rect 551323 587147 551389 587148
rect 551323 586940 551389 586941
rect 551323 586876 551324 586940
rect 551388 586876 551389 586940
rect 551323 586875 551389 586876
rect 551326 586530 551386 586875
rect 550590 581710 550834 581770
rect 550958 586470 551386 586530
rect 550590 577010 550650 581710
rect 550958 578370 551018 586470
rect 551323 586260 551389 586261
rect 551323 586196 551324 586260
rect 551388 586196 551389 586260
rect 551323 586195 551389 586196
rect 551326 582181 551386 586195
rect 551507 582588 551573 582589
rect 551507 582524 551508 582588
rect 551572 582524 551573 582588
rect 551507 582523 551573 582524
rect 551323 582180 551389 582181
rect 551323 582116 551324 582180
rect 551388 582116 551389 582180
rect 551323 582115 551389 582116
rect 551510 578509 551570 582523
rect 551507 578508 551573 578509
rect 551507 578444 551508 578508
rect 551572 578444 551573 578508
rect 551507 578443 551573 578444
rect 550958 578310 551570 578370
rect 551323 578236 551389 578237
rect 551323 578172 551324 578236
rect 551388 578172 551389 578236
rect 551323 578171 551389 578172
rect 551326 577690 551386 578171
rect 550958 577630 551386 577690
rect 550590 576950 550834 577010
rect 550222 575590 550466 575650
rect 550406 569938 550466 575590
rect 550038 569878 550466 569938
rect 550038 562325 550098 569878
rect 550035 562324 550101 562325
rect 550035 562260 550036 562324
rect 550100 562260 550101 562324
rect 550035 562259 550101 562260
rect 550774 560285 550834 576950
rect 550958 560285 551018 577630
rect 551323 577556 551389 577557
rect 551323 577492 551324 577556
rect 551388 577492 551389 577556
rect 551323 577491 551389 577492
rect 551139 563276 551205 563277
rect 551139 563212 551140 563276
rect 551204 563212 551205 563276
rect 551139 563211 551205 563212
rect 550771 560284 550837 560285
rect 550771 560220 550772 560284
rect 550836 560220 550837 560284
rect 550771 560219 550837 560220
rect 550955 560284 551021 560285
rect 550955 560220 550956 560284
rect 551020 560220 551021 560284
rect 550955 560219 551021 560220
rect 551142 560149 551202 563211
rect 551139 560148 551205 560149
rect 551139 560084 551140 560148
rect 551204 560084 551205 560148
rect 551139 560083 551205 560084
rect 550771 560012 550837 560013
rect 550771 559948 550772 560012
rect 550836 559948 550837 560012
rect 550771 559947 550837 559948
rect 550587 548588 550653 548589
rect 550587 548524 550588 548588
rect 550652 548524 550653 548588
rect 550587 548523 550653 548524
rect 550590 538933 550650 548523
rect 550587 538932 550653 538933
rect 550587 538868 550588 538932
rect 550652 538868 550653 538932
rect 550587 538867 550653 538868
rect 549851 534716 549917 534717
rect 549851 534652 549852 534716
rect 549916 534652 549917 534716
rect 549851 534651 549917 534652
rect 546355 531316 546421 531317
rect 546355 531252 546356 531316
rect 546420 531252 546421 531316
rect 546355 531251 546421 531252
rect 550774 530773 550834 559947
rect 550955 555524 551021 555525
rect 550955 555460 550956 555524
rect 551020 555460 551021 555524
rect 550955 555459 551021 555460
rect 550958 532541 551018 555459
rect 551139 543828 551205 543829
rect 551139 543764 551140 543828
rect 551204 543764 551205 543828
rect 551139 543763 551205 543764
rect 551142 543693 551202 543763
rect 551139 543692 551205 543693
rect 551139 543628 551140 543692
rect 551204 543628 551205 543692
rect 551139 543627 551205 543628
rect 550955 532540 551021 532541
rect 550955 532476 550956 532540
rect 551020 532476 551021 532540
rect 550955 532475 551021 532476
rect 551326 531181 551386 577491
rect 551510 569941 551570 578310
rect 551507 569940 551573 569941
rect 551507 569876 551508 569940
rect 551572 569876 551573 569940
rect 551507 569875 551573 569876
rect 551694 569805 551754 595035
rect 551691 569804 551757 569805
rect 551691 569740 551692 569804
rect 551756 569740 551757 569804
rect 551691 569739 551757 569740
rect 551691 562324 551757 562325
rect 551691 562260 551692 562324
rect 551756 562260 551757 562324
rect 551691 562259 551757 562260
rect 551507 560148 551573 560149
rect 551507 560084 551508 560148
rect 551572 560084 551573 560148
rect 551507 560083 551573 560084
rect 551510 543829 551570 560083
rect 551694 548589 551754 562259
rect 551691 548588 551757 548589
rect 551691 548524 551692 548588
rect 551756 548524 551757 548588
rect 551691 548523 551757 548524
rect 551507 543828 551573 543829
rect 551507 543764 551508 543828
rect 551572 543764 551573 543828
rect 551507 543763 551573 543764
rect 551691 543692 551757 543693
rect 551691 543628 551692 543692
rect 551756 543628 551757 543692
rect 551691 543627 551757 543628
rect 551507 538932 551573 538933
rect 551507 538868 551508 538932
rect 551572 538868 551573 538932
rect 551507 538867 551573 538868
rect 551510 532269 551570 538867
rect 551507 532268 551573 532269
rect 551507 532204 551508 532268
rect 551572 532204 551573 532268
rect 551507 532203 551573 532204
rect 551323 531180 551389 531181
rect 551323 531116 551324 531180
rect 551388 531116 551389 531180
rect 551323 531115 551389 531116
rect 551694 531045 551754 543627
rect 551878 531861 551938 634883
rect 552062 533357 552122 651475
rect 552243 648412 552309 648413
rect 552243 648348 552244 648412
rect 552308 648348 552309 648412
rect 552243 648347 552309 648348
rect 552059 533356 552125 533357
rect 552059 533292 552060 533356
rect 552124 533292 552125 533356
rect 552059 533291 552125 533292
rect 552246 532677 552306 648347
rect 552427 647188 552493 647189
rect 552427 647124 552428 647188
rect 552492 647124 552493 647188
rect 552427 647123 552493 647124
rect 552430 533493 552490 647123
rect 552611 644740 552677 644741
rect 552611 644676 552612 644740
rect 552676 644676 552677 644740
rect 552611 644675 552677 644676
rect 552614 533629 552674 644675
rect 552798 545733 552858 654467
rect 552979 587212 553045 587213
rect 552979 587148 552980 587212
rect 553044 587148 553045 587212
rect 552979 587147 553045 587148
rect 552982 582589 553042 587147
rect 552979 582588 553045 582589
rect 552979 582524 552980 582588
rect 553044 582524 553045 582588
rect 552979 582523 553045 582524
rect 552795 545732 552861 545733
rect 552795 545668 552796 545732
rect 552860 545668 552861 545732
rect 552795 545667 552861 545668
rect 552611 533628 552677 533629
rect 552611 533564 552612 533628
rect 552676 533564 552677 533628
rect 552611 533563 552677 533564
rect 552427 533492 552493 533493
rect 552427 533428 552428 533492
rect 552492 533428 552493 533492
rect 552427 533427 552493 533428
rect 552243 532676 552309 532677
rect 552243 532612 552244 532676
rect 552308 532612 552309 532676
rect 552243 532611 552309 532612
rect 553350 531997 553410 658139
rect 553531 656980 553597 656981
rect 553531 656916 553532 656980
rect 553596 656916 553597 656980
rect 553531 656915 553597 656916
rect 553534 532133 553594 656915
rect 553715 655756 553781 655757
rect 553715 655692 553716 655756
rect 553780 655692 553781 655756
rect 553715 655691 553781 655692
rect 553718 532405 553778 655691
rect 553899 650860 553965 650861
rect 553899 650796 553900 650860
rect 553964 650796 553965 650860
rect 553899 650795 553965 650796
rect 553715 532404 553781 532405
rect 553715 532340 553716 532404
rect 553780 532340 553781 532404
rect 553715 532339 553781 532340
rect 553531 532132 553597 532133
rect 553531 532068 553532 532132
rect 553596 532068 553597 532132
rect 553531 532067 553597 532068
rect 553347 531996 553413 531997
rect 553347 531932 553348 531996
rect 553412 531932 553413 531996
rect 553347 531931 553413 531932
rect 551875 531860 551941 531861
rect 551875 531796 551876 531860
rect 551940 531796 551941 531860
rect 551875 531795 551941 531796
rect 551691 531044 551757 531045
rect 551691 530980 551692 531044
rect 551756 530980 551757 531044
rect 551691 530979 551757 530980
rect 550771 530772 550837 530773
rect 550771 530708 550772 530772
rect 550836 530708 550837 530772
rect 550771 530707 550837 530708
rect 553902 530637 553962 650795
rect 554083 643516 554149 643517
rect 554083 643452 554084 643516
rect 554148 643452 554149 643516
rect 554083 643451 554149 643452
rect 554086 530909 554146 643451
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 554083 530908 554149 530909
rect 554083 530844 554084 530908
rect 554148 530844 554149 530908
rect 554083 530843 554149 530844
rect 553899 530636 553965 530637
rect 553899 530572 553900 530636
rect 553964 530572 553965 530636
rect 553899 530571 553965 530572
rect 558804 528912 559404 559898
rect 576804 704838 577404 705800
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 403721 524454 404041 524476
rect 403721 524218 403763 524454
rect 403999 524218 404041 524454
rect 403721 524134 404041 524218
rect 403721 523898 403763 524134
rect 403999 523898 404041 524134
rect 403721 523876 404041 523898
rect 488851 524454 489171 524476
rect 488851 524218 488893 524454
rect 489129 524218 489171 524454
rect 488851 524134 489171 524218
rect 488851 523898 488893 524134
rect 489129 523898 489171 524134
rect 488851 523876 489171 523898
rect 361155 506454 361475 506476
rect 361155 506218 361197 506454
rect 361433 506218 361475 506454
rect 361155 506134 361475 506218
rect 361155 505898 361197 506134
rect 361433 505898 361475 506134
rect 361155 505876 361475 505898
rect 446286 506454 446606 506476
rect 446286 506218 446328 506454
rect 446564 506218 446606 506454
rect 446286 506134 446606 506218
rect 446286 505898 446328 506134
rect 446564 505898 446606 506134
rect 446286 505876 446606 505898
rect 531417 506454 531737 506476
rect 531417 506218 531459 506454
rect 531695 506218 531737 506454
rect 531417 506134 531737 506218
rect 531417 505898 531459 506134
rect 531695 505898 531737 506134
rect 531417 505876 531737 505898
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 324804 474240 325404 502800
rect 342804 488454 343404 502800
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 474240 343404 487898
rect 360804 474240 361404 502800
rect 378804 488454 379404 502800
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 474240 379404 487898
rect 396804 474240 397404 502800
rect 414804 488454 415404 502800
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 317275 428500 317341 428501
rect 317275 428436 317276 428500
rect 317340 428436 317341 428500
rect 317275 428435 317341 428436
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 20483 320788 20549 320789
rect 20483 320724 20484 320788
rect 20548 320724 20549 320788
rect 20483 320723 20549 320724
rect 36804 315600 37404 322800
rect 51579 320788 51645 320789
rect 51579 320724 51580 320788
rect 51644 320724 51645 320788
rect 51579 320723 51645 320724
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 39614 308454 39934 308476
rect 39614 308218 39656 308454
rect 39892 308218 39934 308454
rect 39614 308134 39934 308218
rect 39614 307898 39656 308134
rect 39892 307898 39934 308134
rect 39614 307876 39934 307898
rect 24254 290454 24574 290476
rect 24254 290218 24296 290454
rect 24532 290218 24574 290454
rect 24254 290134 24574 290218
rect 24254 289898 24296 290134
rect 24532 289898 24574 290134
rect 24254 289876 24574 289898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 39614 272454 39934 272476
rect 39614 272218 39656 272454
rect 39892 272218 39934 272454
rect 39614 272134 39934 272218
rect 39614 271898 39656 272134
rect 39892 271898 39934 272134
rect 39614 271876 39934 271898
rect 24254 254454 24574 254476
rect 24254 254218 24296 254454
rect 24532 254218 24574 254454
rect 24254 254134 24574 254218
rect 24254 253898 24296 254134
rect 24532 253898 24574 254134
rect 24254 253876 24574 253898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 51582 236061 51642 320723
rect 54804 315600 55404 322800
rect 72804 315600 73404 322800
rect 90804 315600 91404 322800
rect 108804 315600 109404 322800
rect 70334 308454 70654 308476
rect 70334 308218 70376 308454
rect 70612 308218 70654 308454
rect 70334 308134 70654 308218
rect 70334 307898 70376 308134
rect 70612 307898 70654 308134
rect 70334 307876 70654 307898
rect 101054 308454 101374 308476
rect 101054 308218 101096 308454
rect 101332 308218 101374 308454
rect 101054 308134 101374 308218
rect 101054 307898 101096 308134
rect 101332 307898 101374 308134
rect 101054 307876 101374 307898
rect 126804 308454 127404 322800
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 54974 290454 55294 290476
rect 54974 290218 55016 290454
rect 55252 290218 55294 290454
rect 54974 290134 55294 290218
rect 54974 289898 55016 290134
rect 55252 289898 55294 290134
rect 54974 289876 55294 289898
rect 85694 290454 86014 290476
rect 85694 290218 85736 290454
rect 85972 290218 86014 290454
rect 85694 290134 86014 290218
rect 85694 289898 85736 290134
rect 85972 289898 86014 290134
rect 85694 289876 86014 289898
rect 70334 272454 70654 272476
rect 70334 272218 70376 272454
rect 70612 272218 70654 272454
rect 70334 272134 70654 272218
rect 70334 271898 70376 272134
rect 70612 271898 70654 272134
rect 70334 271876 70654 271898
rect 101054 272454 101374 272476
rect 101054 272218 101096 272454
rect 101332 272218 101374 272454
rect 101054 272134 101374 272218
rect 101054 271898 101096 272134
rect 101332 271898 101374 272134
rect 101054 271876 101374 271898
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 54974 254454 55294 254476
rect 54974 254218 55016 254454
rect 55252 254218 55294 254454
rect 54974 254134 55294 254218
rect 54974 253898 55016 254134
rect 55252 253898 55294 254134
rect 54974 253876 55294 253898
rect 85694 254454 86014 254476
rect 85694 254218 85736 254454
rect 85972 254218 86014 254454
rect 85694 254134 86014 254218
rect 85694 253898 85736 254134
rect 85972 253898 86014 254134
rect 85694 253876 86014 253898
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 51579 236060 51645 236061
rect 51579 235996 51580 236060
rect 51644 235996 51645 236060
rect 51579 235995 51645 235996
rect 18804 219708 19404 235898
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 36804 219708 37404 234000
rect 54804 219708 55404 234000
rect 72804 219708 73404 234000
rect 90804 219708 91404 234000
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 108804 218454 109404 234000
rect 126804 221840 127404 235898
rect 144804 290454 145404 322800
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 221840 145404 253898
rect 162804 308454 163404 322800
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 221840 163404 235898
rect 180804 290454 181404 322800
rect 195099 320516 195165 320517
rect 195099 320452 195100 320516
rect 195164 320452 195165 320516
rect 195099 320451 195165 320452
rect 190315 320244 190381 320245
rect 190315 320180 190316 320244
rect 190380 320180 190381 320244
rect 190315 320179 190381 320180
rect 191603 320244 191669 320245
rect 191603 320180 191604 320244
rect 191668 320180 191669 320244
rect 191603 320179 191669 320180
rect 194363 320244 194429 320245
rect 194363 320180 194364 320244
rect 194428 320180 194429 320244
rect 194363 320179 194429 320180
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 181667 254012 181733 254013
rect 181667 253948 181668 254012
rect 181732 253948 181733 254012
rect 181667 253947 181733 253948
rect 180804 221840 181404 253898
rect 181670 253418 181730 253947
rect 190318 229805 190378 320179
rect 191606 233885 191666 320179
rect 192208 290454 192528 290476
rect 192208 290218 192250 290454
rect 192486 290218 192528 290454
rect 192208 290134 192528 290218
rect 192208 289898 192250 290134
rect 192486 289898 192528 290134
rect 192208 289876 192528 289898
rect 192208 254454 192528 254476
rect 192208 254218 192250 254454
rect 192486 254218 192528 254454
rect 192208 254134 192528 254218
rect 192208 253898 192250 254134
rect 192486 253898 192528 254134
rect 192208 253876 192528 253898
rect 194366 235245 194426 320179
rect 194363 235244 194429 235245
rect 194363 235180 194364 235244
rect 194428 235180 194429 235244
rect 194363 235179 194429 235180
rect 191603 233884 191669 233885
rect 191603 233820 191604 233884
rect 191668 233820 191669 233884
rect 191603 233819 191669 233820
rect 190315 229804 190381 229805
rect 190315 229740 190316 229804
rect 190380 229740 190381 229804
rect 190315 229739 190381 229740
rect 195102 228309 195162 320451
rect 196571 320380 196637 320381
rect 196571 320316 196572 320380
rect 196636 320316 196637 320380
rect 196571 320315 196637 320316
rect 196574 232525 196634 320315
rect 198804 315600 199404 322800
rect 214419 322148 214485 322149
rect 214419 322084 214420 322148
rect 214484 322084 214485 322148
rect 214419 322083 214485 322084
rect 208347 319428 208413 319429
rect 208347 319364 208348 319428
rect 208412 319364 208413 319428
rect 208347 319363 208413 319364
rect 207568 308454 207888 308476
rect 207568 308218 207610 308454
rect 207846 308218 207888 308454
rect 207568 308134 207888 308218
rect 207568 307898 207610 308134
rect 207846 307898 207888 308134
rect 207568 307876 207888 307898
rect 207568 272454 207888 272476
rect 207568 272218 207610 272454
rect 207846 272218 207888 272454
rect 207568 272134 207888 272218
rect 207568 271898 207610 272134
rect 207846 271898 207888 272134
rect 207568 271876 207888 271898
rect 196571 232524 196637 232525
rect 196571 232460 196572 232524
rect 196636 232460 196637 232524
rect 196571 232459 196637 232460
rect 195099 228308 195165 228309
rect 195099 228244 195100 228308
rect 195164 228244 195165 228308
rect 195099 228243 195165 228244
rect 198804 221840 199404 234000
rect 208350 223685 208410 319363
rect 208347 223684 208413 223685
rect 208347 223620 208348 223684
rect 208412 223620 208413 223684
rect 208347 223619 208413 223620
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 28768 200454 29088 200476
rect 28768 200218 28810 200454
rect 29046 200218 29088 200454
rect 28768 200134 29088 200218
rect 28768 199898 28810 200134
rect 29046 199898 29088 200134
rect 28768 199876 29088 199898
rect 59488 200454 59808 200476
rect 59488 200218 59530 200454
rect 59766 200218 59808 200454
rect 59488 200134 59808 200218
rect 59488 199898 59530 200134
rect 59766 199898 59808 200134
rect 59488 199876 59808 199898
rect 90208 200454 90528 200476
rect 90208 200218 90250 200454
rect 90486 200218 90528 200454
rect 90208 200134 90528 200218
rect 90208 199898 90250 200134
rect 90486 199898 90528 200134
rect 90208 199876 90528 199898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 13408 182454 13728 182476
rect 13408 182218 13450 182454
rect 13686 182218 13728 182454
rect 13408 182134 13728 182218
rect 13408 181898 13450 182134
rect 13686 181898 13728 182134
rect 13408 181876 13728 181898
rect 44128 182454 44448 182476
rect 44128 182218 44170 182454
rect 44406 182218 44448 182454
rect 44128 182134 44448 182218
rect 44128 181898 44170 182134
rect 44406 181898 44448 182134
rect 44128 181876 44448 181898
rect 74848 182454 75168 182476
rect 74848 182218 74890 182454
rect 75126 182218 75168 182454
rect 74848 182134 75168 182218
rect 74848 181898 74890 182134
rect 75126 181898 75168 182134
rect 74848 181876 75168 181898
rect 108804 182454 109404 217898
rect 123808 218454 124128 218476
rect 123808 218218 123850 218454
rect 124086 218218 124128 218454
rect 123808 218134 124128 218218
rect 123808 217898 123850 218134
rect 124086 217898 124128 218134
rect 123808 217876 124128 217898
rect 154528 218454 154848 218476
rect 154528 218218 154570 218454
rect 154806 218218 154848 218454
rect 154528 218134 154848 218218
rect 154528 217898 154570 218134
rect 154806 217898 154848 218134
rect 154528 217876 154848 217898
rect 185248 218454 185568 218476
rect 185248 218218 185290 218454
rect 185526 218218 185568 218454
rect 185248 218134 185568 218218
rect 185248 217898 185290 218134
rect 185526 217898 185568 218134
rect 185248 217876 185568 217898
rect 139168 200454 139488 200476
rect 139168 200218 139210 200454
rect 139446 200218 139488 200454
rect 139168 200134 139488 200218
rect 139168 199898 139210 200134
rect 139446 199898 139488 200134
rect 139168 199876 139488 199898
rect 169888 200454 170208 200476
rect 169888 200218 169930 200454
rect 170166 200218 170208 200454
rect 169888 200134 170208 200218
rect 169888 199898 169930 200134
rect 170166 199898 170208 200134
rect 169888 199876 170208 199898
rect 200608 200454 200928 200476
rect 200608 200218 200650 200454
rect 200886 200218 200928 200454
rect 200608 200134 200928 200218
rect 200608 199898 200650 200134
rect 200886 199898 200928 200134
rect 200608 199876 200928 199898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 28768 164454 29088 164476
rect 28768 164218 28810 164454
rect 29046 164218 29088 164454
rect 28768 164134 29088 164218
rect 28768 163898 28810 164134
rect 29046 163898 29088 164134
rect 28768 163876 29088 163898
rect 59488 164454 59808 164476
rect 59488 164218 59530 164454
rect 59766 164218 59808 164454
rect 59488 164134 59808 164218
rect 59488 163898 59530 164134
rect 59766 163898 59808 164134
rect 59488 163876 59808 163898
rect 90208 164454 90528 164476
rect 90208 164218 90250 164454
rect 90486 164218 90528 164454
rect 90208 164134 90528 164218
rect 90208 163898 90250 164134
rect 90486 163898 90528 164134
rect 90208 163876 90528 163898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 13408 146454 13728 146476
rect 13408 146218 13450 146454
rect 13686 146218 13728 146454
rect 13408 146134 13728 146218
rect 13408 145898 13450 146134
rect 13686 145898 13728 146134
rect 13408 145876 13728 145898
rect 44128 146454 44448 146476
rect 44128 146218 44170 146454
rect 44406 146218 44448 146454
rect 44128 146134 44448 146218
rect 44128 145898 44170 146134
rect 44406 145898 44448 146134
rect 44128 145876 44448 145898
rect 74848 146454 75168 146476
rect 74848 146218 74890 146454
rect 75126 146218 75168 146454
rect 74848 146134 75168 146218
rect 74848 145898 74890 146134
rect 75126 145898 75168 146134
rect 74848 145876 75168 145898
rect 108804 146454 109404 181898
rect 123808 182454 124128 182476
rect 123808 182218 123850 182454
rect 124086 182218 124128 182454
rect 123808 182134 124128 182218
rect 123808 181898 123850 182134
rect 124086 181898 124128 182134
rect 123808 181876 124128 181898
rect 154528 182454 154848 182476
rect 154528 182218 154570 182454
rect 154806 182218 154848 182454
rect 154528 182134 154848 182218
rect 154528 181898 154570 182134
rect 154806 181898 154848 182134
rect 154528 181876 154848 181898
rect 185248 182454 185568 182476
rect 185248 182218 185290 182454
rect 185526 182218 185568 182454
rect 185248 182134 185568 182218
rect 185248 181898 185290 182134
rect 185526 181898 185568 182134
rect 185248 181876 185568 181898
rect 139168 164454 139488 164476
rect 139168 164218 139210 164454
rect 139446 164218 139488 164454
rect 139168 164134 139488 164218
rect 139168 163898 139210 164134
rect 139446 163898 139488 164134
rect 139168 163876 139488 163898
rect 169888 164454 170208 164476
rect 169888 164218 169930 164454
rect 170166 164218 170208 164454
rect 169888 164134 170208 164218
rect 169888 163898 169930 164134
rect 170166 163898 170208 164134
rect 169888 163876 170208 163898
rect 200608 164454 200928 164476
rect 200608 164218 200650 164454
rect 200886 164218 200928 164454
rect 200608 164134 200928 164218
rect 200608 163898 200650 164134
rect 200886 163898 200928 164134
rect 200608 163876 200928 163898
rect 214422 159493 214482 322083
rect 216804 315600 217404 322800
rect 234804 315600 235404 322800
rect 252804 315600 253404 322800
rect 270804 315600 271404 322800
rect 280291 317660 280357 317661
rect 280291 317596 280292 317660
rect 280356 317596 280357 317660
rect 280291 317595 280357 317596
rect 280294 317389 280354 317595
rect 280291 317388 280357 317389
rect 280291 317324 280292 317388
rect 280356 317324 280357 317388
rect 280291 317323 280357 317324
rect 280291 309636 280357 309637
rect 280291 309572 280292 309636
rect 280356 309572 280357 309636
rect 280291 309571 280357 309572
rect 238288 308454 238608 308476
rect 238288 308218 238330 308454
rect 238566 308218 238608 308454
rect 238288 308134 238608 308218
rect 238288 307898 238330 308134
rect 238566 307898 238608 308134
rect 238288 307876 238608 307898
rect 269008 308454 269328 308476
rect 269008 308218 269050 308454
rect 269286 308218 269328 308454
rect 269008 308134 269328 308218
rect 269008 307898 269050 308134
rect 269286 307898 269328 308134
rect 269008 307876 269328 307898
rect 280294 306373 280354 309571
rect 280291 306372 280357 306373
rect 280291 306308 280292 306372
rect 280356 306308 280357 306372
rect 280291 306307 280357 306308
rect 280475 306372 280541 306373
rect 280475 306308 280476 306372
rect 280540 306308 280541 306372
rect 280475 306307 280541 306308
rect 280478 296850 280538 306307
rect 280478 296790 280722 296850
rect 280662 296717 280722 296790
rect 280659 296716 280725 296717
rect 280659 296652 280660 296716
rect 280724 296652 280725 296716
rect 280659 296651 280725 296652
rect 281027 296716 281093 296717
rect 281027 296652 281028 296716
rect 281092 296652 281093 296716
rect 281027 296651 281093 296652
rect 281030 295221 281090 296651
rect 281027 295220 281093 295221
rect 281027 295156 281028 295220
rect 281092 295156 281093 295220
rect 281027 295155 281093 295156
rect 222928 290454 223248 290476
rect 222928 290218 222970 290454
rect 223206 290218 223248 290454
rect 222928 290134 223248 290218
rect 222928 289898 222970 290134
rect 223206 289898 223248 290134
rect 222928 289876 223248 289898
rect 253648 290454 253968 290476
rect 253648 290218 253690 290454
rect 253926 290218 253968 290454
rect 253648 290134 253968 290218
rect 253648 289898 253690 290134
rect 253926 289898 253968 290134
rect 253648 289876 253968 289898
rect 288804 290454 289404 325898
rect 293189 326454 293509 326476
rect 293189 326218 293231 326454
rect 293467 326218 293509 326454
rect 293189 326134 293509 326218
rect 293189 325898 293231 326134
rect 293467 325898 293509 326134
rect 293189 325876 293509 325898
rect 294635 308454 294955 308476
rect 294635 308218 294677 308454
rect 294913 308218 294955 308454
rect 294635 308134 294955 308218
rect 294635 307898 294677 308134
rect 294913 307898 294955 308134
rect 294635 307876 294955 307898
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 280475 277540 280541 277541
rect 280475 277476 280476 277540
rect 280540 277476 280541 277540
rect 280475 277475 280541 277476
rect 280478 273461 280538 277475
rect 280475 273460 280541 273461
rect 280475 273396 280476 273460
rect 280540 273396 280541 273460
rect 280475 273395 280541 273396
rect 280291 273188 280357 273189
rect 280291 273124 280292 273188
rect 280356 273124 280357 273188
rect 280291 273123 280357 273124
rect 238288 272454 238608 272476
rect 238288 272218 238330 272454
rect 238566 272218 238608 272454
rect 238288 272134 238608 272218
rect 238288 271898 238330 272134
rect 238566 271898 238608 272134
rect 238288 271876 238608 271898
rect 269008 272454 269328 272476
rect 269008 272218 269050 272454
rect 269286 272218 269328 272454
rect 269008 272134 269328 272218
rect 269008 271898 269050 272134
rect 269286 271898 269328 272134
rect 269008 271876 269328 271898
rect 280294 259589 280354 273123
rect 280291 259588 280357 259589
rect 280291 259524 280292 259588
rect 280356 259524 280357 259588
rect 280291 259523 280357 259524
rect 280475 259588 280541 259589
rect 280475 259524 280476 259588
rect 280540 259524 280541 259588
rect 280475 259523 280541 259524
rect 222928 254454 223248 254476
rect 222928 254218 222970 254454
rect 223206 254218 223248 254454
rect 222928 254134 223248 254218
rect 222928 253898 222970 254134
rect 223206 253898 223248 254134
rect 222928 253876 223248 253898
rect 253648 254454 253968 254476
rect 253648 254218 253690 254454
rect 253926 254218 253968 254454
rect 253648 254134 253968 254218
rect 253648 253898 253690 254134
rect 253926 253898 253968 254134
rect 279371 254012 279437 254013
rect 279371 253948 279372 254012
rect 279436 253948 279437 254012
rect 279371 253947 279437 253948
rect 253648 253876 253968 253898
rect 279374 252058 279434 253947
rect 280478 251157 280538 259523
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 280475 251156 280541 251157
rect 280475 251092 280476 251156
rect 280540 251092 280541 251156
rect 280475 251091 280541 251092
rect 280659 241636 280725 241637
rect 280659 241572 280660 241636
rect 280724 241572 280725 241636
rect 280659 241571 280725 241572
rect 280662 235245 280722 241571
rect 280659 235244 280725 235245
rect 280659 235180 280660 235244
rect 280724 235180 280725 235244
rect 280659 235179 280725 235180
rect 216804 218454 217404 234000
rect 234804 221680 235404 234000
rect 252804 221680 253404 234000
rect 270804 221680 271404 234000
rect 288804 221680 289404 253898
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 221680 307404 235898
rect 324804 398454 325404 430128
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 342804 416454 343404 430128
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 380454 343404 415898
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 332915 302836 332981 302837
rect 332915 302772 332916 302836
rect 332980 302772 332981 302836
rect 332915 302771 332981 302772
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 221680 325404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 214419 159492 214485 159493
rect 214419 159428 214420 159492
rect 214484 159428 214485 159492
rect 214419 159427 214485 159428
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 18804 99440 19404 127228
rect 32259 125084 32325 125085
rect 32259 125020 32260 125084
rect 32324 125020 32325 125084
rect 32259 125019 32325 125020
rect 28768 92454 29088 92476
rect 28768 92218 28810 92454
rect 29046 92218 29088 92454
rect 28768 92134 29088 92218
rect 28768 91898 28810 92134
rect 29046 91898 29088 92134
rect 28768 91876 29088 91898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 13408 74454 13728 74476
rect 13408 74218 13450 74454
rect 13686 74218 13728 74454
rect 13408 74134 13728 74218
rect 13408 73898 13450 74134
rect 13686 73898 13728 74134
rect 13408 73876 13728 73898
rect 28768 56454 29088 56476
rect 28768 56218 28810 56454
rect 29046 56218 29088 56454
rect 28768 56134 29088 56218
rect 28768 55898 28810 56134
rect 29046 55898 29088 56134
rect 28768 55876 29088 55898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 13408 38454 13728 38476
rect 13408 38218 13450 38454
rect 13686 38218 13728 38454
rect 13408 38134 13728 38218
rect 13408 37898 13450 38134
rect 13686 37898 13728 38134
rect 13408 37876 13728 37898
rect 32262 31789 32322 125019
rect 36804 110454 37404 127228
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 99440 37404 109898
rect 54804 99440 55404 127228
rect 72804 110454 73404 127228
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 99440 73404 109898
rect 90804 99440 91404 127228
rect 108804 110454 109404 145898
rect 123808 146454 124128 146476
rect 123808 146218 123850 146454
rect 124086 146218 124128 146454
rect 123808 146134 124128 146218
rect 123808 145898 123850 146134
rect 124086 145898 124128 146134
rect 123808 145876 124128 145898
rect 154528 146454 154848 146476
rect 154528 146218 154570 146454
rect 154806 146218 154848 146454
rect 154528 146134 154848 146218
rect 154528 145898 154570 146134
rect 154806 145898 154848 146134
rect 154528 145876 154848 145898
rect 185248 146454 185568 146476
rect 185248 146218 185290 146454
rect 185526 146218 185568 146454
rect 185248 146134 185568 146218
rect 185248 145898 185290 146134
rect 185526 145898 185568 146134
rect 185248 145876 185568 145898
rect 216804 146454 217404 181898
rect 234804 164454 235404 175440
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 149680 235404 163898
rect 252804 149680 253404 175440
rect 270804 164454 271404 175440
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 149680 271404 163898
rect 288804 149680 289404 175440
rect 306804 164454 307404 175440
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 149680 307404 163898
rect 324804 149680 325404 175440
rect 332918 173909 332978 302771
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 332915 173908 332981 173909
rect 332915 173844 332916 173908
rect 332980 173844 332981 173908
rect 332915 173843 332981 173844
rect 342804 164454 343404 199898
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 139168 128454 139488 128476
rect 139168 128218 139210 128454
rect 139446 128218 139488 128454
rect 139168 128134 139488 128218
rect 139168 127898 139210 128134
rect 139446 127898 139488 128134
rect 139168 127876 139488 127898
rect 169888 128454 170208 128476
rect 169888 128218 169930 128454
rect 170166 128218 170208 128454
rect 169888 128134 170208 128218
rect 169888 127898 169930 128134
rect 170166 127898 170208 128134
rect 169888 127876 170208 127898
rect 200608 128454 200928 128476
rect 200608 128218 200650 128454
rect 200886 128218 200928 128454
rect 200608 128134 200928 128218
rect 200608 127898 200650 128134
rect 200886 127898 200928 128134
rect 200608 127876 200928 127898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 59488 92454 59808 92476
rect 59488 92218 59530 92454
rect 59766 92218 59808 92454
rect 59488 92134 59808 92218
rect 59488 91898 59530 92134
rect 59766 91898 59808 92134
rect 59488 91876 59808 91898
rect 90208 92454 90528 92476
rect 90208 92218 90250 92454
rect 90486 92218 90528 92454
rect 90208 92134 90528 92218
rect 90208 91898 90250 92134
rect 90486 91898 90528 92134
rect 90208 91876 90528 91898
rect 44128 74454 44448 74476
rect 44128 74218 44170 74454
rect 44406 74218 44448 74454
rect 44128 74134 44448 74218
rect 44128 73898 44170 74134
rect 44406 73898 44448 74134
rect 44128 73876 44448 73898
rect 74848 74454 75168 74476
rect 74848 74218 74890 74454
rect 75126 74218 75168 74454
rect 74848 74134 75168 74218
rect 74848 73898 74890 74134
rect 75126 73898 75168 74134
rect 74848 73876 75168 73898
rect 108804 74454 109404 109898
rect 123808 110454 124128 110476
rect 123808 110218 123850 110454
rect 124086 110218 124128 110454
rect 123808 110134 124128 110218
rect 123808 109898 123850 110134
rect 124086 109898 124128 110134
rect 123808 109876 124128 109898
rect 154528 110454 154848 110476
rect 154528 110218 154570 110454
rect 154806 110218 154848 110454
rect 154528 110134 154848 110218
rect 154528 109898 154570 110134
rect 154806 109898 154848 110134
rect 154528 109876 154848 109898
rect 185248 110454 185568 110476
rect 185248 110218 185290 110454
rect 185526 110218 185568 110454
rect 185248 110134 185568 110218
rect 185248 109898 185290 110134
rect 185526 109898 185568 110134
rect 185248 109876 185568 109898
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 139168 92454 139488 92476
rect 139168 92218 139210 92454
rect 139446 92218 139488 92454
rect 139168 92134 139488 92218
rect 139168 91898 139210 92134
rect 139446 91898 139488 92134
rect 139168 91876 139488 91898
rect 169888 92454 170208 92476
rect 169888 92218 169930 92454
rect 170166 92218 170208 92454
rect 169888 92134 170208 92218
rect 169888 91898 169930 92134
rect 170166 91898 170208 92134
rect 169888 91876 170208 91898
rect 200608 92454 200928 92476
rect 200608 92218 200650 92454
rect 200886 92218 200928 92454
rect 200608 92134 200928 92218
rect 200608 91898 200650 92134
rect 200886 91898 200928 92134
rect 200608 91876 200928 91898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 59488 56454 59808 56476
rect 59488 56218 59530 56454
rect 59766 56218 59808 56454
rect 59488 56134 59808 56218
rect 59488 55898 59530 56134
rect 59766 55898 59808 56134
rect 59488 55876 59808 55898
rect 90208 56454 90528 56476
rect 90208 56218 90250 56454
rect 90486 56218 90528 56454
rect 90208 56134 90528 56218
rect 90208 55898 90250 56134
rect 90486 55898 90528 56134
rect 90208 55876 90528 55898
rect 44128 38454 44448 38476
rect 44128 38218 44170 38454
rect 44406 38218 44448 38454
rect 44128 38134 44448 38218
rect 44128 37898 44170 38134
rect 44406 37898 44448 38134
rect 44128 37876 44448 37898
rect 74848 38454 75168 38476
rect 74848 38218 74890 38454
rect 75126 38218 75168 38454
rect 74848 38134 75168 38218
rect 74848 37898 74890 38134
rect 75126 37898 75168 38134
rect 74848 37876 75168 37898
rect 108804 38454 109404 73898
rect 123808 74454 124128 74476
rect 123808 74218 123850 74454
rect 124086 74218 124128 74454
rect 123808 74134 124128 74218
rect 123808 73898 123850 74134
rect 124086 73898 124128 74134
rect 123808 73876 124128 73898
rect 154528 74454 154848 74476
rect 154528 74218 154570 74454
rect 154806 74218 154848 74454
rect 154528 74134 154848 74218
rect 154528 73898 154570 74134
rect 154806 73898 154848 74134
rect 154528 73876 154848 73898
rect 185248 74454 185568 74476
rect 185248 74218 185290 74454
rect 185526 74218 185568 74454
rect 185248 74134 185568 74218
rect 185248 73898 185290 74134
rect 185526 73898 185568 74134
rect 185248 73876 185568 73898
rect 216804 74454 217404 109898
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 234804 92454 235404 103440
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 81488 235404 91898
rect 252804 81488 253404 103440
rect 270804 92454 271404 103440
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 81488 271404 91898
rect 288804 81488 289404 103440
rect 306804 92454 307404 103440
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 81488 307404 91898
rect 324804 81488 325404 103440
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 139168 56454 139488 56476
rect 139168 56218 139210 56454
rect 139446 56218 139488 56454
rect 139168 56134 139488 56218
rect 139168 55898 139210 56134
rect 139446 55898 139488 56134
rect 139168 55876 139488 55898
rect 169888 56454 170208 56476
rect 169888 56218 169930 56454
rect 170166 56218 170208 56454
rect 169888 56134 170208 56218
rect 169888 55898 169930 56134
rect 170166 55898 170208 56134
rect 169888 55876 170208 55898
rect 200608 56454 200928 56476
rect 200608 56218 200650 56454
rect 200886 56218 200928 56454
rect 200608 56134 200928 56218
rect 200608 55898 200650 56134
rect 200886 55898 200928 56134
rect 200608 55876 200928 55898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 32259 31788 32325 31789
rect 32259 31724 32260 31788
rect 32324 31724 32325 31788
rect 32259 31723 32325 31724
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 18804 20454 19404 31440
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 36804 2454 37404 31440
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 54804 20454 55404 31440
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 72804 2454 73404 31440
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 90804 20454 91404 31440
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 108804 2454 109404 37898
rect 123808 38454 124128 38476
rect 123808 38218 123850 38454
rect 124086 38218 124128 38454
rect 123808 38134 124128 38218
rect 123808 37898 123850 38134
rect 124086 37898 124128 38134
rect 123808 37876 124128 37898
rect 154528 38454 154848 38476
rect 154528 38218 154570 38454
rect 154806 38218 154848 38454
rect 154528 38134 154848 38218
rect 154528 37898 154570 38134
rect 154806 37898 154848 38134
rect 154528 37876 154848 37898
rect 185248 38454 185568 38476
rect 185248 38218 185290 38454
rect 185526 38218 185568 38454
rect 185248 38134 185568 38218
rect 185248 37898 185290 38134
rect 185526 37898 185568 38134
rect 185248 37876 185568 37898
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 126804 20454 127404 31440
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 144804 2454 145404 31440
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 162804 20454 163404 31440
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 180804 2454 181404 31440
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 198804 20454 199404 31440
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 216804 2454 217404 37898
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 234804 20454 235404 31440
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 252804 2454 253404 31440
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 270804 20454 271404 31440
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 288804 2454 289404 31440
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 306804 20454 307404 31440
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 324804 2454 325404 31440
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 360804 398454 361404 430128
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 362454 361404 397898
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 182454 361404 217898
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 378804 416454 379404 430128
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 380454 379404 415898
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 396804 398454 397404 430128
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 362454 397404 397898
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 60928 415404 91898
rect 432804 470454 433404 502800
rect 450804 488454 451404 502800
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 473680 451404 487898
rect 468804 473680 469404 502800
rect 486804 488454 487404 502800
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 473680 487404 487898
rect 504804 473680 505404 502800
rect 522804 488454 523404 502800
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 473680 523404 487898
rect 540804 473680 541404 502800
rect 548379 500716 548445 500717
rect 548379 500652 548380 500716
rect 548444 500652 548445 500716
rect 548379 500651 548445 500652
rect 546539 500444 546605 500445
rect 546539 500380 546540 500444
rect 546604 500380 546605 500444
rect 546539 500379 546605 500380
rect 546542 473517 546602 500379
rect 546539 473516 546605 473517
rect 546539 473452 546540 473516
rect 546604 473452 546605 473516
rect 546539 473451 546605 473452
rect 548382 472378 548442 500651
rect 549851 500580 549917 500581
rect 549851 500516 549852 500580
rect 549916 500516 549917 500580
rect 549851 500515 549917 500516
rect 549854 473058 549914 500515
rect 550587 500308 550653 500309
rect 550587 500244 550588 500308
rect 550652 500244 550653 500308
rect 550587 500243 550653 500244
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 550590 468210 550650 500243
rect 550771 500172 550837 500173
rect 550771 500108 550772 500172
rect 550836 500108 550837 500172
rect 550771 500107 550837 500108
rect 550774 470250 550834 500107
rect 558804 488454 559404 502800
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 553347 475556 553413 475557
rect 553347 475492 553348 475556
rect 553412 475492 553413 475556
rect 553347 475491 553413 475492
rect 552059 475420 552125 475421
rect 552059 475356 552060 475420
rect 552124 475356 552125 475420
rect 552059 475355 552125 475356
rect 552062 471885 552122 475355
rect 552059 471884 552125 471885
rect 552059 471820 552060 471884
rect 552124 471820 552125 471884
rect 552059 471819 552125 471820
rect 550774 470190 552122 470250
rect 552062 470117 552122 470190
rect 552059 470116 552125 470117
rect 552059 470052 552060 470116
rect 552124 470052 552125 470116
rect 552059 470051 552125 470052
rect 552059 468348 552125 468349
rect 552059 468284 552060 468348
rect 552124 468284 552125 468348
rect 552059 468283 552125 468284
rect 552062 468210 552122 468283
rect 550590 468150 552122 468210
rect 553350 464541 553410 475491
rect 553347 464540 553413 464541
rect 553347 464476 553348 464540
rect 553412 464476 553413 464540
rect 553347 464475 553413 464476
rect 554822 460325 554882 472822
rect 555190 461549 555250 472142
rect 555187 461548 555253 461549
rect 555187 461484 555188 461548
rect 555252 461484 555253 461548
rect 555187 461483 555253 461484
rect 554819 460324 554885 460325
rect 554819 460260 554820 460324
rect 554884 460260 554885 460324
rect 554819 460259 554885 460260
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 60928 433404 73898
rect 450804 416454 451404 427440
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 60928 451404 91898
rect 468804 398454 469404 427440
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 60928 469404 73898
rect 486804 416454 487404 427440
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 60928 487404 91898
rect 504804 398454 505404 427440
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 60928 505404 73898
rect 522804 416454 523404 427440
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 60928 523404 91898
rect 540804 398454 541404 427440
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 60928 541404 73898
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 60928 559404 91898
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 433568 56454 433888 56476
rect 433568 56218 433610 56454
rect 433846 56218 433888 56454
rect 433568 56134 433888 56218
rect 433568 55898 433610 56134
rect 433846 55898 433888 56134
rect 433568 55876 433888 55898
rect 464288 56454 464608 56476
rect 464288 56218 464330 56454
rect 464566 56218 464608 56454
rect 464288 56134 464608 56218
rect 464288 55898 464330 56134
rect 464566 55898 464608 56134
rect 464288 55876 464608 55898
rect 495008 56454 495328 56476
rect 495008 56218 495050 56454
rect 495286 56218 495328 56454
rect 495008 56134 495328 56218
rect 495008 55898 495050 56134
rect 495286 55898 495328 56134
rect 495008 55876 495328 55898
rect 525728 56454 526048 56476
rect 525728 56218 525770 56454
rect 526006 56218 526048 56454
rect 525728 56134 526048 56218
rect 525728 55898 525770 56134
rect 526006 55898 526048 56134
rect 525728 55876 526048 55898
rect 556448 56454 556768 56476
rect 556448 56218 556490 56454
rect 556726 56218 556768 56454
rect 556448 56134 556768 56218
rect 556448 55898 556490 56134
rect 556726 55898 556768 56134
rect 556448 55876 556768 55898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 418208 38454 418528 38476
rect 418208 38218 418250 38454
rect 418486 38218 418528 38454
rect 418208 38134 418528 38218
rect 418208 37898 418250 38134
rect 418486 37898 418528 38134
rect 418208 37876 418528 37898
rect 448928 38454 449248 38476
rect 448928 38218 448970 38454
rect 449206 38218 449248 38454
rect 448928 38134 449248 38218
rect 448928 37898 448970 38134
rect 449206 37898 449248 38134
rect 448928 37876 449248 37898
rect 479648 38454 479968 38476
rect 479648 38218 479690 38454
rect 479926 38218 479968 38454
rect 479648 38134 479968 38218
rect 479648 37898 479690 38134
rect 479926 37898 479968 38134
rect 479648 37876 479968 37898
rect 510368 38454 510688 38476
rect 510368 38218 510410 38454
rect 510646 38218 510688 38454
rect 510368 38134 510688 38218
rect 510368 37898 510410 38134
rect 510646 37898 510688 38134
rect 510368 37876 510688 37898
rect 541088 38454 541408 38476
rect 541088 38218 541130 38454
rect 541366 38218 541408 38454
rect 541088 38134 541408 38218
rect 541088 37898 541130 38134
rect 541366 37898 541408 38134
rect 541088 37876 541408 37898
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 433568 20454 433888 20476
rect 433568 20218 433610 20454
rect 433846 20218 433888 20454
rect 433568 20134 433888 20218
rect 433568 19898 433610 20134
rect 433846 19898 433888 20134
rect 433568 19876 433888 19898
rect 464288 20454 464608 20476
rect 464288 20218 464330 20454
rect 464566 20218 464608 20454
rect 464288 20134 464608 20218
rect 464288 19898 464330 20134
rect 464566 19898 464608 20134
rect 464288 19876 464608 19898
rect 495008 20454 495328 20476
rect 495008 20218 495050 20454
rect 495286 20218 495328 20454
rect 495008 20134 495328 20218
rect 495008 19898 495050 20134
rect 495286 19898 495328 20134
rect 495008 19876 495328 19898
rect 525728 20454 526048 20476
rect 525728 20218 525770 20454
rect 526006 20218 526048 20454
rect 525728 20134 526048 20218
rect 525728 19898 525770 20134
rect 526006 19898 526048 20134
rect 525728 19876 526048 19898
rect 556448 20454 556768 20476
rect 556448 20218 556490 20454
rect 556726 20218 556768 20454
rect 556448 20134 556768 20218
rect 556448 19898 556490 20134
rect 556726 19898 556768 20134
rect 556448 19876 556768 19898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 414804 -1286 415404 16320
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 432804 2454 433404 16320
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 450804 -1286 451404 16320
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 468804 2454 469404 16320
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 486804 -1286 487404 16320
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 504804 2454 505404 16320
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 522804 -1286 523404 16320
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 540804 2454 541404 16320
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 558804 -1286 559404 16320
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 587200 -2226 587800 706162
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 588140 -3166 588740 707102
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 589080 -4106 589680 708042
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 590020 -5046 590620 708982
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 590960 -5986 591560 709922
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 591900 -6926 592500 710862
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 22054 615772 22290 615858
rect 22054 615708 22140 615772
rect 22140 615708 22204 615772
rect 22204 615708 22290 615772
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 22054 615622 22290 615708
rect 106142 616982 106378 617218
rect 28862 614942 29098 615178
rect 29414 614942 29650 615178
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 107717 524218 107953 524454
rect 107717 523898 107953 524134
rect 192847 524218 193083 524454
rect 192847 523898 193083 524134
rect 65151 506218 65387 506454
rect 65151 505898 65387 506134
rect 150282 506218 150518 506454
rect 150282 505898 150518 506134
rect 235412 506218 235648 506454
rect 235412 505898 235648 506134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 118654 500852 118890 500938
rect 118654 500788 118740 500852
rect 118740 500788 118804 500852
rect 118804 500788 118890 500852
rect 118654 500702 118890 500788
rect 114606 500172 114842 500258
rect 114606 500108 114692 500172
rect 114692 500108 114756 500172
rect 114756 500108 114842 500172
rect 114606 500022 114842 500108
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 23726 470218 23962 470454
rect 23726 469898 23962 470134
rect 54446 470218 54682 470454
rect 54446 469898 54682 470134
rect 85166 470218 85402 470454
rect 85166 469898 85402 470134
rect 115886 470218 116122 470454
rect 115886 469898 116122 470134
rect 146606 470218 146842 470454
rect 146606 469898 146842 470134
rect 39086 452218 39322 452454
rect 39086 451898 39322 452134
rect 69806 452218 70042 452454
rect 69806 451898 70042 452134
rect 100526 452218 100762 452454
rect 100526 451898 100762 452134
rect 131246 452218 131482 452454
rect 131246 451898 131482 452134
rect 23726 434218 23962 434454
rect 23726 433898 23962 434134
rect 54446 434218 54682 434454
rect 54446 433898 54682 434134
rect 85166 434218 85402 434454
rect 85166 433898 85402 434134
rect 115886 434218 116122 434454
rect 115886 433898 116122 434134
rect 146606 434218 146842 434454
rect 146606 433898 146842 434134
rect 39086 416218 39322 416454
rect 39086 415898 39322 416134
rect 69806 416218 70042 416454
rect 69806 415898 70042 416134
rect 100526 416218 100762 416454
rect 100526 415898 100762 416134
rect 131246 416218 131482 416454
rect 131246 415898 131482 416134
rect 129510 401422 129746 401658
rect 122518 400742 122754 400978
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 38917 380218 39153 380454
rect 38917 379898 39153 380134
rect 56847 380218 57083 380454
rect 56847 379898 57083 380134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 29951 362218 30187 362454
rect 29951 361898 30187 362134
rect 47882 362218 48118 362454
rect 47882 361898 48118 362134
rect 65812 362218 66048 362454
rect 65812 361898 66048 362134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 150118 500022 150354 500258
rect 151774 500702 152010 500938
rect 152694 401422 152930 401658
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 157110 421292 157346 421378
rect 157110 421228 157196 421292
rect 157196 421228 157260 421292
rect 157260 421228 157346 421292
rect 157110 421142 157346 421228
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 153798 400742 154034 400978
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 207656 488218 207892 488454
rect 207656 487898 207892 488134
rect 238376 488218 238612 488454
rect 238376 487898 238612 488134
rect 269096 488218 269332 488454
rect 269096 487898 269332 488134
rect 192296 470218 192532 470454
rect 192296 469898 192532 470134
rect 223016 470218 223252 470454
rect 223016 469898 223252 470134
rect 253736 470218 253972 470454
rect 253736 469898 253972 470134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 207656 452218 207892 452454
rect 207656 451898 207892 452134
rect 238376 452218 238612 452454
rect 238376 451898 238612 452134
rect 269096 452218 269332 452454
rect 269096 451898 269332 452134
rect 192296 434218 192532 434454
rect 192296 433898 192532 434134
rect 223016 434218 223252 434454
rect 223016 433898 223252 434134
rect 253736 434218 253972 434454
rect 253736 433898 253972 434134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 281494 421292 281730 421378
rect 281494 421228 281580 421292
rect 281580 421228 281644 421292
rect 281644 421228 281730 421292
rect 281494 421142 281730 421228
rect 207656 416218 207892 416454
rect 207656 415898 207892 416134
rect 238376 416218 238612 416454
rect 238376 415898 238612 416134
rect 269096 416218 269332 416454
rect 269096 415898 269332 416134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 107717 344218 107953 344454
rect 107717 343898 107953 344134
rect 192847 344218 193083 344454
rect 192847 343898 193083 344134
rect 65151 326218 65387 326454
rect 65151 325898 65387 326134
rect 150282 326218 150518 326454
rect 150282 325898 150518 326134
rect 235412 326218 235648 326454
rect 235412 325898 235648 326134
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 323772 650218 324008 650454
rect 323772 649898 324008 650134
rect 354492 650218 354728 650454
rect 354492 649898 354728 650134
rect 385212 650218 385448 650454
rect 385212 649898 385448 650134
rect 415932 650218 416168 650454
rect 415932 649898 416168 650134
rect 446652 650218 446888 650454
rect 446652 649898 446888 650134
rect 464250 650218 464486 650454
rect 464250 649898 464486 650134
rect 339132 632218 339368 632454
rect 339132 631898 339368 632134
rect 369852 632218 370088 632454
rect 369852 631898 370088 632134
rect 400572 632218 400808 632454
rect 400572 631898 400808 632134
rect 431292 632218 431528 632454
rect 431292 631898 431528 632134
rect 479610 632218 479846 632454
rect 479610 631898 479846 632134
rect 323772 614218 324008 614454
rect 323772 613898 324008 614134
rect 354492 614218 354728 614454
rect 354492 613898 354728 614134
rect 385212 614218 385448 614454
rect 385212 613898 385448 614134
rect 415932 614218 416168 614454
rect 415932 613898 416168 614134
rect 446652 614218 446888 614454
rect 446652 613898 446888 614134
rect 464250 614218 464486 614454
rect 464250 613898 464486 614134
rect 339132 596218 339368 596454
rect 339132 595898 339368 596134
rect 369852 596218 370088 596454
rect 369852 595898 370088 596134
rect 400572 596218 400808 596454
rect 400572 595898 400808 596134
rect 431292 596218 431528 596454
rect 431292 595898 431528 596134
rect 479610 596218 479846 596454
rect 479610 595898 479846 596134
rect 323772 578218 324008 578454
rect 323772 577898 324008 578134
rect 354492 578218 354728 578454
rect 354492 577898 354728 578134
rect 385212 578218 385448 578454
rect 385212 577898 385448 578134
rect 415932 578218 416168 578454
rect 415932 577898 416168 578134
rect 446652 578218 446888 578454
rect 446652 577898 446888 578134
rect 464250 578218 464486 578454
rect 464250 577898 464486 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 494970 650218 495206 650454
rect 494970 649898 495206 650134
rect 525690 650218 525926 650454
rect 525690 649898 525926 650134
rect 510330 632218 510566 632454
rect 510330 631898 510566 632134
rect 541050 632218 541286 632454
rect 541050 631898 541286 632134
rect 494970 614218 495206 614454
rect 494970 613898 495206 614134
rect 525690 614218 525926 614454
rect 525690 613898 525926 614134
rect 510330 596218 510566 596454
rect 510330 595898 510566 596134
rect 541050 596218 541286 596454
rect 541050 595898 541286 596134
rect 494970 578218 495206 578454
rect 494970 577898 495206 578134
rect 525690 578218 525926 578454
rect 525690 577898 525926 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 549398 610862 549634 611098
rect 549398 598622 549634 598858
rect 550686 629222 550922 629458
rect 550134 627862 550370 628098
rect 550686 610862 550922 611098
rect 550686 598622 550922 598858
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 403763 524218 403999 524454
rect 403763 523898 403999 524134
rect 488893 524218 489129 524454
rect 488893 523898 489129 524134
rect 361197 506218 361433 506454
rect 361197 505898 361433 506134
rect 446328 506218 446564 506454
rect 446328 505898 446564 506134
rect 531459 506218 531695 506454
rect 531459 505898 531695 506134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 39656 308218 39892 308454
rect 39656 307898 39892 308134
rect 24296 290218 24532 290454
rect 24296 289898 24532 290134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 39656 272218 39892 272454
rect 39656 271898 39892 272134
rect 24296 254218 24532 254454
rect 24296 253898 24532 254134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 70376 308218 70612 308454
rect 70376 307898 70612 308134
rect 101096 308218 101332 308454
rect 101096 307898 101332 308134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 55016 290218 55252 290454
rect 55016 289898 55252 290134
rect 85736 290218 85972 290454
rect 85736 289898 85972 290134
rect 70376 272218 70612 272454
rect 70376 271898 70612 272134
rect 101096 272218 101332 272454
rect 101096 271898 101332 272134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 55016 254218 55252 254454
rect 55016 253898 55252 254134
rect 85736 254218 85972 254454
rect 85736 253898 85972 254134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 181582 253182 181818 253418
rect 192250 290218 192486 290454
rect 192250 289898 192486 290134
rect 192250 254218 192486 254454
rect 192250 253898 192486 254134
rect 207610 308218 207846 308454
rect 207610 307898 207846 308134
rect 207610 272218 207846 272454
rect 207610 271898 207846 272134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 28810 200218 29046 200454
rect 28810 199898 29046 200134
rect 59530 200218 59766 200454
rect 59530 199898 59766 200134
rect 90250 200218 90486 200454
rect 90250 199898 90486 200134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 13450 182218 13686 182454
rect 13450 181898 13686 182134
rect 44170 182218 44406 182454
rect 44170 181898 44406 182134
rect 74890 182218 75126 182454
rect 74890 181898 75126 182134
rect 123850 218218 124086 218454
rect 123850 217898 124086 218134
rect 154570 218218 154806 218454
rect 154570 217898 154806 218134
rect 185290 218218 185526 218454
rect 185290 217898 185526 218134
rect 139210 200218 139446 200454
rect 139210 199898 139446 200134
rect 169930 200218 170166 200454
rect 169930 199898 170166 200134
rect 200650 200218 200886 200454
rect 200650 199898 200886 200134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 28810 164218 29046 164454
rect 28810 163898 29046 164134
rect 59530 164218 59766 164454
rect 59530 163898 59766 164134
rect 90250 164218 90486 164454
rect 90250 163898 90486 164134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 13450 146218 13686 146454
rect 13450 145898 13686 146134
rect 44170 146218 44406 146454
rect 44170 145898 44406 146134
rect 74890 146218 75126 146454
rect 74890 145898 75126 146134
rect 123850 182218 124086 182454
rect 123850 181898 124086 182134
rect 154570 182218 154806 182454
rect 154570 181898 154806 182134
rect 185290 182218 185526 182454
rect 185290 181898 185526 182134
rect 139210 164218 139446 164454
rect 139210 163898 139446 164134
rect 169930 164218 170166 164454
rect 169930 163898 170166 164134
rect 200650 164218 200886 164454
rect 200650 163898 200886 164134
rect 238330 308218 238566 308454
rect 238330 307898 238566 308134
rect 269050 308218 269286 308454
rect 269050 307898 269286 308134
rect 222970 290218 223206 290454
rect 222970 289898 223206 290134
rect 253690 290218 253926 290454
rect 253690 289898 253926 290134
rect 293231 326218 293467 326454
rect 293231 325898 293467 326134
rect 294677 308218 294913 308454
rect 294677 307898 294913 308134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 238330 272218 238566 272454
rect 238330 271898 238566 272134
rect 269050 272218 269286 272454
rect 269050 271898 269286 272134
rect 222970 254218 223206 254454
rect 222970 253898 223206 254134
rect 253690 254218 253926 254454
rect 253690 253898 253926 254134
rect 279286 251822 279522 252058
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 28810 92218 29046 92454
rect 28810 91898 29046 92134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 13450 74218 13686 74454
rect 13450 73898 13686 74134
rect 28810 56218 29046 56454
rect 28810 55898 29046 56134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 13450 38218 13686 38454
rect 13450 37898 13686 38134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 123850 146218 124086 146454
rect 123850 145898 124086 146134
rect 154570 146218 154806 146454
rect 154570 145898 154806 146134
rect 185290 146218 185526 146454
rect 185290 145898 185526 146134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 139210 128218 139446 128454
rect 139210 127898 139446 128134
rect 169930 128218 170166 128454
rect 169930 127898 170166 128134
rect 200650 128218 200886 128454
rect 200650 127898 200886 128134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 59530 92218 59766 92454
rect 59530 91898 59766 92134
rect 90250 92218 90486 92454
rect 90250 91898 90486 92134
rect 44170 74218 44406 74454
rect 44170 73898 44406 74134
rect 74890 74218 75126 74454
rect 74890 73898 75126 74134
rect 123850 110218 124086 110454
rect 123850 109898 124086 110134
rect 154570 110218 154806 110454
rect 154570 109898 154806 110134
rect 185290 110218 185526 110454
rect 185290 109898 185526 110134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 139210 92218 139446 92454
rect 139210 91898 139446 92134
rect 169930 92218 170166 92454
rect 169930 91898 170166 92134
rect 200650 92218 200886 92454
rect 200650 91898 200886 92134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 59530 56218 59766 56454
rect 59530 55898 59766 56134
rect 90250 56218 90486 56454
rect 90250 55898 90486 56134
rect 44170 38218 44406 38454
rect 44170 37898 44406 38134
rect 74890 38218 75126 38454
rect 74890 37898 75126 38134
rect 123850 74218 124086 74454
rect 123850 73898 124086 74134
rect 154570 74218 154806 74454
rect 154570 73898 154806 74134
rect 185290 74218 185526 74454
rect 185290 73898 185526 74134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 139210 56218 139446 56454
rect 139210 55898 139446 56134
rect 169930 56218 170166 56454
rect 169930 55898 170166 56134
rect 200650 56218 200886 56454
rect 200650 55898 200886 56134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 123850 38218 124086 38454
rect 123850 37898 124086 38134
rect 154570 38218 154806 38454
rect 154570 37898 154806 38134
rect 185290 38218 185526 38454
rect 185290 37898 185526 38134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 549766 472822 550002 473058
rect 548294 472142 548530 472378
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 554734 472822 554970 473058
rect 555102 472142 555338 472378
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 433610 56218 433846 56454
rect 433610 55898 433846 56134
rect 464330 56218 464566 56454
rect 464330 55898 464566 56134
rect 495050 56218 495286 56454
rect 495050 55898 495286 56134
rect 525770 56218 526006 56454
rect 525770 55898 526006 56134
rect 556490 56218 556726 56454
rect 556490 55898 556726 56134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 418250 38218 418486 38454
rect 418250 37898 418486 38134
rect 448970 38218 449206 38454
rect 448970 37898 449206 38134
rect 479690 38218 479926 38454
rect 479690 37898 479926 38134
rect 510410 38218 510646 38454
rect 510410 37898 510646 38134
rect 541130 38218 541366 38454
rect 541130 37898 541366 38134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 433610 20218 433846 20454
rect 433610 19898 433846 20134
rect 464330 20218 464566 20454
rect 464330 19898 464566 20134
rect 495050 20218 495286 20454
rect 495050 19898 495286 20134
rect 525770 20218 526006 20454
rect 525770 19898 526006 20134
rect 556490 20218 556726 20454
rect 556490 19898 556726 20134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 323730 650476 324050 650478
rect 354450 650476 354770 650478
rect 385170 650476 385490 650478
rect 415890 650476 416210 650478
rect 446610 650476 446930 650478
rect 464208 650476 464528 650478
rect 494928 650476 495248 650478
rect 525648 650476 525968 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 323772 650454
rect 324008 650218 354492 650454
rect 354728 650218 385212 650454
rect 385448 650218 415932 650454
rect 416168 650218 446652 650454
rect 446888 650218 464250 650454
rect 464486 650218 494970 650454
rect 495206 650218 525690 650454
rect 525926 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 323772 650134
rect 324008 649898 354492 650134
rect 354728 649898 385212 650134
rect 385448 649898 415932 650134
rect 416168 649898 446652 650134
rect 446888 649898 464250 650134
rect 464486 649898 494970 650134
rect 495206 649898 525690 650134
rect 525926 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 323730 649874 324050 649876
rect 354450 649874 354770 649876
rect 385170 649874 385490 649876
rect 415890 649874 416210 649876
rect 446610 649874 446930 649876
rect 464208 649874 464528 649876
rect 494928 649874 495248 649876
rect 525648 649874 525968 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 339090 632476 339410 632478
rect 369810 632476 370130 632478
rect 400530 632476 400850 632478
rect 431250 632476 431570 632478
rect 479568 632476 479888 632478
rect 510288 632476 510608 632478
rect 541008 632476 541328 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 339132 632454
rect 339368 632218 369852 632454
rect 370088 632218 400572 632454
rect 400808 632218 431292 632454
rect 431528 632218 479610 632454
rect 479846 632218 510330 632454
rect 510566 632218 541050 632454
rect 541286 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 339132 632134
rect 339368 631898 369852 632134
rect 370088 631898 400572 632134
rect 400808 631898 431292 632134
rect 431528 631898 479610 632134
rect 479846 631898 510330 632134
rect 510566 631898 541050 632134
rect 541286 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 339090 631874 339410 631876
rect 369810 631874 370130 631876
rect 400530 631874 400850 631876
rect 431250 631874 431570 631876
rect 479568 631874 479888 631876
rect 510288 631874 510608 631876
rect 541008 631874 541328 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect 550092 629458 550964 629500
rect 550092 629222 550686 629458
rect 550922 629222 550964 629458
rect 550092 629180 550964 629222
rect 550092 628098 550412 629180
rect 550092 627862 550134 628098
rect 550370 627862 550412 628098
rect 550092 627820 550412 627862
rect 35812 616940 45516 617260
rect 35812 615900 36132 616940
rect 22012 615858 36132 615900
rect 22012 615622 22054 615858
rect 22290 615622 36132 615858
rect 22012 615580 36132 615622
rect 45196 615900 45516 616940
rect 55132 616940 64836 617260
rect 55132 615900 55452 616940
rect 45196 615580 55452 615900
rect 64516 615900 64836 616940
rect 74452 616940 84156 617260
rect 74452 615900 74772 616940
rect 64516 615580 74772 615900
rect 83836 615900 84156 616940
rect 86780 617218 106420 617260
rect 86780 616982 106142 617218
rect 106378 616982 106420 617218
rect 86780 616940 106420 616982
rect 86780 615900 87100 616940
rect 83836 615580 87100 615900
rect 28820 615178 29692 615220
rect 28820 614942 28862 615178
rect 29098 614942 29414 615178
rect 29650 614942 29692 615178
rect 28820 614900 29692 614942
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 288804 614476 289404 614478
rect 323730 614476 324050 614478
rect 354450 614476 354770 614478
rect 385170 614476 385490 614478
rect 415890 614476 416210 614478
rect 446610 614476 446930 614478
rect 464208 614476 464528 614478
rect 494928 614476 495248 614478
rect 525648 614476 525968 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 288986 614454
rect 289222 614218 323772 614454
rect 324008 614218 354492 614454
rect 354728 614218 385212 614454
rect 385448 614218 415932 614454
rect 416168 614218 446652 614454
rect 446888 614218 464250 614454
rect 464486 614218 494970 614454
rect 495206 614218 525690 614454
rect 525926 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 288986 614134
rect 289222 613898 323772 614134
rect 324008 613898 354492 614134
rect 354728 613898 385212 614134
rect 385448 613898 415932 614134
rect 416168 613898 446652 614134
rect 446888 613898 464250 614134
rect 464486 613898 494970 614134
rect 495206 613898 525690 614134
rect 525926 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 288804 613874 289404 613876
rect 323730 613874 324050 613876
rect 354450 613874 354770 613876
rect 385170 613874 385490 613876
rect 415890 613874 416210 613876
rect 446610 613874 446930 613876
rect 464208 613874 464528 613876
rect 494928 613874 495248 613876
rect 525648 613874 525968 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect 549356 611098 550964 611140
rect 549356 610862 549398 611098
rect 549634 610862 550686 611098
rect 550922 610862 550964 611098
rect 549356 610820 550964 610862
rect 549356 598858 550964 598900
rect 549356 598622 549398 598858
rect 549634 598622 550686 598858
rect 550922 598622 550964 598858
rect 549356 598580 550964 598622
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 162804 596476 163404 596478
rect 306804 596476 307404 596478
rect 339090 596476 339410 596478
rect 369810 596476 370130 596478
rect 400530 596476 400850 596478
rect 431250 596476 431570 596478
rect 479568 596476 479888 596478
rect 510288 596476 510608 596478
rect 541008 596476 541328 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 162986 596454
rect 163222 596218 306986 596454
rect 307222 596218 339132 596454
rect 339368 596218 369852 596454
rect 370088 596218 400572 596454
rect 400808 596218 431292 596454
rect 431528 596218 479610 596454
rect 479846 596218 510330 596454
rect 510566 596218 541050 596454
rect 541286 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 162986 596134
rect 163222 595898 306986 596134
rect 307222 595898 339132 596134
rect 339368 595898 369852 596134
rect 370088 595898 400572 596134
rect 400808 595898 431292 596134
rect 431528 595898 479610 596134
rect 479846 595898 510330 596134
rect 510566 595898 541050 596134
rect 541286 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 162804 595874 163404 595876
rect 306804 595874 307404 595876
rect 339090 595874 339410 595876
rect 369810 595874 370130 595876
rect 400530 595874 400850 595876
rect 431250 595874 431570 595876
rect 479568 595874 479888 595876
rect 510288 595874 510608 595876
rect 541008 595874 541328 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 288804 578476 289404 578478
rect 323730 578476 324050 578478
rect 354450 578476 354770 578478
rect 385170 578476 385490 578478
rect 415890 578476 416210 578478
rect 446610 578476 446930 578478
rect 464208 578476 464528 578478
rect 494928 578476 495248 578478
rect 525648 578476 525968 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 288986 578454
rect 289222 578218 323772 578454
rect 324008 578218 354492 578454
rect 354728 578218 385212 578454
rect 385448 578218 415932 578454
rect 416168 578218 446652 578454
rect 446888 578218 464250 578454
rect 464486 578218 494970 578454
rect 495206 578218 525690 578454
rect 525926 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 288986 578134
rect 289222 577898 323772 578134
rect 324008 577898 354492 578134
rect 354728 577898 385212 578134
rect 385448 577898 415932 578134
rect 416168 577898 446652 578134
rect 446888 577898 464250 578134
rect 464486 577898 494970 578134
rect 495206 577898 525690 578134
rect 525926 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 288804 577874 289404 577876
rect 323730 577874 324050 577876
rect 354450 577874 354770 577876
rect 385170 577874 385490 577876
rect 415890 577874 416210 577876
rect 446610 577874 446930 577876
rect 464208 577874 464528 577876
rect 494928 577874 495248 577876
rect 525648 577874 525968 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586260 559874 586860 559876
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 107675 524476 107995 524478
rect 192805 524476 193125 524478
rect 306804 524476 307404 524478
rect 403721 524476 404041 524478
rect 488851 524476 489171 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 107717 524454
rect 107953 524218 192847 524454
rect 193083 524218 306986 524454
rect 307222 524218 403763 524454
rect 403999 524218 488893 524454
rect 489129 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 107717 524134
rect 107953 523898 192847 524134
rect 193083 523898 306986 524134
rect 307222 523898 403763 524134
rect 403999 523898 488893 524134
rect 489129 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 107675 523874 107995 523876
rect 192805 523874 193125 523876
rect 306804 523874 307404 523876
rect 403721 523874 404041 523876
rect 488851 523874 489171 523876
rect 586260 523874 586860 523876
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 65109 506476 65429 506478
rect 150240 506476 150560 506478
rect 235370 506476 235690 506478
rect 288804 506476 289404 506478
rect 361155 506476 361475 506478
rect 446286 506476 446606 506478
rect 531417 506476 531737 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 65151 506454
rect 65387 506218 150282 506454
rect 150518 506218 235412 506454
rect 235648 506218 288986 506454
rect 289222 506218 361197 506454
rect 361433 506218 446328 506454
rect 446564 506218 531459 506454
rect 531695 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 65151 506134
rect 65387 505898 150282 506134
rect 150518 505898 235412 506134
rect 235648 505898 288986 506134
rect 289222 505898 361197 506134
rect 361433 505898 446328 506134
rect 446564 505898 531459 506134
rect 531695 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 65109 505874 65429 505876
rect 150240 505874 150560 505876
rect 235370 505874 235690 505876
rect 288804 505874 289404 505876
rect 361155 505874 361475 505876
rect 446286 505874 446606 505876
rect 531417 505874 531737 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect 118612 500938 152052 500980
rect 118612 500702 118654 500938
rect 118890 500702 151774 500938
rect 152010 500702 152052 500938
rect 118612 500660 152052 500702
rect 114564 500258 150396 500300
rect 114564 500022 114606 500258
rect 114842 500022 150118 500258
rect 150354 500022 150396 500258
rect 114564 499980 150396 500022
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 207614 488476 207934 488478
rect 238334 488476 238654 488478
rect 269054 488476 269374 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 207656 488454
rect 207892 488218 238376 488454
rect 238612 488218 269096 488454
rect 269332 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 207656 488134
rect 207892 487898 238376 488134
rect 238612 487898 269096 488134
rect 269332 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 207614 487874 207934 487876
rect 238334 487874 238654 487876
rect 269054 487874 269374 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586260 487874 586860 487876
rect 549724 473058 555012 473100
rect 549724 472822 549766 473058
rect 550002 472822 554734 473058
rect 554970 472822 555012 473058
rect 549724 472780 555012 472822
rect 548252 472378 555380 472420
rect 548252 472142 548294 472378
rect 548530 472142 555102 472378
rect 555338 472142 555380 472378
rect 548252 472100 555380 472142
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 23684 470476 24004 470478
rect 54404 470476 54724 470478
rect 85124 470476 85444 470478
rect 115844 470476 116164 470478
rect 146564 470476 146884 470478
rect 180804 470476 181404 470478
rect 192254 470476 192574 470478
rect 222974 470476 223294 470478
rect 253694 470476 254014 470478
rect 288804 470476 289404 470478
rect 432804 470476 433404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 23726 470454
rect 23962 470218 54446 470454
rect 54682 470218 85166 470454
rect 85402 470218 115886 470454
rect 116122 470218 146606 470454
rect 146842 470218 180986 470454
rect 181222 470218 192296 470454
rect 192532 470218 223016 470454
rect 223252 470218 253736 470454
rect 253972 470218 288986 470454
rect 289222 470218 432986 470454
rect 433222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 23726 470134
rect 23962 469898 54446 470134
rect 54682 469898 85166 470134
rect 85402 469898 115886 470134
rect 116122 469898 146606 470134
rect 146842 469898 180986 470134
rect 181222 469898 192296 470134
rect 192532 469898 223016 470134
rect 223252 469898 253736 470134
rect 253972 469898 288986 470134
rect 289222 469898 432986 470134
rect 433222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 23684 469874 24004 469876
rect 54404 469874 54724 469876
rect 85124 469874 85444 469876
rect 115844 469874 116164 469876
rect 146564 469874 146884 469876
rect 180804 469874 181404 469876
rect 192254 469874 192574 469876
rect 222974 469874 223294 469876
rect 253694 469874 254014 469876
rect 288804 469874 289404 469876
rect 432804 469874 433404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -2936 452476 -2336 452478
rect 39044 452476 39364 452478
rect 69764 452476 70084 452478
rect 100484 452476 100804 452478
rect 131204 452476 131524 452478
rect 162804 452476 163404 452478
rect 207614 452476 207934 452478
rect 238334 452476 238654 452478
rect 269054 452476 269374 452478
rect 306804 452476 307404 452478
rect 414804 452476 415404 452478
rect 558804 452476 559404 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 39086 452454
rect 39322 452218 69806 452454
rect 70042 452218 100526 452454
rect 100762 452218 131246 452454
rect 131482 452218 162986 452454
rect 163222 452218 207656 452454
rect 207892 452218 238376 452454
rect 238612 452218 269096 452454
rect 269332 452218 306986 452454
rect 307222 452218 414986 452454
rect 415222 452218 558986 452454
rect 559222 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 39086 452134
rect 39322 451898 69806 452134
rect 70042 451898 100526 452134
rect 100762 451898 131246 452134
rect 131482 451898 162986 452134
rect 163222 451898 207656 452134
rect 207892 451898 238376 452134
rect 238612 451898 269096 452134
rect 269332 451898 306986 452134
rect 307222 451898 414986 452134
rect 415222 451898 558986 452134
rect 559222 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 39044 451874 39364 451876
rect 69764 451874 70084 451876
rect 100484 451874 100804 451876
rect 131204 451874 131524 451876
rect 162804 451874 163404 451876
rect 207614 451874 207934 451876
rect 238334 451874 238654 451876
rect 269054 451874 269374 451876
rect 306804 451874 307404 451876
rect 414804 451874 415404 451876
rect 558804 451874 559404 451876
rect 586260 451874 586860 451876
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 23684 434476 24004 434478
rect 54404 434476 54724 434478
rect 85124 434476 85444 434478
rect 115844 434476 116164 434478
rect 146564 434476 146884 434478
rect 180804 434476 181404 434478
rect 192254 434476 192574 434478
rect 222974 434476 223294 434478
rect 253694 434476 254014 434478
rect 288804 434476 289404 434478
rect 432804 434476 433404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 23726 434454
rect 23962 434218 54446 434454
rect 54682 434218 85166 434454
rect 85402 434218 115886 434454
rect 116122 434218 146606 434454
rect 146842 434218 180986 434454
rect 181222 434218 192296 434454
rect 192532 434218 223016 434454
rect 223252 434218 253736 434454
rect 253972 434218 288986 434454
rect 289222 434218 432986 434454
rect 433222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 23726 434134
rect 23962 433898 54446 434134
rect 54682 433898 85166 434134
rect 85402 433898 115886 434134
rect 116122 433898 146606 434134
rect 146842 433898 180986 434134
rect 181222 433898 192296 434134
rect 192532 433898 223016 434134
rect 223252 433898 253736 434134
rect 253972 433898 288986 434134
rect 289222 433898 432986 434134
rect 433222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 23684 433874 24004 433876
rect 54404 433874 54724 433876
rect 85124 433874 85444 433876
rect 115844 433874 116164 433876
rect 146564 433874 146884 433876
rect 180804 433874 181404 433876
rect 192254 433874 192574 433876
rect 222974 433874 223294 433876
rect 253694 433874 254014 433876
rect 288804 433874 289404 433876
rect 432804 433874 433404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect 157068 421378 281772 421420
rect 157068 421142 157110 421378
rect 157346 421142 281494 421378
rect 281730 421142 281772 421378
rect 157068 421100 281772 421142
rect -2936 416476 -2336 416478
rect 39044 416476 39364 416478
rect 69764 416476 70084 416478
rect 100484 416476 100804 416478
rect 131204 416476 131524 416478
rect 162804 416476 163404 416478
rect 207614 416476 207934 416478
rect 238334 416476 238654 416478
rect 269054 416476 269374 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 39086 416454
rect 39322 416218 69806 416454
rect 70042 416218 100526 416454
rect 100762 416218 131246 416454
rect 131482 416218 162986 416454
rect 163222 416218 207656 416454
rect 207892 416218 238376 416454
rect 238612 416218 269096 416454
rect 269332 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 39086 416134
rect 39322 415898 69806 416134
rect 70042 415898 100526 416134
rect 100762 415898 131246 416134
rect 131482 415898 162986 416134
rect 163222 415898 207656 416134
rect 207892 415898 238376 416134
rect 238612 415898 269096 416134
rect 269332 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 39044 415874 39364 415876
rect 69764 415874 70084 415876
rect 100484 415874 100804 415876
rect 131204 415874 131524 415876
rect 162804 415874 163404 415876
rect 207614 415874 207934 415876
rect 238334 415874 238654 415876
rect 269054 415874 269374 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586260 415874 586860 415876
rect 129468 401658 152972 401700
rect 129468 401422 129510 401658
rect 129746 401422 152694 401658
rect 152930 401422 152972 401658
rect 129468 401380 152972 401422
rect 122476 400978 154076 401020
rect 122476 400742 122518 400978
rect 122754 400742 153798 400978
rect 154034 400742 154076 400978
rect 122476 400700 154076 400742
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 38875 380476 39195 380478
rect 56805 380476 57125 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 38917 380454
rect 39153 380218 56847 380454
rect 57083 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 38917 380134
rect 39153 379898 56847 380134
rect 57083 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 38875 379874 39195 379876
rect 56805 379874 57125 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 29909 362476 30229 362478
rect 47840 362476 48160 362478
rect 65770 362476 66090 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 29951 362454
rect 30187 362218 47882 362454
rect 48118 362218 65812 362454
rect 66048 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 29951 362134
rect 30187 361898 47882 362134
rect 48118 361898 65812 362134
rect 66048 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 29909 361874 30229 361876
rect 47840 361874 48160 361876
rect 65770 361874 66090 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 107675 344476 107995 344478
rect 192805 344476 193125 344478
rect 306804 344476 307404 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 107717 344454
rect 107953 344218 192847 344454
rect 193083 344218 306986 344454
rect 307222 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 107717 344134
rect 107953 343898 192847 344134
rect 193083 343898 306986 344134
rect 307222 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 107675 343874 107995 343876
rect 192805 343874 193125 343876
rect 306804 343874 307404 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 65109 326476 65429 326478
rect 150240 326476 150560 326478
rect 235370 326476 235690 326478
rect 288804 326476 289404 326478
rect 293189 326476 293509 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 65151 326454
rect 65387 326218 150282 326454
rect 150518 326218 235412 326454
rect 235648 326218 288986 326454
rect 289222 326218 293231 326454
rect 293467 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 65151 326134
rect 65387 325898 150282 326134
rect 150518 325898 235412 326134
rect 235648 325898 288986 326134
rect 289222 325898 293231 326134
rect 293467 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 65109 325874 65429 325876
rect 150240 325874 150560 325876
rect 235370 325874 235690 325876
rect 288804 325874 289404 325876
rect 293189 325874 293509 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 39614 308476 39934 308478
rect 70334 308476 70654 308478
rect 101054 308476 101374 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 207568 308476 207888 308478
rect 238288 308476 238608 308478
rect 269008 308476 269328 308478
rect 294635 308476 294955 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 39656 308454
rect 39892 308218 70376 308454
rect 70612 308218 101096 308454
rect 101332 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 207610 308454
rect 207846 308218 238330 308454
rect 238566 308218 269050 308454
rect 269286 308218 294677 308454
rect 294913 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 39656 308134
rect 39892 307898 70376 308134
rect 70612 307898 101096 308134
rect 101332 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 207610 308134
rect 207846 307898 238330 308134
rect 238566 307898 269050 308134
rect 269286 307898 294677 308134
rect 294913 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 39614 307874 39934 307876
rect 70334 307874 70654 307876
rect 101054 307874 101374 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 207568 307874 207888 307876
rect 238288 307874 238608 307876
rect 269008 307874 269328 307876
rect 294635 307874 294955 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 24254 290476 24574 290478
rect 54974 290476 55294 290478
rect 85694 290476 86014 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 192208 290476 192528 290478
rect 222928 290476 223248 290478
rect 253648 290476 253968 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 24296 290454
rect 24532 290218 55016 290454
rect 55252 290218 85736 290454
rect 85972 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 192250 290454
rect 192486 290218 222970 290454
rect 223206 290218 253690 290454
rect 253926 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 24296 290134
rect 24532 289898 55016 290134
rect 55252 289898 85736 290134
rect 85972 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 192250 290134
rect 192486 289898 222970 290134
rect 223206 289898 253690 290134
rect 253926 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 24254 289874 24574 289876
rect 54974 289874 55294 289876
rect 85694 289874 86014 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 192208 289874 192528 289876
rect 222928 289874 223248 289876
rect 253648 289874 253968 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 39614 272476 39934 272478
rect 70334 272476 70654 272478
rect 101054 272476 101374 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 207568 272476 207888 272478
rect 238288 272476 238608 272478
rect 269008 272476 269328 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 39656 272454
rect 39892 272218 70376 272454
rect 70612 272218 101096 272454
rect 101332 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 207610 272454
rect 207846 272218 238330 272454
rect 238566 272218 269050 272454
rect 269286 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 39656 272134
rect 39892 271898 70376 272134
rect 70612 271898 101096 272134
rect 101332 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 207610 272134
rect 207846 271898 238330 272134
rect 238566 271898 269050 272134
rect 269286 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 39614 271874 39934 271876
rect 70334 271874 70654 271876
rect 101054 271874 101374 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 207568 271874 207888 271876
rect 238288 271874 238608 271876
rect 269008 271874 269328 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586260 271874 586860 271876
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 24254 254476 24574 254478
rect 54974 254476 55294 254478
rect 85694 254476 86014 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 192208 254476 192528 254478
rect 222928 254476 223248 254478
rect 253648 254476 253968 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 24296 254454
rect 24532 254218 55016 254454
rect 55252 254218 85736 254454
rect 85972 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 192250 254454
rect 192486 254218 222970 254454
rect 223206 254218 253690 254454
rect 253926 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 24296 254134
rect 24532 253898 55016 254134
rect 55252 253898 85736 254134
rect 85972 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 192250 254134
rect 192486 253898 222970 254134
rect 223206 253898 253690 254134
rect 253926 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 24254 253874 24574 253876
rect 54974 253874 55294 253876
rect 85694 253874 86014 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 192208 253874 192528 253876
rect 222928 253874 223248 253876
rect 253648 253874 253968 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect 181540 253418 248652 253460
rect 181540 253182 181582 253418
rect 181818 253182 248652 253418
rect 181540 253140 248652 253182
rect 248332 252100 248652 253140
rect 257716 253140 267972 253460
rect 257716 252100 258036 253140
rect 248332 251780 258036 252100
rect 267652 252100 267972 253140
rect 267652 252058 279564 252100
rect 267652 251822 279286 252058
rect 279522 251822 279564 252058
rect 267652 251780 279564 251822
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586260 235874 586860 235876
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 108804 218476 109404 218478
rect 123808 218476 124128 218478
rect 154528 218476 154848 218478
rect 185248 218476 185568 218478
rect 216804 218476 217404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 108986 218454
rect 109222 218218 123850 218454
rect 124086 218218 154570 218454
rect 154806 218218 185290 218454
rect 185526 218218 216986 218454
rect 217222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 108986 218134
rect 109222 217898 123850 218134
rect 124086 217898 154570 218134
rect 154806 217898 185290 218134
rect 185526 217898 216986 218134
rect 217222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 108804 217874 109404 217876
rect 123808 217874 124128 217876
rect 154528 217874 154848 217876
rect 185248 217874 185568 217876
rect 216804 217874 217404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -2936 200476 -2336 200478
rect 28768 200476 29088 200478
rect 59488 200476 59808 200478
rect 90208 200476 90528 200478
rect 139168 200476 139488 200478
rect 169888 200476 170208 200478
rect 200608 200476 200928 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 28810 200454
rect 29046 200218 59530 200454
rect 59766 200218 90250 200454
rect 90486 200218 139210 200454
rect 139446 200218 169930 200454
rect 170166 200218 200650 200454
rect 200886 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 28810 200134
rect 29046 199898 59530 200134
rect 59766 199898 90250 200134
rect 90486 199898 139210 200134
rect 139446 199898 169930 200134
rect 170166 199898 200650 200134
rect 200886 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 28768 199874 29088 199876
rect 59488 199874 59808 199876
rect 90208 199874 90528 199876
rect 139168 199874 139488 199876
rect 169888 199874 170208 199876
rect 200608 199874 200928 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586260 199874 586860 199876
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 13408 182476 13728 182478
rect 44128 182476 44448 182478
rect 74848 182476 75168 182478
rect 108804 182476 109404 182478
rect 123808 182476 124128 182478
rect 154528 182476 154848 182478
rect 185248 182476 185568 182478
rect 216804 182476 217404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 13450 182454
rect 13686 182218 44170 182454
rect 44406 182218 74890 182454
rect 75126 182218 108986 182454
rect 109222 182218 123850 182454
rect 124086 182218 154570 182454
rect 154806 182218 185290 182454
rect 185526 182218 216986 182454
rect 217222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 13450 182134
rect 13686 181898 44170 182134
rect 44406 181898 74890 182134
rect 75126 181898 108986 182134
rect 109222 181898 123850 182134
rect 124086 181898 154570 182134
rect 154806 181898 185290 182134
rect 185526 181898 216986 182134
rect 217222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 13408 181874 13728 181876
rect 44128 181874 44448 181876
rect 74848 181874 75168 181876
rect 108804 181874 109404 181876
rect 123808 181874 124128 181876
rect 154528 181874 154848 181876
rect 185248 181874 185568 181876
rect 216804 181874 217404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -2936 164476 -2336 164478
rect 28768 164476 29088 164478
rect 59488 164476 59808 164478
rect 90208 164476 90528 164478
rect 139168 164476 139488 164478
rect 169888 164476 170208 164478
rect 200608 164476 200928 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 28810 164454
rect 29046 164218 59530 164454
rect 59766 164218 90250 164454
rect 90486 164218 139210 164454
rect 139446 164218 169930 164454
rect 170166 164218 200650 164454
rect 200886 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 28810 164134
rect 29046 163898 59530 164134
rect 59766 163898 90250 164134
rect 90486 163898 139210 164134
rect 139446 163898 169930 164134
rect 170166 163898 200650 164134
rect 200886 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 28768 163874 29088 163876
rect 59488 163874 59808 163876
rect 90208 163874 90528 163876
rect 139168 163874 139488 163876
rect 169888 163874 170208 163876
rect 200608 163874 200928 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586260 163874 586860 163876
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 13408 146476 13728 146478
rect 44128 146476 44448 146478
rect 74848 146476 75168 146478
rect 108804 146476 109404 146478
rect 123808 146476 124128 146478
rect 154528 146476 154848 146478
rect 185248 146476 185568 146478
rect 216804 146476 217404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 13450 146454
rect 13686 146218 44170 146454
rect 44406 146218 74890 146454
rect 75126 146218 108986 146454
rect 109222 146218 123850 146454
rect 124086 146218 154570 146454
rect 154806 146218 185290 146454
rect 185526 146218 216986 146454
rect 217222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 13450 146134
rect 13686 145898 44170 146134
rect 44406 145898 74890 146134
rect 75126 145898 108986 146134
rect 109222 145898 123850 146134
rect 124086 145898 154570 146134
rect 154806 145898 185290 146134
rect 185526 145898 216986 146134
rect 217222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 13408 145874 13728 145876
rect 44128 145874 44448 145876
rect 74848 145874 75168 145876
rect 108804 145874 109404 145876
rect 123808 145874 124128 145876
rect 154528 145874 154848 145876
rect 185248 145874 185568 145876
rect 216804 145874 217404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -2936 128476 -2336 128478
rect 139168 128476 139488 128478
rect 169888 128476 170208 128478
rect 200608 128476 200928 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 139210 128454
rect 139446 128218 169930 128454
rect 170166 128218 200650 128454
rect 200886 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 139210 128134
rect 139446 127898 169930 128134
rect 170166 127898 200650 128134
rect 200886 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 139168 127874 139488 127876
rect 169888 127874 170208 127876
rect 200608 127874 200928 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586260 127874 586860 127876
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 123808 110476 124128 110478
rect 154528 110476 154848 110478
rect 185248 110476 185568 110478
rect 216804 110476 217404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 123850 110454
rect 124086 110218 154570 110454
rect 154806 110218 185290 110454
rect 185526 110218 216986 110454
rect 217222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 123850 110134
rect 124086 109898 154570 110134
rect 154806 109898 185290 110134
rect 185526 109898 216986 110134
rect 217222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 123808 109874 124128 109876
rect 154528 109874 154848 109876
rect 185248 109874 185568 109876
rect 216804 109874 217404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -2936 92476 -2336 92478
rect 28768 92476 29088 92478
rect 59488 92476 59808 92478
rect 90208 92476 90528 92478
rect 139168 92476 139488 92478
rect 169888 92476 170208 92478
rect 200608 92476 200928 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 28810 92454
rect 29046 92218 59530 92454
rect 59766 92218 90250 92454
rect 90486 92218 139210 92454
rect 139446 92218 169930 92454
rect 170166 92218 200650 92454
rect 200886 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 28810 92134
rect 29046 91898 59530 92134
rect 59766 91898 90250 92134
rect 90486 91898 139210 92134
rect 139446 91898 169930 92134
rect 170166 91898 200650 92134
rect 200886 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 28768 91874 29088 91876
rect 59488 91874 59808 91876
rect 90208 91874 90528 91876
rect 139168 91874 139488 91876
rect 169888 91874 170208 91876
rect 200608 91874 200928 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586260 91874 586860 91876
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 13408 74476 13728 74478
rect 44128 74476 44448 74478
rect 74848 74476 75168 74478
rect 108804 74476 109404 74478
rect 123808 74476 124128 74478
rect 154528 74476 154848 74478
rect 185248 74476 185568 74478
rect 216804 74476 217404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 13450 74454
rect 13686 74218 44170 74454
rect 44406 74218 74890 74454
rect 75126 74218 108986 74454
rect 109222 74218 123850 74454
rect 124086 74218 154570 74454
rect 154806 74218 185290 74454
rect 185526 74218 216986 74454
rect 217222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 13450 74134
rect 13686 73898 44170 74134
rect 44406 73898 74890 74134
rect 75126 73898 108986 74134
rect 109222 73898 123850 74134
rect 124086 73898 154570 74134
rect 154806 73898 185290 74134
rect 185526 73898 216986 74134
rect 217222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 13408 73874 13728 73876
rect 44128 73874 44448 73876
rect 74848 73874 75168 73876
rect 108804 73874 109404 73876
rect 123808 73874 124128 73876
rect 154528 73874 154848 73876
rect 185248 73874 185568 73876
rect 216804 73874 217404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -2936 56476 -2336 56478
rect 28768 56476 29088 56478
rect 59488 56476 59808 56478
rect 90208 56476 90528 56478
rect 139168 56476 139488 56478
rect 169888 56476 170208 56478
rect 200608 56476 200928 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 433568 56476 433888 56478
rect 464288 56476 464608 56478
rect 495008 56476 495328 56478
rect 525728 56476 526048 56478
rect 556448 56476 556768 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 28810 56454
rect 29046 56218 59530 56454
rect 59766 56218 90250 56454
rect 90486 56218 139210 56454
rect 139446 56218 169930 56454
rect 170166 56218 200650 56454
rect 200886 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 433610 56454
rect 433846 56218 464330 56454
rect 464566 56218 495050 56454
rect 495286 56218 525770 56454
rect 526006 56218 556490 56454
rect 556726 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 28810 56134
rect 29046 55898 59530 56134
rect 59766 55898 90250 56134
rect 90486 55898 139210 56134
rect 139446 55898 169930 56134
rect 170166 55898 200650 56134
rect 200886 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 433610 56134
rect 433846 55898 464330 56134
rect 464566 55898 495050 56134
rect 495286 55898 525770 56134
rect 526006 55898 556490 56134
rect 556726 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 28768 55874 29088 55876
rect 59488 55874 59808 55876
rect 90208 55874 90528 55876
rect 139168 55874 139488 55876
rect 169888 55874 170208 55876
rect 200608 55874 200928 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 433568 55874 433888 55876
rect 464288 55874 464608 55876
rect 495008 55874 495328 55876
rect 525728 55874 526048 55876
rect 556448 55874 556768 55876
rect 586260 55874 586860 55876
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 13408 38476 13728 38478
rect 44128 38476 44448 38478
rect 74848 38476 75168 38478
rect 108804 38476 109404 38478
rect 123808 38476 124128 38478
rect 154528 38476 154848 38478
rect 185248 38476 185568 38478
rect 216804 38476 217404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 418208 38476 418528 38478
rect 448928 38476 449248 38478
rect 479648 38476 479968 38478
rect 510368 38476 510688 38478
rect 541088 38476 541408 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 13450 38454
rect 13686 38218 44170 38454
rect 44406 38218 74890 38454
rect 75126 38218 108986 38454
rect 109222 38218 123850 38454
rect 124086 38218 154570 38454
rect 154806 38218 185290 38454
rect 185526 38218 216986 38454
rect 217222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 418250 38454
rect 418486 38218 448970 38454
rect 449206 38218 479690 38454
rect 479926 38218 510410 38454
rect 510646 38218 541130 38454
rect 541366 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 13450 38134
rect 13686 37898 44170 38134
rect 44406 37898 74890 38134
rect 75126 37898 108986 38134
rect 109222 37898 123850 38134
rect 124086 37898 154570 38134
rect 154806 37898 185290 38134
rect 185526 37898 216986 38134
rect 217222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 418250 38134
rect 418486 37898 448970 38134
rect 449206 37898 479690 38134
rect 479926 37898 510410 38134
rect 510646 37898 541130 38134
rect 541366 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 13408 37874 13728 37876
rect 44128 37874 44448 37876
rect 74848 37874 75168 37876
rect 108804 37874 109404 37876
rect 123808 37874 124128 37876
rect 154528 37874 154848 37876
rect 185248 37874 185568 37876
rect 216804 37874 217404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 418208 37874 418528 37876
rect 448928 37874 449248 37876
rect 479648 37874 479968 37876
rect 510368 37874 510688 37876
rect 541088 37874 541408 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 433568 20476 433888 20478
rect 464288 20476 464608 20478
rect 495008 20476 495328 20478
rect 525728 20476 526048 20478
rect 556448 20476 556768 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 433610 20454
rect 433846 20218 464330 20454
rect 464566 20218 495050 20454
rect 495286 20218 525770 20454
rect 526006 20218 556490 20454
rect 556726 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 433610 20134
rect 433846 19898 464330 20134
rect 464566 19898 495050 20134
rect 495286 19898 525770 20134
rect 526006 19898 556490 20134
rect 556726 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 433568 19874 433888 19876
rect 464288 19874 464608 19876
rect 495008 19874 495328 19876
rect 525728 19874 526048 19876
rect 556448 19874 556768 19876
rect 586260 19874 586860 19876
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 591900 -7506 592500 -7504
use fd_hd  i_fd0_1
timestamp 1607544406
transform 1 0 230000 0 1 31440
box 0 0 108256 50048
use fd_hs  i_fd0_2
timestamp 1607544406
transform 1 0 230000 0 1 103440
box 0 0 112240 46240
use fd_ms  i_fd0_3
timestamp 1607544406
transform 1 0 230000 0 1 175440
box 0 0 106720 46240
use wb_interface  i_itf0
timestamp 1607544406
transform 1 0 119600 0 1 31440
box 0 0 92000 190400
use tdc_inline_1  i_tdc0_1
timestamp 1607544406
transform 1 0 9200 0 1 31440
box 0 0 82800 68000
use tdc_inline_2  i_tdc0_2
timestamp 1607544406
transform 1 0 9200 0 1 127228
box 0 0 92000 92480
use rescue_top  inst_rescue
timestamp 1607544406
transform 1 0 414000 0 1 16320
box 0 0 147200 44608
use fd_inline_1  i_fd2_2
timestamp 1607544406
transform 1 0 20000 0 -1 384200
box 290 2042 56000 27200
use fd_hd_25_1  i_fd2_3
timestamp 1607544406
transform 1 0 188000 0 -1 402224
box 0 0 94746 44112
use wb_extender  i_itf2
timestamp 1607544406
transform 1 0 21600 0 1 322800
box 474 0 257600 26112
use tdc_inline_3  i_tdc2_0
timestamp 1607544406
transform 1 0 20046 0 1 234000
box 0 2128 92000 81600
use tdc_inline_3  i_tdc2_1
timestamp 1607544406
transform 1 0 188000 0 1 234000
box 0 2128 92000 81600
use zero  b_zero.i_zero
timestamp 1607544406
transform 1 0 290800 0 1 304800
box 0 0 10880 24480
use fd_hs  i_fd3_2
timestamp 1607544406
transform 1 0 28000 0 1 571440
box 0 0 112240 46240
use fd_hd_25_1  i_fd3_3
timestamp 1607544406
transform 1 0 188000 0 -1 618224
box 0 0 94746 44112
use wb_extender  i_itf3
timestamp 1607544406
transform 1 0 21600 0 1 502800
box 474 0 257600 26112
use tdc_hd_cbuf2_x4  i_tdc3_0
timestamp 1607544406
transform 1 0 16000 0 1 400000
box 0 2128 138000 87040
use tdc_inline_3  i_tdc3_1
timestamp 1607544406
transform 1 0 188046 0 1 410000
box 0 2128 92000 81600
use fd_ms  i_fd4_2
timestamp 1607544406
transform -1 0 552720 0 1 427440
box 0 0 106720 46240
use fd_hd_25_1  i_fd4_3
timestamp 1607544406
transform -1 0 410746 0 1 430128
box 0 0 94746 44112
use wb_extender  i_itf4
timestamp 1607544406
transform -1 0 575246 0 -1 528912
box 474 0 257600 26112
use tdc_inline_2  i_tdc4_0
timestamp 1607544406
transform 1 0 460000 0 1 570000
box 0 0 92000 92480
use tdc_hd_cbuf2_x4  i_tdc4_1
timestamp 1607544406
transform 1 0 316046 0 -1 657040
box 0 2128 138000 87040
<< labels >>
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 0 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 1 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 2 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 3 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 4 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 5 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 6 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 7 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 8 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 9 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 10 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 11 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 12 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 13 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 14 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 15 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 16 nsew default tristate
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 17 nsew default input
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 18 nsew default input
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 19 nsew default input
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 20 nsew default input
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 21 nsew default input
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 22 nsew default input
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 23 nsew default input
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 24 nsew default input
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 25 nsew default input
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 26 nsew default input
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 27 nsew default input
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 28 nsew default input
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 29 nsew default input
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 30 nsew default input
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 31 nsew default input
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 32 nsew default input
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 33 nsew default input
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 34 nsew default input
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 35 nsew default input
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 36 nsew default input
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 37 nsew default input
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 38 nsew default input
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 39 nsew default input
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 40 nsew default input
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 41 nsew default input
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 42 nsew default input
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 43 nsew default input
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 44 nsew default input
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 45 nsew default input
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 46 nsew default input
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 47 nsew default input
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 48 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 49 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 50 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 51 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 52 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 53 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 54 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 55 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 56 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 57 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 58 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 59 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 60 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 61 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 62 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 63 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 64 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 65 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 66 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 67 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 68 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 69 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 70 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 71 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 72 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 73 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 74 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 75 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 76 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 77 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 78 nsew default tristate
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 79 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 80 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 81 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 82 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 83 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 84 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 85 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 86 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 87 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 88 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 89 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 90 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 91 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 92 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 93 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 94 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 95 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 96 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 97 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 98 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 99 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 100 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 101 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 102 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 103 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 104 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 105 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 106 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 107 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 108 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 109 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 110 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 111 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 112 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 113 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 114 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 115 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 116 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 117 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 118 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 119 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 120 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 121 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 122 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 123 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 124 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 125 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 126 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 127 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 128 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 129 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 130 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 131 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 132 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 133 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 134 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 135 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 136 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 137 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 138 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 139 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 140 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 141 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 142 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 143 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 638 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 639 nsew default input
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 640 nsew default input
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 641 nsew default input
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 642 nsew default input
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
