VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fd_ms
  CLASS BLOCK ;
  FOREIGN fd_ms ;
  ORIGIN 0.000 0.000 ;
  SIZE 533.600 BY 231.200 ;
  PIN bus_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END bus_in[0]
  PIN bus_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END bus_in[10]
  PIN bus_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END bus_in[11]
  PIN bus_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END bus_in[12]
  PIN bus_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END bus_in[13]
  PIN bus_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END bus_in[14]
  PIN bus_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END bus_in[15]
  PIN bus_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 4.000 96.520 ;
    END
  END bus_in[16]
  PIN bus_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END bus_in[17]
  PIN bus_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END bus_in[18]
  PIN bus_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END bus_in[19]
  PIN bus_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END bus_in[1]
  PIN bus_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END bus_in[20]
  PIN bus_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END bus_in[21]
  PIN bus_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 131.280 4.000 131.880 ;
    END
  END bus_in[22]
  PIN bus_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END bus_in[23]
  PIN bus_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END bus_in[24]
  PIN bus_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END bus_in[25]
  PIN bus_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END bus_in[26]
  PIN bus_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.200 4.000 161.800 ;
    END
  END bus_in[27]
  PIN bus_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END bus_in[28]
  PIN bus_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END bus_in[29]
  PIN bus_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.960 4.000 13.560 ;
    END
  END bus_in[2]
  PIN bus_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END bus_in[30]
  PIN bus_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END bus_in[31]
  PIN bus_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END bus_in[32]
  PIN bus_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END bus_in[33]
  PIN bus_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.680 4.000 203.280 ;
    END
  END bus_in[34]
  PIN bus_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.800 4.000 209.400 ;
    END
  END bus_in[35]
  PIN bus_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 211.520 4.000 212.120 ;
    END
  END bus_in[36]
  PIN bus_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END bus_in[37]
  PIN bus_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END bus_in[38]
  PIN bus_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END bus_in[39]
  PIN bus_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END bus_in[3]
  PIN bus_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END bus_in[40]
  PIN bus_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 226.480 4.000 227.080 ;
    END
  END bus_in[41]
  PIN bus_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END bus_in[4]
  PIN bus_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END bus_in[5]
  PIN bus_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END bus_in[6]
  PIN bus_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END bus_in[7]
  PIN bus_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END bus_in[8]
  PIN bus_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END bus_in[9]
  PIN bus_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END bus_out[0]
  PIN bus_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.280 4.000 63.880 ;
    END
  END bus_out[10]
  PIN bus_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END bus_out[11]
  PIN bus_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END bus_out[12]
  PIN bus_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END bus_out[13]
  PIN bus_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END bus_out[14]
  PIN bus_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END bus_out[15]
  PIN bus_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END bus_out[16]
  PIN bus_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END bus_out[17]
  PIN bus_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 4.000 111.480 ;
    END
  END bus_out[18]
  PIN bus_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END bus_out[19]
  PIN bus_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END bus_out[1]
  PIN bus_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END bus_out[20]
  PIN bus_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.560 4.000 129.160 ;
    END
  END bus_out[21]
  PIN bus_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END bus_out[22]
  PIN bus_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END bus_out[23]
  PIN bus_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END bus_out[24]
  PIN bus_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END bus_out[25]
  PIN bus_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END bus_out[26]
  PIN bus_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END bus_out[27]
  PIN bus_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END bus_out[28]
  PIN bus_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.160 4.000 176.760 ;
    END
  END bus_out[29]
  PIN bus_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END bus_out[2]
  PIN bus_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 181.600 4.000 182.200 ;
    END
  END bus_out[30]
  PIN bus_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.720 4.000 188.320 ;
    END
  END bus_out[31]
  PIN bus_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END bus_out[32]
  PIN bus_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END bus_out[33]
  PIN bus_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END bus_out[34]
  PIN bus_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END bus_out[3]
  PIN bus_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END bus_out[4]
  PIN bus_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END bus_out[5]
  PIN bus_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END bus_out[6]
  PIN bus_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 45.600 4.000 46.200 ;
    END
  END bus_out[7]
  PIN bus_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END bus_out[8]
  PIN bus_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END bus_out[9]
  PIN clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 266.890 0.000 267.170 4.000 ;
    END
  END clk_i
  PIN out1_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END out1_o
  PIN out2_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 529.600 115.640 533.600 116.240 ;
    END
  END out2_o
  PIN rst_n_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 266.890 227.200 267.170 231.200 ;
    END
  END rst_n_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 32.180 528.080 35.180 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 122.180 528.080 125.180 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 528.080 220.405 ;
      LAYER met1 ;
        RECT 5.520 2.080 528.080 220.960 ;
      LAYER met2 ;
        RECT 7.450 226.920 266.610 229.685 ;
        RECT 267.450 226.920 518.130 229.685 ;
        RECT 7.450 4.280 518.130 226.920 ;
        RECT 7.450 1.515 266.610 4.280 ;
        RECT 267.450 1.515 518.130 4.280 ;
      LAYER met3 ;
        RECT 4.400 228.800 529.600 229.665 ;
        RECT 4.000 227.480 529.600 228.800 ;
        RECT 4.400 226.080 529.600 227.480 ;
        RECT 4.000 224.080 529.600 226.080 ;
        RECT 4.400 222.680 529.600 224.080 ;
        RECT 4.000 221.360 529.600 222.680 ;
        RECT 4.400 219.960 529.600 221.360 ;
        RECT 4.000 218.640 529.600 219.960 ;
        RECT 4.400 217.240 529.600 218.640 ;
        RECT 4.000 215.240 529.600 217.240 ;
        RECT 4.400 213.840 529.600 215.240 ;
        RECT 4.000 212.520 529.600 213.840 ;
        RECT 4.400 211.120 529.600 212.520 ;
        RECT 4.000 209.800 529.600 211.120 ;
        RECT 4.400 208.400 529.600 209.800 ;
        RECT 4.000 206.400 529.600 208.400 ;
        RECT 4.400 205.000 529.600 206.400 ;
        RECT 4.000 203.680 529.600 205.000 ;
        RECT 4.400 202.280 529.600 203.680 ;
        RECT 4.000 200.960 529.600 202.280 ;
        RECT 4.400 199.560 529.600 200.960 ;
        RECT 4.000 197.560 529.600 199.560 ;
        RECT 4.400 196.160 529.600 197.560 ;
        RECT 4.000 194.840 529.600 196.160 ;
        RECT 4.400 193.440 529.600 194.840 ;
        RECT 4.000 191.440 529.600 193.440 ;
        RECT 4.400 190.040 529.600 191.440 ;
        RECT 4.000 188.720 529.600 190.040 ;
        RECT 4.400 187.320 529.600 188.720 ;
        RECT 4.000 186.000 529.600 187.320 ;
        RECT 4.400 184.600 529.600 186.000 ;
        RECT 4.000 182.600 529.600 184.600 ;
        RECT 4.400 181.200 529.600 182.600 ;
        RECT 4.000 179.880 529.600 181.200 ;
        RECT 4.400 178.480 529.600 179.880 ;
        RECT 4.000 177.160 529.600 178.480 ;
        RECT 4.400 175.760 529.600 177.160 ;
        RECT 4.000 173.760 529.600 175.760 ;
        RECT 4.400 172.360 529.600 173.760 ;
        RECT 4.000 171.040 529.600 172.360 ;
        RECT 4.400 169.640 529.600 171.040 ;
        RECT 4.000 168.320 529.600 169.640 ;
        RECT 4.400 166.920 529.600 168.320 ;
        RECT 4.000 164.920 529.600 166.920 ;
        RECT 4.400 163.520 529.600 164.920 ;
        RECT 4.000 162.200 529.600 163.520 ;
        RECT 4.400 160.800 529.600 162.200 ;
        RECT 4.000 159.480 529.600 160.800 ;
        RECT 4.400 158.080 529.600 159.480 ;
        RECT 4.000 156.080 529.600 158.080 ;
        RECT 4.400 154.680 529.600 156.080 ;
        RECT 4.000 153.360 529.600 154.680 ;
        RECT 4.400 151.960 529.600 153.360 ;
        RECT 4.000 149.960 529.600 151.960 ;
        RECT 4.400 148.560 529.600 149.960 ;
        RECT 4.000 147.240 529.600 148.560 ;
        RECT 4.400 145.840 529.600 147.240 ;
        RECT 4.000 144.520 529.600 145.840 ;
        RECT 4.400 143.120 529.600 144.520 ;
        RECT 4.000 141.120 529.600 143.120 ;
        RECT 4.400 139.720 529.600 141.120 ;
        RECT 4.000 138.400 529.600 139.720 ;
        RECT 4.400 137.000 529.600 138.400 ;
        RECT 4.000 135.680 529.600 137.000 ;
        RECT 4.400 134.280 529.600 135.680 ;
        RECT 4.000 132.280 529.600 134.280 ;
        RECT 4.400 130.880 529.600 132.280 ;
        RECT 4.000 129.560 529.600 130.880 ;
        RECT 4.400 128.160 529.600 129.560 ;
        RECT 4.000 126.840 529.600 128.160 ;
        RECT 4.400 125.440 529.600 126.840 ;
        RECT 4.000 123.440 529.600 125.440 ;
        RECT 4.400 122.040 529.600 123.440 ;
        RECT 4.000 120.720 529.600 122.040 ;
        RECT 4.400 119.320 529.600 120.720 ;
        RECT 4.000 118.000 529.600 119.320 ;
        RECT 4.400 116.640 529.600 118.000 ;
        RECT 4.400 116.600 529.200 116.640 ;
        RECT 4.000 115.240 529.200 116.600 ;
        RECT 4.000 114.600 529.600 115.240 ;
        RECT 4.400 113.200 529.600 114.600 ;
        RECT 4.000 111.880 529.600 113.200 ;
        RECT 4.400 110.480 529.600 111.880 ;
        RECT 4.000 108.480 529.600 110.480 ;
        RECT 4.400 107.080 529.600 108.480 ;
        RECT 4.000 105.760 529.600 107.080 ;
        RECT 4.400 104.360 529.600 105.760 ;
        RECT 4.000 103.040 529.600 104.360 ;
        RECT 4.400 101.640 529.600 103.040 ;
        RECT 4.000 99.640 529.600 101.640 ;
        RECT 4.400 98.240 529.600 99.640 ;
        RECT 4.000 96.920 529.600 98.240 ;
        RECT 4.400 95.520 529.600 96.920 ;
        RECT 4.000 94.200 529.600 95.520 ;
        RECT 4.400 92.800 529.600 94.200 ;
        RECT 4.000 90.800 529.600 92.800 ;
        RECT 4.400 89.400 529.600 90.800 ;
        RECT 4.000 88.080 529.600 89.400 ;
        RECT 4.400 86.680 529.600 88.080 ;
        RECT 4.000 85.360 529.600 86.680 ;
        RECT 4.400 83.960 529.600 85.360 ;
        RECT 4.000 81.960 529.600 83.960 ;
        RECT 4.400 80.560 529.600 81.960 ;
        RECT 4.000 79.240 529.600 80.560 ;
        RECT 4.400 77.840 529.600 79.240 ;
        RECT 4.000 75.840 529.600 77.840 ;
        RECT 4.400 74.440 529.600 75.840 ;
        RECT 4.000 73.120 529.600 74.440 ;
        RECT 4.400 71.720 529.600 73.120 ;
        RECT 4.000 70.400 529.600 71.720 ;
        RECT 4.400 69.000 529.600 70.400 ;
        RECT 4.000 67.000 529.600 69.000 ;
        RECT 4.400 65.600 529.600 67.000 ;
        RECT 4.000 64.280 529.600 65.600 ;
        RECT 4.400 62.880 529.600 64.280 ;
        RECT 4.000 61.560 529.600 62.880 ;
        RECT 4.400 60.160 529.600 61.560 ;
        RECT 4.000 58.160 529.600 60.160 ;
        RECT 4.400 56.760 529.600 58.160 ;
        RECT 4.000 55.440 529.600 56.760 ;
        RECT 4.400 54.040 529.600 55.440 ;
        RECT 4.000 52.720 529.600 54.040 ;
        RECT 4.400 51.320 529.600 52.720 ;
        RECT 4.000 49.320 529.600 51.320 ;
        RECT 4.400 47.920 529.600 49.320 ;
        RECT 4.000 46.600 529.600 47.920 ;
        RECT 4.400 45.200 529.600 46.600 ;
        RECT 4.000 43.880 529.600 45.200 ;
        RECT 4.400 42.480 529.600 43.880 ;
        RECT 4.000 40.480 529.600 42.480 ;
        RECT 4.400 39.080 529.600 40.480 ;
        RECT 4.000 37.760 529.600 39.080 ;
        RECT 4.400 36.360 529.600 37.760 ;
        RECT 4.000 34.360 529.600 36.360 ;
        RECT 4.400 32.960 529.600 34.360 ;
        RECT 4.000 31.640 529.600 32.960 ;
        RECT 4.400 30.240 529.600 31.640 ;
        RECT 4.000 28.920 529.600 30.240 ;
        RECT 4.400 27.520 529.600 28.920 ;
        RECT 4.000 25.520 529.600 27.520 ;
        RECT 4.400 24.120 529.600 25.520 ;
        RECT 4.000 22.800 529.600 24.120 ;
        RECT 4.400 21.400 529.600 22.800 ;
        RECT 4.000 20.080 529.600 21.400 ;
        RECT 4.400 18.680 529.600 20.080 ;
        RECT 4.000 16.680 529.600 18.680 ;
        RECT 4.400 15.280 529.600 16.680 ;
        RECT 4.000 13.960 529.600 15.280 ;
        RECT 4.400 12.560 529.600 13.960 ;
        RECT 4.000 11.240 529.600 12.560 ;
        RECT 4.400 9.840 529.600 11.240 ;
        RECT 4.000 7.840 529.600 9.840 ;
        RECT 4.400 6.440 529.600 7.840 ;
        RECT 4.000 5.120 529.600 6.440 ;
        RECT 4.400 3.720 529.600 5.120 ;
        RECT 4.000 2.400 529.600 3.720 ;
        RECT 4.400 1.535 529.600 2.400 ;
      LAYER met4 ;
        RECT 21.040 10.640 513.985 220.560 ;
      LAYER met5 ;
        RECT 5.520 126.780 528.080 215.190 ;
        RECT 5.520 36.780 528.080 120.580 ;
  END
END fd_ms
END LIBRARY

