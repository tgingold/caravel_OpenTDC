VERSION 5.7 ;
NOWIREEXTENSIONATPIN ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;
MACRO tdc_inline_2
  CLASS BLOCK ;
  FOREIGN tdc_inline_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 460.000 BY 462.400 ;
  PIN bus_in[0]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 2.760 460.000 3.360 ;
    END
  END bus_in[0]
  PIN bus_in[10]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 123.800 460.000 124.400 ;
    END
  END bus_in[10]
  PIN bus_in[11]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 136.040 460.000 136.640 ;
    END
  END bus_in[11]
  PIN bus_in[12]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 148.280 460.000 148.880 ;
    END
  END bus_in[12]
  PIN bus_in[13]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 160.520 460.000 161.120 ;
    END
  END bus_in[13]
  PIN bus_in[14]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 172.760 460.000 173.360 ;
    END
  END bus_in[14]
  PIN bus_in[15]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 185.000 460.000 185.600 ;
    END
  END bus_in[15]
  PIN bus_in[16]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 197.240 460.000 197.840 ;
    END
  END bus_in[16]
  PIN bus_in[17]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 209.480 460.000 210.080 ;
    END
  END bus_in[17]
  PIN bus_in[18]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 221.720 460.000 222.320 ;
    END
  END bus_in[18]
  PIN bus_in[19]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 233.960 460.000 234.560 ;
    END
  END bus_in[19]
  PIN bus_in[1]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 14.320 460.000 14.920 ;
    END
  END bus_in[1]
  PIN bus_in[20]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 245.520 460.000 246.120 ;
    END
  END bus_in[20]
  PIN bus_in[21]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 257.760 460.000 258.360 ;
    END
  END bus_in[21]
  PIN bus_in[22]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 270.000 460.000 270.600 ;
    END
  END bus_in[22]
  PIN bus_in[23]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 282.240 460.000 282.840 ;
    END
  END bus_in[23]
  PIN bus_in[24]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 294.480 460.000 295.080 ;
    END
  END bus_in[24]
  PIN bus_in[25]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 306.720 460.000 307.320 ;
    END
  END bus_in[25]
  PIN bus_in[26]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 318.960 460.000 319.560 ;
    END
  END bus_in[26]
  PIN bus_in[27]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 331.200 460.000 331.800 ;
    END
  END bus_in[27]
  PIN bus_in[28]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 343.440 460.000 344.040 ;
    END
  END bus_in[28]
  PIN bus_in[29]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 355.000 460.000 355.600 ;
    END
  END bus_in[29]
  PIN bus_in[2]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 26.560 460.000 27.160 ;
    END
  END bus_in[2]
  PIN bus_in[30]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 367.240 460.000 367.840 ;
    END
  END bus_in[30]
  PIN bus_in[31]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 379.480 460.000 380.080 ;
    END
  END bus_in[31]
  PIN bus_in[32]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 391.720 460.000 392.320 ;
    END
  END bus_in[32]
  PIN bus_in[33]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 403.960 460.000 404.560 ;
    END
  END bus_in[33]
  PIN bus_in[34]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 416.200 460.000 416.800 ;
    END
  END bus_in[34]
  PIN bus_in[35]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 428.440 460.000 429.040 ;
    END
  END bus_in[35]
  PIN bus_in[36]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 434.560 460.000 435.160 ;
    END
  END bus_in[36]
  PIN bus_in[37]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 440.680 460.000 441.280 ;
    END
  END bus_in[37]
  PIN bus_in[38]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 446.800 460.000 447.400 ;
    END
  END bus_in[38]
  PIN bus_in[39]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 452.920 460.000 453.520 ;
    END
  END bus_in[39]
  PIN bus_in[3]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 38.800 460.000 39.400 ;
    END
  END bus_in[3]
  PIN bus_in[40]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 459.040 460.000 459.640 ;
    END
  END bus_in[40]
  PIN bus_in[41]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 230.090 458.400 230.370 462.400 ;
    END
  END bus_in[41]
  PIN bus_in[4]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 51.040 460.000 51.640 ;
    END
  END bus_in[4]
  PIN bus_in[5]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 63.280 460.000 63.880 ;
    END
  END bus_in[5]
  PIN bus_in[6]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 75.520 460.000 76.120 ;
    END
  END bus_in[6]
  PIN bus_in[7]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 87.760 460.000 88.360 ;
    END
  END bus_in[7]
  PIN bus_in[8]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 100.000 460.000 100.600 ;
    END
  END bus_in[8]
  PIN bus_in[9]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 456.000 112.240 460.000 112.840 ;
    END
  END bus_in[9]
  PIN bus_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 8.200 460.000 8.800 ;
    END
  END bus_out[0]
  PIN bus_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 129.920 460.000 130.520 ;
    END
  END bus_out[10]
  PIN bus_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 142.160 460.000 142.760 ;
    END
  END bus_out[11]
  PIN bus_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 154.400 460.000 155.000 ;
    END
  END bus_out[12]
  PIN bus_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 166.640 460.000 167.240 ;
    END
  END bus_out[13]
  PIN bus_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 178.880 460.000 179.480 ;
    END
  END bus_out[14]
  PIN bus_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 191.120 460.000 191.720 ;
    END
  END bus_out[15]
  PIN bus_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 203.360 460.000 203.960 ;
    END
  END bus_out[16]
  PIN bus_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 215.600 460.000 216.200 ;
    END
  END bus_out[17]
  PIN bus_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 227.840 460.000 228.440 ;
    END
  END bus_out[18]
  PIN bus_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 239.400 460.000 240.000 ;
    END
  END bus_out[19]
  PIN bus_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 20.440 460.000 21.040 ;
    END
  END bus_out[1]
  PIN bus_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 251.640 460.000 252.240 ;
    END
  END bus_out[20]
  PIN bus_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 263.880 460.000 264.480 ;
    END
  END bus_out[21]
  PIN bus_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 276.120 460.000 276.720 ;
    END
  END bus_out[22]
  PIN bus_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 288.360 460.000 288.960 ;
    END
  END bus_out[23]
  PIN bus_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 300.600 460.000 301.200 ;
    END
  END bus_out[24]
  PIN bus_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 312.840 460.000 313.440 ;
    END
  END bus_out[25]
  PIN bus_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 325.080 460.000 325.680 ;
    END
  END bus_out[26]
  PIN bus_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 337.320 460.000 337.920 ;
    END
  END bus_out[27]
  PIN bus_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 349.560 460.000 350.160 ;
    END
  END bus_out[28]
  PIN bus_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 361.120 460.000 361.720 ;
    END
  END bus_out[29]
  PIN bus_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 32.680 460.000 33.280 ;
    END
  END bus_out[2]
  PIN bus_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 373.360 460.000 373.960 ;
    END
  END bus_out[30]
  PIN bus_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 385.600 460.000 386.200 ;
    END
  END bus_out[31]
  PIN bus_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 397.840 460.000 398.440 ;
    END
  END bus_out[32]
  PIN bus_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 410.080 460.000 410.680 ;
    END
  END bus_out[33]
  PIN bus_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 422.320 460.000 422.920 ;
    END
  END bus_out[34]
  PIN bus_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 44.920 460.000 45.520 ;
    END
  END bus_out[3]
  PIN bus_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 57.160 460.000 57.760 ;
    END
  END bus_out[4]
  PIN bus_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 69.400 460.000 70.000 ;
    END
  END bus_out[5]
  PIN bus_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 81.640 460.000 82.240 ;
    END
  END bus_out[6]
  PIN bus_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 93.880 460.000 94.480 ;
    END
  END bus_out[7]
  PIN bus_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 106.120 460.000 106.720 ;
    END
  END bus_out[8]
  PIN bus_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 456.000 118.360 460.000 118.960 ;
    END
  END bus_out[9]
  PIN clk_i
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 115.090 0.000 115.370 4.000 ;
    END
  END clk_i
  PIN inp_i
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 0.000 231.240 4.000 231.840 ;
    END
  END inp_i
  PIN rst_n_i
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 345.090 0.000 345.370 4.000 ;
    END
  END rst_n_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT 
      LAYER met4 ;
      RECT 174.64 10.64 176.24 451.76 ;
      RECT 328.24 10.64 329.84 451.76 ;
      RECT 21.040 10.640 22.640 451.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT 
      LAYER met4 ;
      RECT 251.44 10.64 253.04 451.76 ;
      RECT 405.04 10.64 406.64 451.76 ;
      RECT 97.840 10.640 99.440 451.760 ;
    END
  END VGND
  OBS 
    LAYER li1 ;
    RECT 5.520 10.795 455.255 451.605 ;
    LAYER met1 ;
    RECT 5.520 10.640 455.330 451.760 ;
    LAYER met2 ;
    RECT 8.840 458.120 229.810 459.525 ;
    RECT 230.650 458.120 455.310 459.525 ;
    RECT 8.840 4.280 455.310 458.120 ;
    RECT 8.840 2.875 114.810 4.280 ;
    RECT 115.650 2.875 344.810 4.280 ;
    RECT 345.650 2.875 455.310 4.280 ;
    LAYER met3 ;
    RECT 4.000 458.640 455.600 459.505 ;
    RECT 4.000 453.920 456.000 458.640 ;
    RECT 4.000 452.520 455.600 453.920 ;
    RECT 4.000 447.800 456.000 452.520 ;
    RECT 4.000 446.400 455.600 447.800 ;
    RECT 4.000 441.680 456.000 446.400 ;
    RECT 4.000 440.280 455.600 441.680 ;
    RECT 4.000 435.560 456.000 440.280 ;
    RECT 4.000 434.160 455.600 435.560 ;
    RECT 4.000 429.440 456.000 434.160 ;
    RECT 4.000 428.040 455.600 429.440 ;
    RECT 4.000 423.320 456.000 428.040 ;
    RECT 4.000 421.920 455.600 423.320 ;
    RECT 4.000 417.200 456.000 421.920 ;
    RECT 4.000 415.800 455.600 417.200 ;
    RECT 4.000 411.080 456.000 415.800 ;
    RECT 4.000 409.680 455.600 411.080 ;
    RECT 4.000 404.960 456.000 409.680 ;
    RECT 4.000 403.560 455.600 404.960 ;
    RECT 4.000 398.840 456.000 403.560 ;
    RECT 4.000 397.440 455.600 398.840 ;
    RECT 4.000 392.720 456.000 397.440 ;
    RECT 4.000 391.320 455.600 392.720 ;
    RECT 4.000 386.600 456.000 391.320 ;
    RECT 4.000 385.200 455.600 386.600 ;
    RECT 4.000 380.480 456.000 385.200 ;
    RECT 4.000 379.080 455.600 380.480 ;
    RECT 4.000 374.360 456.000 379.080 ;
    RECT 4.000 372.960 455.600 374.360 ;
    RECT 4.000 368.240 456.000 372.960 ;
    RECT 4.000 366.840 455.600 368.240 ;
    RECT 4.000 362.120 456.000 366.840 ;
    RECT 4.000 360.720 455.600 362.120 ;
    RECT 4.000 356.000 456.000 360.720 ;
    RECT 4.000 354.600 455.600 356.000 ;
    RECT 4.000 350.560 456.000 354.600 ;
    RECT 4.000 349.160 455.600 350.560 ;
    RECT 4.000 344.440 456.000 349.160 ;
    RECT 4.000 343.040 455.600 344.440 ;
    RECT 4.000 338.320 456.000 343.040 ;
    RECT 4.000 336.920 455.600 338.320 ;
    RECT 4.000 332.200 456.000 336.920 ;
    RECT 4.000 330.800 455.600 332.200 ;
    RECT 4.000 326.080 456.000 330.800 ;
    RECT 4.000 324.680 455.600 326.080 ;
    RECT 4.000 319.960 456.000 324.680 ;
    RECT 4.000 318.560 455.600 319.960 ;
    RECT 4.000 313.840 456.000 318.560 ;
    RECT 4.000 312.440 455.600 313.840 ;
    RECT 4.000 307.720 456.000 312.440 ;
    RECT 4.000 306.320 455.600 307.720 ;
    RECT 4.000 301.600 456.000 306.320 ;
    RECT 4.000 300.200 455.600 301.600 ;
    RECT 4.000 295.480 456.000 300.200 ;
    RECT 4.000 294.080 455.600 295.480 ;
    RECT 4.000 289.360 456.000 294.080 ;
    RECT 4.000 287.960 455.600 289.360 ;
    RECT 4.000 283.240 456.000 287.960 ;
    RECT 4.000 281.840 455.600 283.240 ;
    RECT 4.000 277.120 456.000 281.840 ;
    RECT 4.000 275.720 455.600 277.120 ;
    RECT 4.000 271.000 456.000 275.720 ;
    RECT 4.000 269.600 455.600 271.000 ;
    RECT 4.000 264.880 456.000 269.600 ;
    RECT 4.000 263.480 455.600 264.880 ;
    RECT 4.000 258.760 456.000 263.480 ;
    RECT 4.000 257.360 455.600 258.760 ;
    RECT 4.000 252.640 456.000 257.360 ;
    RECT 4.000 251.240 455.600 252.640 ;
    RECT 4.000 246.520 456.000 251.240 ;
    RECT 4.000 245.120 455.600 246.520 ;
    RECT 4.000 240.400 456.000 245.120 ;
    RECT 4.000 239.000 455.600 240.400 ;
    RECT 4.000 234.960 456.000 239.000 ;
    RECT 4.000 233.560 455.600 234.960 ;
    RECT 4.000 232.240 456.000 233.560 ;
    RECT 4.400 230.840 456.000 232.240 ;
    RECT 4.000 228.840 456.000 230.840 ;
    RECT 4.000 227.440 455.600 228.840 ;
    RECT 4.000 222.720 456.000 227.440 ;
    RECT 4.000 221.320 455.600 222.720 ;
    RECT 4.000 216.600 456.000 221.320 ;
    RECT 4.000 215.200 455.600 216.600 ;
    RECT 4.000 210.480 456.000 215.200 ;
    RECT 4.000 209.080 455.600 210.480 ;
    RECT 4.000 204.360 456.000 209.080 ;
    RECT 4.000 202.960 455.600 204.360 ;
    RECT 4.000 198.240 456.000 202.960 ;
    RECT 4.000 196.840 455.600 198.240 ;
    RECT 4.000 192.120 456.000 196.840 ;
    RECT 4.000 190.720 455.600 192.120 ;
    RECT 4.000 186.000 456.000 190.720 ;
    RECT 4.000 184.600 455.600 186.000 ;
    RECT 4.000 179.880 456.000 184.600 ;
    RECT 4.000 178.480 455.600 179.880 ;
    RECT 4.000 173.760 456.000 178.480 ;
    RECT 4.000 172.360 455.600 173.760 ;
    RECT 4.000 167.640 456.000 172.360 ;
    RECT 4.000 166.240 455.600 167.640 ;
    RECT 4.000 161.520 456.000 166.240 ;
    RECT 4.000 160.120 455.600 161.520 ;
    RECT 4.000 155.400 456.000 160.120 ;
    RECT 4.000 154.000 455.600 155.400 ;
    RECT 4.000 149.280 456.000 154.000 ;
    RECT 4.000 147.880 455.600 149.280 ;
    RECT 4.000 143.160 456.000 147.880 ;
    RECT 4.000 141.760 455.600 143.160 ;
    RECT 4.000 137.040 456.000 141.760 ;
    RECT 4.000 135.640 455.600 137.040 ;
    RECT 4.000 130.920 456.000 135.640 ;
    RECT 4.000 129.520 455.600 130.920 ;
    RECT 4.000 124.800 456.000 129.520 ;
    RECT 4.000 123.400 455.600 124.800 ;
    RECT 4.000 119.360 456.000 123.400 ;
    RECT 4.000 117.960 455.600 119.360 ;
    RECT 4.000 113.240 456.000 117.960 ;
    RECT 4.000 111.840 455.600 113.240 ;
    RECT 4.000 107.120 456.000 111.840 ;
    RECT 4.000 105.720 455.600 107.120 ;
    RECT 4.000 101.000 456.000 105.720 ;
    RECT 4.000 99.600 455.600 101.000 ;
    RECT 4.000 94.880 456.000 99.600 ;
    RECT 4.000 93.480 455.600 94.880 ;
    RECT 4.000 88.760 456.000 93.480 ;
    RECT 4.000 87.360 455.600 88.760 ;
    RECT 4.000 82.640 456.000 87.360 ;
    RECT 4.000 81.240 455.600 82.640 ;
    RECT 4.000 76.520 456.000 81.240 ;
    RECT 4.000 75.120 455.600 76.520 ;
    RECT 4.000 70.400 456.000 75.120 ;
    RECT 4.000 69.000 455.600 70.400 ;
    RECT 4.000 64.280 456.000 69.000 ;
    RECT 4.000 62.880 455.600 64.280 ;
    RECT 4.000 58.160 456.000 62.880 ;
    RECT 4.000 56.760 455.600 58.160 ;
    RECT 4.000 52.040 456.000 56.760 ;
    RECT 4.000 50.640 455.600 52.040 ;
    RECT 4.000 45.920 456.000 50.640 ;
    RECT 4.000 44.520 455.600 45.920 ;
    RECT 4.000 39.800 456.000 44.520 ;
    RECT 4.000 38.400 455.600 39.800 ;
    RECT 4.000 33.680 456.000 38.400 ;
    RECT 4.000 32.280 455.600 33.680 ;
    RECT 4.000 27.560 456.000 32.280 ;
    RECT 4.000 26.160 455.600 27.560 ;
    RECT 4.000 21.440 456.000 26.160 ;
    RECT 4.000 20.040 455.600 21.440 ;
    RECT 4.000 15.320 456.000 20.040 ;
    RECT 4.000 13.920 455.600 15.320 ;
    RECT 4.000 9.200 456.000 13.920 ;
    RECT 4.000 7.800 455.600 9.200 ;
    RECT 4.000 3.760 456.000 7.800 ;
    RECT 4.000 2.895 455.600 3.760 ;
    LAYER met4 ;
    RECT 174.640 10.640 406.640 451.760 ;
  END
END tdc_inline_2
END LIBRARY
