VERSION 5.7 ;
NOWIREEXTENSIONATPIN ON ;
DIVIDERCHAR "/" ;
BUSBITCHARS "[]" ;
MACRO tdc_inline_1
  CLASS BLOCK ;
  FOREIGN tdc_inline_1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 414.000 BY 340.000 ;
  PIN bus_in[0]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 2.080 414.000 2.680 ;
    END
  END bus_in[0]
  PIN bus_in[10]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 91.160 414.000 91.760 ;
    END
  END bus_in[10]
  PIN bus_in[11]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 100.000 414.000 100.600 ;
    END
  END bus_in[11]
  PIN bus_in[12]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 108.840 414.000 109.440 ;
    END
  END bus_in[12]
  PIN bus_in[13]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 118.360 414.000 118.960 ;
    END
  END bus_in[13]
  PIN bus_in[14]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 127.200 414.000 127.800 ;
    END
  END bus_in[14]
  PIN bus_in[15]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 136.040 414.000 136.640 ;
    END
  END bus_in[15]
  PIN bus_in[16]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 144.880 414.000 145.480 ;
    END
  END bus_in[16]
  PIN bus_in[17]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 153.720 414.000 154.320 ;
    END
  END bus_in[17]
  PIN bus_in[18]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 162.560 414.000 163.160 ;
    END
  END bus_in[18]
  PIN bus_in[19]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 172.080 414.000 172.680 ;
    END
  END bus_in[19]
  PIN bus_in[1]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 10.920 414.000 11.520 ;
    END
  END bus_in[1]
  PIN bus_in[20]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 180.920 414.000 181.520 ;
    END
  END bus_in[20]
  PIN bus_in[21]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 189.760 414.000 190.360 ;
    END
  END bus_in[21]
  PIN bus_in[22]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 198.600 414.000 199.200 ;
    END
  END bus_in[22]
  PIN bus_in[23]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 207.440 414.000 208.040 ;
    END
  END bus_in[23]
  PIN bus_in[24]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 216.280 414.000 216.880 ;
    END
  END bus_in[24]
  PIN bus_in[25]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 225.120 414.000 225.720 ;
    END
  END bus_in[25]
  PIN bus_in[26]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 234.640 414.000 235.240 ;
    END
  END bus_in[26]
  PIN bus_in[27]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 243.480 414.000 244.080 ;
    END
  END bus_in[27]
  PIN bus_in[28]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 252.320 414.000 252.920 ;
    END
  END bus_in[28]
  PIN bus_in[29]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 261.160 414.000 261.760 ;
    END
  END bus_in[29]
  PIN bus_in[2]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 19.760 414.000 20.360 ;
    END
  END bus_in[2]
  PIN bus_in[30]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 270.000 414.000 270.600 ;
    END
  END bus_in[30]
  PIN bus_in[31]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 278.840 414.000 279.440 ;
    END
  END bus_in[31]
  PIN bus_in[32]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 288.360 414.000 288.960 ;
    END
  END bus_in[32]
  PIN bus_in[33]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 297.200 414.000 297.800 ;
    END
  END bus_in[33]
  PIN bus_in[34]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 306.040 414.000 306.640 ;
    END
  END bus_in[34]
  PIN bus_in[35]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 314.880 414.000 315.480 ;
    END
  END bus_in[35]
  PIN bus_in[36]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 319.640 414.000 320.240 ;
    END
  END bus_in[36]
  PIN bus_in[37]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 323.720 414.000 324.320 ;
    END
  END bus_in[37]
  PIN bus_in[38]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 328.480 414.000 329.080 ;
    END
  END bus_in[38]
  PIN bus_in[39]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 332.560 414.000 333.160 ;
    END
  END bus_in[39]
  PIN bus_in[3]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 28.600 414.000 29.200 ;
    END
  END bus_in[3]
  PIN bus_in[40]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 337.320 414.000 337.920 ;
    END
  END bus_in[40]
  PIN bus_in[41]
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 207.090 336.000 207.370 340.000 ;
    END
  END bus_in[41]
  PIN bus_in[4]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 37.440 414.000 38.040 ;
    END
  END bus_in[4]
  PIN bus_in[5]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 46.280 414.000 46.880 ;
    END
  END bus_in[5]
  PIN bus_in[6]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 55.120 414.000 55.720 ;
    END
  END bus_in[6]
  PIN bus_in[7]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 64.640 414.000 65.240 ;
    END
  END bus_in[7]
  PIN bus_in[8]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 73.480 414.000 74.080 ;
    END
  END bus_in[8]
  PIN bus_in[9]
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 410.000 82.320 414.000 82.920 ;
    END
  END bus_in[9]
  PIN bus_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 6.160 414.000 6.760 ;
    END
  END bus_out[0]
  PIN bus_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 95.920 414.000 96.520 ;
    END
  END bus_out[10]
  PIN bus_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 104.760 414.000 105.360 ;
    END
  END bus_out[11]
  PIN bus_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 113.600 414.000 114.200 ;
    END
  END bus_out[12]
  PIN bus_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 122.440 414.000 123.040 ;
    END
  END bus_out[13]
  PIN bus_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 131.280 414.000 131.880 ;
    END
  END bus_out[14]
  PIN bus_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 140.120 414.000 140.720 ;
    END
  END bus_out[15]
  PIN bus_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 149.640 414.000 150.240 ;
    END
  END bus_out[16]
  PIN bus_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 158.480 414.000 159.080 ;
    END
  END bus_out[17]
  PIN bus_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 167.320 414.000 167.920 ;
    END
  END bus_out[18]
  PIN bus_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 176.160 414.000 176.760 ;
    END
  END bus_out[19]
  PIN bus_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 15.000 414.000 15.600 ;
    END
  END bus_out[1]
  PIN bus_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 185.000 414.000 185.600 ;
    END
  END bus_out[20]
  PIN bus_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 193.840 414.000 194.440 ;
    END
  END bus_out[21]
  PIN bus_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 203.360 414.000 203.960 ;
    END
  END bus_out[22]
  PIN bus_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 212.200 414.000 212.800 ;
    END
  END bus_out[23]
  PIN bus_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 221.040 414.000 221.640 ;
    END
  END bus_out[24]
  PIN bus_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 229.880 414.000 230.480 ;
    END
  END bus_out[25]
  PIN bus_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 238.720 414.000 239.320 ;
    END
  END bus_out[26]
  PIN bus_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 247.560 414.000 248.160 ;
    END
  END bus_out[27]
  PIN bus_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 257.080 414.000 257.680 ;
    END
  END bus_out[28]
  PIN bus_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 265.920 414.000 266.520 ;
    END
  END bus_out[29]
  PIN bus_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 23.840 414.000 24.440 ;
    END
  END bus_out[2]
  PIN bus_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 274.760 414.000 275.360 ;
    END
  END bus_out[30]
  PIN bus_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 283.600 414.000 284.200 ;
    END
  END bus_out[31]
  PIN bus_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 292.440 414.000 293.040 ;
    END
  END bus_out[32]
  PIN bus_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 301.280 414.000 301.880 ;
    END
  END bus_out[33]
  PIN bus_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 310.120 414.000 310.720 ;
    END
  END bus_out[34]
  PIN bus_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 33.360 414.000 33.960 ;
    END
  END bus_out[3]
  PIN bus_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 42.200 414.000 42.800 ;
    END
  END bus_out[4]
  PIN bus_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 51.040 414.000 51.640 ;
    END
  END bus_out[5]
  PIN bus_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 59.880 414.000 60.480 ;
    END
  END bus_out[6]
  PIN bus_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 68.720 414.000 69.320 ;
    END
  END bus_out[7]
  PIN bus_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 77.560 414.000 78.160 ;
    END
  END bus_out[8]
  PIN bus_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT 
      LAYER met3 ;
      RECT 410.000 87.080 414.000 87.680 ;
    END
  END bus_out[9]
  PIN clk_i
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 103.590 0.000 103.870 4.000 ;
    END
  END clk_i
  PIN inp_i
    DIRECTION INPUT ;
    PORT 
      LAYER met3 ;
      RECT 0.000 170.040 4.000 170.640 ;
    END
  END inp_i
  PIN rst_n_i
    DIRECTION INPUT ;
    PORT 
      LAYER met2 ;
      RECT 310.590 0.000 310.870 4.000 ;
    END
  END rst_n_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT 
      LAYER met4 ;
      RECT 174.64 10.64 176.24 329.36 ;
      RECT 328.24 10.64 329.84 329.36 ;
      RECT 21.040 10.640 22.640 329.360 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT 
      LAYER met4 ;
      RECT 251.44 10.64 253.04 329.36 ;
      RECT 405.04 10.64 406.64 329.36 ;
      RECT 97.840 10.640 99.440 329.360 ;
    END
  END VGND
  OBS 
    LAYER li1 ;
    RECT 5.520 10.795 408.480 329.205 ;
    LAYER met1 ;
    RECT 5.520 10.640 408.480 329.360 ;
    LAYER met2 ;
    RECT 10.680 335.720 206.810 337.805 ;
    RECT 207.650 335.720 407.470 337.805 ;
    RECT 10.680 4.280 407.470 335.720 ;
    RECT 10.680 2.195 103.310 4.280 ;
    RECT 104.150 2.195 310.310 4.280 ;
    RECT 311.150 2.195 407.470 4.280 ;
    LAYER met3 ;
    RECT 4.000 336.920 409.600 337.785 ;
    RECT 4.000 333.560 410.000 336.920 ;
    RECT 4.000 332.160 409.600 333.560 ;
    RECT 4.000 329.480 410.000 332.160 ;
    RECT 4.000 328.080 409.600 329.480 ;
    RECT 4.000 324.720 410.000 328.080 ;
    RECT 4.000 323.320 409.600 324.720 ;
    RECT 4.000 320.640 410.000 323.320 ;
    RECT 4.000 319.240 409.600 320.640 ;
    RECT 4.000 315.880 410.000 319.240 ;
    RECT 4.000 314.480 409.600 315.880 ;
    RECT 4.000 311.120 410.000 314.480 ;
    RECT 4.000 309.720 409.600 311.120 ;
    RECT 4.000 307.040 410.000 309.720 ;
    RECT 4.000 305.640 409.600 307.040 ;
    RECT 4.000 302.280 410.000 305.640 ;
    RECT 4.000 300.880 409.600 302.280 ;
    RECT 4.000 298.200 410.000 300.880 ;
    RECT 4.000 296.800 409.600 298.200 ;
    RECT 4.000 293.440 410.000 296.800 ;
    RECT 4.000 292.040 409.600 293.440 ;
    RECT 4.000 289.360 410.000 292.040 ;
    RECT 4.000 287.960 409.600 289.360 ;
    RECT 4.000 284.600 410.000 287.960 ;
    RECT 4.000 283.200 409.600 284.600 ;
    RECT 4.000 279.840 410.000 283.200 ;
    RECT 4.000 278.440 409.600 279.840 ;
    RECT 4.000 275.760 410.000 278.440 ;
    RECT 4.000 274.360 409.600 275.760 ;
    RECT 4.000 271.000 410.000 274.360 ;
    RECT 4.000 269.600 409.600 271.000 ;
    RECT 4.000 266.920 410.000 269.600 ;
    RECT 4.000 265.520 409.600 266.920 ;
    RECT 4.000 262.160 410.000 265.520 ;
    RECT 4.000 260.760 409.600 262.160 ;
    RECT 4.000 258.080 410.000 260.760 ;
    RECT 4.000 256.680 409.600 258.080 ;
    RECT 4.000 253.320 410.000 256.680 ;
    RECT 4.000 251.920 409.600 253.320 ;
    RECT 4.000 248.560 410.000 251.920 ;
    RECT 4.000 247.160 409.600 248.560 ;
    RECT 4.000 244.480 410.000 247.160 ;
    RECT 4.000 243.080 409.600 244.480 ;
    RECT 4.000 239.720 410.000 243.080 ;
    RECT 4.000 238.320 409.600 239.720 ;
    RECT 4.000 235.640 410.000 238.320 ;
    RECT 4.000 234.240 409.600 235.640 ;
    RECT 4.000 230.880 410.000 234.240 ;
    RECT 4.000 229.480 409.600 230.880 ;
    RECT 4.000 226.120 410.000 229.480 ;
    RECT 4.000 224.720 409.600 226.120 ;
    RECT 4.000 222.040 410.000 224.720 ;
    RECT 4.000 220.640 409.600 222.040 ;
    RECT 4.000 217.280 410.000 220.640 ;
    RECT 4.000 215.880 409.600 217.280 ;
    RECT 4.000 213.200 410.000 215.880 ;
    RECT 4.000 211.800 409.600 213.200 ;
    RECT 4.000 208.440 410.000 211.800 ;
    RECT 4.000 207.040 409.600 208.440 ;
    RECT 4.000 204.360 410.000 207.040 ;
    RECT 4.000 202.960 409.600 204.360 ;
    RECT 4.000 199.600 410.000 202.960 ;
    RECT 4.000 198.200 409.600 199.600 ;
    RECT 4.000 194.840 410.000 198.200 ;
    RECT 4.000 193.440 409.600 194.840 ;
    RECT 4.000 190.760 410.000 193.440 ;
    RECT 4.000 189.360 409.600 190.760 ;
    RECT 4.000 186.000 410.000 189.360 ;
    RECT 4.000 184.600 409.600 186.000 ;
    RECT 4.000 181.920 410.000 184.600 ;
    RECT 4.000 180.520 409.600 181.920 ;
    RECT 4.000 177.160 410.000 180.520 ;
    RECT 4.000 175.760 409.600 177.160 ;
    RECT 4.000 173.080 410.000 175.760 ;
    RECT 4.000 171.680 409.600 173.080 ;
    RECT 4.000 171.040 410.000 171.680 ;
    RECT 4.400 169.640 410.000 171.040 ;
    RECT 4.000 168.320 410.000 169.640 ;
    RECT 4.000 166.920 409.600 168.320 ;
    RECT 4.000 163.560 410.000 166.920 ;
    RECT 4.000 162.160 409.600 163.560 ;
    RECT 4.000 159.480 410.000 162.160 ;
    RECT 4.000 158.080 409.600 159.480 ;
    RECT 4.000 154.720 410.000 158.080 ;
    RECT 4.000 153.320 409.600 154.720 ;
    RECT 4.000 150.640 410.000 153.320 ;
    RECT 4.000 149.240 409.600 150.640 ;
    RECT 4.000 145.880 410.000 149.240 ;
    RECT 4.000 144.480 409.600 145.880 ;
    RECT 4.000 141.120 410.000 144.480 ;
    RECT 4.000 139.720 409.600 141.120 ;
    RECT 4.000 137.040 410.000 139.720 ;
    RECT 4.000 135.640 409.600 137.040 ;
    RECT 4.000 132.280 410.000 135.640 ;
    RECT 4.000 130.880 409.600 132.280 ;
    RECT 4.000 128.200 410.000 130.880 ;
    RECT 4.000 126.800 409.600 128.200 ;
    RECT 4.000 123.440 410.000 126.800 ;
    RECT 4.000 122.040 409.600 123.440 ;
    RECT 4.000 119.360 410.000 122.040 ;
    RECT 4.000 117.960 409.600 119.360 ;
    RECT 4.000 114.600 410.000 117.960 ;
    RECT 4.000 113.200 409.600 114.600 ;
    RECT 4.000 109.840 410.000 113.200 ;
    RECT 4.000 108.440 409.600 109.840 ;
    RECT 4.000 105.760 410.000 108.440 ;
    RECT 4.000 104.360 409.600 105.760 ;
    RECT 4.000 101.000 410.000 104.360 ;
    RECT 4.000 99.600 409.600 101.000 ;
    RECT 4.000 96.920 410.000 99.600 ;
    RECT 4.000 95.520 409.600 96.920 ;
    RECT 4.000 92.160 410.000 95.520 ;
    RECT 4.000 90.760 409.600 92.160 ;
    RECT 4.000 88.080 410.000 90.760 ;
    RECT 4.000 86.680 409.600 88.080 ;
    RECT 4.000 83.320 410.000 86.680 ;
    RECT 4.000 81.920 409.600 83.320 ;
    RECT 4.000 78.560 410.000 81.920 ;
    RECT 4.000 77.160 409.600 78.560 ;
    RECT 4.000 74.480 410.000 77.160 ;
    RECT 4.000 73.080 409.600 74.480 ;
    RECT 4.000 69.720 410.000 73.080 ;
    RECT 4.000 68.320 409.600 69.720 ;
    RECT 4.000 65.640 410.000 68.320 ;
    RECT 4.000 64.240 409.600 65.640 ;
    RECT 4.000 60.880 410.000 64.240 ;
    RECT 4.000 59.480 409.600 60.880 ;
    RECT 4.000 56.120 410.000 59.480 ;
    RECT 4.000 54.720 409.600 56.120 ;
    RECT 4.000 52.040 410.000 54.720 ;
    RECT 4.000 50.640 409.600 52.040 ;
    RECT 4.000 47.280 410.000 50.640 ;
    RECT 4.000 45.880 409.600 47.280 ;
    RECT 4.000 43.200 410.000 45.880 ;
    RECT 4.000 41.800 409.600 43.200 ;
    RECT 4.000 38.440 410.000 41.800 ;
    RECT 4.000 37.040 409.600 38.440 ;
    RECT 4.000 34.360 410.000 37.040 ;
    RECT 4.000 32.960 409.600 34.360 ;
    RECT 4.000 29.600 410.000 32.960 ;
    RECT 4.000 28.200 409.600 29.600 ;
    RECT 4.000 24.840 410.000 28.200 ;
    RECT 4.000 23.440 409.600 24.840 ;
    RECT 4.000 20.760 410.000 23.440 ;
    RECT 4.000 19.360 409.600 20.760 ;
    RECT 4.000 16.000 410.000 19.360 ;
    RECT 4.000 14.600 409.600 16.000 ;
    RECT 4.000 11.920 410.000 14.600 ;
    RECT 4.000 10.520 409.600 11.920 ;
    RECT 4.000 7.160 410.000 10.520 ;
    RECT 4.000 5.760 409.600 7.160 ;
    RECT 4.000 3.080 410.000 5.760 ;
    RECT 4.000 2.215 409.600 3.080 ;
    LAYER met4 ;
    RECT 174.640 10.640 406.640 329.360 ;
  END
END tdc_inline_1
END LIBRARY
