magic
tech sky130A
magscale 1 2
timestamp 1607274944
<< viali >>
rect 1933 22025 1967 22059
rect 2301 21957 2335 21991
rect 2393 21889 2427 21923
rect 3129 21889 3163 21923
rect 2485 21821 2519 21855
rect 3773 21753 3807 21787
rect 1933 21481 1967 21515
rect 2485 21345 2519 21379
rect 2393 21277 2427 21311
rect 3129 21277 3163 21311
rect 2301 21209 2335 21243
rect 3773 21209 3807 21243
rect 3773 20937 3807 20971
rect 3129 20801 3163 20835
rect 1933 20393 1967 20427
rect 2485 20257 2519 20291
rect 4877 20257 4911 20291
rect 2393 20189 2427 20223
rect 3129 20189 3163 20223
rect 4233 20189 4267 20223
rect 3773 20121 3807 20155
rect 2301 20053 2335 20087
rect 4877 19849 4911 19883
rect 3129 19713 3163 19747
rect 3773 19713 3807 19747
rect 4233 19713 4267 19747
rect 1933 19305 1967 19339
rect 2485 19169 2519 19203
rect 4877 19169 4911 19203
rect 7085 19169 7119 19203
rect 2393 19101 2427 19135
rect 3129 19101 3163 19135
rect 4233 19101 4267 19135
rect 5337 19101 5371 19135
rect 6441 19101 6475 19135
rect 3773 19033 3807 19067
rect 5981 19033 6015 19067
rect 2301 18965 2335 18999
rect 7085 18761 7119 18795
rect 3129 18625 3163 18659
rect 3773 18625 3807 18659
rect 4233 18625 4267 18659
rect 4877 18625 4911 18659
rect 5337 18625 5371 18659
rect 5981 18625 6015 18659
rect 6441 18625 6475 18659
rect 1933 18217 1967 18251
rect 2485 18081 2519 18115
rect 4877 18081 4911 18115
rect 7085 18081 7119 18115
rect 8189 18081 8223 18115
rect 10397 18081 10431 18115
rect 2393 18013 2427 18047
rect 3129 18013 3163 18047
rect 4233 18013 4267 18047
rect 5337 18013 5371 18047
rect 6452 18013 6486 18047
rect 7545 18013 7579 18047
rect 8660 18013 8694 18047
rect 9753 18013 9787 18047
rect 10857 18013 10891 18047
rect 3773 17945 3807 17979
rect 5981 17945 6015 17979
rect 9293 17945 9327 17979
rect 11501 17945 11535 17979
rect 2301 17877 2335 17911
rect 11501 17673 11535 17707
rect 3129 17537 3163 17571
rect 3773 17537 3807 17571
rect 4233 17537 4267 17571
rect 4877 17537 4911 17571
rect 5337 17537 5371 17571
rect 5981 17537 6015 17571
rect 6441 17537 6475 17571
rect 7085 17537 7119 17571
rect 7545 17537 7579 17571
rect 8189 17537 8223 17571
rect 8649 17537 8683 17571
rect 9293 17537 9327 17571
rect 9753 17537 9787 17571
rect 10397 17537 10431 17571
rect 10857 17537 10891 17571
rect 1933 17129 1967 17163
rect 2485 16993 2519 17027
rect 4877 16993 4911 17027
rect 7085 16993 7119 17027
rect 8189 16993 8223 17027
rect 10397 16993 10431 17027
rect 11501 16993 11535 17027
rect 13709 16993 13743 17027
rect 15917 16993 15951 17027
rect 18125 16993 18159 17027
rect 20333 16993 20367 17027
rect 3129 16925 3163 16959
rect 4233 16925 4267 16959
rect 5337 16925 5371 16959
rect 6452 16925 6486 16959
rect 7545 16925 7579 16959
rect 8660 16925 8694 16959
rect 9753 16925 9787 16959
rect 10857 16925 10891 16959
rect 11961 16925 11995 16959
rect 13065 16925 13099 16959
rect 14180 16925 14214 16959
rect 15273 16925 15307 16959
rect 16377 16925 16411 16959
rect 17481 16925 17515 16959
rect 18585 16925 18619 16959
rect 19689 16925 19723 16959
rect 2393 16857 2427 16891
rect 3773 16857 3807 16891
rect 5981 16857 6015 16891
rect 9293 16857 9327 16891
rect 12605 16857 12639 16891
rect 14813 16857 14847 16891
rect 17021 16857 17055 16891
rect 19229 16857 19263 16891
rect 2301 16789 2335 16823
rect 20333 16585 20367 16619
rect 3129 16449 3163 16483
rect 3773 16449 3807 16483
rect 4233 16449 4267 16483
rect 4877 16449 4911 16483
rect 5337 16449 5371 16483
rect 5981 16449 6015 16483
rect 6441 16449 6475 16483
rect 7085 16449 7119 16483
rect 7545 16449 7579 16483
rect 8189 16449 8223 16483
rect 8649 16449 8683 16483
rect 9293 16449 9327 16483
rect 9753 16449 9787 16483
rect 10397 16449 10431 16483
rect 10857 16449 10891 16483
rect 11501 16449 11535 16483
rect 11961 16449 11995 16483
rect 12605 16449 12639 16483
rect 13065 16449 13099 16483
rect 13709 16449 13743 16483
rect 14169 16449 14203 16483
rect 14813 16449 14847 16483
rect 15273 16449 15307 16483
rect 15917 16449 15951 16483
rect 16377 16449 16411 16483
rect 17021 16449 17055 16483
rect 17481 16449 17515 16483
rect 18125 16449 18159 16483
rect 18585 16449 18619 16483
rect 19229 16449 19263 16483
rect 19689 16449 19723 16483
rect 1933 15973 1967 16007
rect 2485 15905 2519 15939
rect 4877 15905 4911 15939
rect 7085 15905 7119 15939
rect 9293 15905 9327 15939
rect 10397 15905 10431 15939
rect 11501 15905 11535 15939
rect 13709 15905 13743 15939
rect 15917 15905 15951 15939
rect 18125 15905 18159 15939
rect 20333 15905 20367 15939
rect 2393 15837 2427 15871
rect 3129 15837 3163 15871
rect 4233 15837 4267 15871
rect 5337 15837 5371 15871
rect 6452 15837 6486 15871
rect 7545 15837 7579 15871
rect 8660 15837 8694 15871
rect 9753 15837 9787 15871
rect 10857 15837 10891 15871
rect 11961 15837 11995 15871
rect 13065 15837 13099 15871
rect 14180 15837 14214 15871
rect 15273 15837 15307 15871
rect 16377 15837 16411 15871
rect 17481 15837 17515 15871
rect 18585 15837 18619 15871
rect 19689 15837 19723 15871
rect 3773 15769 3807 15803
rect 5981 15769 6015 15803
rect 8189 15769 8223 15803
rect 12605 15769 12639 15803
rect 14813 15769 14847 15803
rect 17021 15769 17055 15803
rect 19229 15769 19263 15803
rect 2301 15701 2335 15735
rect 20333 15497 20367 15531
rect 3129 15361 3163 15395
rect 3773 15361 3807 15395
rect 4233 15361 4267 15395
rect 4877 15361 4911 15395
rect 5337 15361 5371 15395
rect 5981 15361 6015 15395
rect 6441 15361 6475 15395
rect 7085 15361 7119 15395
rect 7545 15361 7579 15395
rect 8189 15361 8223 15395
rect 8649 15361 8683 15395
rect 9293 15361 9327 15395
rect 9753 15361 9787 15395
rect 10397 15361 10431 15395
rect 10857 15361 10891 15395
rect 11501 15361 11535 15395
rect 11961 15361 11995 15395
rect 12605 15361 12639 15395
rect 13065 15361 13099 15395
rect 13709 15361 13743 15395
rect 14169 15361 14203 15395
rect 14813 15361 14847 15395
rect 15273 15361 15307 15395
rect 15917 15361 15951 15395
rect 16377 15361 16411 15395
rect 17021 15361 17055 15395
rect 17481 15361 17515 15395
rect 18125 15361 18159 15395
rect 18585 15361 18619 15395
rect 19229 15361 19263 15395
rect 19689 15361 19723 15395
rect 3773 14953 3807 14987
rect 5981 14817 6015 14851
rect 8189 14817 8223 14851
rect 11501 14817 11535 14851
rect 13709 14817 13743 14851
rect 15917 14817 15951 14851
rect 18125 14817 18159 14851
rect 20333 14817 20367 14851
rect 3129 14749 3163 14783
rect 4233 14749 4267 14783
rect 5337 14749 5371 14783
rect 6452 14749 6486 14783
rect 7545 14749 7579 14783
rect 8660 14749 8694 14783
rect 9753 14749 9787 14783
rect 10857 14749 10891 14783
rect 11961 14749 11995 14783
rect 13065 14749 13099 14783
rect 14180 14749 14214 14783
rect 15273 14749 15307 14783
rect 16377 14749 16411 14783
rect 17481 14749 17515 14783
rect 18585 14749 18619 14783
rect 19689 14749 19723 14783
rect 4877 14681 4911 14715
rect 7085 14681 7119 14715
rect 9293 14681 9327 14715
rect 10397 14681 10431 14715
rect 12605 14681 12639 14715
rect 14813 14681 14847 14715
rect 17021 14681 17055 14715
rect 19229 14681 19263 14715
rect 20333 14409 20367 14443
rect 3129 14273 3163 14307
rect 3773 14273 3807 14307
rect 4233 14273 4267 14307
rect 4877 14273 4911 14307
rect 5337 14273 5371 14307
rect 5981 14273 6015 14307
rect 6441 14273 6475 14307
rect 7085 14273 7119 14307
rect 7545 14273 7579 14307
rect 8189 14273 8223 14307
rect 8649 14273 8683 14307
rect 9293 14273 9327 14307
rect 9753 14273 9787 14307
rect 10397 14273 10431 14307
rect 10857 14273 10891 14307
rect 11501 14273 11535 14307
rect 11961 14273 11995 14307
rect 12605 14273 12639 14307
rect 13065 14273 13099 14307
rect 13709 14273 13743 14307
rect 14169 14273 14203 14307
rect 14813 14273 14847 14307
rect 15273 14273 15307 14307
rect 15917 14273 15951 14307
rect 16377 14273 16411 14307
rect 17021 14273 17055 14307
rect 17481 14273 17515 14307
rect 18125 14273 18159 14307
rect 18585 14273 18619 14307
rect 19229 14273 19263 14307
rect 19689 14273 19723 14307
rect 1933 13797 1967 13831
rect 2485 13729 2519 13763
rect 4877 13729 4911 13763
rect 7085 13729 7119 13763
rect 8189 13729 8223 13763
rect 10397 13729 10431 13763
rect 11501 13729 11535 13763
rect 13709 13729 13743 13763
rect 15917 13729 15951 13763
rect 18125 13729 18159 13763
rect 20333 13729 20367 13763
rect 3129 13661 3163 13695
rect 4233 13661 4267 13695
rect 5337 13661 5371 13695
rect 6452 13661 6486 13695
rect 7545 13661 7579 13695
rect 8660 13661 8694 13695
rect 9753 13661 9787 13695
rect 10857 13661 10891 13695
rect 11961 13661 11995 13695
rect 13065 13661 13099 13695
rect 14180 13661 14214 13695
rect 15273 13661 15307 13695
rect 16377 13661 16411 13695
rect 17481 13661 17515 13695
rect 18585 13661 18619 13695
rect 19689 13661 19723 13695
rect 2393 13593 2427 13627
rect 3773 13593 3807 13627
rect 5981 13593 6015 13627
rect 9293 13593 9327 13627
rect 12605 13593 12639 13627
rect 14813 13593 14847 13627
rect 17021 13593 17055 13627
rect 19229 13593 19263 13627
rect 2301 13525 2335 13559
rect 20333 13321 20367 13355
rect 3129 13185 3163 13219
rect 3773 13185 3807 13219
rect 4233 13185 4267 13219
rect 4877 13185 4911 13219
rect 5337 13185 5371 13219
rect 5981 13185 6015 13219
rect 6441 13185 6475 13219
rect 7085 13185 7119 13219
rect 7545 13185 7579 13219
rect 8189 13185 8223 13219
rect 8649 13185 8683 13219
rect 9293 13185 9327 13219
rect 9753 13185 9787 13219
rect 10397 13185 10431 13219
rect 10857 13185 10891 13219
rect 11501 13185 11535 13219
rect 11961 13185 11995 13219
rect 12605 13185 12639 13219
rect 13065 13185 13099 13219
rect 13709 13185 13743 13219
rect 14169 13185 14203 13219
rect 14813 13185 14847 13219
rect 15273 13185 15307 13219
rect 15917 13185 15951 13219
rect 16377 13185 16411 13219
rect 17021 13185 17055 13219
rect 17481 13185 17515 13219
rect 18125 13185 18159 13219
rect 18585 13185 18619 13219
rect 19229 13185 19263 13219
rect 19689 13185 19723 13219
rect 3773 12777 3807 12811
rect 5981 12641 6015 12675
rect 9293 12641 9327 12675
rect 10397 12641 10431 12675
rect 11501 12641 11535 12675
rect 13709 12641 13743 12675
rect 15917 12641 15951 12675
rect 18125 12641 18159 12675
rect 20333 12641 20367 12675
rect 3129 12573 3163 12607
rect 4233 12573 4267 12607
rect 5337 12573 5371 12607
rect 6452 12573 6486 12607
rect 7545 12573 7579 12607
rect 8660 12573 8694 12607
rect 9753 12573 9787 12607
rect 10857 12573 10891 12607
rect 11961 12573 11995 12607
rect 13065 12573 13099 12607
rect 14180 12573 14214 12607
rect 15273 12573 15307 12607
rect 16377 12573 16411 12607
rect 17481 12573 17515 12607
rect 18585 12573 18619 12607
rect 19689 12573 19723 12607
rect 4877 12505 4911 12539
rect 7085 12505 7119 12539
rect 8189 12505 8223 12539
rect 12605 12505 12639 12539
rect 14813 12505 14847 12539
rect 17021 12505 17055 12539
rect 19229 12505 19263 12539
rect 20333 12233 20367 12267
rect 3129 12097 3163 12131
rect 3773 12097 3807 12131
rect 4233 12097 4267 12131
rect 4877 12097 4911 12131
rect 5337 12097 5371 12131
rect 5981 12097 6015 12131
rect 6441 12097 6475 12131
rect 7085 12097 7119 12131
rect 7545 12097 7579 12131
rect 8189 12097 8223 12131
rect 8649 12097 8683 12131
rect 9293 12097 9327 12131
rect 9753 12097 9787 12131
rect 10397 12097 10431 12131
rect 10857 12097 10891 12131
rect 11501 12097 11535 12131
rect 11961 12097 11995 12131
rect 12605 12097 12639 12131
rect 13065 12097 13099 12131
rect 13709 12097 13743 12131
rect 14169 12097 14203 12131
rect 14813 12097 14847 12131
rect 15273 12097 15307 12131
rect 15917 12097 15951 12131
rect 16377 12097 16411 12131
rect 17021 12097 17055 12131
rect 17481 12097 17515 12131
rect 18125 12097 18159 12131
rect 18585 12097 18619 12131
rect 19229 12097 19263 12131
rect 19689 12097 19723 12131
rect 3773 11553 3807 11587
rect 4877 11553 4911 11587
rect 7085 11553 7119 11587
rect 8189 11553 8223 11587
rect 10397 11553 10431 11587
rect 12605 11553 12639 11587
rect 14813 11553 14847 11587
rect 17021 11553 17055 11587
rect 19229 11553 19263 11587
rect 3129 11485 3163 11519
rect 4233 11485 4267 11519
rect 5337 11485 5371 11519
rect 6452 11485 6486 11519
rect 7545 11485 7579 11519
rect 8660 11485 8694 11519
rect 9753 11485 9787 11519
rect 10857 11485 10891 11519
rect 11961 11485 11995 11519
rect 13065 11485 13099 11519
rect 14180 11485 14214 11519
rect 15273 11485 15307 11519
rect 16377 11485 16411 11519
rect 17481 11485 17515 11519
rect 18585 11485 18619 11519
rect 19689 11485 19723 11519
rect 5981 11417 6015 11451
rect 9293 11417 9327 11451
rect 11501 11417 11535 11451
rect 13709 11417 13743 11451
rect 15917 11417 15951 11451
rect 18125 11417 18159 11451
rect 20333 11417 20367 11451
rect 20333 11145 20367 11179
rect 3129 11009 3163 11043
rect 3773 11009 3807 11043
rect 4233 11009 4267 11043
rect 4877 11009 4911 11043
rect 5337 11009 5371 11043
rect 5981 11009 6015 11043
rect 6441 11009 6475 11043
rect 7085 11009 7119 11043
rect 7545 11009 7579 11043
rect 8189 11009 8223 11043
rect 8649 11009 8683 11043
rect 9293 11009 9327 11043
rect 9753 11009 9787 11043
rect 10397 11009 10431 11043
rect 10857 11009 10891 11043
rect 11501 11009 11535 11043
rect 11961 11009 11995 11043
rect 12605 11009 12639 11043
rect 13065 11009 13099 11043
rect 13709 11009 13743 11043
rect 14169 11009 14203 11043
rect 14813 11009 14847 11043
rect 15273 11009 15307 11043
rect 15917 11009 15951 11043
rect 16377 11009 16411 11043
rect 17021 11009 17055 11043
rect 17481 11009 17515 11043
rect 18125 11009 18159 11043
rect 18585 11009 18619 11043
rect 19229 11009 19263 11043
rect 19689 11009 19723 11043
rect 3773 10601 3807 10635
rect 4877 10465 4911 10499
rect 7085 10465 7119 10499
rect 9293 10465 9327 10499
rect 10397 10465 10431 10499
rect 11501 10465 11535 10499
rect 13709 10465 13743 10499
rect 17021 10465 17055 10499
rect 19229 10465 19263 10499
rect 3129 10397 3163 10431
rect 4233 10397 4267 10431
rect 5337 10397 5371 10431
rect 6452 10397 6486 10431
rect 7545 10397 7579 10431
rect 8660 10397 8694 10431
rect 9753 10397 9787 10431
rect 10857 10397 10891 10431
rect 11961 10397 11995 10431
rect 13065 10397 13099 10431
rect 14180 10397 14214 10431
rect 15273 10397 15307 10431
rect 16377 10397 16411 10431
rect 17481 10397 17515 10431
rect 18585 10397 18619 10431
rect 19689 10397 19723 10431
rect 5981 10329 6015 10363
rect 8189 10329 8223 10363
rect 12605 10329 12639 10363
rect 14813 10329 14847 10363
rect 15917 10329 15951 10363
rect 18125 10329 18159 10363
rect 20333 10329 20367 10363
rect 20333 10057 20367 10091
rect 3129 9921 3163 9955
rect 3773 9921 3807 9955
rect 4233 9921 4267 9955
rect 4877 9921 4911 9955
rect 5337 9921 5371 9955
rect 5981 9921 6015 9955
rect 6441 9921 6475 9955
rect 7085 9921 7119 9955
rect 7545 9921 7579 9955
rect 8189 9921 8223 9955
rect 8649 9921 8683 9955
rect 9293 9921 9327 9955
rect 9753 9921 9787 9955
rect 10397 9921 10431 9955
rect 10857 9921 10891 9955
rect 11501 9921 11535 9955
rect 11961 9921 11995 9955
rect 12605 9921 12639 9955
rect 13065 9921 13099 9955
rect 13709 9921 13743 9955
rect 14169 9921 14203 9955
rect 14813 9921 14847 9955
rect 15273 9921 15307 9955
rect 15917 9921 15951 9955
rect 16377 9921 16411 9955
rect 17021 9921 17055 9955
rect 17481 9921 17515 9955
rect 18125 9921 18159 9955
rect 18585 9921 18619 9955
rect 19229 9921 19263 9955
rect 19689 9921 19723 9955
rect 2485 9377 2519 9411
rect 5981 9377 6015 9411
rect 8189 9377 8223 9411
rect 10397 9377 10431 9411
rect 11501 9377 11535 9411
rect 13709 9377 13743 9411
rect 17021 9377 17055 9411
rect 19229 9377 19263 9411
rect 3129 9309 3163 9343
rect 4233 9309 4267 9343
rect 5337 9309 5371 9343
rect 6452 9309 6486 9343
rect 7545 9309 7579 9343
rect 8660 9309 8694 9343
rect 9753 9309 9787 9343
rect 10857 9309 10891 9343
rect 11961 9309 11995 9343
rect 13065 9309 13099 9343
rect 14180 9309 14214 9343
rect 15273 9309 15307 9343
rect 16377 9309 16411 9343
rect 17481 9309 17515 9343
rect 18585 9309 18619 9343
rect 19689 9309 19723 9343
rect 2393 9241 2427 9275
rect 3773 9241 3807 9275
rect 4877 9241 4911 9275
rect 7085 9241 7119 9275
rect 9293 9241 9327 9275
rect 12605 9241 12639 9275
rect 14813 9241 14847 9275
rect 15917 9241 15951 9275
rect 18125 9241 18159 9275
rect 20333 9241 20367 9275
rect 1933 9173 1967 9207
rect 2301 9173 2335 9207
rect 20333 8969 20367 9003
rect 3129 8833 3163 8867
rect 3773 8833 3807 8867
rect 4233 8833 4267 8867
rect 4877 8833 4911 8867
rect 5337 8833 5371 8867
rect 5981 8833 6015 8867
rect 6441 8833 6475 8867
rect 7085 8833 7119 8867
rect 7545 8833 7579 8867
rect 8189 8833 8223 8867
rect 8649 8833 8683 8867
rect 9293 8833 9327 8867
rect 9753 8833 9787 8867
rect 10397 8833 10431 8867
rect 10857 8833 10891 8867
rect 11501 8833 11535 8867
rect 11961 8833 11995 8867
rect 12605 8833 12639 8867
rect 13065 8833 13099 8867
rect 13709 8833 13743 8867
rect 14169 8833 14203 8867
rect 14813 8833 14847 8867
rect 15273 8833 15307 8867
rect 15917 8833 15951 8867
rect 16377 8833 16411 8867
rect 17021 8833 17055 8867
rect 17481 8833 17515 8867
rect 18125 8833 18159 8867
rect 18585 8833 18619 8867
rect 19229 8833 19263 8867
rect 19689 8833 19723 8867
rect 3773 8425 3807 8459
rect 4877 8289 4911 8323
rect 7085 8289 7119 8323
rect 9293 8289 9327 8323
rect 10397 8289 10431 8323
rect 11501 8289 11535 8323
rect 13709 8289 13743 8323
rect 15917 8289 15951 8323
rect 18125 8289 18159 8323
rect 20333 8289 20367 8323
rect 3129 8221 3163 8255
rect 4233 8221 4267 8255
rect 5337 8221 5371 8255
rect 6452 8221 6486 8255
rect 7545 8221 7579 8255
rect 8660 8221 8694 8255
rect 9753 8221 9787 8255
rect 10857 8221 10891 8255
rect 11961 8221 11995 8255
rect 13065 8221 13099 8255
rect 14180 8221 14214 8255
rect 15273 8221 15307 8255
rect 16377 8221 16411 8255
rect 17481 8221 17515 8255
rect 18585 8221 18619 8255
rect 19689 8221 19723 8255
rect 5981 8153 6015 8187
rect 8189 8153 8223 8187
rect 12605 8153 12639 8187
rect 14813 8153 14847 8187
rect 17021 8153 17055 8187
rect 19229 8153 19263 8187
rect 20333 7881 20367 7915
rect 3129 7745 3163 7779
rect 3773 7745 3807 7779
rect 4233 7745 4267 7779
rect 4877 7745 4911 7779
rect 5337 7745 5371 7779
rect 5981 7745 6015 7779
rect 6441 7745 6475 7779
rect 7085 7745 7119 7779
rect 7545 7745 7579 7779
rect 8189 7745 8223 7779
rect 8649 7745 8683 7779
rect 9293 7745 9327 7779
rect 9753 7745 9787 7779
rect 10397 7745 10431 7779
rect 10857 7745 10891 7779
rect 11501 7745 11535 7779
rect 11961 7745 11995 7779
rect 12605 7745 12639 7779
rect 13065 7745 13099 7779
rect 13709 7745 13743 7779
rect 14169 7745 14203 7779
rect 14813 7745 14847 7779
rect 15273 7745 15307 7779
rect 15917 7745 15951 7779
rect 16377 7745 16411 7779
rect 17021 7745 17055 7779
rect 17481 7745 17515 7779
rect 18125 7745 18159 7779
rect 18585 7745 18619 7779
rect 19229 7745 19263 7779
rect 19689 7745 19723 7779
rect 3129 7133 3163 7167
rect 3773 7133 3807 7167
rect 4233 7133 4267 7167
rect 5337 7133 5371 7167
rect 6452 7133 6486 7167
rect 7545 7133 7579 7167
rect 8660 7133 8694 7167
rect 9293 7133 9327 7167
rect 9753 7133 9787 7167
rect 10857 7133 10891 7167
rect 11961 7133 11995 7167
rect 13065 7133 13099 7167
rect 14180 7133 14214 7167
rect 15273 7133 15307 7167
rect 16377 7133 16411 7167
rect 17481 7133 17515 7167
rect 18585 7133 18619 7167
rect 19689 7133 19723 7167
rect 4877 7065 4911 7099
rect 7085 7065 7119 7099
rect 11501 7065 11535 7099
rect 13709 7065 13743 7099
rect 15917 7065 15951 7099
rect 18125 7065 18159 7099
rect 20333 7065 20367 7099
rect 5981 6997 6015 7031
rect 8189 6997 8223 7031
rect 10397 6997 10431 7031
rect 12605 6997 12639 7031
rect 14813 6997 14847 7031
rect 17021 6997 17055 7031
rect 19229 6997 19263 7031
rect 20333 6793 20367 6827
rect 3129 6657 3163 6691
rect 3773 6657 3807 6691
rect 4233 6657 4267 6691
rect 4877 6657 4911 6691
rect 5337 6657 5371 6691
rect 5981 6657 6015 6691
rect 6441 6657 6475 6691
rect 7085 6657 7119 6691
rect 7545 6657 7579 6691
rect 8189 6657 8223 6691
rect 8649 6657 8683 6691
rect 9293 6657 9327 6691
rect 9753 6657 9787 6691
rect 10397 6657 10431 6691
rect 10857 6657 10891 6691
rect 11501 6657 11535 6691
rect 11961 6657 11995 6691
rect 12605 6657 12639 6691
rect 13065 6657 13099 6691
rect 13709 6657 13743 6691
rect 14169 6657 14203 6691
rect 14813 6657 14847 6691
rect 15273 6657 15307 6691
rect 15917 6657 15951 6691
rect 16377 6657 16411 6691
rect 17021 6657 17055 6691
rect 17481 6657 17515 6691
rect 18125 6657 18159 6691
rect 18585 6657 18619 6691
rect 19229 6657 19263 6691
rect 19689 6657 19723 6691
rect 3773 6249 3807 6283
rect 7085 6113 7119 6147
rect 9293 6113 9327 6147
rect 10397 6113 10431 6147
rect 11501 6113 11535 6147
rect 13709 6113 13743 6147
rect 15917 6113 15951 6147
rect 18125 6113 18159 6147
rect 20333 6113 20367 6147
rect 3129 6045 3163 6079
rect 4244 6045 4278 6079
rect 5337 6045 5371 6079
rect 6441 6045 6475 6079
rect 7545 6045 7579 6079
rect 8660 6045 8694 6079
rect 9753 6045 9787 6079
rect 10857 6045 10891 6079
rect 11961 6045 11995 6079
rect 13065 6045 13099 6079
rect 14180 6045 14214 6079
rect 15273 6045 15307 6079
rect 16377 6045 16411 6079
rect 17481 6045 17515 6079
rect 18585 6045 18619 6079
rect 19689 6045 19723 6079
rect 4877 5977 4911 6011
rect 5981 5977 6015 6011
rect 8189 5977 8223 6011
rect 12605 5977 12639 6011
rect 14813 5977 14847 6011
rect 17021 5977 17055 6011
rect 19229 5977 19263 6011
rect 20333 5705 20367 5739
rect 3129 5569 3163 5603
rect 3773 5569 3807 5603
rect 4233 5569 4267 5603
rect 4877 5569 4911 5603
rect 5337 5569 5371 5603
rect 5981 5569 6015 5603
rect 6441 5569 6475 5603
rect 7085 5569 7119 5603
rect 7545 5569 7579 5603
rect 8189 5569 8223 5603
rect 8649 5569 8683 5603
rect 9293 5569 9327 5603
rect 9753 5569 9787 5603
rect 10397 5569 10431 5603
rect 10857 5569 10891 5603
rect 11501 5569 11535 5603
rect 11961 5569 11995 5603
rect 12605 5569 12639 5603
rect 13065 5569 13099 5603
rect 13709 5569 13743 5603
rect 14169 5569 14203 5603
rect 14813 5569 14847 5603
rect 15273 5569 15307 5603
rect 15917 5569 15951 5603
rect 16377 5569 16411 5603
rect 17021 5569 17055 5603
rect 17481 5569 17515 5603
rect 18125 5569 18159 5603
rect 18585 5569 18619 5603
rect 19229 5569 19263 5603
rect 19689 5569 19723 5603
rect 3129 4957 3163 4991
rect 3773 4957 3807 4991
rect 4233 4957 4267 4991
rect 5337 4957 5371 4991
rect 6441 4957 6475 4991
rect 7545 4957 7579 4991
rect 8649 4957 8683 4991
rect 9753 4957 9787 4991
rect 10857 4957 10891 4991
rect 11961 4957 11995 4991
rect 13065 4957 13099 4991
rect 14180 4957 14214 4991
rect 15273 4957 15307 4991
rect 16377 4957 16411 4991
rect 17481 4957 17515 4991
rect 18585 4957 18619 4991
rect 19689 4957 19723 4991
rect 7085 4889 7119 4923
rect 9293 4889 9327 4923
rect 11501 4889 11535 4923
rect 13709 4889 13743 4923
rect 15917 4889 15951 4923
rect 18125 4889 18159 4923
rect 20333 4889 20367 4923
rect 4877 4821 4911 4855
rect 5981 4821 6015 4855
rect 8189 4821 8223 4855
rect 10397 4821 10431 4855
rect 12605 4821 12639 4855
rect 14813 4821 14847 4855
rect 17021 4821 17055 4855
rect 19229 4821 19263 4855
rect 20333 4617 20367 4651
rect 3129 4481 3163 4515
rect 3773 4481 3807 4515
rect 4233 4481 4267 4515
rect 4877 4481 4911 4515
rect 5337 4481 5371 4515
rect 5981 4481 6015 4515
rect 6441 4481 6475 4515
rect 7085 4481 7119 4515
rect 7545 4481 7579 4515
rect 8189 4481 8223 4515
rect 8649 4481 8683 4515
rect 9293 4481 9327 4515
rect 9753 4481 9787 4515
rect 10397 4481 10431 4515
rect 10857 4481 10891 4515
rect 11501 4481 11535 4515
rect 11961 4481 11995 4515
rect 12605 4481 12639 4515
rect 13065 4481 13099 4515
rect 13709 4481 13743 4515
rect 14169 4481 14203 4515
rect 14813 4481 14847 4515
rect 15273 4481 15307 4515
rect 15917 4481 15951 4515
rect 16377 4481 16411 4515
rect 17021 4481 17055 4515
rect 17481 4481 17515 4515
rect 18125 4481 18159 4515
rect 18585 4481 18619 4515
rect 19229 4481 19263 4515
rect 19689 4481 19723 4515
rect 3773 4073 3807 4107
rect 7085 3937 7119 3971
rect 9293 3937 9327 3971
rect 10397 3937 10431 3971
rect 11501 3937 11535 3971
rect 13709 3937 13743 3971
rect 15917 3937 15951 3971
rect 18125 3937 18159 3971
rect 20333 3937 20367 3971
rect 3129 3869 3163 3903
rect 4244 3869 4278 3903
rect 5337 3869 5371 3903
rect 6441 3869 6475 3903
rect 7545 3869 7579 3903
rect 8660 3869 8694 3903
rect 9753 3869 9787 3903
rect 10857 3869 10891 3903
rect 11961 3869 11995 3903
rect 13065 3869 13099 3903
rect 14180 3869 14214 3903
rect 15273 3869 15307 3903
rect 16377 3869 16411 3903
rect 17481 3869 17515 3903
rect 18585 3869 18619 3903
rect 19689 3869 19723 3903
rect 4877 3801 4911 3835
rect 5981 3801 6015 3835
rect 8189 3801 8223 3835
rect 12605 3801 12639 3835
rect 14813 3801 14847 3835
rect 17021 3801 17055 3835
rect 19229 3801 19263 3835
rect 20333 3461 20367 3495
rect 3129 3393 3163 3427
rect 3773 3393 3807 3427
rect 4233 3393 4267 3427
rect 4877 3393 4911 3427
rect 5337 3393 5371 3427
rect 5981 3393 6015 3427
rect 6441 3393 6475 3427
rect 7085 3393 7119 3427
rect 7545 3393 7579 3427
rect 8189 3393 8223 3427
rect 8649 3393 8683 3427
rect 9293 3393 9327 3427
rect 9753 3393 9787 3427
rect 10397 3393 10431 3427
rect 10857 3393 10891 3427
rect 11501 3393 11535 3427
rect 11961 3393 11995 3427
rect 12605 3393 12639 3427
rect 13065 3393 13099 3427
rect 13709 3393 13743 3427
rect 14169 3393 14203 3427
rect 14813 3393 14847 3427
rect 15273 3393 15307 3427
rect 15917 3393 15951 3427
rect 16377 3393 16411 3427
rect 17021 3393 17055 3427
rect 17481 3393 17515 3427
rect 18125 3393 18159 3427
rect 18585 3393 18619 3427
rect 19229 3393 19263 3427
rect 19689 3393 19723 3427
rect 3773 2985 3807 3019
rect 5981 2849 6015 2883
rect 8189 2849 8223 2883
rect 10397 2849 10431 2883
rect 12605 2849 12639 2883
rect 14813 2849 14847 2883
rect 17021 2849 17055 2883
rect 19229 2849 19263 2883
rect 3129 2781 3163 2815
rect 4244 2781 4278 2815
rect 5337 2781 5371 2815
rect 6441 2781 6475 2815
rect 7545 2781 7579 2815
rect 8660 2781 8694 2815
rect 9753 2781 9787 2815
rect 10857 2781 10891 2815
rect 11961 2781 11995 2815
rect 13065 2781 13099 2815
rect 14169 2781 14203 2815
rect 15273 2781 15307 2815
rect 16377 2781 16411 2815
rect 17481 2781 17515 2815
rect 18585 2781 18619 2815
rect 19689 2781 19723 2815
rect 4877 2713 4911 2747
rect 7085 2713 7119 2747
rect 9293 2713 9327 2747
rect 11501 2713 11535 2747
rect 13709 2713 13743 2747
rect 18125 2713 18159 2747
rect 20333 2713 20367 2747
rect 15917 2645 15951 2679
rect 20333 2441 20367 2475
rect 3129 2305 3163 2339
rect 3773 2305 3807 2339
rect 4233 2305 4267 2339
rect 4877 2305 4911 2339
rect 5337 2305 5371 2339
rect 5981 2305 6015 2339
rect 6441 2305 6475 2339
rect 7085 2305 7119 2339
rect 7545 2305 7579 2339
rect 8189 2305 8223 2339
rect 8649 2305 8683 2339
rect 9293 2305 9327 2339
rect 9753 2305 9787 2339
rect 10397 2305 10431 2339
rect 10857 2305 10891 2339
rect 11501 2305 11535 2339
rect 11961 2305 11995 2339
rect 12605 2305 12639 2339
rect 13065 2305 13099 2339
rect 13709 2305 13743 2339
rect 14169 2305 14203 2339
rect 14813 2305 14847 2339
rect 15273 2305 15307 2339
rect 15917 2305 15951 2339
rect 16377 2305 16411 2339
rect 17021 2305 17055 2339
rect 17481 2305 17515 2339
rect 18125 2305 18159 2339
rect 18585 2305 18619 2339
rect 19229 2305 19263 2339
rect 19689 2305 19723 2339
rect 3773 1897 3807 1931
rect 7085 1761 7119 1795
rect 9293 1761 9327 1795
rect 10397 1761 10431 1795
rect 11501 1761 11535 1795
rect 13709 1761 13743 1795
rect 15917 1761 15951 1795
rect 18125 1761 18159 1795
rect 20333 1761 20367 1795
rect 3129 1693 3163 1727
rect 4244 1693 4278 1727
rect 5337 1693 5371 1727
rect 6441 1693 6475 1727
rect 7545 1693 7579 1727
rect 8660 1693 8694 1727
rect 9753 1693 9787 1727
rect 10857 1693 10891 1727
rect 11961 1693 11995 1727
rect 13065 1693 13099 1727
rect 14180 1693 14214 1727
rect 15273 1693 15307 1727
rect 16377 1693 16411 1727
rect 17481 1693 17515 1727
rect 18585 1693 18619 1727
rect 19689 1693 19723 1727
rect 4877 1625 4911 1659
rect 5981 1625 6015 1659
rect 8189 1625 8223 1659
rect 12605 1625 12639 1659
rect 14813 1625 14847 1659
rect 17021 1625 17055 1659
rect 19229 1625 19263 1659
rect 20333 1353 20367 1387
rect 3129 1217 3163 1251
rect 3773 1217 3807 1251
rect 4233 1217 4267 1251
rect 4877 1217 4911 1251
rect 5337 1217 5371 1251
rect 5981 1217 6015 1251
rect 6441 1217 6475 1251
rect 7085 1217 7119 1251
rect 7545 1217 7579 1251
rect 8189 1217 8223 1251
rect 8649 1217 8683 1251
rect 9293 1217 9327 1251
rect 9753 1217 9787 1251
rect 10397 1217 10431 1251
rect 10857 1217 10891 1251
rect 11501 1217 11535 1251
rect 11961 1217 11995 1251
rect 12605 1217 12639 1251
rect 13065 1217 13099 1251
rect 13709 1217 13743 1251
rect 14169 1217 14203 1251
rect 14813 1217 14847 1251
rect 15273 1217 15307 1251
rect 15917 1217 15951 1251
rect 16377 1217 16411 1251
rect 17021 1217 17055 1251
rect 17481 1217 17515 1251
rect 18125 1217 18159 1251
rect 18585 1217 18619 1251
rect 19229 1217 19263 1251
rect 19689 1217 19723 1251
<< metal1 >>
rect 1904 22170 20764 22192
rect 1904 22118 4446 22170
rect 4498 22118 4510 22170
rect 4562 22118 4574 22170
rect 4626 22118 4638 22170
rect 4690 22118 9774 22170
rect 9826 22118 9838 22170
rect 9890 22118 9902 22170
rect 9954 22118 9966 22170
rect 10018 22118 15102 22170
rect 15154 22118 15166 22170
rect 15218 22118 15230 22170
rect 15282 22118 15294 22170
rect 15346 22118 20764 22170
rect 1904 22096 20764 22118
rect 1918 22056 1924 22068
rect 1879 22028 1924 22056
rect 1918 22016 1924 22028
rect 1976 22016 1982 22068
rect 2286 21988 2292 22000
rect 2247 21960 2292 21988
rect 2286 21948 2292 21960
rect 2344 21988 2350 22000
rect 2344 21960 2608 21988
rect 2344 21948 2350 21960
rect 2381 21923 2439 21929
rect 2381 21920 2393 21923
rect 2304 21892 2393 21920
rect 2304 21784 2332 21892
rect 2381 21889 2393 21892
rect 2427 21889 2439 21923
rect 2580 21920 2608 21960
rect 3117 21923 3175 21929
rect 3117 21920 3129 21923
rect 2580 21892 3129 21920
rect 2381 21883 2439 21889
rect 3117 21889 3129 21892
rect 3163 21889 3175 21923
rect 3117 21883 3175 21889
rect 2470 21852 2476 21864
rect 2431 21824 2476 21852
rect 2470 21812 2476 21824
rect 2528 21812 2534 21864
rect 3761 21787 3819 21793
rect 3761 21784 3773 21787
rect 2304 21756 3773 21784
rect 3761 21753 3773 21756
rect 3807 21753 3819 21787
rect 3761 21747 3819 21753
rect 1904 21626 20764 21648
rect 1904 21574 7110 21626
rect 7162 21574 7174 21626
rect 7226 21574 7238 21626
rect 7290 21574 7302 21626
rect 7354 21574 12438 21626
rect 12490 21574 12502 21626
rect 12554 21574 12566 21626
rect 12618 21574 12630 21626
rect 12682 21574 17766 21626
rect 17818 21574 17830 21626
rect 17882 21574 17894 21626
rect 17946 21574 17958 21626
rect 18010 21574 20764 21626
rect 1904 21552 20764 21574
rect 1921 21515 1979 21521
rect 1921 21481 1933 21515
rect 1967 21512 1979 21515
rect 2286 21512 2292 21524
rect 1967 21484 2292 21512
rect 1967 21481 1979 21484
rect 1921 21475 1979 21481
rect 2286 21472 2292 21484
rect 2344 21472 2350 21524
rect 2470 21376 2476 21388
rect 2431 21348 2476 21376
rect 2470 21336 2476 21348
rect 2528 21336 2534 21388
rect 2381 21311 2439 21317
rect 2381 21277 2393 21311
rect 2427 21308 2439 21311
rect 3117 21311 3175 21317
rect 2427 21280 2792 21308
rect 2427 21277 2439 21280
rect 2381 21271 2439 21277
rect 2286 21200 2292 21252
rect 2344 21240 2350 21252
rect 2764 21240 2792 21280
rect 3117 21277 3129 21311
rect 3163 21308 3175 21311
rect 3850 21308 3856 21320
rect 3163 21280 3856 21308
rect 3163 21277 3175 21280
rect 3117 21271 3175 21277
rect 3850 21268 3856 21280
rect 3908 21268 3914 21320
rect 3761 21243 3819 21249
rect 3761 21240 3773 21243
rect 2344 21212 2389 21240
rect 2764 21212 3773 21240
rect 2344 21200 2350 21212
rect 3761 21209 3773 21212
rect 3807 21209 3819 21243
rect 3761 21203 3819 21209
rect 1904 21082 20764 21104
rect 1904 21030 4446 21082
rect 4498 21030 4510 21082
rect 4562 21030 4574 21082
rect 4626 21030 4638 21082
rect 4690 21030 9774 21082
rect 9826 21030 9838 21082
rect 9890 21030 9902 21082
rect 9954 21030 9966 21082
rect 10018 21030 15102 21082
rect 15154 21030 15166 21082
rect 15218 21030 15230 21082
rect 15282 21030 15294 21082
rect 15346 21030 20764 21082
rect 1904 21008 20764 21030
rect 3761 20971 3819 20977
rect 3761 20937 3773 20971
rect 3807 20968 3819 20971
rect 3850 20968 3856 20980
rect 3807 20940 3856 20968
rect 3807 20937 3819 20940
rect 3761 20931 3819 20937
rect 3850 20928 3856 20940
rect 3908 20928 3914 20980
rect 2286 20792 2292 20844
rect 2344 20832 2350 20844
rect 3117 20835 3175 20841
rect 3117 20832 3129 20835
rect 2344 20804 3129 20832
rect 2344 20792 2350 20804
rect 3117 20801 3129 20804
rect 3163 20801 3175 20835
rect 3117 20795 3175 20801
rect 1904 20538 20764 20560
rect 1904 20486 7110 20538
rect 7162 20486 7174 20538
rect 7226 20486 7238 20538
rect 7290 20486 7302 20538
rect 7354 20486 12438 20538
rect 12490 20486 12502 20538
rect 12554 20486 12566 20538
rect 12618 20486 12630 20538
rect 12682 20486 17766 20538
rect 17818 20486 17830 20538
rect 17882 20486 17894 20538
rect 17946 20486 17958 20538
rect 18010 20486 20764 20538
rect 1904 20464 20764 20486
rect 1921 20427 1979 20433
rect 1921 20393 1933 20427
rect 1967 20424 1979 20427
rect 2286 20424 2292 20436
rect 1967 20396 2292 20424
rect 1967 20393 1979 20396
rect 1921 20387 1979 20393
rect 2286 20384 2292 20396
rect 2344 20384 2350 20436
rect 2470 20288 2476 20300
rect 2431 20260 2476 20288
rect 2470 20248 2476 20260
rect 2528 20248 2534 20300
rect 4865 20291 4923 20297
rect 4865 20288 4877 20291
rect 3132 20260 4877 20288
rect 3132 20229 3160 20260
rect 4865 20257 4877 20260
rect 4911 20257 4923 20291
rect 4865 20251 4923 20257
rect 2381 20223 2439 20229
rect 2381 20189 2393 20223
rect 2427 20189 2439 20223
rect 2381 20183 2439 20189
rect 3117 20223 3175 20229
rect 3117 20189 3129 20223
rect 3163 20189 3175 20223
rect 4218 20220 4224 20232
rect 4179 20192 4224 20220
rect 3117 20183 3175 20189
rect 2396 20152 2424 20183
rect 4218 20180 4224 20192
rect 4276 20180 4282 20232
rect 3761 20155 3819 20161
rect 3761 20152 3773 20155
rect 2396 20124 3773 20152
rect 3761 20121 3773 20124
rect 3807 20121 3819 20155
rect 3761 20115 3819 20121
rect 2286 20044 2292 20096
rect 2344 20084 2350 20096
rect 2344 20056 2389 20084
rect 2344 20044 2350 20056
rect 1904 19994 20764 20016
rect 1904 19942 4446 19994
rect 4498 19942 4510 19994
rect 4562 19942 4574 19994
rect 4626 19942 4638 19994
rect 4690 19942 9774 19994
rect 9826 19942 9838 19994
rect 9890 19942 9902 19994
rect 9954 19942 9966 19994
rect 10018 19942 15102 19994
rect 15154 19942 15166 19994
rect 15218 19942 15230 19994
rect 15282 19942 15294 19994
rect 15346 19942 20764 19994
rect 1904 19920 20764 19942
rect 4218 19840 4224 19892
rect 4276 19880 4282 19892
rect 4865 19883 4923 19889
rect 4865 19880 4877 19883
rect 4276 19852 4877 19880
rect 4276 19840 4282 19852
rect 4865 19849 4877 19852
rect 4911 19849 4923 19883
rect 4865 19843 4923 19849
rect 2286 19704 2292 19756
rect 2344 19744 2350 19756
rect 3117 19747 3175 19753
rect 3117 19744 3129 19747
rect 2344 19716 3129 19744
rect 2344 19704 2350 19716
rect 3117 19713 3129 19716
rect 3163 19713 3175 19747
rect 3117 19707 3175 19713
rect 3761 19747 3819 19753
rect 3761 19713 3773 19747
rect 3807 19744 3819 19747
rect 4221 19747 4279 19753
rect 4221 19744 4233 19747
rect 3807 19716 4233 19744
rect 3807 19713 3819 19716
rect 3761 19707 3819 19713
rect 4221 19713 4233 19716
rect 4267 19713 4279 19747
rect 4221 19707 4279 19713
rect 1904 19450 20764 19472
rect 1904 19398 7110 19450
rect 7162 19398 7174 19450
rect 7226 19398 7238 19450
rect 7290 19398 7302 19450
rect 7354 19398 12438 19450
rect 12490 19398 12502 19450
rect 12554 19398 12566 19450
rect 12618 19398 12630 19450
rect 12682 19398 17766 19450
rect 17818 19398 17830 19450
rect 17882 19398 17894 19450
rect 17946 19398 17958 19450
rect 18010 19398 20764 19450
rect 1904 19376 20764 19398
rect 1921 19339 1979 19345
rect 1921 19305 1933 19339
rect 1967 19336 1979 19339
rect 2286 19336 2292 19348
rect 1967 19308 2292 19336
rect 1967 19305 1979 19308
rect 1921 19299 1979 19305
rect 2286 19296 2292 19308
rect 2344 19296 2350 19348
rect 2470 19200 2476 19212
rect 2431 19172 2476 19200
rect 2470 19160 2476 19172
rect 2528 19160 2534 19212
rect 4865 19203 4923 19209
rect 4865 19200 4877 19203
rect 3132 19172 4877 19200
rect 3132 19141 3160 19172
rect 4865 19169 4877 19172
rect 4911 19169 4923 19203
rect 7073 19203 7131 19209
rect 7073 19200 7085 19203
rect 4865 19163 4923 19169
rect 5340 19172 7085 19200
rect 5340 19141 5368 19172
rect 7073 19169 7085 19172
rect 7119 19169 7131 19203
rect 7073 19163 7131 19169
rect 2381 19135 2439 19141
rect 2381 19101 2393 19135
rect 2427 19101 2439 19135
rect 2381 19095 2439 19101
rect 3117 19135 3175 19141
rect 3117 19101 3129 19135
rect 3163 19101 3175 19135
rect 3117 19095 3175 19101
rect 4221 19135 4279 19141
rect 4221 19101 4233 19135
rect 4267 19101 4279 19135
rect 4221 19095 4279 19101
rect 5325 19135 5383 19141
rect 5325 19101 5337 19135
rect 5371 19101 5383 19135
rect 5325 19095 5383 19101
rect 6429 19135 6487 19141
rect 6429 19101 6441 19135
rect 6475 19132 6487 19135
rect 6978 19132 6984 19144
rect 6475 19104 6984 19132
rect 6475 19101 6487 19104
rect 6429 19095 6487 19101
rect 2396 19064 2424 19095
rect 3761 19067 3819 19073
rect 3761 19064 3773 19067
rect 2396 19036 3773 19064
rect 3761 19033 3773 19036
rect 3807 19033 3819 19067
rect 4236 19064 4264 19095
rect 6978 19092 6984 19104
rect 7036 19092 7042 19144
rect 5969 19067 6027 19073
rect 5969 19064 5981 19067
rect 4236 19036 5981 19064
rect 3761 19027 3819 19033
rect 5969 19033 5981 19036
rect 6015 19033 6027 19067
rect 5969 19027 6027 19033
rect 2286 18956 2292 19008
rect 2344 18996 2350 19008
rect 2344 18968 2389 18996
rect 2344 18956 2350 18968
rect 1904 18906 20764 18928
rect 1904 18854 4446 18906
rect 4498 18854 4510 18906
rect 4562 18854 4574 18906
rect 4626 18854 4638 18906
rect 4690 18854 9774 18906
rect 9826 18854 9838 18906
rect 9890 18854 9902 18906
rect 9954 18854 9966 18906
rect 10018 18854 15102 18906
rect 15154 18854 15166 18906
rect 15218 18854 15230 18906
rect 15282 18854 15294 18906
rect 15346 18854 20764 18906
rect 1904 18832 20764 18854
rect 6978 18752 6984 18804
rect 7036 18792 7042 18804
rect 7073 18795 7131 18801
rect 7073 18792 7085 18795
rect 7036 18764 7085 18792
rect 7036 18752 7042 18764
rect 7073 18761 7085 18764
rect 7119 18761 7131 18795
rect 7073 18755 7131 18761
rect 2286 18616 2292 18668
rect 2344 18656 2350 18668
rect 3117 18659 3175 18665
rect 3117 18656 3129 18659
rect 2344 18628 3129 18656
rect 2344 18616 2350 18628
rect 3117 18625 3129 18628
rect 3163 18625 3175 18659
rect 3117 18619 3175 18625
rect 3761 18659 3819 18665
rect 3761 18625 3773 18659
rect 3807 18656 3819 18659
rect 4221 18659 4279 18665
rect 4221 18656 4233 18659
rect 3807 18628 4233 18656
rect 3807 18625 3819 18628
rect 3761 18619 3819 18625
rect 4221 18625 4233 18628
rect 4267 18625 4279 18659
rect 4221 18619 4279 18625
rect 4865 18659 4923 18665
rect 4865 18625 4877 18659
rect 4911 18656 4923 18659
rect 5325 18659 5383 18665
rect 5325 18656 5337 18659
rect 4911 18628 5337 18656
rect 4911 18625 4923 18628
rect 4865 18619 4923 18625
rect 5325 18625 5337 18628
rect 5371 18625 5383 18659
rect 5325 18619 5383 18625
rect 5969 18659 6027 18665
rect 5969 18625 5981 18659
rect 6015 18656 6027 18659
rect 6429 18659 6487 18665
rect 6429 18656 6441 18659
rect 6015 18628 6441 18656
rect 6015 18625 6027 18628
rect 5969 18619 6027 18625
rect 6429 18625 6441 18628
rect 6475 18625 6487 18659
rect 6429 18619 6487 18625
rect 1904 18362 20764 18384
rect 1904 18310 7110 18362
rect 7162 18310 7174 18362
rect 7226 18310 7238 18362
rect 7290 18310 7302 18362
rect 7354 18310 12438 18362
rect 12490 18310 12502 18362
rect 12554 18310 12566 18362
rect 12618 18310 12630 18362
rect 12682 18310 17766 18362
rect 17818 18310 17830 18362
rect 17882 18310 17894 18362
rect 17946 18310 17958 18362
rect 18010 18310 20764 18362
rect 1904 18288 20764 18310
rect 1921 18251 1979 18257
rect 1921 18217 1933 18251
rect 1967 18248 1979 18251
rect 2286 18248 2292 18260
rect 1967 18220 2292 18248
rect 1967 18217 1979 18220
rect 1921 18211 1979 18217
rect 2286 18208 2292 18220
rect 2344 18208 2350 18260
rect 2470 18112 2476 18124
rect 2431 18084 2476 18112
rect 2470 18072 2476 18084
rect 2528 18072 2534 18124
rect 4865 18115 4923 18121
rect 4865 18112 4877 18115
rect 3132 18084 4877 18112
rect 3132 18053 3160 18084
rect 4865 18081 4877 18084
rect 4911 18081 4923 18115
rect 7073 18115 7131 18121
rect 7073 18112 7085 18115
rect 4865 18075 4923 18081
rect 5340 18084 7085 18112
rect 5340 18053 5368 18084
rect 7073 18081 7085 18084
rect 7119 18081 7131 18115
rect 8177 18115 8235 18121
rect 8177 18112 8189 18115
rect 7073 18075 7131 18081
rect 7364 18084 8189 18112
rect 2381 18047 2439 18053
rect 2381 18013 2393 18047
rect 2427 18013 2439 18047
rect 2381 18007 2439 18013
rect 3117 18047 3175 18053
rect 3117 18013 3129 18047
rect 3163 18013 3175 18047
rect 3117 18007 3175 18013
rect 4221 18047 4279 18053
rect 4221 18013 4233 18047
rect 4267 18013 4279 18047
rect 4221 18007 4279 18013
rect 5325 18047 5383 18053
rect 5325 18013 5337 18047
rect 5371 18013 5383 18047
rect 5325 18007 5383 18013
rect 6440 18047 6498 18053
rect 6440 18013 6452 18047
rect 6486 18013 6498 18047
rect 6440 18007 6498 18013
rect 2396 17976 2424 18007
rect 3761 17979 3819 17985
rect 3761 17976 3773 17979
rect 2396 17948 3773 17976
rect 3761 17945 3773 17948
rect 3807 17945 3819 17979
rect 4236 17976 4264 18007
rect 5969 17979 6027 17985
rect 5969 17976 5981 17979
rect 4236 17948 5981 17976
rect 3761 17939 3819 17945
rect 5969 17945 5981 17948
rect 6015 17945 6027 17979
rect 6444 17976 6472 18007
rect 7364 17976 7392 18084
rect 8177 18081 8189 18084
rect 8223 18081 8235 18115
rect 10385 18115 10443 18121
rect 10385 18112 10397 18115
rect 8177 18075 8235 18081
rect 8663 18084 10397 18112
rect 8663 18053 8691 18084
rect 10385 18081 10397 18084
rect 10431 18081 10443 18115
rect 10385 18075 10443 18081
rect 7533 18047 7591 18053
rect 7533 18013 7545 18047
rect 7579 18013 7591 18047
rect 7533 18007 7591 18013
rect 8648 18047 8706 18053
rect 8648 18013 8660 18047
rect 8694 18013 8706 18047
rect 8648 18007 8706 18013
rect 9741 18047 9799 18053
rect 9741 18013 9753 18047
rect 9787 18013 9799 18047
rect 10842 18044 10848 18056
rect 10803 18016 10848 18044
rect 9741 18007 9799 18013
rect 6444 17948 7392 17976
rect 7548 17976 7576 18007
rect 9281 17979 9339 17985
rect 9281 17976 9293 17979
rect 7548 17948 9293 17976
rect 5969 17939 6027 17945
rect 9281 17945 9293 17948
rect 9327 17945 9339 17979
rect 9756 17976 9784 18007
rect 10842 18004 10848 18016
rect 10900 18004 10906 18056
rect 11489 17979 11547 17985
rect 11489 17976 11501 17979
rect 9756 17948 11501 17976
rect 9281 17939 9339 17945
rect 11489 17945 11501 17948
rect 11535 17945 11547 17979
rect 11489 17939 11547 17945
rect 2286 17868 2292 17920
rect 2344 17908 2350 17920
rect 2344 17880 2389 17908
rect 2344 17868 2350 17880
rect 1904 17818 20764 17840
rect 1904 17766 4446 17818
rect 4498 17766 4510 17818
rect 4562 17766 4574 17818
rect 4626 17766 4638 17818
rect 4690 17766 9774 17818
rect 9826 17766 9838 17818
rect 9890 17766 9902 17818
rect 9954 17766 9966 17818
rect 10018 17766 15102 17818
rect 15154 17766 15166 17818
rect 15218 17766 15230 17818
rect 15282 17766 15294 17818
rect 15346 17766 20764 17818
rect 1904 17744 20764 17766
rect 10842 17664 10848 17716
rect 10900 17704 10906 17716
rect 11489 17707 11547 17713
rect 11489 17704 11501 17707
rect 10900 17676 11501 17704
rect 10900 17664 10906 17676
rect 11489 17673 11501 17676
rect 11535 17673 11547 17707
rect 11489 17667 11547 17673
rect 2286 17528 2292 17580
rect 2344 17568 2350 17580
rect 3117 17571 3175 17577
rect 3117 17568 3129 17571
rect 2344 17540 3129 17568
rect 2344 17528 2350 17540
rect 3117 17537 3129 17540
rect 3163 17537 3175 17571
rect 3117 17531 3175 17537
rect 3761 17571 3819 17577
rect 3761 17537 3773 17571
rect 3807 17568 3819 17571
rect 4221 17571 4279 17577
rect 4221 17568 4233 17571
rect 3807 17540 4233 17568
rect 3807 17537 3819 17540
rect 3761 17531 3819 17537
rect 4221 17537 4233 17540
rect 4267 17537 4279 17571
rect 4221 17531 4279 17537
rect 4865 17571 4923 17577
rect 4865 17537 4877 17571
rect 4911 17568 4923 17571
rect 5325 17571 5383 17577
rect 5325 17568 5337 17571
rect 4911 17540 5337 17568
rect 4911 17537 4923 17540
rect 4865 17531 4923 17537
rect 5325 17537 5337 17540
rect 5371 17537 5383 17571
rect 5325 17531 5383 17537
rect 5969 17571 6027 17577
rect 5969 17537 5981 17571
rect 6015 17568 6027 17571
rect 6429 17571 6487 17577
rect 6429 17568 6441 17571
rect 6015 17540 6441 17568
rect 6015 17537 6027 17540
rect 5969 17531 6027 17537
rect 6429 17537 6441 17540
rect 6475 17537 6487 17571
rect 6429 17531 6487 17537
rect 7073 17571 7131 17577
rect 7073 17537 7085 17571
rect 7119 17568 7131 17571
rect 7533 17571 7591 17577
rect 7533 17568 7545 17571
rect 7119 17540 7545 17568
rect 7119 17537 7131 17540
rect 7073 17531 7131 17537
rect 7533 17537 7545 17540
rect 7579 17537 7591 17571
rect 7533 17531 7591 17537
rect 8177 17571 8235 17577
rect 8177 17537 8189 17571
rect 8223 17568 8235 17571
rect 8637 17571 8695 17577
rect 8637 17568 8649 17571
rect 8223 17540 8649 17568
rect 8223 17537 8235 17540
rect 8177 17531 8235 17537
rect 8637 17537 8649 17540
rect 8683 17537 8695 17571
rect 8637 17531 8695 17537
rect 9281 17571 9339 17577
rect 9281 17537 9293 17571
rect 9327 17568 9339 17571
rect 9741 17571 9799 17577
rect 9741 17568 9753 17571
rect 9327 17540 9753 17568
rect 9327 17537 9339 17540
rect 9281 17531 9339 17537
rect 9741 17537 9753 17540
rect 9787 17537 9799 17571
rect 9741 17531 9799 17537
rect 10385 17571 10443 17577
rect 10385 17537 10397 17571
rect 10431 17568 10443 17571
rect 10845 17571 10903 17577
rect 10845 17568 10857 17571
rect 10431 17540 10857 17568
rect 10431 17537 10443 17540
rect 10385 17531 10443 17537
rect 10845 17537 10857 17540
rect 10891 17537 10903 17571
rect 10845 17531 10903 17537
rect 1904 17274 20764 17296
rect 1904 17222 7110 17274
rect 7162 17222 7174 17274
rect 7226 17222 7238 17274
rect 7290 17222 7302 17274
rect 7354 17222 12438 17274
rect 12490 17222 12502 17274
rect 12554 17222 12566 17274
rect 12618 17222 12630 17274
rect 12682 17222 17766 17274
rect 17818 17222 17830 17274
rect 17882 17222 17894 17274
rect 17946 17222 17958 17274
rect 18010 17222 20764 17274
rect 1904 17200 20764 17222
rect 1921 17163 1979 17169
rect 1921 17129 1933 17163
rect 1967 17160 1979 17163
rect 2286 17160 2292 17172
rect 1967 17132 2292 17160
rect 1967 17129 1979 17132
rect 1921 17123 1979 17129
rect 2286 17120 2292 17132
rect 2344 17120 2350 17172
rect 2470 17024 2476 17036
rect 2431 16996 2476 17024
rect 2470 16984 2476 16996
rect 2528 16984 2534 17036
rect 4865 17027 4923 17033
rect 4865 17024 4877 17027
rect 3132 16996 4877 17024
rect 3132 16965 3160 16996
rect 4865 16993 4877 16996
rect 4911 16993 4923 17027
rect 7073 17027 7131 17033
rect 7073 17024 7085 17027
rect 4865 16987 4923 16993
rect 5340 16996 7085 17024
rect 5340 16965 5368 16996
rect 7073 16993 7085 16996
rect 7119 16993 7131 17027
rect 8177 17027 8235 17033
rect 8177 17024 8189 17027
rect 7073 16987 7131 16993
rect 7364 16996 8189 17024
rect 3117 16959 3175 16965
rect 3117 16925 3129 16959
rect 3163 16925 3175 16959
rect 3117 16919 3175 16925
rect 4221 16959 4279 16965
rect 4221 16925 4233 16959
rect 4267 16925 4279 16959
rect 4221 16919 4279 16925
rect 5325 16959 5383 16965
rect 5325 16925 5337 16959
rect 5371 16925 5383 16959
rect 5325 16919 5383 16925
rect 6440 16959 6498 16965
rect 6440 16925 6452 16959
rect 6486 16925 6498 16959
rect 6440 16919 6498 16925
rect 2381 16891 2439 16897
rect 2381 16857 2393 16891
rect 2427 16888 2439 16891
rect 3761 16891 3819 16897
rect 3761 16888 3773 16891
rect 2427 16860 3773 16888
rect 2427 16857 2439 16860
rect 2381 16851 2439 16857
rect 3761 16857 3773 16860
rect 3807 16857 3819 16891
rect 4236 16888 4264 16919
rect 5969 16891 6027 16897
rect 5969 16888 5981 16891
rect 4236 16860 5981 16888
rect 3761 16851 3819 16857
rect 5969 16857 5981 16860
rect 6015 16857 6027 16891
rect 6444 16888 6472 16919
rect 7364 16888 7392 16996
rect 8177 16993 8189 16996
rect 8223 16993 8235 17027
rect 10385 17027 10443 17033
rect 10385 17024 10397 17027
rect 8177 16987 8235 16993
rect 8663 16996 10397 17024
rect 8663 16965 8691 16996
rect 10385 16993 10397 16996
rect 10431 16993 10443 17027
rect 11489 17027 11547 17033
rect 11489 17024 11501 17027
rect 10385 16987 10443 16993
rect 10584 16996 11501 17024
rect 7533 16959 7591 16965
rect 7533 16925 7545 16959
rect 7579 16925 7591 16959
rect 7533 16919 7591 16925
rect 8648 16959 8706 16965
rect 8648 16925 8660 16959
rect 8694 16925 8706 16959
rect 8648 16919 8706 16925
rect 9741 16959 9799 16965
rect 9741 16925 9753 16959
rect 9787 16956 9799 16959
rect 10584 16956 10612 16996
rect 11489 16993 11501 16996
rect 11535 16993 11547 17027
rect 13697 17027 13755 17033
rect 13697 17024 13709 17027
rect 11489 16987 11547 16993
rect 11964 16996 13709 17024
rect 11964 16965 11992 16996
rect 13697 16993 13709 16996
rect 13743 16993 13755 17027
rect 15905 17027 15963 17033
rect 15905 17024 15917 17027
rect 13697 16987 13755 16993
rect 14183 16996 15917 17024
rect 14183 16965 14211 16996
rect 15905 16993 15917 16996
rect 15951 16993 15963 17027
rect 18113 17027 18171 17033
rect 18113 17024 18125 17027
rect 15905 16987 15963 16993
rect 16380 16996 18125 17024
rect 16380 16965 16408 16996
rect 18113 16993 18125 16996
rect 18159 16993 18171 17027
rect 20321 17027 20379 17033
rect 20321 17024 20333 17027
rect 18113 16987 18171 16993
rect 18588 16996 20333 17024
rect 18588 16965 18616 16996
rect 20321 16993 20333 16996
rect 20367 16993 20379 17027
rect 20321 16987 20379 16993
rect 9787 16928 10612 16956
rect 10845 16959 10903 16965
rect 9787 16925 9799 16928
rect 9741 16919 9799 16925
rect 10845 16925 10857 16959
rect 10891 16925 10903 16959
rect 10845 16919 10903 16925
rect 11949 16959 12007 16965
rect 11949 16925 11961 16959
rect 11995 16925 12007 16959
rect 11949 16919 12007 16925
rect 13053 16959 13111 16965
rect 13053 16925 13065 16959
rect 13099 16925 13111 16959
rect 13053 16919 13111 16925
rect 14168 16959 14226 16965
rect 14168 16925 14180 16959
rect 14214 16925 14226 16959
rect 14168 16919 14226 16925
rect 15261 16959 15319 16965
rect 15261 16925 15273 16959
rect 15307 16925 15319 16959
rect 15261 16919 15319 16925
rect 16365 16959 16423 16965
rect 16365 16925 16377 16959
rect 16411 16925 16423 16959
rect 16365 16919 16423 16925
rect 17469 16959 17527 16965
rect 17469 16925 17481 16959
rect 17515 16925 17527 16959
rect 17469 16919 17527 16925
rect 18573 16959 18631 16965
rect 18573 16925 18585 16959
rect 18619 16925 18631 16959
rect 18573 16919 18631 16925
rect 19677 16959 19735 16965
rect 19677 16925 19689 16959
rect 19723 16956 19735 16959
rect 20134 16956 20140 16968
rect 19723 16928 20140 16956
rect 19723 16925 19735 16928
rect 19677 16919 19735 16925
rect 6444 16860 7392 16888
rect 7548 16888 7576 16919
rect 9281 16891 9339 16897
rect 9281 16888 9293 16891
rect 7548 16860 9293 16888
rect 5969 16851 6027 16857
rect 9281 16857 9293 16860
rect 9327 16857 9339 16891
rect 10860 16888 10888 16919
rect 12593 16891 12651 16897
rect 12593 16888 12605 16891
rect 10860 16860 12605 16888
rect 9281 16851 9339 16857
rect 12593 16857 12605 16860
rect 12639 16857 12651 16891
rect 13068 16888 13096 16919
rect 14801 16891 14859 16897
rect 14801 16888 14813 16891
rect 13068 16860 14813 16888
rect 12593 16851 12651 16857
rect 14801 16857 14813 16860
rect 14847 16857 14859 16891
rect 15276 16888 15304 16919
rect 17009 16891 17067 16897
rect 17009 16888 17021 16891
rect 15276 16860 17021 16888
rect 14801 16851 14859 16857
rect 17009 16857 17021 16860
rect 17055 16857 17067 16891
rect 17484 16888 17512 16919
rect 20134 16916 20140 16928
rect 20192 16916 20198 16968
rect 19217 16891 19275 16897
rect 19217 16888 19229 16891
rect 17484 16860 19229 16888
rect 17009 16851 17067 16857
rect 19217 16857 19229 16860
rect 19263 16857 19275 16891
rect 19217 16851 19275 16857
rect 2286 16780 2292 16832
rect 2344 16820 2350 16832
rect 2344 16792 2389 16820
rect 2344 16780 2350 16792
rect 1904 16730 20764 16752
rect 1904 16678 4446 16730
rect 4498 16678 4510 16730
rect 4562 16678 4574 16730
rect 4626 16678 4638 16730
rect 4690 16678 9774 16730
rect 9826 16678 9838 16730
rect 9890 16678 9902 16730
rect 9954 16678 9966 16730
rect 10018 16678 15102 16730
rect 15154 16678 15166 16730
rect 15218 16678 15230 16730
rect 15282 16678 15294 16730
rect 15346 16678 20764 16730
rect 1904 16656 20764 16678
rect 20134 16576 20140 16628
rect 20192 16616 20198 16628
rect 20321 16619 20379 16625
rect 20321 16616 20333 16619
rect 20192 16588 20333 16616
rect 20192 16576 20198 16588
rect 20321 16585 20333 16588
rect 20367 16585 20379 16619
rect 20321 16579 20379 16585
rect 2286 16440 2292 16492
rect 2344 16480 2350 16492
rect 2562 16480 2568 16492
rect 2344 16452 2568 16480
rect 2344 16440 2350 16452
rect 2562 16440 2568 16452
rect 2620 16480 2626 16492
rect 3117 16483 3175 16489
rect 3117 16480 3129 16483
rect 2620 16452 3129 16480
rect 2620 16440 2626 16452
rect 3117 16449 3129 16452
rect 3163 16449 3175 16483
rect 3117 16443 3175 16449
rect 3761 16483 3819 16489
rect 3761 16449 3773 16483
rect 3807 16480 3819 16483
rect 4221 16483 4279 16489
rect 4221 16480 4233 16483
rect 3807 16452 4233 16480
rect 3807 16449 3819 16452
rect 3761 16443 3819 16449
rect 4221 16449 4233 16452
rect 4267 16449 4279 16483
rect 4221 16443 4279 16449
rect 4865 16483 4923 16489
rect 4865 16449 4877 16483
rect 4911 16480 4923 16483
rect 5325 16483 5383 16489
rect 5325 16480 5337 16483
rect 4911 16452 5337 16480
rect 4911 16449 4923 16452
rect 4865 16443 4923 16449
rect 5325 16449 5337 16452
rect 5371 16449 5383 16483
rect 5325 16443 5383 16449
rect 5969 16483 6027 16489
rect 5969 16449 5981 16483
rect 6015 16480 6027 16483
rect 6429 16483 6487 16489
rect 6429 16480 6441 16483
rect 6015 16452 6441 16480
rect 6015 16449 6027 16452
rect 5969 16443 6027 16449
rect 6429 16449 6441 16452
rect 6475 16449 6487 16483
rect 6429 16443 6487 16449
rect 7073 16483 7131 16489
rect 7073 16449 7085 16483
rect 7119 16480 7131 16483
rect 7533 16483 7591 16489
rect 7533 16480 7545 16483
rect 7119 16452 7545 16480
rect 7119 16449 7131 16452
rect 7073 16443 7131 16449
rect 7533 16449 7545 16452
rect 7579 16449 7591 16483
rect 7533 16443 7591 16449
rect 8177 16483 8235 16489
rect 8177 16449 8189 16483
rect 8223 16480 8235 16483
rect 8637 16483 8695 16489
rect 8637 16480 8649 16483
rect 8223 16452 8649 16480
rect 8223 16449 8235 16452
rect 8177 16443 8235 16449
rect 8637 16449 8649 16452
rect 8683 16449 8695 16483
rect 8637 16443 8695 16449
rect 9281 16483 9339 16489
rect 9281 16449 9293 16483
rect 9327 16480 9339 16483
rect 9741 16483 9799 16489
rect 9741 16480 9753 16483
rect 9327 16452 9753 16480
rect 9327 16449 9339 16452
rect 9281 16443 9339 16449
rect 9741 16449 9753 16452
rect 9787 16449 9799 16483
rect 9741 16443 9799 16449
rect 10385 16483 10443 16489
rect 10385 16449 10397 16483
rect 10431 16480 10443 16483
rect 10845 16483 10903 16489
rect 10845 16480 10857 16483
rect 10431 16452 10857 16480
rect 10431 16449 10443 16452
rect 10385 16443 10443 16449
rect 10845 16449 10857 16452
rect 10891 16449 10903 16483
rect 10845 16443 10903 16449
rect 11489 16483 11547 16489
rect 11489 16449 11501 16483
rect 11535 16480 11547 16483
rect 11949 16483 12007 16489
rect 11949 16480 11961 16483
rect 11535 16452 11961 16480
rect 11535 16449 11547 16452
rect 11489 16443 11547 16449
rect 11949 16449 11961 16452
rect 11995 16449 12007 16483
rect 11949 16443 12007 16449
rect 12593 16483 12651 16489
rect 12593 16449 12605 16483
rect 12639 16480 12651 16483
rect 13053 16483 13111 16489
rect 13053 16480 13065 16483
rect 12639 16452 13065 16480
rect 12639 16449 12651 16452
rect 12593 16443 12651 16449
rect 13053 16449 13065 16452
rect 13099 16449 13111 16483
rect 13053 16443 13111 16449
rect 13697 16483 13755 16489
rect 13697 16449 13709 16483
rect 13743 16480 13755 16483
rect 14157 16483 14215 16489
rect 14157 16480 14169 16483
rect 13743 16452 14169 16480
rect 13743 16449 13755 16452
rect 13697 16443 13755 16449
rect 14157 16449 14169 16452
rect 14203 16449 14215 16483
rect 14157 16443 14215 16449
rect 14801 16483 14859 16489
rect 14801 16449 14813 16483
rect 14847 16480 14859 16483
rect 15261 16483 15319 16489
rect 15261 16480 15273 16483
rect 14847 16452 15273 16480
rect 14847 16449 14859 16452
rect 14801 16443 14859 16449
rect 15261 16449 15273 16452
rect 15307 16449 15319 16483
rect 15261 16443 15319 16449
rect 15905 16483 15963 16489
rect 15905 16449 15917 16483
rect 15951 16480 15963 16483
rect 16365 16483 16423 16489
rect 16365 16480 16377 16483
rect 15951 16452 16377 16480
rect 15951 16449 15963 16452
rect 15905 16443 15963 16449
rect 16365 16449 16377 16452
rect 16411 16449 16423 16483
rect 16365 16443 16423 16449
rect 17009 16483 17067 16489
rect 17009 16449 17021 16483
rect 17055 16480 17067 16483
rect 17469 16483 17527 16489
rect 17469 16480 17481 16483
rect 17055 16452 17481 16480
rect 17055 16449 17067 16452
rect 17009 16443 17067 16449
rect 17469 16449 17481 16452
rect 17515 16449 17527 16483
rect 17469 16443 17527 16449
rect 18113 16483 18171 16489
rect 18113 16449 18125 16483
rect 18159 16480 18171 16483
rect 18573 16483 18631 16489
rect 18573 16480 18585 16483
rect 18159 16452 18585 16480
rect 18159 16449 18171 16452
rect 18113 16443 18171 16449
rect 18573 16449 18585 16452
rect 18619 16449 18631 16483
rect 18573 16443 18631 16449
rect 19217 16483 19275 16489
rect 19217 16449 19229 16483
rect 19263 16480 19275 16483
rect 19677 16483 19735 16489
rect 19677 16480 19689 16483
rect 19263 16452 19689 16480
rect 19263 16449 19275 16452
rect 19217 16443 19275 16449
rect 19677 16449 19689 16452
rect 19723 16449 19735 16483
rect 19677 16443 19735 16449
rect 1904 16186 20764 16208
rect 1904 16134 7110 16186
rect 7162 16134 7174 16186
rect 7226 16134 7238 16186
rect 7290 16134 7302 16186
rect 7354 16134 12438 16186
rect 12490 16134 12502 16186
rect 12554 16134 12566 16186
rect 12618 16134 12630 16186
rect 12682 16134 17766 16186
rect 17818 16134 17830 16186
rect 17882 16134 17894 16186
rect 17946 16134 17958 16186
rect 18010 16134 20764 16186
rect 1904 16112 20764 16134
rect 1921 16007 1979 16013
rect 1921 15973 1933 16007
rect 1967 16004 1979 16007
rect 2562 16004 2568 16016
rect 1967 15976 2568 16004
rect 1967 15973 1979 15976
rect 1921 15967 1979 15973
rect 2562 15964 2568 15976
rect 2620 15964 2626 16016
rect 2470 15936 2476 15948
rect 2431 15908 2476 15936
rect 2470 15896 2476 15908
rect 2528 15896 2534 15948
rect 4865 15939 4923 15945
rect 4865 15936 4877 15939
rect 3132 15908 4877 15936
rect 3132 15877 3160 15908
rect 4865 15905 4877 15908
rect 4911 15905 4923 15939
rect 7073 15939 7131 15945
rect 7073 15936 7085 15939
rect 4865 15899 4923 15905
rect 5340 15908 7085 15936
rect 5340 15877 5368 15908
rect 7073 15905 7085 15908
rect 7119 15905 7131 15939
rect 9281 15939 9339 15945
rect 9281 15936 9293 15939
rect 7073 15899 7131 15905
rect 7548 15908 9293 15936
rect 7548 15877 7576 15908
rect 9281 15905 9293 15908
rect 9327 15905 9339 15939
rect 10385 15939 10443 15945
rect 10385 15936 10397 15939
rect 9281 15899 9339 15905
rect 9572 15908 10397 15936
rect 2381 15871 2439 15877
rect 2381 15837 2393 15871
rect 2427 15837 2439 15871
rect 2381 15831 2439 15837
rect 3117 15871 3175 15877
rect 3117 15837 3129 15871
rect 3163 15837 3175 15871
rect 3117 15831 3175 15837
rect 4221 15871 4279 15877
rect 4221 15837 4233 15871
rect 4267 15837 4279 15871
rect 4221 15831 4279 15837
rect 5325 15871 5383 15877
rect 5325 15837 5337 15871
rect 5371 15837 5383 15871
rect 5325 15831 5383 15837
rect 6440 15871 6498 15877
rect 6440 15837 6452 15871
rect 6486 15837 6498 15871
rect 6440 15831 6498 15837
rect 7533 15871 7591 15877
rect 7533 15837 7545 15871
rect 7579 15837 7591 15871
rect 7533 15831 7591 15837
rect 8648 15871 8706 15877
rect 8648 15837 8660 15871
rect 8694 15837 8706 15871
rect 8648 15831 8706 15837
rect 2396 15800 2424 15831
rect 3761 15803 3819 15809
rect 3761 15800 3773 15803
rect 2396 15772 3773 15800
rect 3761 15769 3773 15772
rect 3807 15769 3819 15803
rect 4236 15800 4264 15831
rect 5969 15803 6027 15809
rect 5969 15800 5981 15803
rect 4236 15772 5981 15800
rect 3761 15763 3819 15769
rect 5969 15769 5981 15772
rect 6015 15769 6027 15803
rect 6455 15800 6483 15831
rect 8177 15803 8235 15809
rect 8177 15800 8189 15803
rect 6455 15772 8189 15800
rect 5969 15763 6027 15769
rect 8177 15769 8189 15772
rect 8223 15769 8235 15803
rect 8663 15800 8691 15831
rect 9572 15800 9600 15908
rect 10385 15905 10397 15908
rect 10431 15905 10443 15939
rect 11489 15939 11547 15945
rect 11489 15936 11501 15939
rect 10385 15899 10443 15905
rect 10584 15908 11501 15936
rect 9741 15871 9799 15877
rect 9741 15837 9753 15871
rect 9787 15868 9799 15871
rect 10584 15868 10612 15908
rect 11489 15905 11501 15908
rect 11535 15905 11547 15939
rect 13697 15939 13755 15945
rect 13697 15936 13709 15939
rect 11489 15899 11547 15905
rect 11964 15908 13709 15936
rect 11964 15877 11992 15908
rect 13697 15905 13709 15908
rect 13743 15905 13755 15939
rect 15905 15939 15963 15945
rect 15905 15936 15917 15939
rect 13697 15899 13755 15905
rect 14183 15908 15917 15936
rect 14183 15877 14211 15908
rect 15905 15905 15917 15908
rect 15951 15905 15963 15939
rect 18113 15939 18171 15945
rect 18113 15936 18125 15939
rect 15905 15899 15963 15905
rect 16380 15908 18125 15936
rect 16380 15877 16408 15908
rect 18113 15905 18125 15908
rect 18159 15905 18171 15939
rect 20321 15939 20379 15945
rect 20321 15936 20333 15939
rect 18113 15899 18171 15905
rect 18588 15908 20333 15936
rect 18588 15877 18616 15908
rect 20321 15905 20333 15908
rect 20367 15905 20379 15939
rect 20321 15899 20379 15905
rect 9787 15840 10612 15868
rect 10845 15871 10903 15877
rect 9787 15837 9799 15840
rect 9741 15831 9799 15837
rect 10845 15837 10857 15871
rect 10891 15837 10903 15871
rect 10845 15831 10903 15837
rect 11949 15871 12007 15877
rect 11949 15837 11961 15871
rect 11995 15837 12007 15871
rect 11949 15831 12007 15837
rect 13053 15871 13111 15877
rect 13053 15837 13065 15871
rect 13099 15837 13111 15871
rect 13053 15831 13111 15837
rect 14168 15871 14226 15877
rect 14168 15837 14180 15871
rect 14214 15837 14226 15871
rect 14168 15831 14226 15837
rect 15261 15871 15319 15877
rect 15261 15837 15273 15871
rect 15307 15837 15319 15871
rect 15261 15831 15319 15837
rect 16365 15871 16423 15877
rect 16365 15837 16377 15871
rect 16411 15837 16423 15871
rect 16365 15831 16423 15837
rect 17469 15871 17527 15877
rect 17469 15837 17481 15871
rect 17515 15837 17527 15871
rect 17469 15831 17527 15837
rect 18573 15871 18631 15877
rect 18573 15837 18585 15871
rect 18619 15837 18631 15871
rect 19674 15868 19680 15880
rect 19635 15840 19680 15868
rect 18573 15831 18631 15837
rect 8663 15772 9600 15800
rect 10860 15800 10888 15831
rect 12593 15803 12651 15809
rect 12593 15800 12605 15803
rect 10860 15772 12605 15800
rect 8177 15763 8235 15769
rect 12593 15769 12605 15772
rect 12639 15769 12651 15803
rect 13068 15800 13096 15831
rect 14801 15803 14859 15809
rect 14801 15800 14813 15803
rect 13068 15772 14813 15800
rect 12593 15763 12651 15769
rect 14801 15769 14813 15772
rect 14847 15769 14859 15803
rect 15276 15800 15304 15831
rect 17009 15803 17067 15809
rect 17009 15800 17021 15803
rect 15276 15772 17021 15800
rect 14801 15763 14859 15769
rect 17009 15769 17021 15772
rect 17055 15769 17067 15803
rect 17484 15800 17512 15831
rect 19674 15828 19680 15840
rect 19732 15828 19738 15880
rect 19217 15803 19275 15809
rect 19217 15800 19229 15803
rect 17484 15772 19229 15800
rect 17009 15763 17067 15769
rect 19217 15769 19229 15772
rect 19263 15769 19275 15803
rect 19217 15763 19275 15769
rect 2286 15692 2292 15744
rect 2344 15732 2350 15744
rect 2344 15704 2389 15732
rect 2344 15692 2350 15704
rect 1904 15642 20764 15664
rect 1904 15590 4446 15642
rect 4498 15590 4510 15642
rect 4562 15590 4574 15642
rect 4626 15590 4638 15642
rect 4690 15590 9774 15642
rect 9826 15590 9838 15642
rect 9890 15590 9902 15642
rect 9954 15590 9966 15642
rect 10018 15590 15102 15642
rect 15154 15590 15166 15642
rect 15218 15590 15230 15642
rect 15282 15590 15294 15642
rect 15346 15590 20764 15642
rect 1904 15568 20764 15590
rect 19674 15488 19680 15540
rect 19732 15528 19738 15540
rect 20321 15531 20379 15537
rect 20321 15528 20333 15531
rect 19732 15500 20333 15528
rect 19732 15488 19738 15500
rect 20321 15497 20333 15500
rect 20367 15497 20379 15531
rect 20321 15491 20379 15497
rect 3117 15395 3175 15401
rect 3117 15361 3129 15395
rect 3163 15361 3175 15395
rect 3117 15355 3175 15361
rect 3761 15395 3819 15401
rect 3761 15361 3773 15395
rect 3807 15392 3819 15395
rect 4221 15395 4279 15401
rect 4221 15392 4233 15395
rect 3807 15364 4233 15392
rect 3807 15361 3819 15364
rect 3761 15355 3819 15361
rect 4221 15361 4233 15364
rect 4267 15361 4279 15395
rect 4221 15355 4279 15361
rect 4865 15395 4923 15401
rect 4865 15361 4877 15395
rect 4911 15392 4923 15395
rect 5325 15395 5383 15401
rect 5325 15392 5337 15395
rect 4911 15364 5337 15392
rect 4911 15361 4923 15364
rect 4865 15355 4923 15361
rect 5325 15361 5337 15364
rect 5371 15361 5383 15395
rect 5325 15355 5383 15361
rect 5969 15395 6027 15401
rect 5969 15361 5981 15395
rect 6015 15392 6027 15395
rect 6429 15395 6487 15401
rect 6429 15392 6441 15395
rect 6015 15364 6441 15392
rect 6015 15361 6027 15364
rect 5969 15355 6027 15361
rect 6429 15361 6441 15364
rect 6475 15361 6487 15395
rect 6429 15355 6487 15361
rect 7073 15395 7131 15401
rect 7073 15361 7085 15395
rect 7119 15392 7131 15395
rect 7533 15395 7591 15401
rect 7533 15392 7545 15395
rect 7119 15364 7545 15392
rect 7119 15361 7131 15364
rect 7073 15355 7131 15361
rect 7533 15361 7545 15364
rect 7579 15361 7591 15395
rect 7533 15355 7591 15361
rect 8177 15395 8235 15401
rect 8177 15361 8189 15395
rect 8223 15392 8235 15395
rect 8637 15395 8695 15401
rect 8637 15392 8649 15395
rect 8223 15364 8649 15392
rect 8223 15361 8235 15364
rect 8177 15355 8235 15361
rect 8637 15361 8649 15364
rect 8683 15361 8695 15395
rect 8637 15355 8695 15361
rect 9281 15395 9339 15401
rect 9281 15361 9293 15395
rect 9327 15392 9339 15395
rect 9741 15395 9799 15401
rect 9741 15392 9753 15395
rect 9327 15364 9753 15392
rect 9327 15361 9339 15364
rect 9281 15355 9339 15361
rect 9741 15361 9753 15364
rect 9787 15361 9799 15395
rect 9741 15355 9799 15361
rect 10385 15395 10443 15401
rect 10385 15361 10397 15395
rect 10431 15392 10443 15395
rect 10845 15395 10903 15401
rect 10845 15392 10857 15395
rect 10431 15364 10857 15392
rect 10431 15361 10443 15364
rect 10385 15355 10443 15361
rect 10845 15361 10857 15364
rect 10891 15361 10903 15395
rect 10845 15355 10903 15361
rect 11489 15395 11547 15401
rect 11489 15361 11501 15395
rect 11535 15392 11547 15395
rect 11949 15395 12007 15401
rect 11949 15392 11961 15395
rect 11535 15364 11961 15392
rect 11535 15361 11547 15364
rect 11489 15355 11547 15361
rect 11949 15361 11961 15364
rect 11995 15361 12007 15395
rect 11949 15355 12007 15361
rect 12593 15395 12651 15401
rect 12593 15361 12605 15395
rect 12639 15392 12651 15395
rect 13053 15395 13111 15401
rect 13053 15392 13065 15395
rect 12639 15364 13065 15392
rect 12639 15361 12651 15364
rect 12593 15355 12651 15361
rect 13053 15361 13065 15364
rect 13099 15361 13111 15395
rect 13053 15355 13111 15361
rect 13697 15395 13755 15401
rect 13697 15361 13709 15395
rect 13743 15392 13755 15395
rect 14157 15395 14215 15401
rect 14157 15392 14169 15395
rect 13743 15364 14169 15392
rect 13743 15361 13755 15364
rect 13697 15355 13755 15361
rect 14157 15361 14169 15364
rect 14203 15361 14215 15395
rect 14157 15355 14215 15361
rect 14801 15395 14859 15401
rect 14801 15361 14813 15395
rect 14847 15392 14859 15395
rect 15261 15395 15319 15401
rect 15261 15392 15273 15395
rect 14847 15364 15273 15392
rect 14847 15361 14859 15364
rect 14801 15355 14859 15361
rect 15261 15361 15273 15364
rect 15307 15361 15319 15395
rect 15261 15355 15319 15361
rect 15905 15395 15963 15401
rect 15905 15361 15917 15395
rect 15951 15392 15963 15395
rect 16365 15395 16423 15401
rect 16365 15392 16377 15395
rect 15951 15364 16377 15392
rect 15951 15361 15963 15364
rect 15905 15355 15963 15361
rect 16365 15361 16377 15364
rect 16411 15361 16423 15395
rect 16365 15355 16423 15361
rect 17009 15395 17067 15401
rect 17009 15361 17021 15395
rect 17055 15392 17067 15395
rect 17469 15395 17527 15401
rect 17469 15392 17481 15395
rect 17055 15364 17481 15392
rect 17055 15361 17067 15364
rect 17009 15355 17067 15361
rect 17469 15361 17481 15364
rect 17515 15361 17527 15395
rect 17469 15355 17527 15361
rect 18113 15395 18171 15401
rect 18113 15361 18125 15395
rect 18159 15392 18171 15395
rect 18573 15395 18631 15401
rect 18573 15392 18585 15395
rect 18159 15364 18585 15392
rect 18159 15361 18171 15364
rect 18113 15355 18171 15361
rect 18573 15361 18585 15364
rect 18619 15361 18631 15395
rect 18573 15355 18631 15361
rect 19217 15395 19275 15401
rect 19217 15361 19229 15395
rect 19263 15392 19275 15395
rect 19677 15395 19735 15401
rect 19677 15392 19689 15395
rect 19263 15364 19689 15392
rect 19263 15361 19275 15364
rect 19217 15355 19275 15361
rect 19677 15361 19689 15364
rect 19723 15361 19735 15395
rect 19677 15355 19735 15361
rect 3132 15324 3160 15355
rect 3132 15296 3804 15324
rect 3776 15268 3804 15296
rect 3758 15216 3764 15268
rect 3816 15216 3822 15268
rect 1904 15098 20764 15120
rect 1904 15046 7110 15098
rect 7162 15046 7174 15098
rect 7226 15046 7238 15098
rect 7290 15046 7302 15098
rect 7354 15046 12438 15098
rect 12490 15046 12502 15098
rect 12554 15046 12566 15098
rect 12618 15046 12630 15098
rect 12682 15046 17766 15098
rect 17818 15046 17830 15098
rect 17882 15046 17894 15098
rect 17946 15046 17958 15098
rect 18010 15046 20764 15098
rect 1904 15024 20764 15046
rect 3758 14984 3764 14996
rect 3719 14956 3764 14984
rect 3758 14944 3764 14956
rect 3816 14944 3822 14996
rect 5969 14851 6027 14857
rect 5969 14848 5981 14851
rect 4236 14820 5981 14848
rect 4236 14789 4264 14820
rect 5969 14817 5981 14820
rect 6015 14817 6027 14851
rect 8177 14851 8235 14857
rect 8177 14848 8189 14851
rect 5969 14811 6027 14817
rect 6455 14820 8189 14848
rect 6455 14789 6483 14820
rect 8177 14817 8189 14820
rect 8223 14817 8235 14851
rect 11489 14851 11547 14857
rect 11489 14848 11501 14851
rect 8177 14811 8235 14817
rect 8663 14820 9600 14848
rect 8663 14789 8691 14820
rect 3117 14783 3175 14789
rect 3117 14749 3129 14783
rect 3163 14749 3175 14783
rect 3117 14743 3175 14749
rect 4221 14783 4279 14789
rect 4221 14749 4233 14783
rect 4267 14749 4279 14783
rect 4221 14743 4279 14749
rect 5325 14783 5383 14789
rect 5325 14749 5337 14783
rect 5371 14749 5383 14783
rect 5325 14743 5383 14749
rect 6440 14783 6498 14789
rect 6440 14749 6452 14783
rect 6486 14749 6498 14783
rect 6440 14743 6498 14749
rect 7533 14783 7591 14789
rect 7533 14749 7545 14783
rect 7579 14749 7591 14783
rect 7533 14743 7591 14749
rect 8648 14783 8706 14789
rect 8648 14749 8660 14783
rect 8694 14749 8706 14783
rect 8648 14743 8706 14749
rect 3132 14712 3160 14743
rect 4865 14715 4923 14721
rect 4865 14712 4877 14715
rect 3132 14684 4877 14712
rect 4865 14681 4877 14684
rect 4911 14681 4923 14715
rect 5340 14712 5368 14743
rect 7073 14715 7131 14721
rect 7073 14712 7085 14715
rect 5340 14684 7085 14712
rect 4865 14675 4923 14681
rect 7073 14681 7085 14684
rect 7119 14681 7131 14715
rect 7548 14712 7576 14743
rect 9281 14715 9339 14721
rect 9281 14712 9293 14715
rect 7548 14684 9293 14712
rect 7073 14675 7131 14681
rect 9281 14681 9293 14684
rect 9327 14681 9339 14715
rect 9572 14712 9600 14820
rect 9756 14820 11501 14848
rect 9756 14789 9784 14820
rect 11489 14817 11501 14820
rect 11535 14817 11547 14851
rect 13697 14851 13755 14857
rect 13697 14848 13709 14851
rect 11489 14811 11547 14817
rect 11964 14820 13709 14848
rect 11964 14789 11992 14820
rect 13697 14817 13709 14820
rect 13743 14817 13755 14851
rect 15905 14851 15963 14857
rect 15905 14848 15917 14851
rect 13697 14811 13755 14817
rect 14183 14820 15917 14848
rect 14183 14789 14211 14820
rect 15905 14817 15917 14820
rect 15951 14817 15963 14851
rect 18113 14851 18171 14857
rect 18113 14848 18125 14851
rect 15905 14811 15963 14817
rect 16380 14820 18125 14848
rect 16380 14789 16408 14820
rect 18113 14817 18125 14820
rect 18159 14817 18171 14851
rect 20321 14851 20379 14857
rect 20321 14848 20333 14851
rect 18113 14811 18171 14817
rect 18588 14820 20333 14848
rect 18588 14789 18616 14820
rect 20321 14817 20333 14820
rect 20367 14817 20379 14851
rect 20321 14811 20379 14817
rect 9741 14783 9799 14789
rect 9741 14749 9753 14783
rect 9787 14749 9799 14783
rect 9741 14743 9799 14749
rect 10845 14783 10903 14789
rect 10845 14749 10857 14783
rect 10891 14749 10903 14783
rect 10845 14743 10903 14749
rect 11949 14783 12007 14789
rect 11949 14749 11961 14783
rect 11995 14749 12007 14783
rect 11949 14743 12007 14749
rect 13053 14783 13111 14789
rect 13053 14749 13065 14783
rect 13099 14749 13111 14783
rect 13053 14743 13111 14749
rect 14168 14783 14226 14789
rect 14168 14749 14180 14783
rect 14214 14749 14226 14783
rect 14168 14743 14226 14749
rect 15261 14783 15319 14789
rect 15261 14749 15273 14783
rect 15307 14749 15319 14783
rect 15261 14743 15319 14749
rect 16365 14783 16423 14789
rect 16365 14749 16377 14783
rect 16411 14749 16423 14783
rect 16365 14743 16423 14749
rect 17469 14783 17527 14789
rect 17469 14749 17481 14783
rect 17515 14749 17527 14783
rect 17469 14743 17527 14749
rect 18573 14783 18631 14789
rect 18573 14749 18585 14783
rect 18619 14749 18631 14783
rect 18573 14743 18631 14749
rect 19677 14783 19735 14789
rect 19677 14749 19689 14783
rect 19723 14780 19735 14783
rect 20134 14780 20140 14792
rect 19723 14752 20140 14780
rect 19723 14749 19735 14752
rect 19677 14743 19735 14749
rect 10385 14715 10443 14721
rect 10385 14712 10397 14715
rect 9572 14684 10397 14712
rect 9281 14675 9339 14681
rect 10385 14681 10397 14684
rect 10431 14681 10443 14715
rect 10860 14712 10888 14743
rect 12593 14715 12651 14721
rect 12593 14712 12605 14715
rect 10860 14684 12605 14712
rect 10385 14675 10443 14681
rect 12593 14681 12605 14684
rect 12639 14681 12651 14715
rect 13068 14712 13096 14743
rect 14801 14715 14859 14721
rect 14801 14712 14813 14715
rect 13068 14684 14813 14712
rect 12593 14675 12651 14681
rect 14801 14681 14813 14684
rect 14847 14681 14859 14715
rect 15276 14712 15304 14743
rect 17009 14715 17067 14721
rect 17009 14712 17021 14715
rect 15276 14684 17021 14712
rect 14801 14675 14859 14681
rect 17009 14681 17021 14684
rect 17055 14681 17067 14715
rect 17484 14712 17512 14743
rect 20134 14740 20140 14752
rect 20192 14740 20198 14792
rect 19217 14715 19275 14721
rect 19217 14712 19229 14715
rect 17484 14684 19229 14712
rect 17009 14675 17067 14681
rect 19217 14681 19229 14684
rect 19263 14681 19275 14715
rect 19217 14675 19275 14681
rect 1904 14554 20764 14576
rect 1904 14502 4446 14554
rect 4498 14502 4510 14554
rect 4562 14502 4574 14554
rect 4626 14502 4638 14554
rect 4690 14502 9774 14554
rect 9826 14502 9838 14554
rect 9890 14502 9902 14554
rect 9954 14502 9966 14554
rect 10018 14502 15102 14554
rect 15154 14502 15166 14554
rect 15218 14502 15230 14554
rect 15282 14502 15294 14554
rect 15346 14502 20764 14554
rect 1904 14480 20764 14502
rect 20134 14400 20140 14452
rect 20192 14440 20198 14452
rect 20321 14443 20379 14449
rect 20321 14440 20333 14443
rect 20192 14412 20333 14440
rect 20192 14400 20198 14412
rect 20321 14409 20333 14412
rect 20367 14409 20379 14443
rect 20321 14403 20379 14409
rect 2286 14264 2292 14316
rect 2344 14304 2350 14316
rect 3117 14307 3175 14313
rect 3117 14304 3129 14307
rect 2344 14276 3129 14304
rect 2344 14264 2350 14276
rect 3117 14273 3129 14276
rect 3163 14273 3175 14307
rect 3117 14267 3175 14273
rect 3761 14307 3819 14313
rect 3761 14273 3773 14307
rect 3807 14304 3819 14307
rect 4221 14307 4279 14313
rect 4221 14304 4233 14307
rect 3807 14276 4233 14304
rect 3807 14273 3819 14276
rect 3761 14267 3819 14273
rect 4221 14273 4233 14276
rect 4267 14273 4279 14307
rect 4221 14267 4279 14273
rect 4865 14307 4923 14313
rect 4865 14273 4877 14307
rect 4911 14304 4923 14307
rect 5325 14307 5383 14313
rect 5325 14304 5337 14307
rect 4911 14276 5337 14304
rect 4911 14273 4923 14276
rect 4865 14267 4923 14273
rect 5325 14273 5337 14276
rect 5371 14273 5383 14307
rect 5325 14267 5383 14273
rect 5969 14307 6027 14313
rect 5969 14273 5981 14307
rect 6015 14304 6027 14307
rect 6429 14307 6487 14313
rect 6429 14304 6441 14307
rect 6015 14276 6441 14304
rect 6015 14273 6027 14276
rect 5969 14267 6027 14273
rect 6429 14273 6441 14276
rect 6475 14273 6487 14307
rect 6429 14267 6487 14273
rect 7073 14307 7131 14313
rect 7073 14273 7085 14307
rect 7119 14304 7131 14307
rect 7533 14307 7591 14313
rect 7533 14304 7545 14307
rect 7119 14276 7545 14304
rect 7119 14273 7131 14276
rect 7073 14267 7131 14273
rect 7533 14273 7545 14276
rect 7579 14273 7591 14307
rect 7533 14267 7591 14273
rect 8177 14307 8235 14313
rect 8177 14273 8189 14307
rect 8223 14304 8235 14307
rect 8637 14307 8695 14313
rect 8637 14304 8649 14307
rect 8223 14276 8649 14304
rect 8223 14273 8235 14276
rect 8177 14267 8235 14273
rect 8637 14273 8649 14276
rect 8683 14273 8695 14307
rect 8637 14267 8695 14273
rect 9281 14307 9339 14313
rect 9281 14273 9293 14307
rect 9327 14304 9339 14307
rect 9741 14307 9799 14313
rect 9741 14304 9753 14307
rect 9327 14276 9753 14304
rect 9327 14273 9339 14276
rect 9281 14267 9339 14273
rect 9741 14273 9753 14276
rect 9787 14273 9799 14307
rect 9741 14267 9799 14273
rect 10385 14307 10443 14313
rect 10385 14273 10397 14307
rect 10431 14304 10443 14307
rect 10845 14307 10903 14313
rect 10845 14304 10857 14307
rect 10431 14276 10857 14304
rect 10431 14273 10443 14276
rect 10385 14267 10443 14273
rect 10845 14273 10857 14276
rect 10891 14273 10903 14307
rect 10845 14267 10903 14273
rect 11489 14307 11547 14313
rect 11489 14273 11501 14307
rect 11535 14304 11547 14307
rect 11949 14307 12007 14313
rect 11949 14304 11961 14307
rect 11535 14276 11961 14304
rect 11535 14273 11547 14276
rect 11489 14267 11547 14273
rect 11949 14273 11961 14276
rect 11995 14273 12007 14307
rect 11949 14267 12007 14273
rect 12593 14307 12651 14313
rect 12593 14273 12605 14307
rect 12639 14304 12651 14307
rect 13053 14307 13111 14313
rect 13053 14304 13065 14307
rect 12639 14276 13065 14304
rect 12639 14273 12651 14276
rect 12593 14267 12651 14273
rect 13053 14273 13065 14276
rect 13099 14273 13111 14307
rect 13053 14267 13111 14273
rect 13697 14307 13755 14313
rect 13697 14273 13709 14307
rect 13743 14304 13755 14307
rect 14157 14307 14215 14313
rect 14157 14304 14169 14307
rect 13743 14276 14169 14304
rect 13743 14273 13755 14276
rect 13697 14267 13755 14273
rect 14157 14273 14169 14276
rect 14203 14273 14215 14307
rect 14157 14267 14215 14273
rect 14801 14307 14859 14313
rect 14801 14273 14813 14307
rect 14847 14304 14859 14307
rect 15261 14307 15319 14313
rect 15261 14304 15273 14307
rect 14847 14276 15273 14304
rect 14847 14273 14859 14276
rect 14801 14267 14859 14273
rect 15261 14273 15273 14276
rect 15307 14273 15319 14307
rect 15261 14267 15319 14273
rect 15905 14307 15963 14313
rect 15905 14273 15917 14307
rect 15951 14304 15963 14307
rect 16365 14307 16423 14313
rect 16365 14304 16377 14307
rect 15951 14276 16377 14304
rect 15951 14273 15963 14276
rect 15905 14267 15963 14273
rect 16365 14273 16377 14276
rect 16411 14273 16423 14307
rect 16365 14267 16423 14273
rect 17009 14307 17067 14313
rect 17009 14273 17021 14307
rect 17055 14304 17067 14307
rect 17469 14307 17527 14313
rect 17469 14304 17481 14307
rect 17055 14276 17481 14304
rect 17055 14273 17067 14276
rect 17009 14267 17067 14273
rect 17469 14273 17481 14276
rect 17515 14273 17527 14307
rect 17469 14267 17527 14273
rect 18113 14307 18171 14313
rect 18113 14273 18125 14307
rect 18159 14304 18171 14307
rect 18573 14307 18631 14313
rect 18573 14304 18585 14307
rect 18159 14276 18585 14304
rect 18159 14273 18171 14276
rect 18113 14267 18171 14273
rect 18573 14273 18585 14276
rect 18619 14273 18631 14307
rect 18573 14267 18631 14273
rect 19217 14307 19275 14313
rect 19217 14273 19229 14307
rect 19263 14304 19275 14307
rect 19677 14307 19735 14313
rect 19677 14304 19689 14307
rect 19263 14276 19689 14304
rect 19263 14273 19275 14276
rect 19217 14267 19275 14273
rect 19677 14273 19689 14276
rect 19723 14273 19735 14307
rect 19677 14267 19735 14273
rect 1904 14010 20764 14032
rect 1904 13958 7110 14010
rect 7162 13958 7174 14010
rect 7226 13958 7238 14010
rect 7290 13958 7302 14010
rect 7354 13958 12438 14010
rect 12490 13958 12502 14010
rect 12554 13958 12566 14010
rect 12618 13958 12630 14010
rect 12682 13958 17766 14010
rect 17818 13958 17830 14010
rect 17882 13958 17894 14010
rect 17946 13958 17958 14010
rect 18010 13958 20764 14010
rect 1904 13936 20764 13958
rect 1921 13831 1979 13837
rect 1921 13797 1933 13831
rect 1967 13828 1979 13831
rect 2286 13828 2292 13840
rect 1967 13800 2292 13828
rect 1967 13797 1979 13800
rect 1921 13791 1979 13797
rect 2286 13788 2292 13800
rect 2344 13788 2350 13840
rect 2470 13760 2476 13772
rect 2431 13732 2476 13760
rect 2470 13720 2476 13732
rect 2528 13720 2534 13772
rect 4865 13763 4923 13769
rect 4865 13760 4877 13763
rect 3132 13732 4877 13760
rect 3132 13701 3160 13732
rect 4865 13729 4877 13732
rect 4911 13729 4923 13763
rect 7073 13763 7131 13769
rect 7073 13760 7085 13763
rect 4865 13723 4923 13729
rect 5340 13732 7085 13760
rect 5340 13701 5368 13732
rect 7073 13729 7085 13732
rect 7119 13729 7131 13763
rect 8177 13763 8235 13769
rect 8177 13760 8189 13763
rect 7073 13723 7131 13729
rect 7364 13732 8189 13760
rect 3117 13695 3175 13701
rect 3117 13661 3129 13695
rect 3163 13661 3175 13695
rect 3117 13655 3175 13661
rect 4221 13695 4279 13701
rect 4221 13661 4233 13695
rect 4267 13661 4279 13695
rect 4221 13655 4279 13661
rect 5325 13695 5383 13701
rect 5325 13661 5337 13695
rect 5371 13661 5383 13695
rect 5325 13655 5383 13661
rect 6440 13695 6498 13701
rect 6440 13661 6452 13695
rect 6486 13661 6498 13695
rect 6440 13655 6498 13661
rect 2381 13627 2439 13633
rect 2381 13593 2393 13627
rect 2427 13624 2439 13627
rect 3761 13627 3819 13633
rect 3761 13624 3773 13627
rect 2427 13596 3773 13624
rect 2427 13593 2439 13596
rect 2381 13587 2439 13593
rect 3761 13593 3773 13596
rect 3807 13593 3819 13627
rect 4236 13624 4264 13655
rect 5969 13627 6027 13633
rect 5969 13624 5981 13627
rect 4236 13596 5981 13624
rect 3761 13587 3819 13593
rect 5969 13593 5981 13596
rect 6015 13593 6027 13627
rect 6455 13624 6483 13655
rect 7364 13624 7392 13732
rect 8177 13729 8189 13732
rect 8223 13729 8235 13763
rect 10385 13763 10443 13769
rect 10385 13760 10397 13763
rect 8177 13723 8235 13729
rect 8652 13732 10397 13760
rect 8652 13701 8680 13732
rect 10385 13729 10397 13732
rect 10431 13729 10443 13763
rect 11489 13763 11547 13769
rect 11489 13760 11501 13763
rect 10385 13723 10443 13729
rect 10584 13732 11501 13760
rect 7533 13695 7591 13701
rect 7533 13661 7545 13695
rect 7579 13661 7591 13695
rect 7533 13655 7591 13661
rect 8648 13695 8706 13701
rect 8648 13661 8660 13695
rect 8694 13661 8706 13695
rect 8648 13655 8706 13661
rect 9741 13695 9799 13701
rect 9741 13661 9753 13695
rect 9787 13692 9799 13695
rect 10584 13692 10612 13732
rect 11489 13729 11501 13732
rect 11535 13729 11547 13763
rect 13697 13763 13755 13769
rect 13697 13760 13709 13763
rect 11489 13723 11547 13729
rect 11964 13732 13709 13760
rect 11964 13701 11992 13732
rect 13697 13729 13709 13732
rect 13743 13729 13755 13763
rect 15905 13763 15963 13769
rect 15905 13760 15917 13763
rect 13697 13723 13755 13729
rect 14172 13732 15917 13760
rect 14172 13701 14200 13732
rect 15905 13729 15917 13732
rect 15951 13729 15963 13763
rect 18113 13763 18171 13769
rect 18113 13760 18125 13763
rect 15905 13723 15963 13729
rect 16380 13732 18125 13760
rect 16380 13701 16408 13732
rect 18113 13729 18125 13732
rect 18159 13729 18171 13763
rect 20321 13763 20379 13769
rect 20321 13760 20333 13763
rect 18113 13723 18171 13729
rect 18588 13732 20333 13760
rect 18588 13701 18616 13732
rect 20321 13729 20333 13732
rect 20367 13729 20379 13763
rect 20321 13723 20379 13729
rect 9787 13664 10612 13692
rect 10845 13695 10903 13701
rect 9787 13661 9799 13664
rect 9741 13655 9799 13661
rect 10845 13661 10857 13695
rect 10891 13661 10903 13695
rect 10845 13655 10903 13661
rect 11949 13695 12007 13701
rect 11949 13661 11961 13695
rect 11995 13661 12007 13695
rect 11949 13655 12007 13661
rect 13053 13695 13111 13701
rect 13053 13661 13065 13695
rect 13099 13661 13111 13695
rect 13053 13655 13111 13661
rect 14168 13695 14226 13701
rect 14168 13661 14180 13695
rect 14214 13661 14226 13695
rect 14168 13655 14226 13661
rect 15261 13695 15319 13701
rect 15261 13661 15273 13695
rect 15307 13661 15319 13695
rect 15261 13655 15319 13661
rect 16365 13695 16423 13701
rect 16365 13661 16377 13695
rect 16411 13661 16423 13695
rect 16365 13655 16423 13661
rect 17469 13695 17527 13701
rect 17469 13661 17481 13695
rect 17515 13661 17527 13695
rect 17469 13655 17527 13661
rect 18573 13695 18631 13701
rect 18573 13661 18585 13695
rect 18619 13661 18631 13695
rect 19674 13692 19680 13704
rect 19635 13664 19680 13692
rect 18573 13655 18631 13661
rect 6455 13596 7392 13624
rect 7548 13624 7576 13655
rect 9281 13627 9339 13633
rect 9281 13624 9293 13627
rect 7548 13596 9293 13624
rect 5969 13587 6027 13593
rect 9281 13593 9293 13596
rect 9327 13593 9339 13627
rect 10860 13624 10888 13655
rect 12593 13627 12651 13633
rect 12593 13624 12605 13627
rect 10860 13596 12605 13624
rect 9281 13587 9339 13593
rect 12593 13593 12605 13596
rect 12639 13593 12651 13627
rect 13068 13624 13096 13655
rect 14801 13627 14859 13633
rect 14801 13624 14813 13627
rect 13068 13596 14813 13624
rect 12593 13587 12651 13593
rect 14801 13593 14813 13596
rect 14847 13593 14859 13627
rect 15276 13624 15304 13655
rect 17009 13627 17067 13633
rect 17009 13624 17021 13627
rect 15276 13596 17021 13624
rect 14801 13587 14859 13593
rect 17009 13593 17021 13596
rect 17055 13593 17067 13627
rect 17484 13624 17512 13655
rect 19674 13652 19680 13664
rect 19732 13652 19738 13704
rect 19217 13627 19275 13633
rect 19217 13624 19229 13627
rect 17484 13596 19229 13624
rect 17009 13587 17067 13593
rect 19217 13593 19229 13596
rect 19263 13593 19275 13627
rect 19217 13587 19275 13593
rect 2286 13516 2292 13568
rect 2344 13556 2350 13568
rect 2344 13528 2389 13556
rect 2344 13516 2350 13528
rect 1904 13466 20764 13488
rect 1904 13414 4446 13466
rect 4498 13414 4510 13466
rect 4562 13414 4574 13466
rect 4626 13414 4638 13466
rect 4690 13414 9774 13466
rect 9826 13414 9838 13466
rect 9890 13414 9902 13466
rect 9954 13414 9966 13466
rect 10018 13414 15102 13466
rect 15154 13414 15166 13466
rect 15218 13414 15230 13466
rect 15282 13414 15294 13466
rect 15346 13414 20764 13466
rect 1904 13392 20764 13414
rect 19674 13312 19680 13364
rect 19732 13352 19738 13364
rect 20321 13355 20379 13361
rect 20321 13352 20333 13355
rect 19732 13324 20333 13352
rect 19732 13312 19738 13324
rect 20321 13321 20333 13324
rect 20367 13321 20379 13355
rect 20321 13315 20379 13321
rect 3117 13219 3175 13225
rect 3117 13185 3129 13219
rect 3163 13185 3175 13219
rect 3117 13179 3175 13185
rect 3761 13219 3819 13225
rect 3761 13185 3773 13219
rect 3807 13216 3819 13219
rect 4221 13219 4279 13225
rect 4221 13216 4233 13219
rect 3807 13188 4233 13216
rect 3807 13185 3819 13188
rect 3761 13179 3819 13185
rect 4221 13185 4233 13188
rect 4267 13185 4279 13219
rect 4221 13179 4279 13185
rect 4865 13219 4923 13225
rect 4865 13185 4877 13219
rect 4911 13216 4923 13219
rect 5325 13219 5383 13225
rect 5325 13216 5337 13219
rect 4911 13188 5337 13216
rect 4911 13185 4923 13188
rect 4865 13179 4923 13185
rect 5325 13185 5337 13188
rect 5371 13185 5383 13219
rect 5325 13179 5383 13185
rect 5969 13219 6027 13225
rect 5969 13185 5981 13219
rect 6015 13216 6027 13219
rect 6429 13219 6487 13225
rect 6429 13216 6441 13219
rect 6015 13188 6441 13216
rect 6015 13185 6027 13188
rect 5969 13179 6027 13185
rect 6429 13185 6441 13188
rect 6475 13185 6487 13219
rect 6429 13179 6487 13185
rect 7073 13219 7131 13225
rect 7073 13185 7085 13219
rect 7119 13216 7131 13219
rect 7533 13219 7591 13225
rect 7533 13216 7545 13219
rect 7119 13188 7545 13216
rect 7119 13185 7131 13188
rect 7073 13179 7131 13185
rect 7533 13185 7545 13188
rect 7579 13185 7591 13219
rect 7533 13179 7591 13185
rect 8177 13219 8235 13225
rect 8177 13185 8189 13219
rect 8223 13216 8235 13219
rect 8637 13219 8695 13225
rect 8637 13216 8649 13219
rect 8223 13188 8649 13216
rect 8223 13185 8235 13188
rect 8177 13179 8235 13185
rect 8637 13185 8649 13188
rect 8683 13185 8695 13219
rect 8637 13179 8695 13185
rect 9281 13219 9339 13225
rect 9281 13185 9293 13219
rect 9327 13216 9339 13219
rect 9741 13219 9799 13225
rect 9741 13216 9753 13219
rect 9327 13188 9753 13216
rect 9327 13185 9339 13188
rect 9281 13179 9339 13185
rect 9741 13185 9753 13188
rect 9787 13185 9799 13219
rect 9741 13179 9799 13185
rect 10385 13219 10443 13225
rect 10385 13185 10397 13219
rect 10431 13216 10443 13219
rect 10845 13219 10903 13225
rect 10845 13216 10857 13219
rect 10431 13188 10857 13216
rect 10431 13185 10443 13188
rect 10385 13179 10443 13185
rect 10845 13185 10857 13188
rect 10891 13185 10903 13219
rect 10845 13179 10903 13185
rect 11489 13219 11547 13225
rect 11489 13185 11501 13219
rect 11535 13216 11547 13219
rect 11949 13219 12007 13225
rect 11949 13216 11961 13219
rect 11535 13188 11961 13216
rect 11535 13185 11547 13188
rect 11489 13179 11547 13185
rect 11949 13185 11961 13188
rect 11995 13185 12007 13219
rect 11949 13179 12007 13185
rect 12593 13219 12651 13225
rect 12593 13185 12605 13219
rect 12639 13216 12651 13219
rect 13053 13219 13111 13225
rect 13053 13216 13065 13219
rect 12639 13188 13065 13216
rect 12639 13185 12651 13188
rect 12593 13179 12651 13185
rect 13053 13185 13065 13188
rect 13099 13185 13111 13219
rect 13053 13179 13111 13185
rect 13697 13219 13755 13225
rect 13697 13185 13709 13219
rect 13743 13216 13755 13219
rect 14157 13219 14215 13225
rect 14157 13216 14169 13219
rect 13743 13188 14169 13216
rect 13743 13185 13755 13188
rect 13697 13179 13755 13185
rect 14157 13185 14169 13188
rect 14203 13185 14215 13219
rect 14157 13179 14215 13185
rect 14801 13219 14859 13225
rect 14801 13185 14813 13219
rect 14847 13216 14859 13219
rect 15261 13219 15319 13225
rect 15261 13216 15273 13219
rect 14847 13188 15273 13216
rect 14847 13185 14859 13188
rect 14801 13179 14859 13185
rect 15261 13185 15273 13188
rect 15307 13185 15319 13219
rect 15261 13179 15319 13185
rect 15905 13219 15963 13225
rect 15905 13185 15917 13219
rect 15951 13216 15963 13219
rect 16365 13219 16423 13225
rect 16365 13216 16377 13219
rect 15951 13188 16377 13216
rect 15951 13185 15963 13188
rect 15905 13179 15963 13185
rect 16365 13185 16377 13188
rect 16411 13185 16423 13219
rect 16365 13179 16423 13185
rect 17009 13219 17067 13225
rect 17009 13185 17021 13219
rect 17055 13216 17067 13219
rect 17469 13219 17527 13225
rect 17469 13216 17481 13219
rect 17055 13188 17481 13216
rect 17055 13185 17067 13188
rect 17009 13179 17067 13185
rect 17469 13185 17481 13188
rect 17515 13185 17527 13219
rect 17469 13179 17527 13185
rect 18113 13219 18171 13225
rect 18113 13185 18125 13219
rect 18159 13216 18171 13219
rect 18573 13219 18631 13225
rect 18573 13216 18585 13219
rect 18159 13188 18585 13216
rect 18159 13185 18171 13188
rect 18113 13179 18171 13185
rect 18573 13185 18585 13188
rect 18619 13185 18631 13219
rect 18573 13179 18631 13185
rect 19217 13219 19275 13225
rect 19217 13185 19229 13219
rect 19263 13216 19275 13219
rect 19677 13219 19735 13225
rect 19677 13216 19689 13219
rect 19263 13188 19689 13216
rect 19263 13185 19275 13188
rect 19217 13179 19275 13185
rect 19677 13185 19689 13188
rect 19723 13185 19735 13219
rect 19677 13179 19735 13185
rect 3132 13148 3160 13179
rect 3132 13120 3804 13148
rect 3776 13092 3804 13120
rect 3758 13040 3764 13092
rect 3816 13040 3822 13092
rect 1904 12922 20764 12944
rect 1904 12870 7110 12922
rect 7162 12870 7174 12922
rect 7226 12870 7238 12922
rect 7290 12870 7302 12922
rect 7354 12870 12438 12922
rect 12490 12870 12502 12922
rect 12554 12870 12566 12922
rect 12618 12870 12630 12922
rect 12682 12870 17766 12922
rect 17818 12870 17830 12922
rect 17882 12870 17894 12922
rect 17946 12870 17958 12922
rect 18010 12870 20764 12922
rect 1904 12848 20764 12870
rect 3758 12808 3764 12820
rect 3719 12780 3764 12808
rect 3758 12768 3764 12780
rect 3816 12768 3822 12820
rect 5969 12675 6027 12681
rect 5969 12672 5981 12675
rect 4236 12644 5981 12672
rect 4236 12613 4264 12644
rect 5969 12641 5981 12644
rect 6015 12641 6027 12675
rect 9281 12675 9339 12681
rect 9281 12672 9293 12675
rect 5969 12635 6027 12641
rect 6455 12644 7392 12672
rect 6455 12613 6483 12644
rect 3117 12607 3175 12613
rect 3117 12573 3129 12607
rect 3163 12573 3175 12607
rect 3117 12567 3175 12573
rect 4221 12607 4279 12613
rect 4221 12573 4233 12607
rect 4267 12573 4279 12607
rect 4221 12567 4279 12573
rect 5325 12607 5383 12613
rect 5325 12573 5337 12607
rect 5371 12573 5383 12607
rect 5325 12567 5383 12573
rect 6440 12607 6498 12613
rect 6440 12573 6452 12607
rect 6486 12573 6498 12607
rect 6440 12567 6498 12573
rect 3132 12536 3160 12567
rect 4865 12539 4923 12545
rect 4865 12536 4877 12539
rect 3132 12508 4877 12536
rect 4865 12505 4877 12508
rect 4911 12505 4923 12539
rect 5340 12536 5368 12567
rect 7073 12539 7131 12545
rect 7073 12536 7085 12539
rect 5340 12508 7085 12536
rect 4865 12499 4923 12505
rect 7073 12505 7085 12508
rect 7119 12505 7131 12539
rect 7364 12536 7392 12644
rect 7548 12644 9293 12672
rect 7548 12613 7576 12644
rect 9281 12641 9293 12644
rect 9327 12641 9339 12675
rect 10385 12675 10443 12681
rect 10385 12672 10397 12675
rect 9281 12635 9339 12641
rect 9572 12644 10397 12672
rect 7533 12607 7591 12613
rect 7533 12573 7545 12607
rect 7579 12573 7591 12607
rect 7533 12567 7591 12573
rect 8648 12607 8706 12613
rect 8648 12573 8660 12607
rect 8694 12573 8706 12607
rect 8648 12567 8706 12573
rect 8177 12539 8235 12545
rect 8177 12536 8189 12539
rect 7364 12508 8189 12536
rect 7073 12499 7131 12505
rect 8177 12505 8189 12508
rect 8223 12505 8235 12539
rect 8652 12536 8680 12567
rect 9572 12536 9600 12644
rect 10385 12641 10397 12644
rect 10431 12641 10443 12675
rect 11489 12675 11547 12681
rect 11489 12672 11501 12675
rect 10385 12635 10443 12641
rect 10584 12644 11501 12672
rect 9741 12607 9799 12613
rect 9741 12573 9753 12607
rect 9787 12604 9799 12607
rect 10584 12604 10612 12644
rect 11489 12641 11501 12644
rect 11535 12641 11547 12675
rect 13697 12675 13755 12681
rect 13697 12672 13709 12675
rect 11489 12635 11547 12641
rect 11964 12644 13709 12672
rect 11964 12613 11992 12644
rect 13697 12641 13709 12644
rect 13743 12641 13755 12675
rect 15905 12675 15963 12681
rect 15905 12672 15917 12675
rect 13697 12635 13755 12641
rect 14172 12644 15917 12672
rect 14172 12613 14200 12644
rect 15905 12641 15917 12644
rect 15951 12641 15963 12675
rect 18113 12675 18171 12681
rect 18113 12672 18125 12675
rect 15905 12635 15963 12641
rect 16380 12644 18125 12672
rect 16380 12613 16408 12644
rect 18113 12641 18125 12644
rect 18159 12641 18171 12675
rect 20321 12675 20379 12681
rect 20321 12672 20333 12675
rect 18113 12635 18171 12641
rect 18588 12644 20333 12672
rect 18588 12613 18616 12644
rect 20321 12641 20333 12644
rect 20367 12641 20379 12675
rect 20321 12635 20379 12641
rect 9787 12576 10612 12604
rect 10845 12607 10903 12613
rect 9787 12573 9799 12576
rect 9741 12567 9799 12573
rect 10845 12573 10857 12607
rect 10891 12573 10903 12607
rect 10845 12567 10903 12573
rect 11949 12607 12007 12613
rect 11949 12573 11961 12607
rect 11995 12573 12007 12607
rect 11949 12567 12007 12573
rect 13053 12607 13111 12613
rect 13053 12573 13065 12607
rect 13099 12573 13111 12607
rect 13053 12567 13111 12573
rect 14168 12607 14226 12613
rect 14168 12573 14180 12607
rect 14214 12573 14226 12607
rect 14168 12567 14226 12573
rect 15261 12607 15319 12613
rect 15261 12573 15273 12607
rect 15307 12573 15319 12607
rect 15261 12567 15319 12573
rect 16365 12607 16423 12613
rect 16365 12573 16377 12607
rect 16411 12573 16423 12607
rect 16365 12567 16423 12573
rect 17469 12607 17527 12613
rect 17469 12573 17481 12607
rect 17515 12573 17527 12607
rect 17469 12567 17527 12573
rect 18573 12607 18631 12613
rect 18573 12573 18585 12607
rect 18619 12573 18631 12607
rect 18573 12567 18631 12573
rect 19677 12607 19735 12613
rect 19677 12573 19689 12607
rect 19723 12604 19735 12607
rect 20134 12604 20140 12616
rect 19723 12576 20140 12604
rect 19723 12573 19735 12576
rect 19677 12567 19735 12573
rect 8652 12508 9600 12536
rect 10860 12536 10888 12567
rect 12593 12539 12651 12545
rect 12593 12536 12605 12539
rect 10860 12508 12605 12536
rect 8177 12499 8235 12505
rect 12593 12505 12605 12508
rect 12639 12505 12651 12539
rect 13068 12536 13096 12567
rect 14801 12539 14859 12545
rect 14801 12536 14813 12539
rect 13068 12508 14813 12536
rect 12593 12499 12651 12505
rect 14801 12505 14813 12508
rect 14847 12505 14859 12539
rect 15276 12536 15304 12567
rect 17009 12539 17067 12545
rect 17009 12536 17021 12539
rect 15276 12508 17021 12536
rect 14801 12499 14859 12505
rect 17009 12505 17021 12508
rect 17055 12505 17067 12539
rect 17484 12536 17512 12567
rect 20134 12564 20140 12576
rect 20192 12564 20198 12616
rect 19217 12539 19275 12545
rect 19217 12536 19229 12539
rect 17484 12508 19229 12536
rect 17009 12499 17067 12505
rect 19217 12505 19229 12508
rect 19263 12505 19275 12539
rect 19217 12499 19275 12505
rect 1904 12378 20764 12400
rect 1904 12326 4446 12378
rect 4498 12326 4510 12378
rect 4562 12326 4574 12378
rect 4626 12326 4638 12378
rect 4690 12326 9774 12378
rect 9826 12326 9838 12378
rect 9890 12326 9902 12378
rect 9954 12326 9966 12378
rect 10018 12326 15102 12378
rect 15154 12326 15166 12378
rect 15218 12326 15230 12378
rect 15282 12326 15294 12378
rect 15346 12326 20764 12378
rect 1904 12304 20764 12326
rect 20134 12224 20140 12276
rect 20192 12264 20198 12276
rect 20321 12267 20379 12273
rect 20321 12264 20333 12267
rect 20192 12236 20333 12264
rect 20192 12224 20198 12236
rect 20321 12233 20333 12236
rect 20367 12233 20379 12267
rect 20321 12227 20379 12233
rect 3117 12131 3175 12137
rect 3117 12097 3129 12131
rect 3163 12097 3175 12131
rect 3117 12091 3175 12097
rect 3761 12131 3819 12137
rect 3761 12097 3773 12131
rect 3807 12128 3819 12131
rect 4221 12131 4279 12137
rect 4221 12128 4233 12131
rect 3807 12100 4233 12128
rect 3807 12097 3819 12100
rect 3761 12091 3819 12097
rect 4221 12097 4233 12100
rect 4267 12097 4279 12131
rect 4221 12091 4279 12097
rect 4865 12131 4923 12137
rect 4865 12097 4877 12131
rect 4911 12128 4923 12131
rect 5325 12131 5383 12137
rect 5325 12128 5337 12131
rect 4911 12100 5337 12128
rect 4911 12097 4923 12100
rect 4865 12091 4923 12097
rect 5325 12097 5337 12100
rect 5371 12097 5383 12131
rect 5325 12091 5383 12097
rect 5969 12131 6027 12137
rect 5969 12097 5981 12131
rect 6015 12128 6027 12131
rect 6429 12131 6487 12137
rect 6429 12128 6441 12131
rect 6015 12100 6441 12128
rect 6015 12097 6027 12100
rect 5969 12091 6027 12097
rect 6429 12097 6441 12100
rect 6475 12097 6487 12131
rect 6429 12091 6487 12097
rect 7073 12131 7131 12137
rect 7073 12097 7085 12131
rect 7119 12128 7131 12131
rect 7533 12131 7591 12137
rect 7533 12128 7545 12131
rect 7119 12100 7545 12128
rect 7119 12097 7131 12100
rect 7073 12091 7131 12097
rect 7533 12097 7545 12100
rect 7579 12097 7591 12131
rect 7533 12091 7591 12097
rect 8177 12131 8235 12137
rect 8177 12097 8189 12131
rect 8223 12128 8235 12131
rect 8637 12131 8695 12137
rect 8637 12128 8649 12131
rect 8223 12100 8649 12128
rect 8223 12097 8235 12100
rect 8177 12091 8235 12097
rect 8637 12097 8649 12100
rect 8683 12097 8695 12131
rect 8637 12091 8695 12097
rect 9281 12131 9339 12137
rect 9281 12097 9293 12131
rect 9327 12128 9339 12131
rect 9741 12131 9799 12137
rect 9741 12128 9753 12131
rect 9327 12100 9753 12128
rect 9327 12097 9339 12100
rect 9281 12091 9339 12097
rect 9741 12097 9753 12100
rect 9787 12097 9799 12131
rect 9741 12091 9799 12097
rect 10385 12131 10443 12137
rect 10385 12097 10397 12131
rect 10431 12128 10443 12131
rect 10845 12131 10903 12137
rect 10845 12128 10857 12131
rect 10431 12100 10857 12128
rect 10431 12097 10443 12100
rect 10385 12091 10443 12097
rect 10845 12097 10857 12100
rect 10891 12097 10903 12131
rect 10845 12091 10903 12097
rect 11489 12131 11547 12137
rect 11489 12097 11501 12131
rect 11535 12128 11547 12131
rect 11949 12131 12007 12137
rect 11949 12128 11961 12131
rect 11535 12100 11961 12128
rect 11535 12097 11547 12100
rect 11489 12091 11547 12097
rect 11949 12097 11961 12100
rect 11995 12097 12007 12131
rect 11949 12091 12007 12097
rect 12593 12131 12651 12137
rect 12593 12097 12605 12131
rect 12639 12128 12651 12131
rect 13053 12131 13111 12137
rect 13053 12128 13065 12131
rect 12639 12100 13065 12128
rect 12639 12097 12651 12100
rect 12593 12091 12651 12097
rect 13053 12097 13065 12100
rect 13099 12097 13111 12131
rect 13053 12091 13111 12097
rect 13697 12131 13755 12137
rect 13697 12097 13709 12131
rect 13743 12128 13755 12131
rect 14157 12131 14215 12137
rect 14157 12128 14169 12131
rect 13743 12100 14169 12128
rect 13743 12097 13755 12100
rect 13697 12091 13755 12097
rect 14157 12097 14169 12100
rect 14203 12097 14215 12131
rect 14157 12091 14215 12097
rect 14801 12131 14859 12137
rect 14801 12097 14813 12131
rect 14847 12128 14859 12131
rect 15261 12131 15319 12137
rect 15261 12128 15273 12131
rect 14847 12100 15273 12128
rect 14847 12097 14859 12100
rect 14801 12091 14859 12097
rect 15261 12097 15273 12100
rect 15307 12097 15319 12131
rect 15261 12091 15319 12097
rect 15905 12131 15963 12137
rect 15905 12097 15917 12131
rect 15951 12128 15963 12131
rect 16365 12131 16423 12137
rect 16365 12128 16377 12131
rect 15951 12100 16377 12128
rect 15951 12097 15963 12100
rect 15905 12091 15963 12097
rect 16365 12097 16377 12100
rect 16411 12097 16423 12131
rect 16365 12091 16423 12097
rect 17009 12131 17067 12137
rect 17009 12097 17021 12131
rect 17055 12128 17067 12131
rect 17469 12131 17527 12137
rect 17469 12128 17481 12131
rect 17055 12100 17481 12128
rect 17055 12097 17067 12100
rect 17009 12091 17067 12097
rect 17469 12097 17481 12100
rect 17515 12097 17527 12131
rect 17469 12091 17527 12097
rect 18113 12131 18171 12137
rect 18113 12097 18125 12131
rect 18159 12128 18171 12131
rect 18573 12131 18631 12137
rect 18573 12128 18585 12131
rect 18159 12100 18585 12128
rect 18159 12097 18171 12100
rect 18113 12091 18171 12097
rect 18573 12097 18585 12100
rect 18619 12097 18631 12131
rect 18573 12091 18631 12097
rect 19217 12131 19275 12137
rect 19217 12097 19229 12131
rect 19263 12128 19275 12131
rect 19677 12131 19735 12137
rect 19677 12128 19689 12131
rect 19263 12100 19689 12128
rect 19263 12097 19275 12100
rect 19217 12091 19275 12097
rect 19677 12097 19689 12100
rect 19723 12097 19735 12131
rect 19677 12091 19735 12097
rect 3132 11992 3160 12091
rect 3758 11992 3764 12004
rect 3132 11964 3764 11992
rect 3758 11952 3764 11964
rect 3816 11952 3822 12004
rect 1904 11834 20764 11856
rect 1904 11782 7110 11834
rect 7162 11782 7174 11834
rect 7226 11782 7238 11834
rect 7290 11782 7302 11834
rect 7354 11782 12438 11834
rect 12490 11782 12502 11834
rect 12554 11782 12566 11834
rect 12618 11782 12630 11834
rect 12682 11782 17766 11834
rect 17818 11782 17830 11834
rect 17882 11782 17894 11834
rect 17946 11782 17958 11834
rect 18010 11782 20764 11834
rect 1904 11760 20764 11782
rect 3758 11584 3764 11596
rect 3719 11556 3764 11584
rect 3758 11544 3764 11556
rect 3816 11544 3822 11596
rect 4865 11587 4923 11593
rect 4865 11584 4877 11587
rect 3960 11556 4877 11584
rect 3117 11519 3175 11525
rect 3117 11485 3129 11519
rect 3163 11516 3175 11519
rect 3960 11516 3988 11556
rect 4865 11553 4877 11556
rect 4911 11553 4923 11587
rect 7073 11587 7131 11593
rect 7073 11584 7085 11587
rect 4865 11547 4923 11553
rect 5340 11556 7085 11584
rect 5340 11525 5368 11556
rect 7073 11553 7085 11556
rect 7119 11553 7131 11587
rect 8177 11587 8235 11593
rect 8177 11584 8189 11587
rect 7073 11547 7131 11553
rect 7364 11556 8189 11584
rect 3163 11488 3988 11516
rect 4221 11519 4279 11525
rect 3163 11485 3175 11488
rect 3117 11479 3175 11485
rect 4221 11485 4233 11519
rect 4267 11485 4279 11519
rect 4221 11479 4279 11485
rect 5325 11519 5383 11525
rect 5325 11485 5337 11519
rect 5371 11485 5383 11519
rect 5325 11479 5383 11485
rect 6440 11519 6498 11525
rect 6440 11485 6452 11519
rect 6486 11485 6498 11519
rect 6440 11479 6498 11485
rect 4236 11448 4264 11479
rect 5969 11451 6027 11457
rect 5969 11448 5981 11451
rect 4236 11420 5981 11448
rect 5969 11417 5981 11420
rect 6015 11417 6027 11451
rect 6444 11448 6472 11479
rect 7364 11448 7392 11556
rect 8177 11553 8189 11556
rect 8223 11553 8235 11587
rect 10385 11587 10443 11593
rect 10385 11584 10397 11587
rect 8177 11547 8235 11553
rect 8652 11556 10397 11584
rect 8652 11525 8680 11556
rect 10385 11553 10397 11556
rect 10431 11553 10443 11587
rect 12593 11587 12651 11593
rect 12593 11584 12605 11587
rect 10385 11547 10443 11553
rect 10860 11556 12605 11584
rect 10860 11525 10888 11556
rect 12593 11553 12605 11556
rect 12639 11553 12651 11587
rect 14801 11587 14859 11593
rect 14801 11584 14813 11587
rect 12593 11547 12651 11553
rect 13068 11556 14813 11584
rect 13068 11525 13096 11556
rect 14801 11553 14813 11556
rect 14847 11553 14859 11587
rect 17009 11587 17067 11593
rect 17009 11584 17021 11587
rect 14801 11547 14859 11553
rect 15276 11556 17021 11584
rect 15276 11525 15304 11556
rect 17009 11553 17021 11556
rect 17055 11553 17067 11587
rect 19217 11587 19275 11593
rect 19217 11584 19229 11587
rect 17009 11547 17067 11553
rect 17484 11556 19229 11584
rect 17484 11525 17512 11556
rect 19217 11553 19229 11556
rect 19263 11553 19275 11587
rect 19217 11547 19275 11553
rect 7533 11519 7591 11525
rect 7533 11485 7545 11519
rect 7579 11485 7591 11519
rect 7533 11479 7591 11485
rect 8648 11519 8706 11525
rect 8648 11485 8660 11519
rect 8694 11485 8706 11519
rect 8648 11479 8706 11485
rect 9741 11519 9799 11525
rect 9741 11485 9753 11519
rect 9787 11485 9799 11519
rect 9741 11479 9799 11485
rect 10845 11519 10903 11525
rect 10845 11485 10857 11519
rect 10891 11485 10903 11519
rect 10845 11479 10903 11485
rect 11949 11519 12007 11525
rect 11949 11485 11961 11519
rect 11995 11485 12007 11519
rect 11949 11479 12007 11485
rect 13053 11519 13111 11525
rect 13053 11485 13065 11519
rect 13099 11485 13111 11519
rect 13053 11479 13111 11485
rect 14168 11519 14226 11525
rect 14168 11485 14180 11519
rect 14214 11485 14226 11519
rect 14168 11479 14226 11485
rect 15261 11519 15319 11525
rect 15261 11485 15273 11519
rect 15307 11485 15319 11519
rect 15261 11479 15319 11485
rect 16365 11519 16423 11525
rect 16365 11485 16377 11519
rect 16411 11485 16423 11519
rect 16365 11479 16423 11485
rect 17469 11519 17527 11525
rect 17469 11485 17481 11519
rect 17515 11485 17527 11519
rect 17469 11479 17527 11485
rect 18573 11519 18631 11525
rect 18573 11485 18585 11519
rect 18619 11485 18631 11519
rect 19674 11516 19680 11528
rect 19635 11488 19680 11516
rect 18573 11479 18631 11485
rect 6444 11420 7392 11448
rect 7548 11448 7576 11479
rect 9281 11451 9339 11457
rect 9281 11448 9293 11451
rect 7548 11420 9293 11448
rect 5969 11411 6027 11417
rect 9281 11417 9293 11420
rect 9327 11417 9339 11451
rect 9756 11448 9784 11479
rect 11489 11451 11547 11457
rect 11489 11448 11501 11451
rect 9756 11420 11501 11448
rect 9281 11411 9339 11417
rect 11489 11417 11501 11420
rect 11535 11417 11547 11451
rect 11964 11448 11992 11479
rect 13697 11451 13755 11457
rect 13697 11448 13709 11451
rect 11964 11420 13709 11448
rect 11489 11411 11547 11417
rect 13697 11417 13709 11420
rect 13743 11417 13755 11451
rect 14172 11448 14200 11479
rect 15905 11451 15963 11457
rect 15905 11448 15917 11451
rect 14172 11420 15917 11448
rect 13697 11411 13755 11417
rect 15905 11417 15917 11420
rect 15951 11417 15963 11451
rect 16380 11448 16408 11479
rect 18113 11451 18171 11457
rect 18113 11448 18125 11451
rect 16380 11420 18125 11448
rect 15905 11411 15963 11417
rect 18113 11417 18125 11420
rect 18159 11417 18171 11451
rect 18588 11448 18616 11479
rect 19674 11476 19680 11488
rect 19732 11476 19738 11528
rect 20321 11451 20379 11457
rect 20321 11448 20333 11451
rect 18588 11420 20333 11448
rect 18113 11411 18171 11417
rect 20321 11417 20333 11420
rect 20367 11417 20379 11451
rect 20321 11411 20379 11417
rect 1904 11290 20764 11312
rect 1904 11238 4446 11290
rect 4498 11238 4510 11290
rect 4562 11238 4574 11290
rect 4626 11238 4638 11290
rect 4690 11238 9774 11290
rect 9826 11238 9838 11290
rect 9890 11238 9902 11290
rect 9954 11238 9966 11290
rect 10018 11238 15102 11290
rect 15154 11238 15166 11290
rect 15218 11238 15230 11290
rect 15282 11238 15294 11290
rect 15346 11238 20764 11290
rect 1904 11216 20764 11238
rect 19674 11136 19680 11188
rect 19732 11176 19738 11188
rect 20321 11179 20379 11185
rect 20321 11176 20333 11179
rect 19732 11148 20333 11176
rect 19732 11136 19738 11148
rect 20321 11145 20333 11148
rect 20367 11145 20379 11179
rect 20321 11139 20379 11145
rect 3117 11043 3175 11049
rect 3117 11009 3129 11043
rect 3163 11009 3175 11043
rect 3117 11003 3175 11009
rect 3761 11043 3819 11049
rect 3761 11009 3773 11043
rect 3807 11040 3819 11043
rect 4221 11043 4279 11049
rect 4221 11040 4233 11043
rect 3807 11012 4233 11040
rect 3807 11009 3819 11012
rect 3761 11003 3819 11009
rect 4221 11009 4233 11012
rect 4267 11009 4279 11043
rect 4221 11003 4279 11009
rect 4865 11043 4923 11049
rect 4865 11009 4877 11043
rect 4911 11040 4923 11043
rect 5325 11043 5383 11049
rect 5325 11040 5337 11043
rect 4911 11012 5337 11040
rect 4911 11009 4923 11012
rect 4865 11003 4923 11009
rect 5325 11009 5337 11012
rect 5371 11009 5383 11043
rect 5325 11003 5383 11009
rect 5969 11043 6027 11049
rect 5969 11009 5981 11043
rect 6015 11040 6027 11043
rect 6429 11043 6487 11049
rect 6429 11040 6441 11043
rect 6015 11012 6441 11040
rect 6015 11009 6027 11012
rect 5969 11003 6027 11009
rect 6429 11009 6441 11012
rect 6475 11009 6487 11043
rect 6429 11003 6487 11009
rect 7073 11043 7131 11049
rect 7073 11009 7085 11043
rect 7119 11040 7131 11043
rect 7533 11043 7591 11049
rect 7533 11040 7545 11043
rect 7119 11012 7545 11040
rect 7119 11009 7131 11012
rect 7073 11003 7131 11009
rect 7533 11009 7545 11012
rect 7579 11009 7591 11043
rect 7533 11003 7591 11009
rect 8177 11043 8235 11049
rect 8177 11009 8189 11043
rect 8223 11040 8235 11043
rect 8637 11043 8695 11049
rect 8637 11040 8649 11043
rect 8223 11012 8649 11040
rect 8223 11009 8235 11012
rect 8177 11003 8235 11009
rect 8637 11009 8649 11012
rect 8683 11009 8695 11043
rect 8637 11003 8695 11009
rect 9281 11043 9339 11049
rect 9281 11009 9293 11043
rect 9327 11040 9339 11043
rect 9741 11043 9799 11049
rect 9741 11040 9753 11043
rect 9327 11012 9753 11040
rect 9327 11009 9339 11012
rect 9281 11003 9339 11009
rect 9741 11009 9753 11012
rect 9787 11009 9799 11043
rect 9741 11003 9799 11009
rect 10385 11043 10443 11049
rect 10385 11009 10397 11043
rect 10431 11040 10443 11043
rect 10845 11043 10903 11049
rect 10845 11040 10857 11043
rect 10431 11012 10857 11040
rect 10431 11009 10443 11012
rect 10385 11003 10443 11009
rect 10845 11009 10857 11012
rect 10891 11009 10903 11043
rect 10845 11003 10903 11009
rect 11489 11043 11547 11049
rect 11489 11009 11501 11043
rect 11535 11040 11547 11043
rect 11949 11043 12007 11049
rect 11949 11040 11961 11043
rect 11535 11012 11961 11040
rect 11535 11009 11547 11012
rect 11489 11003 11547 11009
rect 11949 11009 11961 11012
rect 11995 11009 12007 11043
rect 11949 11003 12007 11009
rect 12593 11043 12651 11049
rect 12593 11009 12605 11043
rect 12639 11040 12651 11043
rect 13053 11043 13111 11049
rect 13053 11040 13065 11043
rect 12639 11012 13065 11040
rect 12639 11009 12651 11012
rect 12593 11003 12651 11009
rect 13053 11009 13065 11012
rect 13099 11009 13111 11043
rect 13053 11003 13111 11009
rect 13697 11043 13755 11049
rect 13697 11009 13709 11043
rect 13743 11040 13755 11043
rect 14157 11043 14215 11049
rect 14157 11040 14169 11043
rect 13743 11012 14169 11040
rect 13743 11009 13755 11012
rect 13697 11003 13755 11009
rect 14157 11009 14169 11012
rect 14203 11009 14215 11043
rect 14157 11003 14215 11009
rect 14801 11043 14859 11049
rect 14801 11009 14813 11043
rect 14847 11040 14859 11043
rect 15261 11043 15319 11049
rect 15261 11040 15273 11043
rect 14847 11012 15273 11040
rect 14847 11009 14859 11012
rect 14801 11003 14859 11009
rect 15261 11009 15273 11012
rect 15307 11009 15319 11043
rect 15261 11003 15319 11009
rect 15905 11043 15963 11049
rect 15905 11009 15917 11043
rect 15951 11040 15963 11043
rect 16365 11043 16423 11049
rect 16365 11040 16377 11043
rect 15951 11012 16377 11040
rect 15951 11009 15963 11012
rect 15905 11003 15963 11009
rect 16365 11009 16377 11012
rect 16411 11009 16423 11043
rect 16365 11003 16423 11009
rect 17009 11043 17067 11049
rect 17009 11009 17021 11043
rect 17055 11040 17067 11043
rect 17469 11043 17527 11049
rect 17469 11040 17481 11043
rect 17055 11012 17481 11040
rect 17055 11009 17067 11012
rect 17009 11003 17067 11009
rect 17469 11009 17481 11012
rect 17515 11009 17527 11043
rect 17469 11003 17527 11009
rect 18113 11043 18171 11049
rect 18113 11009 18125 11043
rect 18159 11040 18171 11043
rect 18573 11043 18631 11049
rect 18573 11040 18585 11043
rect 18159 11012 18585 11040
rect 18159 11009 18171 11012
rect 18113 11003 18171 11009
rect 18573 11009 18585 11012
rect 18619 11009 18631 11043
rect 18573 11003 18631 11009
rect 19217 11043 19275 11049
rect 19217 11009 19229 11043
rect 19263 11040 19275 11043
rect 19677 11043 19735 11049
rect 19677 11040 19689 11043
rect 19263 11012 19689 11040
rect 19263 11009 19275 11012
rect 19217 11003 19275 11009
rect 19677 11009 19689 11012
rect 19723 11009 19735 11043
rect 19677 11003 19735 11009
rect 3132 10904 3160 11003
rect 3758 10904 3764 10916
rect 3132 10876 3764 10904
rect 3758 10864 3764 10876
rect 3816 10864 3822 10916
rect 1904 10746 20764 10768
rect 1904 10694 7110 10746
rect 7162 10694 7174 10746
rect 7226 10694 7238 10746
rect 7290 10694 7302 10746
rect 7354 10694 12438 10746
rect 12490 10694 12502 10746
rect 12554 10694 12566 10746
rect 12618 10694 12630 10746
rect 12682 10694 17766 10746
rect 17818 10694 17830 10746
rect 17882 10694 17894 10746
rect 17946 10694 17958 10746
rect 18010 10694 20764 10746
rect 1904 10672 20764 10694
rect 3758 10632 3764 10644
rect 3719 10604 3764 10632
rect 3758 10592 3764 10604
rect 3816 10592 3822 10644
rect 4865 10499 4923 10505
rect 4865 10496 4877 10499
rect 3132 10468 4877 10496
rect 3132 10437 3160 10468
rect 4865 10465 4877 10468
rect 4911 10465 4923 10499
rect 7073 10499 7131 10505
rect 7073 10496 7085 10499
rect 4865 10459 4923 10465
rect 5340 10468 7085 10496
rect 5340 10437 5368 10468
rect 7073 10465 7085 10468
rect 7119 10465 7131 10499
rect 9281 10499 9339 10505
rect 9281 10496 9293 10499
rect 7073 10459 7131 10465
rect 7548 10468 9293 10496
rect 7548 10437 7576 10468
rect 9281 10465 9293 10468
rect 9327 10465 9339 10499
rect 10385 10499 10443 10505
rect 10385 10496 10397 10499
rect 9281 10459 9339 10465
rect 9572 10468 10397 10496
rect 3117 10431 3175 10437
rect 3117 10397 3129 10431
rect 3163 10397 3175 10431
rect 3117 10391 3175 10397
rect 4221 10431 4279 10437
rect 4221 10397 4233 10431
rect 4267 10397 4279 10431
rect 4221 10391 4279 10397
rect 5325 10431 5383 10437
rect 5325 10397 5337 10431
rect 5371 10397 5383 10431
rect 5325 10391 5383 10397
rect 6440 10431 6498 10437
rect 6440 10397 6452 10431
rect 6486 10397 6498 10431
rect 6440 10391 6498 10397
rect 7533 10431 7591 10437
rect 7533 10397 7545 10431
rect 7579 10397 7591 10431
rect 7533 10391 7591 10397
rect 8648 10431 8706 10437
rect 8648 10397 8660 10431
rect 8694 10397 8706 10431
rect 8648 10391 8706 10397
rect 4236 10360 4264 10391
rect 5969 10363 6027 10369
rect 5969 10360 5981 10363
rect 4236 10332 5981 10360
rect 5969 10329 5981 10332
rect 6015 10329 6027 10363
rect 6444 10360 6472 10391
rect 8177 10363 8235 10369
rect 8177 10360 8189 10363
rect 6444 10332 8189 10360
rect 5969 10323 6027 10329
rect 8177 10329 8189 10332
rect 8223 10329 8235 10363
rect 8652 10360 8680 10391
rect 9572 10360 9600 10468
rect 10385 10465 10397 10468
rect 10431 10465 10443 10499
rect 11489 10499 11547 10505
rect 11489 10496 11501 10499
rect 10385 10459 10443 10465
rect 10584 10468 11501 10496
rect 9741 10431 9799 10437
rect 9741 10397 9753 10431
rect 9787 10428 9799 10431
rect 10584 10428 10612 10468
rect 11489 10465 11501 10468
rect 11535 10465 11547 10499
rect 13697 10499 13755 10505
rect 13697 10496 13709 10499
rect 11489 10459 11547 10465
rect 11964 10468 13709 10496
rect 11964 10437 11992 10468
rect 13697 10465 13709 10468
rect 13743 10465 13755 10499
rect 17009 10499 17067 10505
rect 17009 10496 17021 10499
rect 13697 10459 13755 10465
rect 14172 10468 15212 10496
rect 14172 10437 14200 10468
rect 9787 10400 10612 10428
rect 10845 10431 10903 10437
rect 9787 10397 9799 10400
rect 9741 10391 9799 10397
rect 10845 10397 10857 10431
rect 10891 10397 10903 10431
rect 10845 10391 10903 10397
rect 11949 10431 12007 10437
rect 11949 10397 11961 10431
rect 11995 10397 12007 10431
rect 11949 10391 12007 10397
rect 13053 10431 13111 10437
rect 13053 10397 13065 10431
rect 13099 10397 13111 10431
rect 13053 10391 13111 10397
rect 14168 10431 14226 10437
rect 14168 10397 14180 10431
rect 14214 10397 14226 10431
rect 14168 10391 14226 10397
rect 8652 10332 9600 10360
rect 10860 10360 10888 10391
rect 12593 10363 12651 10369
rect 12593 10360 12605 10363
rect 10860 10332 12605 10360
rect 8177 10323 8235 10329
rect 12593 10329 12605 10332
rect 12639 10329 12651 10363
rect 13068 10360 13096 10391
rect 14801 10363 14859 10369
rect 14801 10360 14813 10363
rect 13068 10332 14813 10360
rect 12593 10323 12651 10329
rect 14801 10329 14813 10332
rect 14847 10329 14859 10363
rect 15184 10360 15212 10468
rect 15276 10468 17021 10496
rect 15276 10437 15304 10468
rect 17009 10465 17021 10468
rect 17055 10465 17067 10499
rect 19217 10499 19275 10505
rect 19217 10496 19229 10499
rect 17009 10459 17067 10465
rect 17484 10468 19229 10496
rect 17484 10437 17512 10468
rect 19217 10465 19229 10468
rect 19263 10465 19275 10499
rect 19217 10459 19275 10465
rect 15261 10431 15319 10437
rect 15261 10397 15273 10431
rect 15307 10397 15319 10431
rect 15261 10391 15319 10397
rect 16365 10431 16423 10437
rect 16365 10397 16377 10431
rect 16411 10397 16423 10431
rect 16365 10391 16423 10397
rect 17469 10431 17527 10437
rect 17469 10397 17481 10431
rect 17515 10397 17527 10431
rect 17469 10391 17527 10397
rect 18573 10431 18631 10437
rect 18573 10397 18585 10431
rect 18619 10397 18631 10431
rect 18573 10391 18631 10397
rect 19677 10431 19735 10437
rect 19677 10397 19689 10431
rect 19723 10428 19735 10431
rect 20134 10428 20140 10440
rect 19723 10400 20140 10428
rect 19723 10397 19735 10400
rect 19677 10391 19735 10397
rect 15905 10363 15963 10369
rect 15905 10360 15917 10363
rect 15184 10332 15917 10360
rect 14801 10323 14859 10329
rect 15905 10329 15917 10332
rect 15951 10329 15963 10363
rect 16380 10360 16408 10391
rect 18113 10363 18171 10369
rect 18113 10360 18125 10363
rect 16380 10332 18125 10360
rect 15905 10323 15963 10329
rect 18113 10329 18125 10332
rect 18159 10329 18171 10363
rect 18588 10360 18616 10391
rect 20134 10388 20140 10400
rect 20192 10388 20198 10440
rect 20321 10363 20379 10369
rect 20321 10360 20333 10363
rect 18588 10332 20333 10360
rect 18113 10323 18171 10329
rect 20321 10329 20333 10332
rect 20367 10329 20379 10363
rect 20321 10323 20379 10329
rect 1904 10202 20764 10224
rect 1904 10150 4446 10202
rect 4498 10150 4510 10202
rect 4562 10150 4574 10202
rect 4626 10150 4638 10202
rect 4690 10150 9774 10202
rect 9826 10150 9838 10202
rect 9890 10150 9902 10202
rect 9954 10150 9966 10202
rect 10018 10150 15102 10202
rect 15154 10150 15166 10202
rect 15218 10150 15230 10202
rect 15282 10150 15294 10202
rect 15346 10150 20764 10202
rect 1904 10128 20764 10150
rect 20134 10048 20140 10100
rect 20192 10088 20198 10100
rect 20321 10091 20379 10097
rect 20321 10088 20333 10091
rect 20192 10060 20333 10088
rect 20192 10048 20198 10060
rect 20321 10057 20333 10060
rect 20367 10057 20379 10091
rect 20321 10051 20379 10057
rect 2286 9912 2292 9964
rect 2344 9952 2350 9964
rect 3117 9955 3175 9961
rect 3117 9952 3129 9955
rect 2344 9924 3129 9952
rect 2344 9912 2350 9924
rect 3117 9921 3129 9924
rect 3163 9921 3175 9955
rect 3117 9915 3175 9921
rect 3761 9955 3819 9961
rect 3761 9921 3773 9955
rect 3807 9952 3819 9955
rect 4221 9955 4279 9961
rect 4221 9952 4233 9955
rect 3807 9924 4233 9952
rect 3807 9921 3819 9924
rect 3761 9915 3819 9921
rect 4221 9921 4233 9924
rect 4267 9921 4279 9955
rect 4221 9915 4279 9921
rect 4865 9955 4923 9961
rect 4865 9921 4877 9955
rect 4911 9952 4923 9955
rect 5325 9955 5383 9961
rect 5325 9952 5337 9955
rect 4911 9924 5337 9952
rect 4911 9921 4923 9924
rect 4865 9915 4923 9921
rect 5325 9921 5337 9924
rect 5371 9921 5383 9955
rect 5325 9915 5383 9921
rect 5969 9955 6027 9961
rect 5969 9921 5981 9955
rect 6015 9952 6027 9955
rect 6429 9955 6487 9961
rect 6429 9952 6441 9955
rect 6015 9924 6441 9952
rect 6015 9921 6027 9924
rect 5969 9915 6027 9921
rect 6429 9921 6441 9924
rect 6475 9921 6487 9955
rect 6429 9915 6487 9921
rect 7073 9955 7131 9961
rect 7073 9921 7085 9955
rect 7119 9952 7131 9955
rect 7533 9955 7591 9961
rect 7533 9952 7545 9955
rect 7119 9924 7545 9952
rect 7119 9921 7131 9924
rect 7073 9915 7131 9921
rect 7533 9921 7545 9924
rect 7579 9921 7591 9955
rect 7533 9915 7591 9921
rect 8177 9955 8235 9961
rect 8177 9921 8189 9955
rect 8223 9952 8235 9955
rect 8637 9955 8695 9961
rect 8637 9952 8649 9955
rect 8223 9924 8649 9952
rect 8223 9921 8235 9924
rect 8177 9915 8235 9921
rect 8637 9921 8649 9924
rect 8683 9921 8695 9955
rect 8637 9915 8695 9921
rect 9281 9955 9339 9961
rect 9281 9921 9293 9955
rect 9327 9952 9339 9955
rect 9741 9955 9799 9961
rect 9741 9952 9753 9955
rect 9327 9924 9753 9952
rect 9327 9921 9339 9924
rect 9281 9915 9339 9921
rect 9741 9921 9753 9924
rect 9787 9921 9799 9955
rect 9741 9915 9799 9921
rect 10385 9955 10443 9961
rect 10385 9921 10397 9955
rect 10431 9952 10443 9955
rect 10845 9955 10903 9961
rect 10845 9952 10857 9955
rect 10431 9924 10857 9952
rect 10431 9921 10443 9924
rect 10385 9915 10443 9921
rect 10845 9921 10857 9924
rect 10891 9921 10903 9955
rect 10845 9915 10903 9921
rect 11489 9955 11547 9961
rect 11489 9921 11501 9955
rect 11535 9952 11547 9955
rect 11949 9955 12007 9961
rect 11949 9952 11961 9955
rect 11535 9924 11961 9952
rect 11535 9921 11547 9924
rect 11489 9915 11547 9921
rect 11949 9921 11961 9924
rect 11995 9921 12007 9955
rect 11949 9915 12007 9921
rect 12593 9955 12651 9961
rect 12593 9921 12605 9955
rect 12639 9952 12651 9955
rect 13053 9955 13111 9961
rect 13053 9952 13065 9955
rect 12639 9924 13065 9952
rect 12639 9921 12651 9924
rect 12593 9915 12651 9921
rect 13053 9921 13065 9924
rect 13099 9921 13111 9955
rect 13053 9915 13111 9921
rect 13697 9955 13755 9961
rect 13697 9921 13709 9955
rect 13743 9952 13755 9955
rect 14157 9955 14215 9961
rect 14157 9952 14169 9955
rect 13743 9924 14169 9952
rect 13743 9921 13755 9924
rect 13697 9915 13755 9921
rect 14157 9921 14169 9924
rect 14203 9921 14215 9955
rect 14157 9915 14215 9921
rect 14801 9955 14859 9961
rect 14801 9921 14813 9955
rect 14847 9952 14859 9955
rect 15261 9955 15319 9961
rect 15261 9952 15273 9955
rect 14847 9924 15273 9952
rect 14847 9921 14859 9924
rect 14801 9915 14859 9921
rect 15261 9921 15273 9924
rect 15307 9921 15319 9955
rect 15261 9915 15319 9921
rect 15905 9955 15963 9961
rect 15905 9921 15917 9955
rect 15951 9952 15963 9955
rect 16365 9955 16423 9961
rect 16365 9952 16377 9955
rect 15951 9924 16377 9952
rect 15951 9921 15963 9924
rect 15905 9915 15963 9921
rect 16365 9921 16377 9924
rect 16411 9921 16423 9955
rect 16365 9915 16423 9921
rect 17009 9955 17067 9961
rect 17009 9921 17021 9955
rect 17055 9952 17067 9955
rect 17469 9955 17527 9961
rect 17469 9952 17481 9955
rect 17055 9924 17481 9952
rect 17055 9921 17067 9924
rect 17009 9915 17067 9921
rect 17469 9921 17481 9924
rect 17515 9921 17527 9955
rect 17469 9915 17527 9921
rect 18113 9955 18171 9961
rect 18113 9921 18125 9955
rect 18159 9952 18171 9955
rect 18573 9955 18631 9961
rect 18573 9952 18585 9955
rect 18159 9924 18585 9952
rect 18159 9921 18171 9924
rect 18113 9915 18171 9921
rect 18573 9921 18585 9924
rect 18619 9921 18631 9955
rect 18573 9915 18631 9921
rect 19217 9955 19275 9961
rect 19217 9921 19229 9955
rect 19263 9952 19275 9955
rect 19677 9955 19735 9961
rect 19677 9952 19689 9955
rect 19263 9924 19689 9952
rect 19263 9921 19275 9924
rect 19217 9915 19275 9921
rect 19677 9921 19689 9924
rect 19723 9921 19735 9955
rect 19677 9915 19735 9921
rect 1904 9658 20764 9680
rect 1904 9606 7110 9658
rect 7162 9606 7174 9658
rect 7226 9606 7238 9658
rect 7290 9606 7302 9658
rect 7354 9606 12438 9658
rect 12490 9606 12502 9658
rect 12554 9606 12566 9658
rect 12618 9606 12630 9658
rect 12682 9606 17766 9658
rect 17818 9606 17830 9658
rect 17882 9606 17894 9658
rect 17946 9606 17958 9658
rect 18010 9606 20764 9658
rect 1904 9584 20764 9606
rect 2470 9408 2476 9420
rect 2431 9380 2476 9408
rect 2470 9368 2476 9380
rect 2528 9368 2534 9420
rect 5969 9411 6027 9417
rect 5969 9408 5981 9411
rect 4236 9380 5981 9408
rect 2286 9300 2292 9352
rect 2344 9300 2350 9352
rect 4236 9349 4264 9380
rect 5969 9377 5981 9380
rect 6015 9377 6027 9411
rect 8177 9411 8235 9417
rect 8177 9408 8189 9411
rect 5969 9371 6027 9377
rect 6444 9380 8189 9408
rect 6444 9349 6472 9380
rect 8177 9377 8189 9380
rect 8223 9377 8235 9411
rect 10385 9411 10443 9417
rect 10385 9408 10397 9411
rect 8177 9371 8235 9377
rect 8652 9380 10397 9408
rect 8652 9349 8680 9380
rect 10385 9377 10397 9380
rect 10431 9377 10443 9411
rect 11489 9411 11547 9417
rect 11489 9408 11501 9411
rect 10385 9371 10443 9377
rect 10584 9380 11501 9408
rect 3117 9343 3175 9349
rect 3117 9309 3129 9343
rect 3163 9340 3175 9343
rect 4221 9343 4279 9349
rect 3163 9312 3896 9340
rect 3163 9309 3175 9312
rect 3117 9303 3175 9309
rect 2304 9272 2332 9300
rect 1936 9244 2332 9272
rect 2381 9275 2439 9281
rect 1936 9213 1964 9244
rect 2381 9241 2393 9275
rect 2427 9272 2439 9275
rect 3761 9275 3819 9281
rect 3761 9272 3773 9275
rect 2427 9244 3773 9272
rect 2427 9241 2439 9244
rect 2381 9235 2439 9241
rect 3761 9241 3773 9244
rect 3807 9241 3819 9275
rect 3868 9272 3896 9312
rect 4221 9309 4233 9343
rect 4267 9309 4279 9343
rect 4221 9303 4279 9309
rect 5325 9343 5383 9349
rect 5325 9309 5337 9343
rect 5371 9309 5383 9343
rect 5325 9303 5383 9309
rect 6440 9343 6498 9349
rect 6440 9309 6452 9343
rect 6486 9309 6498 9343
rect 6440 9303 6498 9309
rect 7533 9343 7591 9349
rect 7533 9309 7545 9343
rect 7579 9309 7591 9343
rect 7533 9303 7591 9309
rect 8648 9343 8706 9349
rect 8648 9309 8660 9343
rect 8694 9309 8706 9343
rect 8648 9303 8706 9309
rect 9741 9343 9799 9349
rect 9741 9309 9753 9343
rect 9787 9340 9799 9343
rect 10584 9340 10612 9380
rect 11489 9377 11501 9380
rect 11535 9377 11547 9411
rect 13697 9411 13755 9417
rect 13697 9408 13709 9411
rect 11489 9371 11547 9377
rect 11964 9380 13709 9408
rect 11964 9349 11992 9380
rect 13697 9377 13709 9380
rect 13743 9377 13755 9411
rect 17009 9411 17067 9417
rect 17009 9408 17021 9411
rect 13697 9371 13755 9377
rect 14172 9380 14936 9408
rect 14172 9349 14200 9380
rect 9787 9312 10612 9340
rect 10845 9343 10903 9349
rect 9787 9309 9799 9312
rect 9741 9303 9799 9309
rect 10845 9309 10857 9343
rect 10891 9309 10903 9343
rect 10845 9303 10903 9309
rect 11949 9343 12007 9349
rect 11949 9309 11961 9343
rect 11995 9309 12007 9343
rect 11949 9303 12007 9309
rect 13053 9343 13111 9349
rect 13053 9309 13065 9343
rect 13099 9309 13111 9343
rect 13053 9303 13111 9309
rect 14168 9343 14226 9349
rect 14168 9309 14180 9343
rect 14214 9309 14226 9343
rect 14168 9303 14226 9309
rect 4865 9275 4923 9281
rect 4865 9272 4877 9275
rect 3868 9244 4877 9272
rect 3761 9235 3819 9241
rect 4865 9241 4877 9244
rect 4911 9241 4923 9275
rect 5340 9272 5368 9303
rect 7073 9275 7131 9281
rect 7073 9272 7085 9275
rect 5340 9244 7085 9272
rect 4865 9235 4923 9241
rect 7073 9241 7085 9244
rect 7119 9241 7131 9275
rect 7548 9272 7576 9303
rect 9281 9275 9339 9281
rect 9281 9272 9293 9275
rect 7548 9244 9293 9272
rect 7073 9235 7131 9241
rect 9281 9241 9293 9244
rect 9327 9241 9339 9275
rect 10860 9272 10888 9303
rect 12593 9275 12651 9281
rect 12593 9272 12605 9275
rect 10860 9244 12605 9272
rect 9281 9235 9339 9241
rect 12593 9241 12605 9244
rect 12639 9241 12651 9275
rect 13068 9272 13096 9303
rect 14801 9275 14859 9281
rect 14801 9272 14813 9275
rect 13068 9244 14813 9272
rect 12593 9235 12651 9241
rect 14801 9241 14813 9244
rect 14847 9241 14859 9275
rect 14908 9272 14936 9380
rect 15276 9380 17021 9408
rect 15276 9349 15304 9380
rect 17009 9377 17021 9380
rect 17055 9377 17067 9411
rect 19217 9411 19275 9417
rect 19217 9408 19229 9411
rect 17009 9371 17067 9377
rect 17484 9380 19229 9408
rect 17484 9349 17512 9380
rect 19217 9377 19229 9380
rect 19263 9377 19275 9411
rect 19217 9371 19275 9377
rect 15261 9343 15319 9349
rect 15261 9309 15273 9343
rect 15307 9309 15319 9343
rect 15261 9303 15319 9309
rect 16365 9343 16423 9349
rect 16365 9309 16377 9343
rect 16411 9309 16423 9343
rect 16365 9303 16423 9309
rect 17469 9343 17527 9349
rect 17469 9309 17481 9343
rect 17515 9309 17527 9343
rect 17469 9303 17527 9309
rect 18573 9343 18631 9349
rect 18573 9309 18585 9343
rect 18619 9309 18631 9343
rect 19674 9340 19680 9352
rect 19635 9312 19680 9340
rect 18573 9303 18631 9309
rect 15905 9275 15963 9281
rect 15905 9272 15917 9275
rect 14908 9244 15917 9272
rect 14801 9235 14859 9241
rect 15905 9241 15917 9244
rect 15951 9241 15963 9275
rect 16380 9272 16408 9303
rect 18113 9275 18171 9281
rect 18113 9272 18125 9275
rect 16380 9244 18125 9272
rect 15905 9235 15963 9241
rect 18113 9241 18125 9244
rect 18159 9241 18171 9275
rect 18588 9272 18616 9303
rect 19674 9300 19680 9312
rect 19732 9300 19738 9352
rect 20321 9275 20379 9281
rect 20321 9272 20333 9275
rect 18588 9244 20333 9272
rect 18113 9235 18171 9241
rect 20321 9241 20333 9244
rect 20367 9241 20379 9275
rect 20321 9235 20379 9241
rect 1921 9207 1979 9213
rect 1921 9173 1933 9207
rect 1967 9173 1979 9207
rect 1921 9167 1979 9173
rect 2286 9164 2292 9216
rect 2344 9204 2350 9216
rect 2344 9176 2389 9204
rect 2344 9164 2350 9176
rect 1904 9114 20764 9136
rect 1904 9062 4446 9114
rect 4498 9062 4510 9114
rect 4562 9062 4574 9114
rect 4626 9062 4638 9114
rect 4690 9062 9774 9114
rect 9826 9062 9838 9114
rect 9890 9062 9902 9114
rect 9954 9062 9966 9114
rect 10018 9062 15102 9114
rect 15154 9062 15166 9114
rect 15218 9062 15230 9114
rect 15282 9062 15294 9114
rect 15346 9062 20764 9114
rect 1904 9040 20764 9062
rect 19674 8960 19680 9012
rect 19732 9000 19738 9012
rect 20321 9003 20379 9009
rect 20321 9000 20333 9003
rect 19732 8972 20333 9000
rect 19732 8960 19738 8972
rect 20321 8969 20333 8972
rect 20367 8969 20379 9003
rect 20321 8963 20379 8969
rect 3117 8867 3175 8873
rect 3117 8833 3129 8867
rect 3163 8833 3175 8867
rect 3117 8827 3175 8833
rect 3761 8867 3819 8873
rect 3761 8833 3773 8867
rect 3807 8864 3819 8867
rect 4221 8867 4279 8873
rect 4221 8864 4233 8867
rect 3807 8836 4233 8864
rect 3807 8833 3819 8836
rect 3761 8827 3819 8833
rect 4221 8833 4233 8836
rect 4267 8833 4279 8867
rect 4221 8827 4279 8833
rect 4865 8867 4923 8873
rect 4865 8833 4877 8867
rect 4911 8864 4923 8867
rect 5325 8867 5383 8873
rect 5325 8864 5337 8867
rect 4911 8836 5337 8864
rect 4911 8833 4923 8836
rect 4865 8827 4923 8833
rect 5325 8833 5337 8836
rect 5371 8833 5383 8867
rect 5325 8827 5383 8833
rect 5969 8867 6027 8873
rect 5969 8833 5981 8867
rect 6015 8864 6027 8867
rect 6429 8867 6487 8873
rect 6429 8864 6441 8867
rect 6015 8836 6441 8864
rect 6015 8833 6027 8836
rect 5969 8827 6027 8833
rect 6429 8833 6441 8836
rect 6475 8833 6487 8867
rect 6429 8827 6487 8833
rect 7073 8867 7131 8873
rect 7073 8833 7085 8867
rect 7119 8864 7131 8867
rect 7533 8867 7591 8873
rect 7533 8864 7545 8867
rect 7119 8836 7545 8864
rect 7119 8833 7131 8836
rect 7073 8827 7131 8833
rect 7533 8833 7545 8836
rect 7579 8833 7591 8867
rect 7533 8827 7591 8833
rect 8177 8867 8235 8873
rect 8177 8833 8189 8867
rect 8223 8864 8235 8867
rect 8637 8867 8695 8873
rect 8637 8864 8649 8867
rect 8223 8836 8649 8864
rect 8223 8833 8235 8836
rect 8177 8827 8235 8833
rect 8637 8833 8649 8836
rect 8683 8833 8695 8867
rect 8637 8827 8695 8833
rect 9281 8867 9339 8873
rect 9281 8833 9293 8867
rect 9327 8864 9339 8867
rect 9741 8867 9799 8873
rect 9741 8864 9753 8867
rect 9327 8836 9753 8864
rect 9327 8833 9339 8836
rect 9281 8827 9339 8833
rect 9741 8833 9753 8836
rect 9787 8833 9799 8867
rect 9741 8827 9799 8833
rect 10385 8867 10443 8873
rect 10385 8833 10397 8867
rect 10431 8864 10443 8867
rect 10845 8867 10903 8873
rect 10845 8864 10857 8867
rect 10431 8836 10857 8864
rect 10431 8833 10443 8836
rect 10385 8827 10443 8833
rect 10845 8833 10857 8836
rect 10891 8833 10903 8867
rect 10845 8827 10903 8833
rect 11489 8867 11547 8873
rect 11489 8833 11501 8867
rect 11535 8864 11547 8867
rect 11949 8867 12007 8873
rect 11949 8864 11961 8867
rect 11535 8836 11961 8864
rect 11535 8833 11547 8836
rect 11489 8827 11547 8833
rect 11949 8833 11961 8836
rect 11995 8833 12007 8867
rect 11949 8827 12007 8833
rect 12593 8867 12651 8873
rect 12593 8833 12605 8867
rect 12639 8864 12651 8867
rect 13053 8867 13111 8873
rect 13053 8864 13065 8867
rect 12639 8836 13065 8864
rect 12639 8833 12651 8836
rect 12593 8827 12651 8833
rect 13053 8833 13065 8836
rect 13099 8833 13111 8867
rect 13053 8827 13111 8833
rect 13697 8867 13755 8873
rect 13697 8833 13709 8867
rect 13743 8864 13755 8867
rect 14157 8867 14215 8873
rect 14157 8864 14169 8867
rect 13743 8836 14169 8864
rect 13743 8833 13755 8836
rect 13697 8827 13755 8833
rect 14157 8833 14169 8836
rect 14203 8833 14215 8867
rect 14157 8827 14215 8833
rect 14801 8867 14859 8873
rect 14801 8833 14813 8867
rect 14847 8864 14859 8867
rect 15261 8867 15319 8873
rect 15261 8864 15273 8867
rect 14847 8836 15273 8864
rect 14847 8833 14859 8836
rect 14801 8827 14859 8833
rect 15261 8833 15273 8836
rect 15307 8833 15319 8867
rect 15261 8827 15319 8833
rect 15905 8867 15963 8873
rect 15905 8833 15917 8867
rect 15951 8864 15963 8867
rect 16365 8867 16423 8873
rect 16365 8864 16377 8867
rect 15951 8836 16377 8864
rect 15951 8833 15963 8836
rect 15905 8827 15963 8833
rect 16365 8833 16377 8836
rect 16411 8833 16423 8867
rect 16365 8827 16423 8833
rect 17009 8867 17067 8873
rect 17009 8833 17021 8867
rect 17055 8864 17067 8867
rect 17469 8867 17527 8873
rect 17469 8864 17481 8867
rect 17055 8836 17481 8864
rect 17055 8833 17067 8836
rect 17009 8827 17067 8833
rect 17469 8833 17481 8836
rect 17515 8833 17527 8867
rect 17469 8827 17527 8833
rect 18113 8867 18171 8873
rect 18113 8833 18125 8867
rect 18159 8864 18171 8867
rect 18573 8867 18631 8873
rect 18573 8864 18585 8867
rect 18159 8836 18585 8864
rect 18159 8833 18171 8836
rect 18113 8827 18171 8833
rect 18573 8833 18585 8836
rect 18619 8833 18631 8867
rect 18573 8827 18631 8833
rect 19217 8867 19275 8873
rect 19217 8833 19229 8867
rect 19263 8864 19275 8867
rect 19677 8867 19735 8873
rect 19677 8864 19689 8867
rect 19263 8836 19689 8864
rect 19263 8833 19275 8836
rect 19217 8827 19275 8833
rect 19677 8833 19689 8836
rect 19723 8833 19735 8867
rect 19677 8827 19735 8833
rect 3132 8728 3160 8827
rect 3758 8728 3764 8740
rect 3132 8700 3764 8728
rect 3758 8688 3764 8700
rect 3816 8688 3822 8740
rect 1904 8570 20764 8592
rect 1904 8518 7110 8570
rect 7162 8518 7174 8570
rect 7226 8518 7238 8570
rect 7290 8518 7302 8570
rect 7354 8518 12438 8570
rect 12490 8518 12502 8570
rect 12554 8518 12566 8570
rect 12618 8518 12630 8570
rect 12682 8518 17766 8570
rect 17818 8518 17830 8570
rect 17882 8518 17894 8570
rect 17946 8518 17958 8570
rect 18010 8518 20764 8570
rect 1904 8496 20764 8518
rect 3758 8456 3764 8468
rect 3719 8428 3764 8456
rect 3758 8416 3764 8428
rect 3816 8416 3822 8468
rect 4865 8323 4923 8329
rect 4865 8320 4877 8323
rect 3132 8292 4877 8320
rect 3132 8261 3160 8292
rect 4865 8289 4877 8292
rect 4911 8289 4923 8323
rect 7073 8323 7131 8329
rect 7073 8320 7085 8323
rect 4865 8283 4923 8289
rect 5340 8292 7085 8320
rect 5340 8261 5368 8292
rect 7073 8289 7085 8292
rect 7119 8289 7131 8323
rect 9281 8323 9339 8329
rect 9281 8320 9293 8323
rect 7073 8283 7131 8289
rect 7548 8292 9293 8320
rect 7548 8261 7576 8292
rect 9281 8289 9293 8292
rect 9327 8289 9339 8323
rect 10385 8323 10443 8329
rect 10385 8320 10397 8323
rect 9281 8283 9339 8289
rect 9572 8292 10397 8320
rect 3117 8255 3175 8261
rect 3117 8221 3129 8255
rect 3163 8221 3175 8255
rect 3117 8215 3175 8221
rect 4221 8255 4279 8261
rect 4221 8221 4233 8255
rect 4267 8221 4279 8255
rect 4221 8215 4279 8221
rect 5325 8255 5383 8261
rect 5325 8221 5337 8255
rect 5371 8221 5383 8255
rect 5325 8215 5383 8221
rect 6440 8255 6498 8261
rect 6440 8221 6452 8255
rect 6486 8221 6498 8255
rect 6440 8215 6498 8221
rect 7533 8255 7591 8261
rect 7533 8221 7545 8255
rect 7579 8221 7591 8255
rect 7533 8215 7591 8221
rect 8648 8255 8706 8261
rect 8648 8221 8660 8255
rect 8694 8221 8706 8255
rect 8648 8215 8706 8221
rect 4236 8184 4264 8215
rect 5969 8187 6027 8193
rect 5969 8184 5981 8187
rect 4236 8156 5981 8184
rect 5969 8153 5981 8156
rect 6015 8153 6027 8187
rect 6444 8184 6472 8215
rect 8177 8187 8235 8193
rect 8177 8184 8189 8187
rect 6444 8156 8189 8184
rect 5969 8147 6027 8153
rect 8177 8153 8189 8156
rect 8223 8153 8235 8187
rect 8652 8184 8680 8215
rect 9572 8184 9600 8292
rect 10385 8289 10397 8292
rect 10431 8289 10443 8323
rect 11489 8323 11547 8329
rect 11489 8320 11501 8323
rect 10385 8283 10443 8289
rect 10584 8292 11501 8320
rect 9741 8255 9799 8261
rect 9741 8221 9753 8255
rect 9787 8252 9799 8255
rect 10584 8252 10612 8292
rect 11489 8289 11501 8292
rect 11535 8289 11547 8323
rect 13697 8323 13755 8329
rect 13697 8320 13709 8323
rect 11489 8283 11547 8289
rect 11964 8292 13709 8320
rect 11964 8261 11992 8292
rect 13697 8289 13709 8292
rect 13743 8289 13755 8323
rect 15905 8323 15963 8329
rect 15905 8320 15917 8323
rect 13697 8283 13755 8289
rect 14172 8292 15917 8320
rect 14172 8261 14200 8292
rect 15905 8289 15917 8292
rect 15951 8289 15963 8323
rect 18113 8323 18171 8329
rect 18113 8320 18125 8323
rect 15905 8283 15963 8289
rect 16380 8292 18125 8320
rect 16380 8261 16408 8292
rect 18113 8289 18125 8292
rect 18159 8289 18171 8323
rect 20321 8323 20379 8329
rect 20321 8320 20333 8323
rect 18113 8283 18171 8289
rect 18588 8292 20333 8320
rect 18588 8261 18616 8292
rect 20321 8289 20333 8292
rect 20367 8289 20379 8323
rect 20321 8283 20379 8289
rect 9787 8224 10612 8252
rect 10845 8255 10903 8261
rect 9787 8221 9799 8224
rect 9741 8215 9799 8221
rect 10845 8221 10857 8255
rect 10891 8221 10903 8255
rect 10845 8215 10903 8221
rect 11949 8255 12007 8261
rect 11949 8221 11961 8255
rect 11995 8221 12007 8255
rect 11949 8215 12007 8221
rect 13053 8255 13111 8261
rect 13053 8221 13065 8255
rect 13099 8221 13111 8255
rect 13053 8215 13111 8221
rect 14168 8255 14226 8261
rect 14168 8221 14180 8255
rect 14214 8221 14226 8255
rect 14168 8215 14226 8221
rect 15261 8255 15319 8261
rect 15261 8221 15273 8255
rect 15307 8221 15319 8255
rect 15261 8215 15319 8221
rect 16365 8255 16423 8261
rect 16365 8221 16377 8255
rect 16411 8221 16423 8255
rect 16365 8215 16423 8221
rect 17469 8255 17527 8261
rect 17469 8221 17481 8255
rect 17515 8221 17527 8255
rect 17469 8215 17527 8221
rect 18573 8255 18631 8261
rect 18573 8221 18585 8255
rect 18619 8221 18631 8255
rect 18573 8215 18631 8221
rect 19677 8255 19735 8261
rect 19677 8221 19689 8255
rect 19723 8252 19735 8255
rect 20134 8252 20140 8264
rect 19723 8224 20140 8252
rect 19723 8221 19735 8224
rect 19677 8215 19735 8221
rect 8652 8156 9600 8184
rect 10860 8184 10888 8215
rect 12593 8187 12651 8193
rect 12593 8184 12605 8187
rect 10860 8156 12605 8184
rect 8177 8147 8235 8153
rect 12593 8153 12605 8156
rect 12639 8153 12651 8187
rect 13068 8184 13096 8215
rect 14801 8187 14859 8193
rect 14801 8184 14813 8187
rect 13068 8156 14813 8184
rect 12593 8147 12651 8153
rect 14801 8153 14813 8156
rect 14847 8153 14859 8187
rect 15276 8184 15304 8215
rect 17009 8187 17067 8193
rect 17009 8184 17021 8187
rect 15276 8156 17021 8184
rect 14801 8147 14859 8153
rect 17009 8153 17021 8156
rect 17055 8153 17067 8187
rect 17484 8184 17512 8215
rect 20134 8212 20140 8224
rect 20192 8212 20198 8264
rect 19217 8187 19275 8193
rect 19217 8184 19229 8187
rect 17484 8156 19229 8184
rect 17009 8147 17067 8153
rect 19217 8153 19229 8156
rect 19263 8153 19275 8187
rect 19217 8147 19275 8153
rect 1904 8026 20764 8048
rect 1904 7974 4446 8026
rect 4498 7974 4510 8026
rect 4562 7974 4574 8026
rect 4626 7974 4638 8026
rect 4690 7974 9774 8026
rect 9826 7974 9838 8026
rect 9890 7974 9902 8026
rect 9954 7974 9966 8026
rect 10018 7974 15102 8026
rect 15154 7974 15166 8026
rect 15218 7974 15230 8026
rect 15282 7974 15294 8026
rect 15346 7974 20764 8026
rect 1904 7952 20764 7974
rect 20134 7872 20140 7924
rect 20192 7912 20198 7924
rect 20321 7915 20379 7921
rect 20321 7912 20333 7915
rect 20192 7884 20333 7912
rect 20192 7872 20198 7884
rect 20321 7881 20333 7884
rect 20367 7881 20379 7915
rect 20321 7875 20379 7881
rect 3117 7779 3175 7785
rect 3117 7745 3129 7779
rect 3163 7745 3175 7779
rect 3117 7739 3175 7745
rect 3761 7779 3819 7785
rect 3761 7745 3773 7779
rect 3807 7776 3819 7779
rect 4221 7779 4279 7785
rect 4221 7776 4233 7779
rect 3807 7748 4233 7776
rect 3807 7745 3819 7748
rect 3761 7739 3819 7745
rect 4221 7745 4233 7748
rect 4267 7745 4279 7779
rect 4221 7739 4279 7745
rect 4865 7779 4923 7785
rect 4865 7745 4877 7779
rect 4911 7776 4923 7779
rect 5325 7779 5383 7785
rect 5325 7776 5337 7779
rect 4911 7748 5337 7776
rect 4911 7745 4923 7748
rect 4865 7739 4923 7745
rect 5325 7745 5337 7748
rect 5371 7745 5383 7779
rect 5325 7739 5383 7745
rect 5969 7779 6027 7785
rect 5969 7745 5981 7779
rect 6015 7776 6027 7779
rect 6429 7779 6487 7785
rect 6429 7776 6441 7779
rect 6015 7748 6441 7776
rect 6015 7745 6027 7748
rect 5969 7739 6027 7745
rect 6429 7745 6441 7748
rect 6475 7745 6487 7779
rect 6429 7739 6487 7745
rect 7073 7779 7131 7785
rect 7073 7745 7085 7779
rect 7119 7776 7131 7779
rect 7533 7779 7591 7785
rect 7533 7776 7545 7779
rect 7119 7748 7545 7776
rect 7119 7745 7131 7748
rect 7073 7739 7131 7745
rect 7533 7745 7545 7748
rect 7579 7745 7591 7779
rect 7533 7739 7591 7745
rect 8177 7779 8235 7785
rect 8177 7745 8189 7779
rect 8223 7776 8235 7779
rect 8637 7779 8695 7785
rect 8637 7776 8649 7779
rect 8223 7748 8649 7776
rect 8223 7745 8235 7748
rect 8177 7739 8235 7745
rect 8637 7745 8649 7748
rect 8683 7745 8695 7779
rect 8637 7739 8695 7745
rect 9281 7779 9339 7785
rect 9281 7745 9293 7779
rect 9327 7776 9339 7779
rect 9741 7779 9799 7785
rect 9741 7776 9753 7779
rect 9327 7748 9753 7776
rect 9327 7745 9339 7748
rect 9281 7739 9339 7745
rect 9741 7745 9753 7748
rect 9787 7745 9799 7779
rect 9741 7739 9799 7745
rect 10385 7779 10443 7785
rect 10385 7745 10397 7779
rect 10431 7776 10443 7779
rect 10845 7779 10903 7785
rect 10845 7776 10857 7779
rect 10431 7748 10857 7776
rect 10431 7745 10443 7748
rect 10385 7739 10443 7745
rect 10845 7745 10857 7748
rect 10891 7745 10903 7779
rect 10845 7739 10903 7745
rect 11489 7779 11547 7785
rect 11489 7745 11501 7779
rect 11535 7776 11547 7779
rect 11949 7779 12007 7785
rect 11949 7776 11961 7779
rect 11535 7748 11961 7776
rect 11535 7745 11547 7748
rect 11489 7739 11547 7745
rect 11949 7745 11961 7748
rect 11995 7745 12007 7779
rect 11949 7739 12007 7745
rect 12593 7779 12651 7785
rect 12593 7745 12605 7779
rect 12639 7776 12651 7779
rect 13053 7779 13111 7785
rect 13053 7776 13065 7779
rect 12639 7748 13065 7776
rect 12639 7745 12651 7748
rect 12593 7739 12651 7745
rect 13053 7745 13065 7748
rect 13099 7745 13111 7779
rect 13053 7739 13111 7745
rect 13697 7779 13755 7785
rect 13697 7745 13709 7779
rect 13743 7776 13755 7779
rect 14157 7779 14215 7785
rect 14157 7776 14169 7779
rect 13743 7748 14169 7776
rect 13743 7745 13755 7748
rect 13697 7739 13755 7745
rect 14157 7745 14169 7748
rect 14203 7745 14215 7779
rect 14157 7739 14215 7745
rect 14801 7779 14859 7785
rect 14801 7745 14813 7779
rect 14847 7776 14859 7779
rect 15261 7779 15319 7785
rect 15261 7776 15273 7779
rect 14847 7748 15273 7776
rect 14847 7745 14859 7748
rect 14801 7739 14859 7745
rect 15261 7745 15273 7748
rect 15307 7745 15319 7779
rect 15261 7739 15319 7745
rect 15905 7779 15963 7785
rect 15905 7745 15917 7779
rect 15951 7776 15963 7779
rect 16365 7779 16423 7785
rect 16365 7776 16377 7779
rect 15951 7748 16377 7776
rect 15951 7745 15963 7748
rect 15905 7739 15963 7745
rect 16365 7745 16377 7748
rect 16411 7745 16423 7779
rect 16365 7739 16423 7745
rect 17009 7779 17067 7785
rect 17009 7745 17021 7779
rect 17055 7776 17067 7779
rect 17469 7779 17527 7785
rect 17469 7776 17481 7779
rect 17055 7748 17481 7776
rect 17055 7745 17067 7748
rect 17009 7739 17067 7745
rect 17469 7745 17481 7748
rect 17515 7745 17527 7779
rect 17469 7739 17527 7745
rect 18113 7779 18171 7785
rect 18113 7745 18125 7779
rect 18159 7776 18171 7779
rect 18573 7779 18631 7785
rect 18573 7776 18585 7779
rect 18159 7748 18585 7776
rect 18159 7745 18171 7748
rect 18113 7739 18171 7745
rect 18573 7745 18585 7748
rect 18619 7745 18631 7779
rect 18573 7739 18631 7745
rect 19217 7779 19275 7785
rect 19217 7745 19229 7779
rect 19263 7776 19275 7779
rect 19677 7779 19735 7785
rect 19677 7776 19689 7779
rect 19263 7748 19689 7776
rect 19263 7745 19275 7748
rect 19217 7739 19275 7745
rect 19677 7745 19689 7748
rect 19723 7745 19735 7779
rect 19677 7739 19735 7745
rect 3132 7640 3160 7739
rect 3758 7640 3764 7652
rect 3132 7612 3764 7640
rect 3758 7600 3764 7612
rect 3816 7600 3822 7652
rect 1904 7482 20764 7504
rect 1904 7430 7110 7482
rect 7162 7430 7174 7482
rect 7226 7430 7238 7482
rect 7290 7430 7302 7482
rect 7354 7430 12438 7482
rect 12490 7430 12502 7482
rect 12554 7430 12566 7482
rect 12618 7430 12630 7482
rect 12682 7430 17766 7482
rect 17818 7430 17830 7482
rect 17882 7430 17894 7482
rect 17946 7430 17958 7482
rect 18010 7430 20764 7482
rect 1904 7408 20764 7430
rect 6352 7204 6564 7232
rect 3117 7167 3175 7173
rect 3117 7133 3129 7167
rect 3163 7133 3175 7167
rect 3758 7164 3764 7176
rect 3719 7136 3764 7164
rect 3117 7127 3175 7133
rect 3132 7096 3160 7127
rect 3758 7124 3764 7136
rect 3816 7124 3822 7176
rect 4221 7167 4279 7173
rect 4221 7133 4233 7167
rect 4267 7164 4279 7167
rect 5325 7167 5383 7173
rect 4267 7136 5092 7164
rect 4267 7133 4279 7136
rect 4221 7127 4279 7133
rect 4865 7099 4923 7105
rect 4865 7096 4877 7099
rect 3132 7068 4877 7096
rect 4865 7065 4877 7068
rect 4911 7065 4923 7099
rect 4865 7059 4923 7065
rect 5064 7028 5092 7136
rect 5325 7133 5337 7167
rect 5371 7164 5383 7167
rect 6352 7164 6380 7204
rect 5371 7136 6380 7164
rect 6440 7167 6498 7173
rect 5371 7133 5383 7136
rect 5325 7127 5383 7133
rect 6440 7133 6452 7167
rect 6486 7133 6498 7167
rect 6440 7127 6498 7133
rect 5969 7031 6027 7037
rect 5969 7028 5981 7031
rect 5064 7000 5981 7028
rect 5969 6997 5981 7000
rect 6015 6997 6027 7031
rect 6444 7028 6472 7127
rect 6536 7096 6564 7204
rect 8560 7204 8772 7232
rect 7533 7167 7591 7173
rect 7533 7133 7545 7167
rect 7579 7164 7591 7167
rect 8560 7164 8588 7204
rect 7579 7136 8588 7164
rect 8648 7167 8706 7173
rect 7579 7133 7591 7136
rect 7533 7127 7591 7133
rect 8648 7133 8660 7167
rect 8694 7133 8706 7167
rect 8744 7164 8772 7204
rect 9281 7167 9339 7173
rect 9281 7164 9293 7167
rect 8744 7136 9293 7164
rect 8648 7127 8706 7133
rect 9281 7133 9293 7136
rect 9327 7133 9339 7167
rect 9281 7127 9339 7133
rect 9741 7167 9799 7173
rect 9741 7133 9753 7167
rect 9787 7133 9799 7167
rect 9741 7127 9799 7133
rect 10845 7167 10903 7173
rect 10845 7133 10857 7167
rect 10891 7164 10903 7167
rect 11949 7167 12007 7173
rect 10891 7136 11716 7164
rect 10891 7133 10903 7136
rect 10845 7127 10903 7133
rect 7073 7099 7131 7105
rect 7073 7096 7085 7099
rect 6536 7068 7085 7096
rect 7073 7065 7085 7068
rect 7119 7065 7131 7099
rect 7073 7059 7131 7065
rect 8177 7031 8235 7037
rect 8177 7028 8189 7031
rect 6444 7000 8189 7028
rect 5969 6991 6027 6997
rect 8177 6997 8189 7000
rect 8223 6997 8235 7031
rect 8652 7028 8680 7127
rect 9756 7096 9784 7127
rect 11489 7099 11547 7105
rect 11489 7096 11501 7099
rect 9756 7068 11501 7096
rect 11489 7065 11501 7068
rect 11535 7065 11547 7099
rect 11489 7059 11547 7065
rect 10385 7031 10443 7037
rect 10385 7028 10397 7031
rect 8652 7000 10397 7028
rect 8177 6991 8235 6997
rect 10385 6997 10397 7000
rect 10431 6997 10443 7031
rect 11688 7028 11716 7136
rect 11949 7133 11961 7167
rect 11995 7133 12007 7167
rect 11949 7127 12007 7133
rect 13053 7167 13111 7173
rect 13053 7133 13065 7167
rect 13099 7164 13111 7167
rect 14168 7167 14226 7173
rect 13099 7136 13924 7164
rect 13099 7133 13111 7136
rect 13053 7127 13111 7133
rect 11964 7096 11992 7127
rect 13697 7099 13755 7105
rect 13697 7096 13709 7099
rect 11964 7068 13709 7096
rect 13697 7065 13709 7068
rect 13743 7065 13755 7099
rect 13697 7059 13755 7065
rect 12593 7031 12651 7037
rect 12593 7028 12605 7031
rect 11688 7000 12605 7028
rect 10385 6991 10443 6997
rect 12593 6997 12605 7000
rect 12639 6997 12651 7031
rect 13896 7028 13924 7136
rect 14168 7133 14180 7167
rect 14214 7133 14226 7167
rect 14168 7127 14226 7133
rect 15261 7167 15319 7173
rect 15261 7133 15273 7167
rect 15307 7164 15319 7167
rect 16365 7167 16423 7173
rect 15307 7136 16132 7164
rect 15307 7133 15319 7136
rect 15261 7127 15319 7133
rect 14172 7096 14200 7127
rect 15905 7099 15963 7105
rect 15905 7096 15917 7099
rect 14172 7068 15917 7096
rect 15905 7065 15917 7068
rect 15951 7065 15963 7099
rect 15905 7059 15963 7065
rect 14801 7031 14859 7037
rect 14801 7028 14813 7031
rect 13896 7000 14813 7028
rect 12593 6991 12651 6997
rect 14801 6997 14813 7000
rect 14847 6997 14859 7031
rect 16104 7028 16132 7136
rect 16365 7133 16377 7167
rect 16411 7133 16423 7167
rect 16365 7127 16423 7133
rect 17469 7167 17527 7173
rect 17469 7133 17481 7167
rect 17515 7164 17527 7167
rect 18573 7167 18631 7173
rect 17515 7136 18340 7164
rect 17515 7133 17527 7136
rect 17469 7127 17527 7133
rect 16380 7096 16408 7127
rect 18113 7099 18171 7105
rect 18113 7096 18125 7099
rect 16380 7068 18125 7096
rect 18113 7065 18125 7068
rect 18159 7065 18171 7099
rect 18113 7059 18171 7065
rect 17009 7031 17067 7037
rect 17009 7028 17021 7031
rect 16104 7000 17021 7028
rect 14801 6991 14859 6997
rect 17009 6997 17021 7000
rect 17055 6997 17067 7031
rect 18312 7028 18340 7136
rect 18573 7133 18585 7167
rect 18619 7133 18631 7167
rect 19674 7164 19680 7176
rect 19635 7136 19680 7164
rect 18573 7127 18631 7133
rect 18588 7096 18616 7127
rect 19674 7124 19680 7136
rect 19732 7124 19738 7176
rect 20321 7099 20379 7105
rect 20321 7096 20333 7099
rect 18588 7068 20333 7096
rect 20321 7065 20333 7068
rect 20367 7065 20379 7099
rect 20321 7059 20379 7065
rect 19217 7031 19275 7037
rect 19217 7028 19229 7031
rect 18312 7000 19229 7028
rect 17009 6991 17067 6997
rect 19217 6997 19229 7000
rect 19263 6997 19275 7031
rect 19217 6991 19275 6997
rect 1904 6938 20764 6960
rect 1904 6886 4446 6938
rect 4498 6886 4510 6938
rect 4562 6886 4574 6938
rect 4626 6886 4638 6938
rect 4690 6886 9774 6938
rect 9826 6886 9838 6938
rect 9890 6886 9902 6938
rect 9954 6886 9966 6938
rect 10018 6886 15102 6938
rect 15154 6886 15166 6938
rect 15218 6886 15230 6938
rect 15282 6886 15294 6938
rect 15346 6886 20764 6938
rect 1904 6864 20764 6886
rect 19674 6784 19680 6836
rect 19732 6824 19738 6836
rect 20321 6827 20379 6833
rect 20321 6824 20333 6827
rect 19732 6796 20333 6824
rect 19732 6784 19738 6796
rect 20321 6793 20333 6796
rect 20367 6793 20379 6827
rect 20321 6787 20379 6793
rect 3117 6691 3175 6697
rect 3117 6657 3129 6691
rect 3163 6657 3175 6691
rect 3117 6651 3175 6657
rect 3761 6691 3819 6697
rect 3761 6657 3773 6691
rect 3807 6688 3819 6691
rect 4221 6691 4279 6697
rect 4221 6688 4233 6691
rect 3807 6660 4233 6688
rect 3807 6657 3819 6660
rect 3761 6651 3819 6657
rect 4221 6657 4233 6660
rect 4267 6657 4279 6691
rect 4221 6651 4279 6657
rect 4865 6691 4923 6697
rect 4865 6657 4877 6691
rect 4911 6688 4923 6691
rect 5325 6691 5383 6697
rect 5325 6688 5337 6691
rect 4911 6660 5337 6688
rect 4911 6657 4923 6660
rect 4865 6651 4923 6657
rect 5325 6657 5337 6660
rect 5371 6657 5383 6691
rect 5325 6651 5383 6657
rect 5969 6691 6027 6697
rect 5969 6657 5981 6691
rect 6015 6688 6027 6691
rect 6429 6691 6487 6697
rect 6429 6688 6441 6691
rect 6015 6660 6441 6688
rect 6015 6657 6027 6660
rect 5969 6651 6027 6657
rect 6429 6657 6441 6660
rect 6475 6657 6487 6691
rect 6429 6651 6487 6657
rect 7073 6691 7131 6697
rect 7073 6657 7085 6691
rect 7119 6688 7131 6691
rect 7533 6691 7591 6697
rect 7533 6688 7545 6691
rect 7119 6660 7545 6688
rect 7119 6657 7131 6660
rect 7073 6651 7131 6657
rect 7533 6657 7545 6660
rect 7579 6657 7591 6691
rect 7533 6651 7591 6657
rect 8177 6691 8235 6697
rect 8177 6657 8189 6691
rect 8223 6688 8235 6691
rect 8637 6691 8695 6697
rect 8637 6688 8649 6691
rect 8223 6660 8649 6688
rect 8223 6657 8235 6660
rect 8177 6651 8235 6657
rect 8637 6657 8649 6660
rect 8683 6657 8695 6691
rect 8637 6651 8695 6657
rect 9281 6691 9339 6697
rect 9281 6657 9293 6691
rect 9327 6688 9339 6691
rect 9741 6691 9799 6697
rect 9741 6688 9753 6691
rect 9327 6660 9753 6688
rect 9327 6657 9339 6660
rect 9281 6651 9339 6657
rect 9741 6657 9753 6660
rect 9787 6657 9799 6691
rect 9741 6651 9799 6657
rect 10385 6691 10443 6697
rect 10385 6657 10397 6691
rect 10431 6688 10443 6691
rect 10845 6691 10903 6697
rect 10845 6688 10857 6691
rect 10431 6660 10857 6688
rect 10431 6657 10443 6660
rect 10385 6651 10443 6657
rect 10845 6657 10857 6660
rect 10891 6657 10903 6691
rect 10845 6651 10903 6657
rect 11489 6691 11547 6697
rect 11489 6657 11501 6691
rect 11535 6688 11547 6691
rect 11949 6691 12007 6697
rect 11949 6688 11961 6691
rect 11535 6660 11961 6688
rect 11535 6657 11547 6660
rect 11489 6651 11547 6657
rect 11949 6657 11961 6660
rect 11995 6657 12007 6691
rect 11949 6651 12007 6657
rect 12593 6691 12651 6697
rect 12593 6657 12605 6691
rect 12639 6688 12651 6691
rect 13053 6691 13111 6697
rect 13053 6688 13065 6691
rect 12639 6660 13065 6688
rect 12639 6657 12651 6660
rect 12593 6651 12651 6657
rect 13053 6657 13065 6660
rect 13099 6657 13111 6691
rect 13053 6651 13111 6657
rect 13697 6691 13755 6697
rect 13697 6657 13709 6691
rect 13743 6688 13755 6691
rect 14157 6691 14215 6697
rect 14157 6688 14169 6691
rect 13743 6660 14169 6688
rect 13743 6657 13755 6660
rect 13697 6651 13755 6657
rect 14157 6657 14169 6660
rect 14203 6657 14215 6691
rect 14157 6651 14215 6657
rect 14801 6691 14859 6697
rect 14801 6657 14813 6691
rect 14847 6688 14859 6691
rect 15261 6691 15319 6697
rect 15261 6688 15273 6691
rect 14847 6660 15273 6688
rect 14847 6657 14859 6660
rect 14801 6651 14859 6657
rect 15261 6657 15273 6660
rect 15307 6657 15319 6691
rect 15261 6651 15319 6657
rect 15905 6691 15963 6697
rect 15905 6657 15917 6691
rect 15951 6688 15963 6691
rect 16365 6691 16423 6697
rect 16365 6688 16377 6691
rect 15951 6660 16377 6688
rect 15951 6657 15963 6660
rect 15905 6651 15963 6657
rect 16365 6657 16377 6660
rect 16411 6657 16423 6691
rect 16365 6651 16423 6657
rect 17009 6691 17067 6697
rect 17009 6657 17021 6691
rect 17055 6688 17067 6691
rect 17469 6691 17527 6697
rect 17469 6688 17481 6691
rect 17055 6660 17481 6688
rect 17055 6657 17067 6660
rect 17009 6651 17067 6657
rect 17469 6657 17481 6660
rect 17515 6657 17527 6691
rect 17469 6651 17527 6657
rect 18113 6691 18171 6697
rect 18113 6657 18125 6691
rect 18159 6688 18171 6691
rect 18573 6691 18631 6697
rect 18573 6688 18585 6691
rect 18159 6660 18585 6688
rect 18159 6657 18171 6660
rect 18113 6651 18171 6657
rect 18573 6657 18585 6660
rect 18619 6657 18631 6691
rect 18573 6651 18631 6657
rect 19217 6691 19275 6697
rect 19217 6657 19229 6691
rect 19263 6688 19275 6691
rect 19677 6691 19735 6697
rect 19677 6688 19689 6691
rect 19263 6660 19689 6688
rect 19263 6657 19275 6660
rect 19217 6651 19275 6657
rect 19677 6657 19689 6660
rect 19723 6657 19735 6691
rect 19677 6651 19735 6657
rect 3132 6552 3160 6651
rect 3758 6552 3764 6564
rect 3132 6524 3764 6552
rect 3758 6512 3764 6524
rect 3816 6512 3822 6564
rect 1904 6394 20764 6416
rect 1904 6342 7110 6394
rect 7162 6342 7174 6394
rect 7226 6342 7238 6394
rect 7290 6342 7302 6394
rect 7354 6342 12438 6394
rect 12490 6342 12502 6394
rect 12554 6342 12566 6394
rect 12618 6342 12630 6394
rect 12682 6342 17766 6394
rect 17818 6342 17830 6394
rect 17882 6342 17894 6394
rect 17946 6342 17958 6394
rect 18010 6342 20764 6394
rect 1904 6320 20764 6342
rect 3758 6280 3764 6292
rect 3719 6252 3764 6280
rect 3758 6240 3764 6252
rect 3816 6240 3822 6292
rect 7073 6147 7131 6153
rect 7073 6144 7085 6147
rect 4236 6116 5276 6144
rect 4236 6085 4264 6116
rect 3117 6079 3175 6085
rect 3117 6045 3129 6079
rect 3163 6045 3175 6079
rect 3117 6039 3175 6045
rect 4232 6079 4290 6085
rect 4232 6045 4244 6079
rect 4278 6045 4290 6079
rect 4232 6039 4290 6045
rect 3132 6008 3160 6039
rect 4865 6011 4923 6017
rect 4865 6008 4877 6011
rect 3132 5980 4877 6008
rect 4865 5977 4877 5980
rect 4911 5977 4923 6011
rect 5248 6008 5276 6116
rect 5340 6116 7085 6144
rect 5340 6085 5368 6116
rect 7073 6113 7085 6116
rect 7119 6113 7131 6147
rect 9281 6147 9339 6153
rect 9281 6144 9293 6147
rect 7073 6107 7131 6113
rect 7548 6116 9293 6144
rect 7548 6085 7576 6116
rect 9281 6113 9293 6116
rect 9327 6113 9339 6147
rect 10385 6147 10443 6153
rect 10385 6144 10397 6147
rect 9281 6107 9339 6113
rect 9572 6116 10397 6144
rect 5325 6079 5383 6085
rect 5325 6045 5337 6079
rect 5371 6045 5383 6079
rect 5325 6039 5383 6045
rect 6429 6079 6487 6085
rect 6429 6045 6441 6079
rect 6475 6045 6487 6079
rect 6429 6039 6487 6045
rect 7533 6079 7591 6085
rect 7533 6045 7545 6079
rect 7579 6045 7591 6079
rect 7533 6039 7591 6045
rect 8648 6079 8706 6085
rect 8648 6045 8660 6079
rect 8694 6045 8706 6079
rect 8648 6039 8706 6045
rect 5969 6011 6027 6017
rect 5969 6008 5981 6011
rect 5248 5980 5981 6008
rect 4865 5971 4923 5977
rect 5969 5977 5981 5980
rect 6015 5977 6027 6011
rect 6444 6008 6472 6039
rect 8177 6011 8235 6017
rect 8177 6008 8189 6011
rect 6444 5980 8189 6008
rect 5969 5971 6027 5977
rect 8177 5977 8189 5980
rect 8223 5977 8235 6011
rect 8652 6008 8680 6039
rect 9572 6008 9600 6116
rect 10385 6113 10397 6116
rect 10431 6113 10443 6147
rect 11489 6147 11547 6153
rect 11489 6144 11501 6147
rect 10385 6107 10443 6113
rect 10584 6116 11501 6144
rect 9741 6079 9799 6085
rect 9741 6045 9753 6079
rect 9787 6076 9799 6079
rect 10584 6076 10612 6116
rect 11489 6113 11501 6116
rect 11535 6113 11547 6147
rect 13697 6147 13755 6153
rect 13697 6144 13709 6147
rect 11489 6107 11547 6113
rect 11964 6116 13709 6144
rect 11964 6085 11992 6116
rect 13697 6113 13709 6116
rect 13743 6113 13755 6147
rect 15905 6147 15963 6153
rect 15905 6144 15917 6147
rect 13697 6107 13755 6113
rect 14172 6116 15917 6144
rect 14172 6085 14200 6116
rect 15905 6113 15917 6116
rect 15951 6113 15963 6147
rect 18113 6147 18171 6153
rect 18113 6144 18125 6147
rect 15905 6107 15963 6113
rect 16380 6116 18125 6144
rect 16380 6085 16408 6116
rect 18113 6113 18125 6116
rect 18159 6113 18171 6147
rect 20321 6147 20379 6153
rect 20321 6144 20333 6147
rect 18113 6107 18171 6113
rect 18588 6116 20333 6144
rect 18588 6085 18616 6116
rect 20321 6113 20333 6116
rect 20367 6113 20379 6147
rect 20321 6107 20379 6113
rect 9787 6048 10612 6076
rect 10845 6079 10903 6085
rect 9787 6045 9799 6048
rect 9741 6039 9799 6045
rect 10845 6045 10857 6079
rect 10891 6045 10903 6079
rect 10845 6039 10903 6045
rect 11949 6079 12007 6085
rect 11949 6045 11961 6079
rect 11995 6045 12007 6079
rect 11949 6039 12007 6045
rect 13053 6079 13111 6085
rect 13053 6045 13065 6079
rect 13099 6045 13111 6079
rect 13053 6039 13111 6045
rect 14168 6079 14226 6085
rect 14168 6045 14180 6079
rect 14214 6045 14226 6079
rect 14168 6039 14226 6045
rect 15261 6079 15319 6085
rect 15261 6045 15273 6079
rect 15307 6045 15319 6079
rect 15261 6039 15319 6045
rect 16365 6079 16423 6085
rect 16365 6045 16377 6079
rect 16411 6045 16423 6079
rect 16365 6039 16423 6045
rect 17469 6079 17527 6085
rect 17469 6045 17481 6079
rect 17515 6045 17527 6079
rect 17469 6039 17527 6045
rect 18573 6079 18631 6085
rect 18573 6045 18585 6079
rect 18619 6045 18631 6079
rect 18573 6039 18631 6045
rect 19677 6079 19735 6085
rect 19677 6045 19689 6079
rect 19723 6076 19735 6079
rect 20134 6076 20140 6088
rect 19723 6048 20140 6076
rect 19723 6045 19735 6048
rect 19677 6039 19735 6045
rect 8652 5980 9600 6008
rect 10860 6008 10888 6039
rect 12593 6011 12651 6017
rect 12593 6008 12605 6011
rect 10860 5980 12605 6008
rect 8177 5971 8235 5977
rect 12593 5977 12605 5980
rect 12639 5977 12651 6011
rect 13068 6008 13096 6039
rect 14801 6011 14859 6017
rect 14801 6008 14813 6011
rect 13068 5980 14813 6008
rect 12593 5971 12651 5977
rect 14801 5977 14813 5980
rect 14847 5977 14859 6011
rect 15276 6008 15304 6039
rect 17009 6011 17067 6017
rect 17009 6008 17021 6011
rect 15276 5980 17021 6008
rect 14801 5971 14859 5977
rect 17009 5977 17021 5980
rect 17055 5977 17067 6011
rect 17484 6008 17512 6039
rect 20134 6036 20140 6048
rect 20192 6036 20198 6088
rect 19217 6011 19275 6017
rect 19217 6008 19229 6011
rect 17484 5980 19229 6008
rect 17009 5971 17067 5977
rect 19217 5977 19229 5980
rect 19263 5977 19275 6011
rect 19217 5971 19275 5977
rect 1904 5850 20764 5872
rect 1904 5798 4446 5850
rect 4498 5798 4510 5850
rect 4562 5798 4574 5850
rect 4626 5798 4638 5850
rect 4690 5798 9774 5850
rect 9826 5798 9838 5850
rect 9890 5798 9902 5850
rect 9954 5798 9966 5850
rect 10018 5798 15102 5850
rect 15154 5798 15166 5850
rect 15218 5798 15230 5850
rect 15282 5798 15294 5850
rect 15346 5798 20764 5850
rect 1904 5776 20764 5798
rect 20134 5696 20140 5748
rect 20192 5736 20198 5748
rect 20321 5739 20379 5745
rect 20321 5736 20333 5739
rect 20192 5708 20333 5736
rect 20192 5696 20198 5708
rect 20321 5705 20333 5708
rect 20367 5705 20379 5739
rect 20321 5699 20379 5705
rect 3117 5603 3175 5609
rect 3117 5569 3129 5603
rect 3163 5569 3175 5603
rect 3117 5563 3175 5569
rect 3761 5603 3819 5609
rect 3761 5569 3773 5603
rect 3807 5600 3819 5603
rect 4221 5603 4279 5609
rect 4221 5600 4233 5603
rect 3807 5572 4233 5600
rect 3807 5569 3819 5572
rect 3761 5563 3819 5569
rect 4221 5569 4233 5572
rect 4267 5569 4279 5603
rect 4221 5563 4279 5569
rect 4865 5603 4923 5609
rect 4865 5569 4877 5603
rect 4911 5600 4923 5603
rect 5325 5603 5383 5609
rect 5325 5600 5337 5603
rect 4911 5572 5337 5600
rect 4911 5569 4923 5572
rect 4865 5563 4923 5569
rect 5325 5569 5337 5572
rect 5371 5569 5383 5603
rect 5325 5563 5383 5569
rect 5969 5603 6027 5609
rect 5969 5569 5981 5603
rect 6015 5600 6027 5603
rect 6429 5603 6487 5609
rect 6429 5600 6441 5603
rect 6015 5572 6441 5600
rect 6015 5569 6027 5572
rect 5969 5563 6027 5569
rect 6429 5569 6441 5572
rect 6475 5569 6487 5603
rect 6429 5563 6487 5569
rect 7073 5603 7131 5609
rect 7073 5569 7085 5603
rect 7119 5600 7131 5603
rect 7533 5603 7591 5609
rect 7533 5600 7545 5603
rect 7119 5572 7545 5600
rect 7119 5569 7131 5572
rect 7073 5563 7131 5569
rect 7533 5569 7545 5572
rect 7579 5569 7591 5603
rect 7533 5563 7591 5569
rect 8177 5603 8235 5609
rect 8177 5569 8189 5603
rect 8223 5600 8235 5603
rect 8637 5603 8695 5609
rect 8637 5600 8649 5603
rect 8223 5572 8649 5600
rect 8223 5569 8235 5572
rect 8177 5563 8235 5569
rect 8637 5569 8649 5572
rect 8683 5569 8695 5603
rect 8637 5563 8695 5569
rect 9281 5603 9339 5609
rect 9281 5569 9293 5603
rect 9327 5600 9339 5603
rect 9741 5603 9799 5609
rect 9741 5600 9753 5603
rect 9327 5572 9753 5600
rect 9327 5569 9339 5572
rect 9281 5563 9339 5569
rect 9741 5569 9753 5572
rect 9787 5569 9799 5603
rect 9741 5563 9799 5569
rect 10385 5603 10443 5609
rect 10385 5569 10397 5603
rect 10431 5600 10443 5603
rect 10845 5603 10903 5609
rect 10845 5600 10857 5603
rect 10431 5572 10857 5600
rect 10431 5569 10443 5572
rect 10385 5563 10443 5569
rect 10845 5569 10857 5572
rect 10891 5569 10903 5603
rect 10845 5563 10903 5569
rect 11489 5603 11547 5609
rect 11489 5569 11501 5603
rect 11535 5600 11547 5603
rect 11949 5603 12007 5609
rect 11949 5600 11961 5603
rect 11535 5572 11961 5600
rect 11535 5569 11547 5572
rect 11489 5563 11547 5569
rect 11949 5569 11961 5572
rect 11995 5569 12007 5603
rect 11949 5563 12007 5569
rect 12593 5603 12651 5609
rect 12593 5569 12605 5603
rect 12639 5600 12651 5603
rect 13053 5603 13111 5609
rect 13053 5600 13065 5603
rect 12639 5572 13065 5600
rect 12639 5569 12651 5572
rect 12593 5563 12651 5569
rect 13053 5569 13065 5572
rect 13099 5569 13111 5603
rect 13053 5563 13111 5569
rect 13697 5603 13755 5609
rect 13697 5569 13709 5603
rect 13743 5600 13755 5603
rect 14157 5603 14215 5609
rect 14157 5600 14169 5603
rect 13743 5572 14169 5600
rect 13743 5569 13755 5572
rect 13697 5563 13755 5569
rect 14157 5569 14169 5572
rect 14203 5569 14215 5603
rect 14157 5563 14215 5569
rect 14801 5603 14859 5609
rect 14801 5569 14813 5603
rect 14847 5600 14859 5603
rect 15261 5603 15319 5609
rect 15261 5600 15273 5603
rect 14847 5572 15273 5600
rect 14847 5569 14859 5572
rect 14801 5563 14859 5569
rect 15261 5569 15273 5572
rect 15307 5569 15319 5603
rect 15261 5563 15319 5569
rect 15905 5603 15963 5609
rect 15905 5569 15917 5603
rect 15951 5600 15963 5603
rect 16365 5603 16423 5609
rect 16365 5600 16377 5603
rect 15951 5572 16377 5600
rect 15951 5569 15963 5572
rect 15905 5563 15963 5569
rect 16365 5569 16377 5572
rect 16411 5569 16423 5603
rect 16365 5563 16423 5569
rect 17009 5603 17067 5609
rect 17009 5569 17021 5603
rect 17055 5600 17067 5603
rect 17469 5603 17527 5609
rect 17469 5600 17481 5603
rect 17055 5572 17481 5600
rect 17055 5569 17067 5572
rect 17009 5563 17067 5569
rect 17469 5569 17481 5572
rect 17515 5569 17527 5603
rect 17469 5563 17527 5569
rect 18113 5603 18171 5609
rect 18113 5569 18125 5603
rect 18159 5600 18171 5603
rect 18573 5603 18631 5609
rect 18573 5600 18585 5603
rect 18159 5572 18585 5600
rect 18159 5569 18171 5572
rect 18113 5563 18171 5569
rect 18573 5569 18585 5572
rect 18619 5569 18631 5603
rect 18573 5563 18631 5569
rect 19217 5603 19275 5609
rect 19217 5569 19229 5603
rect 19263 5600 19275 5603
rect 19677 5603 19735 5609
rect 19677 5600 19689 5603
rect 19263 5572 19689 5600
rect 19263 5569 19275 5572
rect 19217 5563 19275 5569
rect 19677 5569 19689 5572
rect 19723 5569 19735 5603
rect 19677 5563 19735 5569
rect 3132 5464 3160 5563
rect 3758 5464 3764 5476
rect 3132 5436 3764 5464
rect 3758 5424 3764 5436
rect 3816 5424 3822 5476
rect 1904 5306 20764 5328
rect 1904 5254 7110 5306
rect 7162 5254 7174 5306
rect 7226 5254 7238 5306
rect 7290 5254 7302 5306
rect 7354 5254 12438 5306
rect 12490 5254 12502 5306
rect 12554 5254 12566 5306
rect 12618 5254 12630 5306
rect 12682 5254 17766 5306
rect 17818 5254 17830 5306
rect 17882 5254 17894 5306
rect 17946 5254 17958 5306
rect 18010 5254 20764 5306
rect 1904 5232 20764 5254
rect 3117 4991 3175 4997
rect 3117 4957 3129 4991
rect 3163 4957 3175 4991
rect 3758 4988 3764 5000
rect 3719 4960 3764 4988
rect 3117 4951 3175 4957
rect 3132 4852 3160 4951
rect 3758 4948 3764 4960
rect 3816 4948 3822 5000
rect 4221 4991 4279 4997
rect 4221 4957 4233 4991
rect 4267 4988 4279 4991
rect 5325 4991 5383 4997
rect 4267 4960 5276 4988
rect 4267 4957 4279 4960
rect 4221 4951 4279 4957
rect 4865 4855 4923 4861
rect 4865 4852 4877 4855
rect 3132 4824 4877 4852
rect 4865 4821 4877 4824
rect 4911 4821 4923 4855
rect 5248 4852 5276 4960
rect 5325 4957 5337 4991
rect 5371 4957 5383 4991
rect 5325 4951 5383 4957
rect 6429 4991 6487 4997
rect 6429 4957 6441 4991
rect 6475 4988 6487 4991
rect 7533 4991 7591 4997
rect 6475 4960 7300 4988
rect 6475 4957 6487 4960
rect 6429 4951 6487 4957
rect 5340 4920 5368 4951
rect 7073 4923 7131 4929
rect 7073 4920 7085 4923
rect 5340 4892 7085 4920
rect 7073 4889 7085 4892
rect 7119 4889 7131 4923
rect 7073 4883 7131 4889
rect 5969 4855 6027 4861
rect 5969 4852 5981 4855
rect 5248 4824 5981 4852
rect 4865 4815 4923 4821
rect 5969 4821 5981 4824
rect 6015 4821 6027 4855
rect 7272 4852 7300 4960
rect 7533 4957 7545 4991
rect 7579 4957 7591 4991
rect 7533 4951 7591 4957
rect 8637 4991 8695 4997
rect 8637 4957 8649 4991
rect 8683 4988 8695 4991
rect 9741 4991 9799 4997
rect 8683 4960 9692 4988
rect 8683 4957 8695 4960
rect 8637 4951 8695 4957
rect 7548 4920 7576 4951
rect 9281 4923 9339 4929
rect 9281 4920 9293 4923
rect 7548 4892 9293 4920
rect 9281 4889 9293 4892
rect 9327 4889 9339 4923
rect 9281 4883 9339 4889
rect 8177 4855 8235 4861
rect 8177 4852 8189 4855
rect 7272 4824 8189 4852
rect 5969 4815 6027 4821
rect 8177 4821 8189 4824
rect 8223 4821 8235 4855
rect 9664 4852 9692 4960
rect 9741 4957 9753 4991
rect 9787 4988 9799 4991
rect 10845 4991 10903 4997
rect 9787 4960 10612 4988
rect 9787 4957 9799 4960
rect 9741 4951 9799 4957
rect 10584 4920 10612 4960
rect 10845 4957 10857 4991
rect 10891 4988 10903 4991
rect 11949 4991 12007 4997
rect 10891 4960 11716 4988
rect 10891 4957 10903 4960
rect 10845 4951 10903 4957
rect 11489 4923 11547 4929
rect 11489 4920 11501 4923
rect 10584 4892 11501 4920
rect 11489 4889 11501 4892
rect 11535 4889 11547 4923
rect 11489 4883 11547 4889
rect 10385 4855 10443 4861
rect 10385 4852 10397 4855
rect 9664 4824 10397 4852
rect 8177 4815 8235 4821
rect 10385 4821 10397 4824
rect 10431 4821 10443 4855
rect 11688 4852 11716 4960
rect 11949 4957 11961 4991
rect 11995 4957 12007 4991
rect 11949 4951 12007 4957
rect 13053 4991 13111 4997
rect 13053 4957 13065 4991
rect 13099 4988 13111 4991
rect 14168 4991 14226 4997
rect 13099 4960 13924 4988
rect 13099 4957 13111 4960
rect 13053 4951 13111 4957
rect 11964 4920 11992 4951
rect 13697 4923 13755 4929
rect 13697 4920 13709 4923
rect 11964 4892 13709 4920
rect 13697 4889 13709 4892
rect 13743 4889 13755 4923
rect 13697 4883 13755 4889
rect 12593 4855 12651 4861
rect 12593 4852 12605 4855
rect 11688 4824 12605 4852
rect 10385 4815 10443 4821
rect 12593 4821 12605 4824
rect 12639 4821 12651 4855
rect 13896 4852 13924 4960
rect 14168 4957 14180 4991
rect 14214 4957 14226 4991
rect 14168 4951 14226 4957
rect 15261 4991 15319 4997
rect 15261 4957 15273 4991
rect 15307 4988 15319 4991
rect 16365 4991 16423 4997
rect 15307 4960 16132 4988
rect 15307 4957 15319 4960
rect 15261 4951 15319 4957
rect 14172 4920 14200 4951
rect 15905 4923 15963 4929
rect 15905 4920 15917 4923
rect 14172 4892 15917 4920
rect 15905 4889 15917 4892
rect 15951 4889 15963 4923
rect 15905 4883 15963 4889
rect 14801 4855 14859 4861
rect 14801 4852 14813 4855
rect 13896 4824 14813 4852
rect 12593 4815 12651 4821
rect 14801 4821 14813 4824
rect 14847 4821 14859 4855
rect 16104 4852 16132 4960
rect 16365 4957 16377 4991
rect 16411 4957 16423 4991
rect 16365 4951 16423 4957
rect 17469 4991 17527 4997
rect 17469 4957 17481 4991
rect 17515 4988 17527 4991
rect 18573 4991 18631 4997
rect 17515 4960 18340 4988
rect 17515 4957 17527 4960
rect 17469 4951 17527 4957
rect 16380 4920 16408 4951
rect 18113 4923 18171 4929
rect 18113 4920 18125 4923
rect 16380 4892 18125 4920
rect 18113 4889 18125 4892
rect 18159 4889 18171 4923
rect 18113 4883 18171 4889
rect 17009 4855 17067 4861
rect 17009 4852 17021 4855
rect 16104 4824 17021 4852
rect 14801 4815 14859 4821
rect 17009 4821 17021 4824
rect 17055 4821 17067 4855
rect 18312 4852 18340 4960
rect 18573 4957 18585 4991
rect 18619 4957 18631 4991
rect 19674 4988 19680 5000
rect 19635 4960 19680 4988
rect 18573 4951 18631 4957
rect 18588 4920 18616 4951
rect 19674 4948 19680 4960
rect 19732 4948 19738 5000
rect 20321 4923 20379 4929
rect 20321 4920 20333 4923
rect 18588 4892 20333 4920
rect 20321 4889 20333 4892
rect 20367 4889 20379 4923
rect 20321 4883 20379 4889
rect 19217 4855 19275 4861
rect 19217 4852 19229 4855
rect 18312 4824 19229 4852
rect 17009 4815 17067 4821
rect 19217 4821 19229 4824
rect 19263 4821 19275 4855
rect 19217 4815 19275 4821
rect 1904 4762 20764 4784
rect 1904 4710 4446 4762
rect 4498 4710 4510 4762
rect 4562 4710 4574 4762
rect 4626 4710 4638 4762
rect 4690 4710 9774 4762
rect 9826 4710 9838 4762
rect 9890 4710 9902 4762
rect 9954 4710 9966 4762
rect 10018 4710 15102 4762
rect 15154 4710 15166 4762
rect 15218 4710 15230 4762
rect 15282 4710 15294 4762
rect 15346 4710 20764 4762
rect 1904 4688 20764 4710
rect 19674 4608 19680 4660
rect 19732 4648 19738 4660
rect 20321 4651 20379 4657
rect 20321 4648 20333 4651
rect 19732 4620 20333 4648
rect 19732 4608 19738 4620
rect 20321 4617 20333 4620
rect 20367 4617 20379 4651
rect 20321 4611 20379 4617
rect 3117 4515 3175 4521
rect 3117 4481 3129 4515
rect 3163 4481 3175 4515
rect 3117 4475 3175 4481
rect 3761 4515 3819 4521
rect 3761 4481 3773 4515
rect 3807 4512 3819 4515
rect 4221 4515 4279 4521
rect 4221 4512 4233 4515
rect 3807 4484 4233 4512
rect 3807 4481 3819 4484
rect 3761 4475 3819 4481
rect 4221 4481 4233 4484
rect 4267 4481 4279 4515
rect 4221 4475 4279 4481
rect 4865 4515 4923 4521
rect 4865 4481 4877 4515
rect 4911 4512 4923 4515
rect 5325 4515 5383 4521
rect 5325 4512 5337 4515
rect 4911 4484 5337 4512
rect 4911 4481 4923 4484
rect 4865 4475 4923 4481
rect 5325 4481 5337 4484
rect 5371 4481 5383 4515
rect 5325 4475 5383 4481
rect 5969 4515 6027 4521
rect 5969 4481 5981 4515
rect 6015 4512 6027 4515
rect 6429 4515 6487 4521
rect 6429 4512 6441 4515
rect 6015 4484 6441 4512
rect 6015 4481 6027 4484
rect 5969 4475 6027 4481
rect 6429 4481 6441 4484
rect 6475 4481 6487 4515
rect 6429 4475 6487 4481
rect 7073 4515 7131 4521
rect 7073 4481 7085 4515
rect 7119 4512 7131 4515
rect 7533 4515 7591 4521
rect 7533 4512 7545 4515
rect 7119 4484 7545 4512
rect 7119 4481 7131 4484
rect 7073 4475 7131 4481
rect 7533 4481 7545 4484
rect 7579 4481 7591 4515
rect 7533 4475 7591 4481
rect 8177 4515 8235 4521
rect 8177 4481 8189 4515
rect 8223 4512 8235 4515
rect 8637 4515 8695 4521
rect 8637 4512 8649 4515
rect 8223 4484 8649 4512
rect 8223 4481 8235 4484
rect 8177 4475 8235 4481
rect 8637 4481 8649 4484
rect 8683 4481 8695 4515
rect 8637 4475 8695 4481
rect 9281 4515 9339 4521
rect 9281 4481 9293 4515
rect 9327 4512 9339 4515
rect 9741 4515 9799 4521
rect 9741 4512 9753 4515
rect 9327 4484 9753 4512
rect 9327 4481 9339 4484
rect 9281 4475 9339 4481
rect 9741 4481 9753 4484
rect 9787 4481 9799 4515
rect 9741 4475 9799 4481
rect 10385 4515 10443 4521
rect 10385 4481 10397 4515
rect 10431 4512 10443 4515
rect 10845 4515 10903 4521
rect 10845 4512 10857 4515
rect 10431 4484 10857 4512
rect 10431 4481 10443 4484
rect 10385 4475 10443 4481
rect 10845 4481 10857 4484
rect 10891 4481 10903 4515
rect 10845 4475 10903 4481
rect 11489 4515 11547 4521
rect 11489 4481 11501 4515
rect 11535 4512 11547 4515
rect 11949 4515 12007 4521
rect 11949 4512 11961 4515
rect 11535 4484 11961 4512
rect 11535 4481 11547 4484
rect 11489 4475 11547 4481
rect 11949 4481 11961 4484
rect 11995 4481 12007 4515
rect 11949 4475 12007 4481
rect 12593 4515 12651 4521
rect 12593 4481 12605 4515
rect 12639 4512 12651 4515
rect 13053 4515 13111 4521
rect 13053 4512 13065 4515
rect 12639 4484 13065 4512
rect 12639 4481 12651 4484
rect 12593 4475 12651 4481
rect 13053 4481 13065 4484
rect 13099 4481 13111 4515
rect 13053 4475 13111 4481
rect 13697 4515 13755 4521
rect 13697 4481 13709 4515
rect 13743 4512 13755 4515
rect 14157 4515 14215 4521
rect 14157 4512 14169 4515
rect 13743 4484 14169 4512
rect 13743 4481 13755 4484
rect 13697 4475 13755 4481
rect 14157 4481 14169 4484
rect 14203 4481 14215 4515
rect 14157 4475 14215 4481
rect 14801 4515 14859 4521
rect 14801 4481 14813 4515
rect 14847 4512 14859 4515
rect 15261 4515 15319 4521
rect 15261 4512 15273 4515
rect 14847 4484 15273 4512
rect 14847 4481 14859 4484
rect 14801 4475 14859 4481
rect 15261 4481 15273 4484
rect 15307 4481 15319 4515
rect 15261 4475 15319 4481
rect 15905 4515 15963 4521
rect 15905 4481 15917 4515
rect 15951 4512 15963 4515
rect 16365 4515 16423 4521
rect 16365 4512 16377 4515
rect 15951 4484 16377 4512
rect 15951 4481 15963 4484
rect 15905 4475 15963 4481
rect 16365 4481 16377 4484
rect 16411 4481 16423 4515
rect 16365 4475 16423 4481
rect 17009 4515 17067 4521
rect 17009 4481 17021 4515
rect 17055 4512 17067 4515
rect 17469 4515 17527 4521
rect 17469 4512 17481 4515
rect 17055 4484 17481 4512
rect 17055 4481 17067 4484
rect 17009 4475 17067 4481
rect 17469 4481 17481 4484
rect 17515 4481 17527 4515
rect 17469 4475 17527 4481
rect 18113 4515 18171 4521
rect 18113 4481 18125 4515
rect 18159 4512 18171 4515
rect 18573 4515 18631 4521
rect 18573 4512 18585 4515
rect 18159 4484 18585 4512
rect 18159 4481 18171 4484
rect 18113 4475 18171 4481
rect 18573 4481 18585 4484
rect 18619 4481 18631 4515
rect 18573 4475 18631 4481
rect 19217 4515 19275 4521
rect 19217 4481 19229 4515
rect 19263 4512 19275 4515
rect 19677 4515 19735 4521
rect 19677 4512 19689 4515
rect 19263 4484 19689 4512
rect 19263 4481 19275 4484
rect 19217 4475 19275 4481
rect 19677 4481 19689 4484
rect 19723 4481 19735 4515
rect 19677 4475 19735 4481
rect 3132 4376 3160 4475
rect 3758 4376 3764 4388
rect 3132 4348 3764 4376
rect 3758 4336 3764 4348
rect 3816 4336 3822 4388
rect 1904 4218 20764 4240
rect 1904 4166 7110 4218
rect 7162 4166 7174 4218
rect 7226 4166 7238 4218
rect 7290 4166 7302 4218
rect 7354 4166 12438 4218
rect 12490 4166 12502 4218
rect 12554 4166 12566 4218
rect 12618 4166 12630 4218
rect 12682 4166 17766 4218
rect 17818 4166 17830 4218
rect 17882 4166 17894 4218
rect 17946 4166 17958 4218
rect 18010 4166 20764 4218
rect 1904 4144 20764 4166
rect 3758 4104 3764 4116
rect 3719 4076 3764 4104
rect 3758 4064 3764 4076
rect 3816 4064 3822 4116
rect 7073 3971 7131 3977
rect 7073 3968 7085 3971
rect 4236 3940 5276 3968
rect 4236 3909 4264 3940
rect 3117 3903 3175 3909
rect 3117 3869 3129 3903
rect 3163 3869 3175 3903
rect 3117 3863 3175 3869
rect 4232 3903 4290 3909
rect 4232 3869 4244 3903
rect 4278 3869 4290 3903
rect 4232 3863 4290 3869
rect 3132 3832 3160 3863
rect 4865 3835 4923 3841
rect 4865 3832 4877 3835
rect 3132 3804 4877 3832
rect 4865 3801 4877 3804
rect 4911 3801 4923 3835
rect 5248 3832 5276 3940
rect 5340 3940 7085 3968
rect 5340 3909 5368 3940
rect 7073 3937 7085 3940
rect 7119 3937 7131 3971
rect 9281 3971 9339 3977
rect 9281 3968 9293 3971
rect 7073 3931 7131 3937
rect 7548 3940 9293 3968
rect 7548 3909 7576 3940
rect 9281 3937 9293 3940
rect 9327 3937 9339 3971
rect 10385 3971 10443 3977
rect 10385 3968 10397 3971
rect 9281 3931 9339 3937
rect 9572 3940 10397 3968
rect 5325 3903 5383 3909
rect 5325 3869 5337 3903
rect 5371 3869 5383 3903
rect 5325 3863 5383 3869
rect 6429 3903 6487 3909
rect 6429 3869 6441 3903
rect 6475 3869 6487 3903
rect 6429 3863 6487 3869
rect 7533 3903 7591 3909
rect 7533 3869 7545 3903
rect 7579 3869 7591 3903
rect 7533 3863 7591 3869
rect 8648 3903 8706 3909
rect 8648 3869 8660 3903
rect 8694 3869 8706 3903
rect 8648 3863 8706 3869
rect 5969 3835 6027 3841
rect 5969 3832 5981 3835
rect 5248 3804 5981 3832
rect 4865 3795 4923 3801
rect 5969 3801 5981 3804
rect 6015 3801 6027 3835
rect 6444 3832 6472 3863
rect 8177 3835 8235 3841
rect 8177 3832 8189 3835
rect 6444 3804 8189 3832
rect 5969 3795 6027 3801
rect 8177 3801 8189 3804
rect 8223 3801 8235 3835
rect 8652 3832 8680 3863
rect 9572 3832 9600 3940
rect 10385 3937 10397 3940
rect 10431 3937 10443 3971
rect 11489 3971 11547 3977
rect 11489 3968 11501 3971
rect 10385 3931 10443 3937
rect 10584 3940 11501 3968
rect 9741 3903 9799 3909
rect 9741 3869 9753 3903
rect 9787 3900 9799 3903
rect 10584 3900 10612 3940
rect 11489 3937 11501 3940
rect 11535 3937 11547 3971
rect 13697 3971 13755 3977
rect 13697 3968 13709 3971
rect 11489 3931 11547 3937
rect 11964 3940 13709 3968
rect 11964 3909 11992 3940
rect 13697 3937 13709 3940
rect 13743 3937 13755 3971
rect 15905 3971 15963 3977
rect 15905 3968 15917 3971
rect 13697 3931 13755 3937
rect 14172 3940 15917 3968
rect 14172 3909 14200 3940
rect 15905 3937 15917 3940
rect 15951 3937 15963 3971
rect 18113 3971 18171 3977
rect 18113 3968 18125 3971
rect 15905 3931 15963 3937
rect 16380 3940 18125 3968
rect 16380 3909 16408 3940
rect 18113 3937 18125 3940
rect 18159 3937 18171 3971
rect 20321 3971 20379 3977
rect 20321 3968 20333 3971
rect 18113 3931 18171 3937
rect 18588 3940 20333 3968
rect 18588 3909 18616 3940
rect 20321 3937 20333 3940
rect 20367 3937 20379 3971
rect 20321 3931 20379 3937
rect 9787 3872 10612 3900
rect 10845 3903 10903 3909
rect 9787 3869 9799 3872
rect 9741 3863 9799 3869
rect 10845 3869 10857 3903
rect 10891 3869 10903 3903
rect 10845 3863 10903 3869
rect 11949 3903 12007 3909
rect 11949 3869 11961 3903
rect 11995 3869 12007 3903
rect 11949 3863 12007 3869
rect 13053 3903 13111 3909
rect 13053 3869 13065 3903
rect 13099 3869 13111 3903
rect 13053 3863 13111 3869
rect 14168 3903 14226 3909
rect 14168 3869 14180 3903
rect 14214 3869 14226 3903
rect 14168 3863 14226 3869
rect 15261 3903 15319 3909
rect 15261 3869 15273 3903
rect 15307 3869 15319 3903
rect 15261 3863 15319 3869
rect 16365 3903 16423 3909
rect 16365 3869 16377 3903
rect 16411 3869 16423 3903
rect 16365 3863 16423 3869
rect 17469 3903 17527 3909
rect 17469 3869 17481 3903
rect 17515 3869 17527 3903
rect 17469 3863 17527 3869
rect 18573 3903 18631 3909
rect 18573 3869 18585 3903
rect 18619 3869 18631 3903
rect 18573 3863 18631 3869
rect 19677 3903 19735 3909
rect 19677 3869 19689 3903
rect 19723 3900 19735 3903
rect 20226 3900 20232 3912
rect 19723 3872 20232 3900
rect 19723 3869 19735 3872
rect 19677 3863 19735 3869
rect 8652 3804 9600 3832
rect 10860 3832 10888 3863
rect 12593 3835 12651 3841
rect 12593 3832 12605 3835
rect 10860 3804 12605 3832
rect 8177 3795 8235 3801
rect 12593 3801 12605 3804
rect 12639 3801 12651 3835
rect 13068 3832 13096 3863
rect 14801 3835 14859 3841
rect 14801 3832 14813 3835
rect 13068 3804 14813 3832
rect 12593 3795 12651 3801
rect 14801 3801 14813 3804
rect 14847 3801 14859 3835
rect 15276 3832 15304 3863
rect 17009 3835 17067 3841
rect 17009 3832 17021 3835
rect 15276 3804 17021 3832
rect 14801 3795 14859 3801
rect 17009 3801 17021 3804
rect 17055 3801 17067 3835
rect 17484 3832 17512 3863
rect 20226 3860 20232 3872
rect 20284 3860 20290 3912
rect 19217 3835 19275 3841
rect 19217 3832 19229 3835
rect 17484 3804 19229 3832
rect 17009 3795 17067 3801
rect 19217 3801 19229 3804
rect 19263 3801 19275 3835
rect 19217 3795 19275 3801
rect 1904 3674 20764 3696
rect 1904 3622 4446 3674
rect 4498 3622 4510 3674
rect 4562 3622 4574 3674
rect 4626 3622 4638 3674
rect 4690 3622 9774 3674
rect 9826 3622 9838 3674
rect 9890 3622 9902 3674
rect 9954 3622 9966 3674
rect 10018 3622 15102 3674
rect 15154 3622 15166 3674
rect 15218 3622 15230 3674
rect 15282 3622 15294 3674
rect 15346 3622 20764 3674
rect 1904 3600 20764 3622
rect 20226 3452 20232 3504
rect 20284 3492 20290 3504
rect 20321 3495 20379 3501
rect 20321 3492 20333 3495
rect 20284 3464 20333 3492
rect 20284 3452 20290 3464
rect 20321 3461 20333 3464
rect 20367 3461 20379 3495
rect 20321 3455 20379 3461
rect 3117 3427 3175 3433
rect 3117 3393 3129 3427
rect 3163 3393 3175 3427
rect 3117 3387 3175 3393
rect 3761 3427 3819 3433
rect 3761 3393 3773 3427
rect 3807 3424 3819 3427
rect 4221 3427 4279 3433
rect 4221 3424 4233 3427
rect 3807 3396 4233 3424
rect 3807 3393 3819 3396
rect 3761 3387 3819 3393
rect 4221 3393 4233 3396
rect 4267 3393 4279 3427
rect 4221 3387 4279 3393
rect 4865 3427 4923 3433
rect 4865 3393 4877 3427
rect 4911 3424 4923 3427
rect 5325 3427 5383 3433
rect 5325 3424 5337 3427
rect 4911 3396 5337 3424
rect 4911 3393 4923 3396
rect 4865 3387 4923 3393
rect 5325 3393 5337 3396
rect 5371 3393 5383 3427
rect 5325 3387 5383 3393
rect 5969 3427 6027 3433
rect 5969 3393 5981 3427
rect 6015 3424 6027 3427
rect 6429 3427 6487 3433
rect 6429 3424 6441 3427
rect 6015 3396 6441 3424
rect 6015 3393 6027 3396
rect 5969 3387 6027 3393
rect 6429 3393 6441 3396
rect 6475 3393 6487 3427
rect 6429 3387 6487 3393
rect 7073 3427 7131 3433
rect 7073 3393 7085 3427
rect 7119 3424 7131 3427
rect 7533 3427 7591 3433
rect 7533 3424 7545 3427
rect 7119 3396 7545 3424
rect 7119 3393 7131 3396
rect 7073 3387 7131 3393
rect 7533 3393 7545 3396
rect 7579 3393 7591 3427
rect 7533 3387 7591 3393
rect 8177 3427 8235 3433
rect 8177 3393 8189 3427
rect 8223 3424 8235 3427
rect 8637 3427 8695 3433
rect 8637 3424 8649 3427
rect 8223 3396 8649 3424
rect 8223 3393 8235 3396
rect 8177 3387 8235 3393
rect 8637 3393 8649 3396
rect 8683 3393 8695 3427
rect 8637 3387 8695 3393
rect 9281 3427 9339 3433
rect 9281 3393 9293 3427
rect 9327 3424 9339 3427
rect 9741 3427 9799 3433
rect 9741 3424 9753 3427
rect 9327 3396 9753 3424
rect 9327 3393 9339 3396
rect 9281 3387 9339 3393
rect 9741 3393 9753 3396
rect 9787 3393 9799 3427
rect 9741 3387 9799 3393
rect 10385 3427 10443 3433
rect 10385 3393 10397 3427
rect 10431 3424 10443 3427
rect 10845 3427 10903 3433
rect 10845 3424 10857 3427
rect 10431 3396 10857 3424
rect 10431 3393 10443 3396
rect 10385 3387 10443 3393
rect 10845 3393 10857 3396
rect 10891 3393 10903 3427
rect 10845 3387 10903 3393
rect 11489 3427 11547 3433
rect 11489 3393 11501 3427
rect 11535 3424 11547 3427
rect 11949 3427 12007 3433
rect 11949 3424 11961 3427
rect 11535 3396 11961 3424
rect 11535 3393 11547 3396
rect 11489 3387 11547 3393
rect 11949 3393 11961 3396
rect 11995 3393 12007 3427
rect 11949 3387 12007 3393
rect 12593 3427 12651 3433
rect 12593 3393 12605 3427
rect 12639 3424 12651 3427
rect 13053 3427 13111 3433
rect 13053 3424 13065 3427
rect 12639 3396 13065 3424
rect 12639 3393 12651 3396
rect 12593 3387 12651 3393
rect 13053 3393 13065 3396
rect 13099 3393 13111 3427
rect 13053 3387 13111 3393
rect 13697 3427 13755 3433
rect 13697 3393 13709 3427
rect 13743 3424 13755 3427
rect 14157 3427 14215 3433
rect 14157 3424 14169 3427
rect 13743 3396 14169 3424
rect 13743 3393 13755 3396
rect 13697 3387 13755 3393
rect 14157 3393 14169 3396
rect 14203 3393 14215 3427
rect 14157 3387 14215 3393
rect 14801 3427 14859 3433
rect 14801 3393 14813 3427
rect 14847 3424 14859 3427
rect 15261 3427 15319 3433
rect 15261 3424 15273 3427
rect 14847 3396 15273 3424
rect 14847 3393 14859 3396
rect 14801 3387 14859 3393
rect 15261 3393 15273 3396
rect 15307 3393 15319 3427
rect 15261 3387 15319 3393
rect 15905 3427 15963 3433
rect 15905 3393 15917 3427
rect 15951 3424 15963 3427
rect 16365 3427 16423 3433
rect 16365 3424 16377 3427
rect 15951 3396 16377 3424
rect 15951 3393 15963 3396
rect 15905 3387 15963 3393
rect 16365 3393 16377 3396
rect 16411 3393 16423 3427
rect 16365 3387 16423 3393
rect 17009 3427 17067 3433
rect 17009 3393 17021 3427
rect 17055 3424 17067 3427
rect 17469 3427 17527 3433
rect 17469 3424 17481 3427
rect 17055 3396 17481 3424
rect 17055 3393 17067 3396
rect 17009 3387 17067 3393
rect 17469 3393 17481 3396
rect 17515 3393 17527 3427
rect 17469 3387 17527 3393
rect 18113 3427 18171 3433
rect 18113 3393 18125 3427
rect 18159 3424 18171 3427
rect 18573 3427 18631 3433
rect 18573 3424 18585 3427
rect 18159 3396 18585 3424
rect 18159 3393 18171 3396
rect 18113 3387 18171 3393
rect 18573 3393 18585 3396
rect 18619 3393 18631 3427
rect 18573 3387 18631 3393
rect 19217 3427 19275 3433
rect 19217 3393 19229 3427
rect 19263 3424 19275 3427
rect 19677 3427 19735 3433
rect 19677 3424 19689 3427
rect 19263 3396 19689 3424
rect 19263 3393 19275 3396
rect 19217 3387 19275 3393
rect 19677 3393 19689 3396
rect 19723 3393 19735 3427
rect 19677 3387 19735 3393
rect 3132 3288 3160 3387
rect 3758 3288 3764 3300
rect 3132 3260 3764 3288
rect 3758 3248 3764 3260
rect 3816 3248 3822 3300
rect 1904 3130 20764 3152
rect 1904 3078 7110 3130
rect 7162 3078 7174 3130
rect 7226 3078 7238 3130
rect 7290 3078 7302 3130
rect 7354 3078 12438 3130
rect 12490 3078 12502 3130
rect 12554 3078 12566 3130
rect 12618 3078 12630 3130
rect 12682 3078 17766 3130
rect 17818 3078 17830 3130
rect 17882 3078 17894 3130
rect 17946 3078 17958 3130
rect 18010 3078 20764 3130
rect 1904 3056 20764 3078
rect 3758 3016 3764 3028
rect 3719 2988 3764 3016
rect 3758 2976 3764 2988
rect 3816 2976 3822 3028
rect 5969 2883 6027 2889
rect 5969 2880 5981 2883
rect 4236 2852 5981 2880
rect 4236 2821 4264 2852
rect 5969 2849 5981 2852
rect 6015 2849 6027 2883
rect 8177 2883 8235 2889
rect 8177 2880 8189 2883
rect 5969 2843 6027 2849
rect 6444 2852 8189 2880
rect 6444 2821 6472 2852
rect 8177 2849 8189 2852
rect 8223 2849 8235 2883
rect 10385 2883 10443 2889
rect 10385 2880 10397 2883
rect 8177 2843 8235 2849
rect 8652 2852 10397 2880
rect 8652 2821 8680 2852
rect 10385 2849 10397 2852
rect 10431 2849 10443 2883
rect 12593 2883 12651 2889
rect 12593 2880 12605 2883
rect 10385 2843 10443 2849
rect 10860 2852 12605 2880
rect 10860 2821 10888 2852
rect 12593 2849 12605 2852
rect 12639 2849 12651 2883
rect 14801 2883 14859 2889
rect 14801 2880 14813 2883
rect 12593 2843 12651 2849
rect 13068 2852 14813 2880
rect 13068 2821 13096 2852
rect 14801 2849 14813 2852
rect 14847 2849 14859 2883
rect 17009 2883 17067 2889
rect 17009 2880 17021 2883
rect 14801 2843 14859 2849
rect 15276 2852 17021 2880
rect 3117 2815 3175 2821
rect 3117 2781 3129 2815
rect 3163 2812 3175 2815
rect 4232 2815 4290 2821
rect 3163 2784 3804 2812
rect 3163 2781 3175 2784
rect 3117 2775 3175 2781
rect 3776 2744 3804 2784
rect 4232 2781 4244 2815
rect 4278 2781 4290 2815
rect 4232 2775 4290 2781
rect 5325 2815 5383 2821
rect 5325 2781 5337 2815
rect 5371 2812 5383 2815
rect 6429 2815 6487 2821
rect 5371 2784 6196 2812
rect 5371 2781 5383 2784
rect 5325 2775 5383 2781
rect 4865 2747 4923 2753
rect 4865 2744 4877 2747
rect 3776 2716 4877 2744
rect 4865 2713 4877 2716
rect 4911 2713 4923 2747
rect 6168 2744 6196 2784
rect 6429 2781 6441 2815
rect 6475 2781 6487 2815
rect 6429 2775 6487 2781
rect 7533 2815 7591 2821
rect 7533 2781 7545 2815
rect 7579 2812 7591 2815
rect 8648 2815 8706 2821
rect 7579 2784 8404 2812
rect 7579 2781 7591 2784
rect 7533 2775 7591 2781
rect 7073 2747 7131 2753
rect 7073 2744 7085 2747
rect 6168 2716 7085 2744
rect 4865 2707 4923 2713
rect 7073 2713 7085 2716
rect 7119 2713 7131 2747
rect 8376 2744 8404 2784
rect 8648 2781 8660 2815
rect 8694 2781 8706 2815
rect 8648 2775 8706 2781
rect 9741 2815 9799 2821
rect 9741 2781 9753 2815
rect 9787 2812 9799 2815
rect 10845 2815 10903 2821
rect 9787 2784 10612 2812
rect 9787 2781 9799 2784
rect 9741 2775 9799 2781
rect 9281 2747 9339 2753
rect 9281 2744 9293 2747
rect 8376 2716 9293 2744
rect 7073 2707 7131 2713
rect 9281 2713 9293 2716
rect 9327 2713 9339 2747
rect 10584 2744 10612 2784
rect 10845 2781 10857 2815
rect 10891 2781 10903 2815
rect 10845 2775 10903 2781
rect 11949 2815 12007 2821
rect 11949 2781 11961 2815
rect 11995 2812 12007 2815
rect 13053 2815 13111 2821
rect 11995 2784 12820 2812
rect 11995 2781 12007 2784
rect 11949 2775 12007 2781
rect 11489 2747 11547 2753
rect 11489 2744 11501 2747
rect 10584 2716 11501 2744
rect 9281 2707 9339 2713
rect 11489 2713 11501 2716
rect 11535 2713 11547 2747
rect 12792 2744 12820 2784
rect 13053 2781 13065 2815
rect 13099 2781 13111 2815
rect 13053 2775 13111 2781
rect 14157 2815 14215 2821
rect 14157 2781 14169 2815
rect 14203 2812 14215 2815
rect 14982 2812 14988 2824
rect 14203 2784 14988 2812
rect 14203 2781 14215 2784
rect 14157 2775 14215 2781
rect 14982 2772 14988 2784
rect 15040 2772 15046 2824
rect 15276 2821 15304 2852
rect 17009 2849 17021 2852
rect 17055 2849 17067 2883
rect 19217 2883 19275 2889
rect 19217 2880 19229 2883
rect 17009 2843 17067 2849
rect 17484 2852 19229 2880
rect 17484 2821 17512 2852
rect 19217 2849 19229 2852
rect 19263 2849 19275 2883
rect 19217 2843 19275 2849
rect 15261 2815 15319 2821
rect 15261 2781 15273 2815
rect 15307 2781 15319 2815
rect 15261 2775 15319 2781
rect 16365 2815 16423 2821
rect 16365 2781 16377 2815
rect 16411 2812 16423 2815
rect 17469 2815 17527 2821
rect 16411 2784 17236 2812
rect 16411 2781 16423 2784
rect 16365 2775 16423 2781
rect 13697 2747 13755 2753
rect 13697 2744 13709 2747
rect 12792 2716 13709 2744
rect 11489 2707 11547 2713
rect 13697 2713 13709 2716
rect 13743 2713 13755 2747
rect 17208 2744 17236 2784
rect 17469 2781 17481 2815
rect 17515 2781 17527 2815
rect 17469 2775 17527 2781
rect 18573 2815 18631 2821
rect 18573 2781 18585 2815
rect 18619 2812 18631 2815
rect 19677 2815 19735 2821
rect 18619 2784 19260 2812
rect 18619 2781 18631 2784
rect 18573 2775 18631 2781
rect 18113 2747 18171 2753
rect 18113 2744 18125 2747
rect 17208 2716 18125 2744
rect 13697 2707 13755 2713
rect 18113 2713 18125 2716
rect 18159 2713 18171 2747
rect 19232 2744 19260 2784
rect 19677 2781 19689 2815
rect 19723 2812 19735 2815
rect 20134 2812 20140 2824
rect 19723 2784 20140 2812
rect 19723 2781 19735 2784
rect 19677 2775 19735 2781
rect 20134 2772 20140 2784
rect 20192 2772 20198 2824
rect 20321 2747 20379 2753
rect 20321 2744 20333 2747
rect 19232 2716 20333 2744
rect 18113 2707 18171 2713
rect 20321 2713 20333 2716
rect 20367 2713 20379 2747
rect 20321 2707 20379 2713
rect 14982 2636 14988 2688
rect 15040 2676 15046 2688
rect 15905 2679 15963 2685
rect 15905 2676 15917 2679
rect 15040 2648 15917 2676
rect 15040 2636 15046 2648
rect 15905 2645 15917 2648
rect 15951 2645 15963 2679
rect 15905 2639 15963 2645
rect 1904 2586 20764 2608
rect 1904 2534 4446 2586
rect 4498 2534 4510 2586
rect 4562 2534 4574 2586
rect 4626 2534 4638 2586
rect 4690 2534 9774 2586
rect 9826 2534 9838 2586
rect 9890 2534 9902 2586
rect 9954 2534 9966 2586
rect 10018 2534 15102 2586
rect 15154 2534 15166 2586
rect 15218 2534 15230 2586
rect 15282 2534 15294 2586
rect 15346 2534 20764 2586
rect 1904 2512 20764 2534
rect 20134 2432 20140 2484
rect 20192 2472 20198 2484
rect 20321 2475 20379 2481
rect 20321 2472 20333 2475
rect 20192 2444 20333 2472
rect 20192 2432 20198 2444
rect 20321 2441 20333 2444
rect 20367 2441 20379 2475
rect 20321 2435 20379 2441
rect 3117 2339 3175 2345
rect 3117 2305 3129 2339
rect 3163 2305 3175 2339
rect 3117 2299 3175 2305
rect 3761 2339 3819 2345
rect 3761 2305 3773 2339
rect 3807 2336 3819 2339
rect 4221 2339 4279 2345
rect 4221 2336 4233 2339
rect 3807 2308 4233 2336
rect 3807 2305 3819 2308
rect 3761 2299 3819 2305
rect 4221 2305 4233 2308
rect 4267 2305 4279 2339
rect 4221 2299 4279 2305
rect 4865 2339 4923 2345
rect 4865 2305 4877 2339
rect 4911 2336 4923 2339
rect 5325 2339 5383 2345
rect 5325 2336 5337 2339
rect 4911 2308 5337 2336
rect 4911 2305 4923 2308
rect 4865 2299 4923 2305
rect 5325 2305 5337 2308
rect 5371 2305 5383 2339
rect 5325 2299 5383 2305
rect 5969 2339 6027 2345
rect 5969 2305 5981 2339
rect 6015 2336 6027 2339
rect 6429 2339 6487 2345
rect 6429 2336 6441 2339
rect 6015 2308 6441 2336
rect 6015 2305 6027 2308
rect 5969 2299 6027 2305
rect 6429 2305 6441 2308
rect 6475 2305 6487 2339
rect 6429 2299 6487 2305
rect 7073 2339 7131 2345
rect 7073 2305 7085 2339
rect 7119 2336 7131 2339
rect 7533 2339 7591 2345
rect 7533 2336 7545 2339
rect 7119 2308 7545 2336
rect 7119 2305 7131 2308
rect 7073 2299 7131 2305
rect 7533 2305 7545 2308
rect 7579 2305 7591 2339
rect 7533 2299 7591 2305
rect 8177 2339 8235 2345
rect 8177 2305 8189 2339
rect 8223 2336 8235 2339
rect 8637 2339 8695 2345
rect 8637 2336 8649 2339
rect 8223 2308 8649 2336
rect 8223 2305 8235 2308
rect 8177 2299 8235 2305
rect 8637 2305 8649 2308
rect 8683 2305 8695 2339
rect 8637 2299 8695 2305
rect 9281 2339 9339 2345
rect 9281 2305 9293 2339
rect 9327 2336 9339 2339
rect 9741 2339 9799 2345
rect 9741 2336 9753 2339
rect 9327 2308 9753 2336
rect 9327 2305 9339 2308
rect 9281 2299 9339 2305
rect 9741 2305 9753 2308
rect 9787 2305 9799 2339
rect 9741 2299 9799 2305
rect 10385 2339 10443 2345
rect 10385 2305 10397 2339
rect 10431 2336 10443 2339
rect 10845 2339 10903 2345
rect 10845 2336 10857 2339
rect 10431 2308 10857 2336
rect 10431 2305 10443 2308
rect 10385 2299 10443 2305
rect 10845 2305 10857 2308
rect 10891 2305 10903 2339
rect 10845 2299 10903 2305
rect 11489 2339 11547 2345
rect 11489 2305 11501 2339
rect 11535 2336 11547 2339
rect 11949 2339 12007 2345
rect 11949 2336 11961 2339
rect 11535 2308 11961 2336
rect 11535 2305 11547 2308
rect 11489 2299 11547 2305
rect 11949 2305 11961 2308
rect 11995 2305 12007 2339
rect 11949 2299 12007 2305
rect 12593 2339 12651 2345
rect 12593 2305 12605 2339
rect 12639 2336 12651 2339
rect 13053 2339 13111 2345
rect 13053 2336 13065 2339
rect 12639 2308 13065 2336
rect 12639 2305 12651 2308
rect 12593 2299 12651 2305
rect 13053 2305 13065 2308
rect 13099 2305 13111 2339
rect 13053 2299 13111 2305
rect 13697 2339 13755 2345
rect 13697 2305 13709 2339
rect 13743 2336 13755 2339
rect 14157 2339 14215 2345
rect 14157 2336 14169 2339
rect 13743 2308 14169 2336
rect 13743 2305 13755 2308
rect 13697 2299 13755 2305
rect 14157 2305 14169 2308
rect 14203 2305 14215 2339
rect 14157 2299 14215 2305
rect 14801 2339 14859 2345
rect 14801 2305 14813 2339
rect 14847 2336 14859 2339
rect 15261 2339 15319 2345
rect 15261 2336 15273 2339
rect 14847 2308 15273 2336
rect 14847 2305 14859 2308
rect 14801 2299 14859 2305
rect 15261 2305 15273 2308
rect 15307 2305 15319 2339
rect 15261 2299 15319 2305
rect 15905 2339 15963 2345
rect 15905 2305 15917 2339
rect 15951 2336 15963 2339
rect 16365 2339 16423 2345
rect 16365 2336 16377 2339
rect 15951 2308 16377 2336
rect 15951 2305 15963 2308
rect 15905 2299 15963 2305
rect 16365 2305 16377 2308
rect 16411 2305 16423 2339
rect 16365 2299 16423 2305
rect 17009 2339 17067 2345
rect 17009 2305 17021 2339
rect 17055 2336 17067 2339
rect 17469 2339 17527 2345
rect 17469 2336 17481 2339
rect 17055 2308 17481 2336
rect 17055 2305 17067 2308
rect 17009 2299 17067 2305
rect 17469 2305 17481 2308
rect 17515 2305 17527 2339
rect 17469 2299 17527 2305
rect 18113 2339 18171 2345
rect 18113 2305 18125 2339
rect 18159 2336 18171 2339
rect 18573 2339 18631 2345
rect 18573 2336 18585 2339
rect 18159 2308 18585 2336
rect 18159 2305 18171 2308
rect 18113 2299 18171 2305
rect 18573 2305 18585 2308
rect 18619 2305 18631 2339
rect 18573 2299 18631 2305
rect 19217 2339 19275 2345
rect 19217 2305 19229 2339
rect 19263 2336 19275 2339
rect 19677 2339 19735 2345
rect 19677 2336 19689 2339
rect 19263 2308 19689 2336
rect 19263 2305 19275 2308
rect 19217 2299 19275 2305
rect 19677 2305 19689 2308
rect 19723 2305 19735 2339
rect 19677 2299 19735 2305
rect 3132 2200 3160 2299
rect 3758 2200 3764 2212
rect 3132 2172 3764 2200
rect 3758 2160 3764 2172
rect 3816 2160 3822 2212
rect 1904 2042 20764 2064
rect 1904 1990 7110 2042
rect 7162 1990 7174 2042
rect 7226 1990 7238 2042
rect 7290 1990 7302 2042
rect 7354 1990 12438 2042
rect 12490 1990 12502 2042
rect 12554 1990 12566 2042
rect 12618 1990 12630 2042
rect 12682 1990 17766 2042
rect 17818 1990 17830 2042
rect 17882 1990 17894 2042
rect 17946 1990 17958 2042
rect 18010 1990 20764 2042
rect 1904 1968 20764 1990
rect 3758 1928 3764 1940
rect 3719 1900 3764 1928
rect 3758 1888 3764 1900
rect 3816 1888 3822 1940
rect 7073 1795 7131 1801
rect 7073 1792 7085 1795
rect 4236 1764 5276 1792
rect 4236 1733 4264 1764
rect 3117 1727 3175 1733
rect 3117 1693 3129 1727
rect 3163 1693 3175 1727
rect 3117 1687 3175 1693
rect 4232 1727 4290 1733
rect 4232 1693 4244 1727
rect 4278 1693 4290 1727
rect 4232 1687 4290 1693
rect 3132 1656 3160 1687
rect 4865 1659 4923 1665
rect 4865 1656 4877 1659
rect 3132 1628 4877 1656
rect 4865 1625 4877 1628
rect 4911 1625 4923 1659
rect 5248 1656 5276 1764
rect 5340 1764 7085 1792
rect 5340 1733 5368 1764
rect 7073 1761 7085 1764
rect 7119 1761 7131 1795
rect 9281 1795 9339 1801
rect 9281 1792 9293 1795
rect 7073 1755 7131 1761
rect 7548 1764 9293 1792
rect 7548 1733 7576 1764
rect 9281 1761 9293 1764
rect 9327 1761 9339 1795
rect 10385 1795 10443 1801
rect 10385 1792 10397 1795
rect 9281 1755 9339 1761
rect 9572 1764 10397 1792
rect 5325 1727 5383 1733
rect 5325 1693 5337 1727
rect 5371 1693 5383 1727
rect 5325 1687 5383 1693
rect 6429 1727 6487 1733
rect 6429 1693 6441 1727
rect 6475 1693 6487 1727
rect 6429 1687 6487 1693
rect 7533 1727 7591 1733
rect 7533 1693 7545 1727
rect 7579 1693 7591 1727
rect 7533 1687 7591 1693
rect 8648 1727 8706 1733
rect 8648 1693 8660 1727
rect 8694 1693 8706 1727
rect 8648 1687 8706 1693
rect 5969 1659 6027 1665
rect 5969 1656 5981 1659
rect 5248 1628 5981 1656
rect 4865 1619 4923 1625
rect 5969 1625 5981 1628
rect 6015 1625 6027 1659
rect 6444 1656 6472 1687
rect 8177 1659 8235 1665
rect 8177 1656 8189 1659
rect 6444 1628 8189 1656
rect 5969 1619 6027 1625
rect 8177 1625 8189 1628
rect 8223 1625 8235 1659
rect 8652 1656 8680 1687
rect 9572 1656 9600 1764
rect 10385 1761 10397 1764
rect 10431 1761 10443 1795
rect 11489 1795 11547 1801
rect 11489 1792 11501 1795
rect 10385 1755 10443 1761
rect 10584 1764 11501 1792
rect 9741 1727 9799 1733
rect 9741 1693 9753 1727
rect 9787 1724 9799 1727
rect 10584 1724 10612 1764
rect 11489 1761 11501 1764
rect 11535 1761 11547 1795
rect 13697 1795 13755 1801
rect 13697 1792 13709 1795
rect 11489 1755 11547 1761
rect 11964 1764 13709 1792
rect 11964 1733 11992 1764
rect 13697 1761 13709 1764
rect 13743 1761 13755 1795
rect 15905 1795 15963 1801
rect 15905 1792 15917 1795
rect 13697 1755 13755 1761
rect 14172 1764 15917 1792
rect 14172 1733 14200 1764
rect 15905 1761 15917 1764
rect 15951 1761 15963 1795
rect 18113 1795 18171 1801
rect 18113 1792 18125 1795
rect 15905 1755 15963 1761
rect 16380 1764 18125 1792
rect 16380 1733 16408 1764
rect 18113 1761 18125 1764
rect 18159 1761 18171 1795
rect 20321 1795 20379 1801
rect 20321 1792 20333 1795
rect 18113 1755 18171 1761
rect 18588 1764 20333 1792
rect 18588 1733 18616 1764
rect 20321 1761 20333 1764
rect 20367 1761 20379 1795
rect 20321 1755 20379 1761
rect 9787 1696 10612 1724
rect 10845 1727 10903 1733
rect 9787 1693 9799 1696
rect 9741 1687 9799 1693
rect 10845 1693 10857 1727
rect 10891 1693 10903 1727
rect 10845 1687 10903 1693
rect 11949 1727 12007 1733
rect 11949 1693 11961 1727
rect 11995 1693 12007 1727
rect 11949 1687 12007 1693
rect 13053 1727 13111 1733
rect 13053 1693 13065 1727
rect 13099 1693 13111 1727
rect 13053 1687 13111 1693
rect 14168 1727 14226 1733
rect 14168 1693 14180 1727
rect 14214 1693 14226 1727
rect 14168 1687 14226 1693
rect 15261 1727 15319 1733
rect 15261 1693 15273 1727
rect 15307 1693 15319 1727
rect 15261 1687 15319 1693
rect 16365 1727 16423 1733
rect 16365 1693 16377 1727
rect 16411 1693 16423 1727
rect 16365 1687 16423 1693
rect 17469 1727 17527 1733
rect 17469 1693 17481 1727
rect 17515 1693 17527 1727
rect 17469 1687 17527 1693
rect 18573 1727 18631 1733
rect 18573 1693 18585 1727
rect 18619 1693 18631 1727
rect 18573 1687 18631 1693
rect 19677 1727 19735 1733
rect 19677 1693 19689 1727
rect 19723 1724 19735 1727
rect 20134 1724 20140 1736
rect 19723 1696 20140 1724
rect 19723 1693 19735 1696
rect 19677 1687 19735 1693
rect 8652 1628 9600 1656
rect 10860 1656 10888 1687
rect 12593 1659 12651 1665
rect 12593 1656 12605 1659
rect 10860 1628 12605 1656
rect 8177 1619 8235 1625
rect 12593 1625 12605 1628
rect 12639 1625 12651 1659
rect 13068 1656 13096 1687
rect 14801 1659 14859 1665
rect 14801 1656 14813 1659
rect 13068 1628 14813 1656
rect 12593 1619 12651 1625
rect 14801 1625 14813 1628
rect 14847 1625 14859 1659
rect 15276 1656 15304 1687
rect 17009 1659 17067 1665
rect 17009 1656 17021 1659
rect 15276 1628 17021 1656
rect 14801 1619 14859 1625
rect 17009 1625 17021 1628
rect 17055 1625 17067 1659
rect 17484 1656 17512 1687
rect 20134 1684 20140 1696
rect 20192 1684 20198 1736
rect 19217 1659 19275 1665
rect 19217 1656 19229 1659
rect 17484 1628 19229 1656
rect 17009 1619 17067 1625
rect 19217 1625 19229 1628
rect 19263 1625 19275 1659
rect 19217 1619 19275 1625
rect 1904 1498 20764 1520
rect 1904 1446 4446 1498
rect 4498 1446 4510 1498
rect 4562 1446 4574 1498
rect 4626 1446 4638 1498
rect 4690 1446 9774 1498
rect 9826 1446 9838 1498
rect 9890 1446 9902 1498
rect 9954 1446 9966 1498
rect 10018 1446 15102 1498
rect 15154 1446 15166 1498
rect 15218 1446 15230 1498
rect 15282 1446 15294 1498
rect 15346 1446 20764 1498
rect 1904 1424 20764 1446
rect 20134 1344 20140 1396
rect 20192 1384 20198 1396
rect 20321 1387 20379 1393
rect 20321 1384 20333 1387
rect 20192 1356 20333 1384
rect 20192 1344 20198 1356
rect 20321 1353 20333 1356
rect 20367 1353 20379 1387
rect 20321 1347 20379 1353
rect 2930 1208 2936 1260
rect 2988 1248 2994 1260
rect 3117 1251 3175 1257
rect 3117 1248 3129 1251
rect 2988 1220 3129 1248
rect 2988 1208 2994 1220
rect 3117 1217 3129 1220
rect 3163 1217 3175 1251
rect 3117 1211 3175 1217
rect 3761 1251 3819 1257
rect 3761 1217 3773 1251
rect 3807 1248 3819 1251
rect 4221 1251 4279 1257
rect 4221 1248 4233 1251
rect 3807 1220 4233 1248
rect 3807 1217 3819 1220
rect 3761 1211 3819 1217
rect 4221 1217 4233 1220
rect 4267 1217 4279 1251
rect 4221 1211 4279 1217
rect 4865 1251 4923 1257
rect 4865 1217 4877 1251
rect 4911 1248 4923 1251
rect 5325 1251 5383 1257
rect 5325 1248 5337 1251
rect 4911 1220 5337 1248
rect 4911 1217 4923 1220
rect 4865 1211 4923 1217
rect 5325 1217 5337 1220
rect 5371 1217 5383 1251
rect 5325 1211 5383 1217
rect 5969 1251 6027 1257
rect 5969 1217 5981 1251
rect 6015 1248 6027 1251
rect 6429 1251 6487 1257
rect 6429 1248 6441 1251
rect 6015 1220 6441 1248
rect 6015 1217 6027 1220
rect 5969 1211 6027 1217
rect 6429 1217 6441 1220
rect 6475 1217 6487 1251
rect 6429 1211 6487 1217
rect 7073 1251 7131 1257
rect 7073 1217 7085 1251
rect 7119 1248 7131 1251
rect 7533 1251 7591 1257
rect 7533 1248 7545 1251
rect 7119 1220 7545 1248
rect 7119 1217 7131 1220
rect 7073 1211 7131 1217
rect 7533 1217 7545 1220
rect 7579 1217 7591 1251
rect 7533 1211 7591 1217
rect 8177 1251 8235 1257
rect 8177 1217 8189 1251
rect 8223 1248 8235 1251
rect 8637 1251 8695 1257
rect 8637 1248 8649 1251
rect 8223 1220 8649 1248
rect 8223 1217 8235 1220
rect 8177 1211 8235 1217
rect 8637 1217 8649 1220
rect 8683 1217 8695 1251
rect 8637 1211 8695 1217
rect 9281 1251 9339 1257
rect 9281 1217 9293 1251
rect 9327 1248 9339 1251
rect 9741 1251 9799 1257
rect 9741 1248 9753 1251
rect 9327 1220 9753 1248
rect 9327 1217 9339 1220
rect 9281 1211 9339 1217
rect 9741 1217 9753 1220
rect 9787 1217 9799 1251
rect 9741 1211 9799 1217
rect 10385 1251 10443 1257
rect 10385 1217 10397 1251
rect 10431 1248 10443 1251
rect 10845 1251 10903 1257
rect 10845 1248 10857 1251
rect 10431 1220 10857 1248
rect 10431 1217 10443 1220
rect 10385 1211 10443 1217
rect 10845 1217 10857 1220
rect 10891 1217 10903 1251
rect 10845 1211 10903 1217
rect 11489 1251 11547 1257
rect 11489 1217 11501 1251
rect 11535 1248 11547 1251
rect 11949 1251 12007 1257
rect 11949 1248 11961 1251
rect 11535 1220 11961 1248
rect 11535 1217 11547 1220
rect 11489 1211 11547 1217
rect 11949 1217 11961 1220
rect 11995 1217 12007 1251
rect 11949 1211 12007 1217
rect 12593 1251 12651 1257
rect 12593 1217 12605 1251
rect 12639 1248 12651 1251
rect 13053 1251 13111 1257
rect 13053 1248 13065 1251
rect 12639 1220 13065 1248
rect 12639 1217 12651 1220
rect 12593 1211 12651 1217
rect 13053 1217 13065 1220
rect 13099 1217 13111 1251
rect 13053 1211 13111 1217
rect 13697 1251 13755 1257
rect 13697 1217 13709 1251
rect 13743 1248 13755 1251
rect 14157 1251 14215 1257
rect 14157 1248 14169 1251
rect 13743 1220 14169 1248
rect 13743 1217 13755 1220
rect 13697 1211 13755 1217
rect 14157 1217 14169 1220
rect 14203 1217 14215 1251
rect 14157 1211 14215 1217
rect 14801 1251 14859 1257
rect 14801 1217 14813 1251
rect 14847 1248 14859 1251
rect 15261 1251 15319 1257
rect 15261 1248 15273 1251
rect 14847 1220 15273 1248
rect 14847 1217 14859 1220
rect 14801 1211 14859 1217
rect 15261 1217 15273 1220
rect 15307 1217 15319 1251
rect 15261 1211 15319 1217
rect 15905 1251 15963 1257
rect 15905 1217 15917 1251
rect 15951 1248 15963 1251
rect 16365 1251 16423 1257
rect 16365 1248 16377 1251
rect 15951 1220 16377 1248
rect 15951 1217 15963 1220
rect 15905 1211 15963 1217
rect 16365 1217 16377 1220
rect 16411 1217 16423 1251
rect 16365 1211 16423 1217
rect 17009 1251 17067 1257
rect 17009 1217 17021 1251
rect 17055 1248 17067 1251
rect 17469 1251 17527 1257
rect 17469 1248 17481 1251
rect 17055 1220 17481 1248
rect 17055 1217 17067 1220
rect 17009 1211 17067 1217
rect 17469 1217 17481 1220
rect 17515 1217 17527 1251
rect 17469 1211 17527 1217
rect 18113 1251 18171 1257
rect 18113 1217 18125 1251
rect 18159 1248 18171 1251
rect 18573 1251 18631 1257
rect 18573 1248 18585 1251
rect 18159 1220 18585 1248
rect 18159 1217 18171 1220
rect 18113 1211 18171 1217
rect 18573 1217 18585 1220
rect 18619 1217 18631 1251
rect 18573 1211 18631 1217
rect 19217 1251 19275 1257
rect 19217 1217 19229 1251
rect 19263 1248 19275 1251
rect 19677 1251 19735 1257
rect 19677 1248 19689 1251
rect 19263 1220 19689 1248
rect 19263 1217 19275 1220
rect 19217 1211 19275 1217
rect 19677 1217 19689 1220
rect 19723 1217 19735 1251
rect 19677 1211 19735 1217
rect 1904 954 20764 976
rect 1904 902 7110 954
rect 7162 902 7174 954
rect 7226 902 7238 954
rect 7290 902 7302 954
rect 7354 902 12438 954
rect 12490 902 12502 954
rect 12554 902 12566 954
rect 12618 902 12630 954
rect 12682 902 17766 954
rect 17818 902 17830 954
rect 17882 902 17894 954
rect 17946 902 17958 954
rect 18010 902 20764 954
rect 1904 880 20764 902
<< via1 >>
rect 4446 22118 4498 22170
rect 4510 22118 4562 22170
rect 4574 22118 4626 22170
rect 4638 22118 4690 22170
rect 9774 22118 9826 22170
rect 9838 22118 9890 22170
rect 9902 22118 9954 22170
rect 9966 22118 10018 22170
rect 15102 22118 15154 22170
rect 15166 22118 15218 22170
rect 15230 22118 15282 22170
rect 15294 22118 15346 22170
rect 1924 22059 1976 22068
rect 1924 22025 1933 22059
rect 1933 22025 1967 22059
rect 1967 22025 1976 22059
rect 1924 22016 1976 22025
rect 2292 21991 2344 22000
rect 2292 21957 2301 21991
rect 2301 21957 2335 21991
rect 2335 21957 2344 21991
rect 2292 21948 2344 21957
rect 2476 21855 2528 21864
rect 2476 21821 2485 21855
rect 2485 21821 2519 21855
rect 2519 21821 2528 21855
rect 2476 21812 2528 21821
rect 7110 21574 7162 21626
rect 7174 21574 7226 21626
rect 7238 21574 7290 21626
rect 7302 21574 7354 21626
rect 12438 21574 12490 21626
rect 12502 21574 12554 21626
rect 12566 21574 12618 21626
rect 12630 21574 12682 21626
rect 17766 21574 17818 21626
rect 17830 21574 17882 21626
rect 17894 21574 17946 21626
rect 17958 21574 18010 21626
rect 2292 21472 2344 21524
rect 2476 21379 2528 21388
rect 2476 21345 2485 21379
rect 2485 21345 2519 21379
rect 2519 21345 2528 21379
rect 2476 21336 2528 21345
rect 2292 21243 2344 21252
rect 2292 21209 2301 21243
rect 2301 21209 2335 21243
rect 2335 21209 2344 21243
rect 3856 21268 3908 21320
rect 2292 21200 2344 21209
rect 4446 21030 4498 21082
rect 4510 21030 4562 21082
rect 4574 21030 4626 21082
rect 4638 21030 4690 21082
rect 9774 21030 9826 21082
rect 9838 21030 9890 21082
rect 9902 21030 9954 21082
rect 9966 21030 10018 21082
rect 15102 21030 15154 21082
rect 15166 21030 15218 21082
rect 15230 21030 15282 21082
rect 15294 21030 15346 21082
rect 3856 20928 3908 20980
rect 2292 20792 2344 20844
rect 7110 20486 7162 20538
rect 7174 20486 7226 20538
rect 7238 20486 7290 20538
rect 7302 20486 7354 20538
rect 12438 20486 12490 20538
rect 12502 20486 12554 20538
rect 12566 20486 12618 20538
rect 12630 20486 12682 20538
rect 17766 20486 17818 20538
rect 17830 20486 17882 20538
rect 17894 20486 17946 20538
rect 17958 20486 18010 20538
rect 2292 20384 2344 20436
rect 2476 20291 2528 20300
rect 2476 20257 2485 20291
rect 2485 20257 2519 20291
rect 2519 20257 2528 20291
rect 2476 20248 2528 20257
rect 4224 20223 4276 20232
rect 4224 20189 4233 20223
rect 4233 20189 4267 20223
rect 4267 20189 4276 20223
rect 4224 20180 4276 20189
rect 2292 20087 2344 20096
rect 2292 20053 2301 20087
rect 2301 20053 2335 20087
rect 2335 20053 2344 20087
rect 2292 20044 2344 20053
rect 4446 19942 4498 19994
rect 4510 19942 4562 19994
rect 4574 19942 4626 19994
rect 4638 19942 4690 19994
rect 9774 19942 9826 19994
rect 9838 19942 9890 19994
rect 9902 19942 9954 19994
rect 9966 19942 10018 19994
rect 15102 19942 15154 19994
rect 15166 19942 15218 19994
rect 15230 19942 15282 19994
rect 15294 19942 15346 19994
rect 4224 19840 4276 19892
rect 2292 19704 2344 19756
rect 7110 19398 7162 19450
rect 7174 19398 7226 19450
rect 7238 19398 7290 19450
rect 7302 19398 7354 19450
rect 12438 19398 12490 19450
rect 12502 19398 12554 19450
rect 12566 19398 12618 19450
rect 12630 19398 12682 19450
rect 17766 19398 17818 19450
rect 17830 19398 17882 19450
rect 17894 19398 17946 19450
rect 17958 19398 18010 19450
rect 2292 19296 2344 19348
rect 2476 19203 2528 19212
rect 2476 19169 2485 19203
rect 2485 19169 2519 19203
rect 2519 19169 2528 19203
rect 2476 19160 2528 19169
rect 6984 19092 7036 19144
rect 2292 18999 2344 19008
rect 2292 18965 2301 18999
rect 2301 18965 2335 18999
rect 2335 18965 2344 18999
rect 2292 18956 2344 18965
rect 4446 18854 4498 18906
rect 4510 18854 4562 18906
rect 4574 18854 4626 18906
rect 4638 18854 4690 18906
rect 9774 18854 9826 18906
rect 9838 18854 9890 18906
rect 9902 18854 9954 18906
rect 9966 18854 10018 18906
rect 15102 18854 15154 18906
rect 15166 18854 15218 18906
rect 15230 18854 15282 18906
rect 15294 18854 15346 18906
rect 6984 18752 7036 18804
rect 2292 18616 2344 18668
rect 7110 18310 7162 18362
rect 7174 18310 7226 18362
rect 7238 18310 7290 18362
rect 7302 18310 7354 18362
rect 12438 18310 12490 18362
rect 12502 18310 12554 18362
rect 12566 18310 12618 18362
rect 12630 18310 12682 18362
rect 17766 18310 17818 18362
rect 17830 18310 17882 18362
rect 17894 18310 17946 18362
rect 17958 18310 18010 18362
rect 2292 18208 2344 18260
rect 2476 18115 2528 18124
rect 2476 18081 2485 18115
rect 2485 18081 2519 18115
rect 2519 18081 2528 18115
rect 2476 18072 2528 18081
rect 10848 18047 10900 18056
rect 10848 18013 10857 18047
rect 10857 18013 10891 18047
rect 10891 18013 10900 18047
rect 10848 18004 10900 18013
rect 2292 17911 2344 17920
rect 2292 17877 2301 17911
rect 2301 17877 2335 17911
rect 2335 17877 2344 17911
rect 2292 17868 2344 17877
rect 4446 17766 4498 17818
rect 4510 17766 4562 17818
rect 4574 17766 4626 17818
rect 4638 17766 4690 17818
rect 9774 17766 9826 17818
rect 9838 17766 9890 17818
rect 9902 17766 9954 17818
rect 9966 17766 10018 17818
rect 15102 17766 15154 17818
rect 15166 17766 15218 17818
rect 15230 17766 15282 17818
rect 15294 17766 15346 17818
rect 10848 17664 10900 17716
rect 2292 17528 2344 17580
rect 7110 17222 7162 17274
rect 7174 17222 7226 17274
rect 7238 17222 7290 17274
rect 7302 17222 7354 17274
rect 12438 17222 12490 17274
rect 12502 17222 12554 17274
rect 12566 17222 12618 17274
rect 12630 17222 12682 17274
rect 17766 17222 17818 17274
rect 17830 17222 17882 17274
rect 17894 17222 17946 17274
rect 17958 17222 18010 17274
rect 2292 17120 2344 17172
rect 2476 17027 2528 17036
rect 2476 16993 2485 17027
rect 2485 16993 2519 17027
rect 2519 16993 2528 17027
rect 2476 16984 2528 16993
rect 20140 16916 20192 16968
rect 2292 16823 2344 16832
rect 2292 16789 2301 16823
rect 2301 16789 2335 16823
rect 2335 16789 2344 16823
rect 2292 16780 2344 16789
rect 4446 16678 4498 16730
rect 4510 16678 4562 16730
rect 4574 16678 4626 16730
rect 4638 16678 4690 16730
rect 9774 16678 9826 16730
rect 9838 16678 9890 16730
rect 9902 16678 9954 16730
rect 9966 16678 10018 16730
rect 15102 16678 15154 16730
rect 15166 16678 15218 16730
rect 15230 16678 15282 16730
rect 15294 16678 15346 16730
rect 20140 16576 20192 16628
rect 2292 16440 2344 16492
rect 2568 16440 2620 16492
rect 7110 16134 7162 16186
rect 7174 16134 7226 16186
rect 7238 16134 7290 16186
rect 7302 16134 7354 16186
rect 12438 16134 12490 16186
rect 12502 16134 12554 16186
rect 12566 16134 12618 16186
rect 12630 16134 12682 16186
rect 17766 16134 17818 16186
rect 17830 16134 17882 16186
rect 17894 16134 17946 16186
rect 17958 16134 18010 16186
rect 2568 15964 2620 16016
rect 2476 15939 2528 15948
rect 2476 15905 2485 15939
rect 2485 15905 2519 15939
rect 2519 15905 2528 15939
rect 2476 15896 2528 15905
rect 19680 15871 19732 15880
rect 19680 15837 19689 15871
rect 19689 15837 19723 15871
rect 19723 15837 19732 15871
rect 19680 15828 19732 15837
rect 2292 15735 2344 15744
rect 2292 15701 2301 15735
rect 2301 15701 2335 15735
rect 2335 15701 2344 15735
rect 2292 15692 2344 15701
rect 4446 15590 4498 15642
rect 4510 15590 4562 15642
rect 4574 15590 4626 15642
rect 4638 15590 4690 15642
rect 9774 15590 9826 15642
rect 9838 15590 9890 15642
rect 9902 15590 9954 15642
rect 9966 15590 10018 15642
rect 15102 15590 15154 15642
rect 15166 15590 15218 15642
rect 15230 15590 15282 15642
rect 15294 15590 15346 15642
rect 19680 15488 19732 15540
rect 3764 15216 3816 15268
rect 7110 15046 7162 15098
rect 7174 15046 7226 15098
rect 7238 15046 7290 15098
rect 7302 15046 7354 15098
rect 12438 15046 12490 15098
rect 12502 15046 12554 15098
rect 12566 15046 12618 15098
rect 12630 15046 12682 15098
rect 17766 15046 17818 15098
rect 17830 15046 17882 15098
rect 17894 15046 17946 15098
rect 17958 15046 18010 15098
rect 3764 14987 3816 14996
rect 3764 14953 3773 14987
rect 3773 14953 3807 14987
rect 3807 14953 3816 14987
rect 3764 14944 3816 14953
rect 20140 14740 20192 14792
rect 4446 14502 4498 14554
rect 4510 14502 4562 14554
rect 4574 14502 4626 14554
rect 4638 14502 4690 14554
rect 9774 14502 9826 14554
rect 9838 14502 9890 14554
rect 9902 14502 9954 14554
rect 9966 14502 10018 14554
rect 15102 14502 15154 14554
rect 15166 14502 15218 14554
rect 15230 14502 15282 14554
rect 15294 14502 15346 14554
rect 20140 14400 20192 14452
rect 2292 14264 2344 14316
rect 7110 13958 7162 14010
rect 7174 13958 7226 14010
rect 7238 13958 7290 14010
rect 7302 13958 7354 14010
rect 12438 13958 12490 14010
rect 12502 13958 12554 14010
rect 12566 13958 12618 14010
rect 12630 13958 12682 14010
rect 17766 13958 17818 14010
rect 17830 13958 17882 14010
rect 17894 13958 17946 14010
rect 17958 13958 18010 14010
rect 2292 13788 2344 13840
rect 2476 13763 2528 13772
rect 2476 13729 2485 13763
rect 2485 13729 2519 13763
rect 2519 13729 2528 13763
rect 2476 13720 2528 13729
rect 19680 13695 19732 13704
rect 19680 13661 19689 13695
rect 19689 13661 19723 13695
rect 19723 13661 19732 13695
rect 19680 13652 19732 13661
rect 2292 13559 2344 13568
rect 2292 13525 2301 13559
rect 2301 13525 2335 13559
rect 2335 13525 2344 13559
rect 2292 13516 2344 13525
rect 4446 13414 4498 13466
rect 4510 13414 4562 13466
rect 4574 13414 4626 13466
rect 4638 13414 4690 13466
rect 9774 13414 9826 13466
rect 9838 13414 9890 13466
rect 9902 13414 9954 13466
rect 9966 13414 10018 13466
rect 15102 13414 15154 13466
rect 15166 13414 15218 13466
rect 15230 13414 15282 13466
rect 15294 13414 15346 13466
rect 19680 13312 19732 13364
rect 3764 13040 3816 13092
rect 7110 12870 7162 12922
rect 7174 12870 7226 12922
rect 7238 12870 7290 12922
rect 7302 12870 7354 12922
rect 12438 12870 12490 12922
rect 12502 12870 12554 12922
rect 12566 12870 12618 12922
rect 12630 12870 12682 12922
rect 17766 12870 17818 12922
rect 17830 12870 17882 12922
rect 17894 12870 17946 12922
rect 17958 12870 18010 12922
rect 3764 12811 3816 12820
rect 3764 12777 3773 12811
rect 3773 12777 3807 12811
rect 3807 12777 3816 12811
rect 3764 12768 3816 12777
rect 20140 12564 20192 12616
rect 4446 12326 4498 12378
rect 4510 12326 4562 12378
rect 4574 12326 4626 12378
rect 4638 12326 4690 12378
rect 9774 12326 9826 12378
rect 9838 12326 9890 12378
rect 9902 12326 9954 12378
rect 9966 12326 10018 12378
rect 15102 12326 15154 12378
rect 15166 12326 15218 12378
rect 15230 12326 15282 12378
rect 15294 12326 15346 12378
rect 20140 12224 20192 12276
rect 3764 11952 3816 12004
rect 7110 11782 7162 11834
rect 7174 11782 7226 11834
rect 7238 11782 7290 11834
rect 7302 11782 7354 11834
rect 12438 11782 12490 11834
rect 12502 11782 12554 11834
rect 12566 11782 12618 11834
rect 12630 11782 12682 11834
rect 17766 11782 17818 11834
rect 17830 11782 17882 11834
rect 17894 11782 17946 11834
rect 17958 11782 18010 11834
rect 3764 11587 3816 11596
rect 3764 11553 3773 11587
rect 3773 11553 3807 11587
rect 3807 11553 3816 11587
rect 3764 11544 3816 11553
rect 19680 11519 19732 11528
rect 19680 11485 19689 11519
rect 19689 11485 19723 11519
rect 19723 11485 19732 11519
rect 19680 11476 19732 11485
rect 4446 11238 4498 11290
rect 4510 11238 4562 11290
rect 4574 11238 4626 11290
rect 4638 11238 4690 11290
rect 9774 11238 9826 11290
rect 9838 11238 9890 11290
rect 9902 11238 9954 11290
rect 9966 11238 10018 11290
rect 15102 11238 15154 11290
rect 15166 11238 15218 11290
rect 15230 11238 15282 11290
rect 15294 11238 15346 11290
rect 19680 11136 19732 11188
rect 3764 10864 3816 10916
rect 7110 10694 7162 10746
rect 7174 10694 7226 10746
rect 7238 10694 7290 10746
rect 7302 10694 7354 10746
rect 12438 10694 12490 10746
rect 12502 10694 12554 10746
rect 12566 10694 12618 10746
rect 12630 10694 12682 10746
rect 17766 10694 17818 10746
rect 17830 10694 17882 10746
rect 17894 10694 17946 10746
rect 17958 10694 18010 10746
rect 3764 10635 3816 10644
rect 3764 10601 3773 10635
rect 3773 10601 3807 10635
rect 3807 10601 3816 10635
rect 3764 10592 3816 10601
rect 20140 10388 20192 10440
rect 4446 10150 4498 10202
rect 4510 10150 4562 10202
rect 4574 10150 4626 10202
rect 4638 10150 4690 10202
rect 9774 10150 9826 10202
rect 9838 10150 9890 10202
rect 9902 10150 9954 10202
rect 9966 10150 10018 10202
rect 15102 10150 15154 10202
rect 15166 10150 15218 10202
rect 15230 10150 15282 10202
rect 15294 10150 15346 10202
rect 20140 10048 20192 10100
rect 2292 9912 2344 9964
rect 7110 9606 7162 9658
rect 7174 9606 7226 9658
rect 7238 9606 7290 9658
rect 7302 9606 7354 9658
rect 12438 9606 12490 9658
rect 12502 9606 12554 9658
rect 12566 9606 12618 9658
rect 12630 9606 12682 9658
rect 17766 9606 17818 9658
rect 17830 9606 17882 9658
rect 17894 9606 17946 9658
rect 17958 9606 18010 9658
rect 2476 9411 2528 9420
rect 2476 9377 2485 9411
rect 2485 9377 2519 9411
rect 2519 9377 2528 9411
rect 2476 9368 2528 9377
rect 2292 9300 2344 9352
rect 19680 9343 19732 9352
rect 19680 9309 19689 9343
rect 19689 9309 19723 9343
rect 19723 9309 19732 9343
rect 19680 9300 19732 9309
rect 2292 9207 2344 9216
rect 2292 9173 2301 9207
rect 2301 9173 2335 9207
rect 2335 9173 2344 9207
rect 2292 9164 2344 9173
rect 4446 9062 4498 9114
rect 4510 9062 4562 9114
rect 4574 9062 4626 9114
rect 4638 9062 4690 9114
rect 9774 9062 9826 9114
rect 9838 9062 9890 9114
rect 9902 9062 9954 9114
rect 9966 9062 10018 9114
rect 15102 9062 15154 9114
rect 15166 9062 15218 9114
rect 15230 9062 15282 9114
rect 15294 9062 15346 9114
rect 19680 8960 19732 9012
rect 3764 8688 3816 8740
rect 7110 8518 7162 8570
rect 7174 8518 7226 8570
rect 7238 8518 7290 8570
rect 7302 8518 7354 8570
rect 12438 8518 12490 8570
rect 12502 8518 12554 8570
rect 12566 8518 12618 8570
rect 12630 8518 12682 8570
rect 17766 8518 17818 8570
rect 17830 8518 17882 8570
rect 17894 8518 17946 8570
rect 17958 8518 18010 8570
rect 3764 8459 3816 8468
rect 3764 8425 3773 8459
rect 3773 8425 3807 8459
rect 3807 8425 3816 8459
rect 3764 8416 3816 8425
rect 20140 8212 20192 8264
rect 4446 7974 4498 8026
rect 4510 7974 4562 8026
rect 4574 7974 4626 8026
rect 4638 7974 4690 8026
rect 9774 7974 9826 8026
rect 9838 7974 9890 8026
rect 9902 7974 9954 8026
rect 9966 7974 10018 8026
rect 15102 7974 15154 8026
rect 15166 7974 15218 8026
rect 15230 7974 15282 8026
rect 15294 7974 15346 8026
rect 20140 7872 20192 7924
rect 3764 7600 3816 7652
rect 7110 7430 7162 7482
rect 7174 7430 7226 7482
rect 7238 7430 7290 7482
rect 7302 7430 7354 7482
rect 12438 7430 12490 7482
rect 12502 7430 12554 7482
rect 12566 7430 12618 7482
rect 12630 7430 12682 7482
rect 17766 7430 17818 7482
rect 17830 7430 17882 7482
rect 17894 7430 17946 7482
rect 17958 7430 18010 7482
rect 3764 7167 3816 7176
rect 3764 7133 3773 7167
rect 3773 7133 3807 7167
rect 3807 7133 3816 7167
rect 3764 7124 3816 7133
rect 19680 7167 19732 7176
rect 19680 7133 19689 7167
rect 19689 7133 19723 7167
rect 19723 7133 19732 7167
rect 19680 7124 19732 7133
rect 4446 6886 4498 6938
rect 4510 6886 4562 6938
rect 4574 6886 4626 6938
rect 4638 6886 4690 6938
rect 9774 6886 9826 6938
rect 9838 6886 9890 6938
rect 9902 6886 9954 6938
rect 9966 6886 10018 6938
rect 15102 6886 15154 6938
rect 15166 6886 15218 6938
rect 15230 6886 15282 6938
rect 15294 6886 15346 6938
rect 19680 6784 19732 6836
rect 3764 6512 3816 6564
rect 7110 6342 7162 6394
rect 7174 6342 7226 6394
rect 7238 6342 7290 6394
rect 7302 6342 7354 6394
rect 12438 6342 12490 6394
rect 12502 6342 12554 6394
rect 12566 6342 12618 6394
rect 12630 6342 12682 6394
rect 17766 6342 17818 6394
rect 17830 6342 17882 6394
rect 17894 6342 17946 6394
rect 17958 6342 18010 6394
rect 3764 6283 3816 6292
rect 3764 6249 3773 6283
rect 3773 6249 3807 6283
rect 3807 6249 3816 6283
rect 3764 6240 3816 6249
rect 20140 6036 20192 6088
rect 4446 5798 4498 5850
rect 4510 5798 4562 5850
rect 4574 5798 4626 5850
rect 4638 5798 4690 5850
rect 9774 5798 9826 5850
rect 9838 5798 9890 5850
rect 9902 5798 9954 5850
rect 9966 5798 10018 5850
rect 15102 5798 15154 5850
rect 15166 5798 15218 5850
rect 15230 5798 15282 5850
rect 15294 5798 15346 5850
rect 20140 5696 20192 5748
rect 3764 5424 3816 5476
rect 7110 5254 7162 5306
rect 7174 5254 7226 5306
rect 7238 5254 7290 5306
rect 7302 5254 7354 5306
rect 12438 5254 12490 5306
rect 12502 5254 12554 5306
rect 12566 5254 12618 5306
rect 12630 5254 12682 5306
rect 17766 5254 17818 5306
rect 17830 5254 17882 5306
rect 17894 5254 17946 5306
rect 17958 5254 18010 5306
rect 3764 4991 3816 5000
rect 3764 4957 3773 4991
rect 3773 4957 3807 4991
rect 3807 4957 3816 4991
rect 3764 4948 3816 4957
rect 19680 4991 19732 5000
rect 19680 4957 19689 4991
rect 19689 4957 19723 4991
rect 19723 4957 19732 4991
rect 19680 4948 19732 4957
rect 4446 4710 4498 4762
rect 4510 4710 4562 4762
rect 4574 4710 4626 4762
rect 4638 4710 4690 4762
rect 9774 4710 9826 4762
rect 9838 4710 9890 4762
rect 9902 4710 9954 4762
rect 9966 4710 10018 4762
rect 15102 4710 15154 4762
rect 15166 4710 15218 4762
rect 15230 4710 15282 4762
rect 15294 4710 15346 4762
rect 19680 4608 19732 4660
rect 3764 4336 3816 4388
rect 7110 4166 7162 4218
rect 7174 4166 7226 4218
rect 7238 4166 7290 4218
rect 7302 4166 7354 4218
rect 12438 4166 12490 4218
rect 12502 4166 12554 4218
rect 12566 4166 12618 4218
rect 12630 4166 12682 4218
rect 17766 4166 17818 4218
rect 17830 4166 17882 4218
rect 17894 4166 17946 4218
rect 17958 4166 18010 4218
rect 3764 4107 3816 4116
rect 3764 4073 3773 4107
rect 3773 4073 3807 4107
rect 3807 4073 3816 4107
rect 3764 4064 3816 4073
rect 20232 3860 20284 3912
rect 4446 3622 4498 3674
rect 4510 3622 4562 3674
rect 4574 3622 4626 3674
rect 4638 3622 4690 3674
rect 9774 3622 9826 3674
rect 9838 3622 9890 3674
rect 9902 3622 9954 3674
rect 9966 3622 10018 3674
rect 15102 3622 15154 3674
rect 15166 3622 15218 3674
rect 15230 3622 15282 3674
rect 15294 3622 15346 3674
rect 20232 3452 20284 3504
rect 3764 3248 3816 3300
rect 7110 3078 7162 3130
rect 7174 3078 7226 3130
rect 7238 3078 7290 3130
rect 7302 3078 7354 3130
rect 12438 3078 12490 3130
rect 12502 3078 12554 3130
rect 12566 3078 12618 3130
rect 12630 3078 12682 3130
rect 17766 3078 17818 3130
rect 17830 3078 17882 3130
rect 17894 3078 17946 3130
rect 17958 3078 18010 3130
rect 3764 3019 3816 3028
rect 3764 2985 3773 3019
rect 3773 2985 3807 3019
rect 3807 2985 3816 3019
rect 3764 2976 3816 2985
rect 14988 2772 15040 2824
rect 20140 2772 20192 2824
rect 14988 2636 15040 2688
rect 4446 2534 4498 2586
rect 4510 2534 4562 2586
rect 4574 2534 4626 2586
rect 4638 2534 4690 2586
rect 9774 2534 9826 2586
rect 9838 2534 9890 2586
rect 9902 2534 9954 2586
rect 9966 2534 10018 2586
rect 15102 2534 15154 2586
rect 15166 2534 15218 2586
rect 15230 2534 15282 2586
rect 15294 2534 15346 2586
rect 20140 2432 20192 2484
rect 3764 2160 3816 2212
rect 7110 1990 7162 2042
rect 7174 1990 7226 2042
rect 7238 1990 7290 2042
rect 7302 1990 7354 2042
rect 12438 1990 12490 2042
rect 12502 1990 12554 2042
rect 12566 1990 12618 2042
rect 12630 1990 12682 2042
rect 17766 1990 17818 2042
rect 17830 1990 17882 2042
rect 17894 1990 17946 2042
rect 17958 1990 18010 2042
rect 3764 1931 3816 1940
rect 3764 1897 3773 1931
rect 3773 1897 3807 1931
rect 3807 1897 3816 1931
rect 3764 1888 3816 1897
rect 20140 1684 20192 1736
rect 4446 1446 4498 1498
rect 4510 1446 4562 1498
rect 4574 1446 4626 1498
rect 4638 1446 4690 1498
rect 9774 1446 9826 1498
rect 9838 1446 9890 1498
rect 9902 1446 9954 1498
rect 9966 1446 10018 1498
rect 15102 1446 15154 1498
rect 15166 1446 15218 1498
rect 15230 1446 15282 1498
rect 15294 1446 15346 1498
rect 20140 1344 20192 1396
rect 2936 1208 2988 1260
rect 7110 902 7162 954
rect 7174 902 7226 954
rect 7238 902 7290 954
rect 7302 902 7354 954
rect 12438 902 12490 954
rect 12502 902 12554 954
rect 12566 902 12618 954
rect 12630 902 12682 954
rect 17766 902 17818 954
rect 17830 902 17882 954
rect 17894 902 17946 954
rect 17958 902 18010 954
<< metal2 >>
rect 1922 22376 1978 22385
rect 1922 22311 1978 22320
rect 1936 22074 1964 22311
rect 4420 22172 4716 22192
rect 4476 22170 4500 22172
rect 4556 22170 4580 22172
rect 4636 22170 4660 22172
rect 4498 22118 4500 22170
rect 4562 22118 4574 22170
rect 4636 22118 4638 22170
rect 4476 22116 4500 22118
rect 4556 22116 4580 22118
rect 4636 22116 4660 22118
rect 4420 22096 4716 22116
rect 9748 22172 10044 22192
rect 9804 22170 9828 22172
rect 9884 22170 9908 22172
rect 9964 22170 9988 22172
rect 9826 22118 9828 22170
rect 9890 22118 9902 22170
rect 9964 22118 9966 22170
rect 9804 22116 9828 22118
rect 9884 22116 9908 22118
rect 9964 22116 9988 22118
rect 9748 22096 10044 22116
rect 15076 22172 15372 22192
rect 15132 22170 15156 22172
rect 15212 22170 15236 22172
rect 15292 22170 15316 22172
rect 15154 22118 15156 22170
rect 15218 22118 15230 22170
rect 15292 22118 15294 22170
rect 15132 22116 15156 22118
rect 15212 22116 15236 22118
rect 15292 22116 15316 22118
rect 15076 22096 15372 22116
rect 1924 22068 1976 22074
rect 1924 22010 1976 22016
rect 2292 22000 2344 22006
rect 2292 21942 2344 21948
rect 2304 21530 2332 21942
rect 2476 21864 2528 21870
rect 2474 21832 2476 21841
rect 2528 21832 2530 21841
rect 2474 21767 2530 21776
rect 7084 21628 7380 21648
rect 7140 21626 7164 21628
rect 7220 21626 7244 21628
rect 7300 21626 7324 21628
rect 7162 21574 7164 21626
rect 7226 21574 7238 21626
rect 7300 21574 7302 21626
rect 7140 21572 7164 21574
rect 7220 21572 7244 21574
rect 7300 21572 7324 21574
rect 7084 21552 7380 21572
rect 12412 21628 12708 21648
rect 12468 21626 12492 21628
rect 12548 21626 12572 21628
rect 12628 21626 12652 21628
rect 12490 21574 12492 21626
rect 12554 21574 12566 21626
rect 12628 21574 12630 21626
rect 12468 21572 12492 21574
rect 12548 21572 12572 21574
rect 12628 21572 12652 21574
rect 12412 21552 12708 21572
rect 17740 21628 18036 21648
rect 17796 21626 17820 21628
rect 17876 21626 17900 21628
rect 17956 21626 17980 21628
rect 17818 21574 17820 21626
rect 17882 21574 17894 21626
rect 17956 21574 17958 21626
rect 17796 21572 17820 21574
rect 17876 21572 17900 21574
rect 17956 21572 17980 21574
rect 17740 21552 18036 21572
rect 2292 21524 2344 21530
rect 2292 21466 2344 21472
rect 2476 21388 2528 21394
rect 2476 21330 2528 21336
rect 2488 21297 2516 21330
rect 3856 21320 3908 21326
rect 2474 21288 2530 21297
rect 2292 21252 2344 21258
rect 3856 21262 3908 21268
rect 2474 21223 2530 21232
rect 2292 21194 2344 21200
rect 2304 20850 2332 21194
rect 3868 20986 3896 21262
rect 4420 21084 4716 21104
rect 4476 21082 4500 21084
rect 4556 21082 4580 21084
rect 4636 21082 4660 21084
rect 4498 21030 4500 21082
rect 4562 21030 4574 21082
rect 4636 21030 4638 21082
rect 4476 21028 4500 21030
rect 4556 21028 4580 21030
rect 4636 21028 4660 21030
rect 4420 21008 4716 21028
rect 9748 21084 10044 21104
rect 9804 21082 9828 21084
rect 9884 21082 9908 21084
rect 9964 21082 9988 21084
rect 9826 21030 9828 21082
rect 9890 21030 9902 21082
rect 9964 21030 9966 21082
rect 9804 21028 9828 21030
rect 9884 21028 9908 21030
rect 9964 21028 9988 21030
rect 9748 21008 10044 21028
rect 15076 21084 15372 21104
rect 15132 21082 15156 21084
rect 15212 21082 15236 21084
rect 15292 21082 15316 21084
rect 15154 21030 15156 21082
rect 15218 21030 15230 21082
rect 15292 21030 15294 21082
rect 15132 21028 15156 21030
rect 15212 21028 15236 21030
rect 15292 21028 15316 21030
rect 15076 21008 15372 21028
rect 3856 20980 3908 20986
rect 3856 20922 3908 20928
rect 2292 20844 2344 20850
rect 2292 20786 2344 20792
rect 2304 20442 2332 20786
rect 7084 20540 7380 20560
rect 7140 20538 7164 20540
rect 7220 20538 7244 20540
rect 7300 20538 7324 20540
rect 7162 20486 7164 20538
rect 7226 20486 7238 20538
rect 7300 20486 7302 20538
rect 7140 20484 7164 20486
rect 7220 20484 7244 20486
rect 7300 20484 7324 20486
rect 7084 20464 7380 20484
rect 12412 20540 12708 20560
rect 12468 20538 12492 20540
rect 12548 20538 12572 20540
rect 12628 20538 12652 20540
rect 12490 20486 12492 20538
rect 12554 20486 12566 20538
rect 12628 20486 12630 20538
rect 12468 20484 12492 20486
rect 12548 20484 12572 20486
rect 12628 20484 12652 20486
rect 12412 20464 12708 20484
rect 17740 20540 18036 20560
rect 17796 20538 17820 20540
rect 17876 20538 17900 20540
rect 17956 20538 17980 20540
rect 17818 20486 17820 20538
rect 17882 20486 17894 20538
rect 17956 20486 17958 20538
rect 17796 20484 17820 20486
rect 17876 20484 17900 20486
rect 17956 20484 17980 20486
rect 17740 20464 18036 20484
rect 2292 20436 2344 20442
rect 2292 20378 2344 20384
rect 2476 20300 2528 20306
rect 2476 20242 2528 20248
rect 2488 20209 2516 20242
rect 4224 20232 4276 20238
rect 2474 20200 2530 20209
rect 4224 20174 4276 20180
rect 2474 20135 2530 20144
rect 2292 20096 2344 20102
rect 2292 20038 2344 20044
rect 2304 19762 2332 20038
rect 4236 19898 4264 20174
rect 4420 19996 4716 20016
rect 4476 19994 4500 19996
rect 4556 19994 4580 19996
rect 4636 19994 4660 19996
rect 4498 19942 4500 19994
rect 4562 19942 4574 19994
rect 4636 19942 4638 19994
rect 4476 19940 4500 19942
rect 4556 19940 4580 19942
rect 4636 19940 4660 19942
rect 4420 19920 4716 19940
rect 9748 19996 10044 20016
rect 9804 19994 9828 19996
rect 9884 19994 9908 19996
rect 9964 19994 9988 19996
rect 9826 19942 9828 19994
rect 9890 19942 9902 19994
rect 9964 19942 9966 19994
rect 9804 19940 9828 19942
rect 9884 19940 9908 19942
rect 9964 19940 9988 19942
rect 9748 19920 10044 19940
rect 15076 19996 15372 20016
rect 15132 19994 15156 19996
rect 15212 19994 15236 19996
rect 15292 19994 15316 19996
rect 15154 19942 15156 19994
rect 15218 19942 15230 19994
rect 15292 19942 15294 19994
rect 15132 19940 15156 19942
rect 15212 19940 15236 19942
rect 15292 19940 15316 19942
rect 15076 19920 15372 19940
rect 4224 19892 4276 19898
rect 4224 19834 4276 19840
rect 2292 19756 2344 19762
rect 2292 19698 2344 19704
rect 2304 19354 2332 19698
rect 7084 19452 7380 19472
rect 7140 19450 7164 19452
rect 7220 19450 7244 19452
rect 7300 19450 7324 19452
rect 7162 19398 7164 19450
rect 7226 19398 7238 19450
rect 7300 19398 7302 19450
rect 7140 19396 7164 19398
rect 7220 19396 7244 19398
rect 7300 19396 7324 19398
rect 7084 19376 7380 19396
rect 12412 19452 12708 19472
rect 12468 19450 12492 19452
rect 12548 19450 12572 19452
rect 12628 19450 12652 19452
rect 12490 19398 12492 19450
rect 12554 19398 12566 19450
rect 12628 19398 12630 19450
rect 12468 19396 12492 19398
rect 12548 19396 12572 19398
rect 12628 19396 12652 19398
rect 12412 19376 12708 19396
rect 17740 19452 18036 19472
rect 17796 19450 17820 19452
rect 17876 19450 17900 19452
rect 17956 19450 17980 19452
rect 17818 19398 17820 19450
rect 17882 19398 17894 19450
rect 17956 19398 17958 19450
rect 17796 19396 17820 19398
rect 17876 19396 17900 19398
rect 17956 19396 17980 19398
rect 17740 19376 18036 19396
rect 2292 19348 2344 19354
rect 2292 19290 2344 19296
rect 2476 19212 2528 19218
rect 2476 19154 2528 19160
rect 2488 19121 2516 19154
rect 6984 19144 7036 19150
rect 2474 19112 2530 19121
rect 6984 19086 7036 19092
rect 2474 19047 2530 19056
rect 2292 19008 2344 19014
rect 2292 18950 2344 18956
rect 2304 18674 2332 18950
rect 4420 18908 4716 18928
rect 4476 18906 4500 18908
rect 4556 18906 4580 18908
rect 4636 18906 4660 18908
rect 4498 18854 4500 18906
rect 4562 18854 4574 18906
rect 4636 18854 4638 18906
rect 4476 18852 4500 18854
rect 4556 18852 4580 18854
rect 4636 18852 4660 18854
rect 4420 18832 4716 18852
rect 6996 18810 7024 19086
rect 9748 18908 10044 18928
rect 9804 18906 9828 18908
rect 9884 18906 9908 18908
rect 9964 18906 9988 18908
rect 9826 18854 9828 18906
rect 9890 18854 9902 18906
rect 9964 18854 9966 18906
rect 9804 18852 9828 18854
rect 9884 18852 9908 18854
rect 9964 18852 9988 18854
rect 9748 18832 10044 18852
rect 15076 18908 15372 18928
rect 15132 18906 15156 18908
rect 15212 18906 15236 18908
rect 15292 18906 15316 18908
rect 15154 18854 15156 18906
rect 15218 18854 15230 18906
rect 15292 18854 15294 18906
rect 15132 18852 15156 18854
rect 15212 18852 15236 18854
rect 15292 18852 15316 18854
rect 15076 18832 15372 18852
rect 6984 18804 7036 18810
rect 6984 18746 7036 18752
rect 2292 18668 2344 18674
rect 2292 18610 2344 18616
rect 2304 18266 2332 18610
rect 7084 18364 7380 18384
rect 7140 18362 7164 18364
rect 7220 18362 7244 18364
rect 7300 18362 7324 18364
rect 7162 18310 7164 18362
rect 7226 18310 7238 18362
rect 7300 18310 7302 18362
rect 7140 18308 7164 18310
rect 7220 18308 7244 18310
rect 7300 18308 7324 18310
rect 7084 18288 7380 18308
rect 12412 18364 12708 18384
rect 12468 18362 12492 18364
rect 12548 18362 12572 18364
rect 12628 18362 12652 18364
rect 12490 18310 12492 18362
rect 12554 18310 12566 18362
rect 12628 18310 12630 18362
rect 12468 18308 12492 18310
rect 12548 18308 12572 18310
rect 12628 18308 12652 18310
rect 12412 18288 12708 18308
rect 17740 18364 18036 18384
rect 17796 18362 17820 18364
rect 17876 18362 17900 18364
rect 17956 18362 17980 18364
rect 17818 18310 17820 18362
rect 17882 18310 17894 18362
rect 17956 18310 17958 18362
rect 17796 18308 17820 18310
rect 17876 18308 17900 18310
rect 17956 18308 17980 18310
rect 17740 18288 18036 18308
rect 2292 18260 2344 18266
rect 2292 18202 2344 18208
rect 2476 18124 2528 18130
rect 2476 18066 2528 18072
rect 2488 18033 2516 18066
rect 10848 18056 10900 18062
rect 2474 18024 2530 18033
rect 10848 17998 10900 18004
rect 2474 17959 2530 17968
rect 2292 17920 2344 17926
rect 2292 17862 2344 17868
rect 2304 17586 2332 17862
rect 4420 17820 4716 17840
rect 4476 17818 4500 17820
rect 4556 17818 4580 17820
rect 4636 17818 4660 17820
rect 4498 17766 4500 17818
rect 4562 17766 4574 17818
rect 4636 17766 4638 17818
rect 4476 17764 4500 17766
rect 4556 17764 4580 17766
rect 4636 17764 4660 17766
rect 4420 17744 4716 17764
rect 9748 17820 10044 17840
rect 9804 17818 9828 17820
rect 9884 17818 9908 17820
rect 9964 17818 9988 17820
rect 9826 17766 9828 17818
rect 9890 17766 9902 17818
rect 9964 17766 9966 17818
rect 9804 17764 9828 17766
rect 9884 17764 9908 17766
rect 9964 17764 9988 17766
rect 9748 17744 10044 17764
rect 10860 17722 10888 17998
rect 15076 17820 15372 17840
rect 15132 17818 15156 17820
rect 15212 17818 15236 17820
rect 15292 17818 15316 17820
rect 15154 17766 15156 17818
rect 15218 17766 15230 17818
rect 15292 17766 15294 17818
rect 15132 17764 15156 17766
rect 15212 17764 15236 17766
rect 15292 17764 15316 17766
rect 15076 17744 15372 17764
rect 10848 17716 10900 17722
rect 10848 17658 10900 17664
rect 2292 17580 2344 17586
rect 2292 17522 2344 17528
rect 2304 17178 2332 17522
rect 7084 17276 7380 17296
rect 7140 17274 7164 17276
rect 7220 17274 7244 17276
rect 7300 17274 7324 17276
rect 7162 17222 7164 17274
rect 7226 17222 7238 17274
rect 7300 17222 7302 17274
rect 7140 17220 7164 17222
rect 7220 17220 7244 17222
rect 7300 17220 7324 17222
rect 7084 17200 7380 17220
rect 12412 17276 12708 17296
rect 12468 17274 12492 17276
rect 12548 17274 12572 17276
rect 12628 17274 12652 17276
rect 12490 17222 12492 17274
rect 12554 17222 12566 17274
rect 12628 17222 12630 17274
rect 12468 17220 12492 17222
rect 12548 17220 12572 17222
rect 12628 17220 12652 17222
rect 12412 17200 12708 17220
rect 17740 17276 18036 17296
rect 17796 17274 17820 17276
rect 17876 17274 17900 17276
rect 17956 17274 17980 17276
rect 17818 17222 17820 17274
rect 17882 17222 17894 17274
rect 17956 17222 17958 17274
rect 17796 17220 17820 17222
rect 17876 17220 17900 17222
rect 17956 17220 17980 17222
rect 17740 17200 18036 17220
rect 2292 17172 2344 17178
rect 2292 17114 2344 17120
rect 2476 17036 2528 17042
rect 2476 16978 2528 16984
rect 2292 16832 2344 16838
rect 2292 16774 2344 16780
rect 2304 16498 2332 16774
rect 2488 16673 2516 16978
rect 20140 16968 20192 16974
rect 20140 16910 20192 16916
rect 4420 16732 4716 16752
rect 4476 16730 4500 16732
rect 4556 16730 4580 16732
rect 4636 16730 4660 16732
rect 4498 16678 4500 16730
rect 4562 16678 4574 16730
rect 4636 16678 4638 16730
rect 4476 16676 4500 16678
rect 4556 16676 4580 16678
rect 4636 16676 4660 16678
rect 2474 16664 2530 16673
rect 4420 16656 4716 16676
rect 9748 16732 10044 16752
rect 9804 16730 9828 16732
rect 9884 16730 9908 16732
rect 9964 16730 9988 16732
rect 9826 16678 9828 16730
rect 9890 16678 9902 16730
rect 9964 16678 9966 16730
rect 9804 16676 9828 16678
rect 9884 16676 9908 16678
rect 9964 16676 9988 16678
rect 9748 16656 10044 16676
rect 15076 16732 15372 16752
rect 15132 16730 15156 16732
rect 15212 16730 15236 16732
rect 15292 16730 15316 16732
rect 15154 16678 15156 16730
rect 15218 16678 15230 16730
rect 15292 16678 15294 16730
rect 15132 16676 15156 16678
rect 15212 16676 15236 16678
rect 15292 16676 15316 16678
rect 15076 16656 15372 16676
rect 20152 16634 20180 16910
rect 2474 16599 2530 16608
rect 20140 16628 20192 16634
rect 20140 16570 20192 16576
rect 2292 16492 2344 16498
rect 2292 16434 2344 16440
rect 2568 16492 2620 16498
rect 2568 16434 2620 16440
rect 2580 16022 2608 16434
rect 7084 16188 7380 16208
rect 7140 16186 7164 16188
rect 7220 16186 7244 16188
rect 7300 16186 7324 16188
rect 7162 16134 7164 16186
rect 7226 16134 7238 16186
rect 7300 16134 7302 16186
rect 7140 16132 7164 16134
rect 7220 16132 7244 16134
rect 7300 16132 7324 16134
rect 7084 16112 7380 16132
rect 12412 16188 12708 16208
rect 12468 16186 12492 16188
rect 12548 16186 12572 16188
rect 12628 16186 12652 16188
rect 12490 16134 12492 16186
rect 12554 16134 12566 16186
rect 12628 16134 12630 16186
rect 12468 16132 12492 16134
rect 12548 16132 12572 16134
rect 12628 16132 12652 16134
rect 12412 16112 12708 16132
rect 17740 16188 18036 16208
rect 17796 16186 17820 16188
rect 17876 16186 17900 16188
rect 17956 16186 17980 16188
rect 17818 16134 17820 16186
rect 17882 16134 17894 16186
rect 17956 16134 17958 16186
rect 17796 16132 17820 16134
rect 17876 16132 17900 16134
rect 17956 16132 17980 16134
rect 17740 16112 18036 16132
rect 2568 16016 2620 16022
rect 2568 15958 2620 15964
rect 2476 15948 2528 15954
rect 2476 15890 2528 15896
rect 2488 15857 2516 15890
rect 19680 15880 19732 15886
rect 2474 15848 2530 15857
rect 19680 15822 19732 15828
rect 2474 15783 2530 15792
rect 2292 15744 2344 15750
rect 2292 15686 2344 15692
rect 2304 14322 2332 15686
rect 4420 15644 4716 15664
rect 4476 15642 4500 15644
rect 4556 15642 4580 15644
rect 4636 15642 4660 15644
rect 4498 15590 4500 15642
rect 4562 15590 4574 15642
rect 4636 15590 4638 15642
rect 4476 15588 4500 15590
rect 4556 15588 4580 15590
rect 4636 15588 4660 15590
rect 4420 15568 4716 15588
rect 9748 15644 10044 15664
rect 9804 15642 9828 15644
rect 9884 15642 9908 15644
rect 9964 15642 9988 15644
rect 9826 15590 9828 15642
rect 9890 15590 9902 15642
rect 9964 15590 9966 15642
rect 9804 15588 9828 15590
rect 9884 15588 9908 15590
rect 9964 15588 9988 15590
rect 9748 15568 10044 15588
rect 15076 15644 15372 15664
rect 15132 15642 15156 15644
rect 15212 15642 15236 15644
rect 15292 15642 15316 15644
rect 15154 15590 15156 15642
rect 15218 15590 15230 15642
rect 15292 15590 15294 15642
rect 15132 15588 15156 15590
rect 15212 15588 15236 15590
rect 15292 15588 15316 15590
rect 15076 15568 15372 15588
rect 19692 15546 19720 15822
rect 19680 15540 19732 15546
rect 19680 15482 19732 15488
rect 3764 15268 3816 15274
rect 3764 15210 3816 15216
rect 3776 15002 3804 15210
rect 7084 15100 7380 15120
rect 7140 15098 7164 15100
rect 7220 15098 7244 15100
rect 7300 15098 7324 15100
rect 7162 15046 7164 15098
rect 7226 15046 7238 15098
rect 7300 15046 7302 15098
rect 7140 15044 7164 15046
rect 7220 15044 7244 15046
rect 7300 15044 7324 15046
rect 7084 15024 7380 15044
rect 12412 15100 12708 15120
rect 12468 15098 12492 15100
rect 12548 15098 12572 15100
rect 12628 15098 12652 15100
rect 12490 15046 12492 15098
rect 12554 15046 12566 15098
rect 12628 15046 12630 15098
rect 12468 15044 12492 15046
rect 12548 15044 12572 15046
rect 12628 15044 12652 15046
rect 12412 15024 12708 15044
rect 17740 15100 18036 15120
rect 17796 15098 17820 15100
rect 17876 15098 17900 15100
rect 17956 15098 17980 15100
rect 17818 15046 17820 15098
rect 17882 15046 17894 15098
rect 17956 15046 17958 15098
rect 17796 15044 17820 15046
rect 17876 15044 17900 15046
rect 17956 15044 17980 15046
rect 17740 15024 18036 15044
rect 3764 14996 3816 15002
rect 3764 14938 3816 14944
rect 20140 14792 20192 14798
rect 20140 14734 20192 14740
rect 4420 14556 4716 14576
rect 4476 14554 4500 14556
rect 4556 14554 4580 14556
rect 4636 14554 4660 14556
rect 4498 14502 4500 14554
rect 4562 14502 4574 14554
rect 4636 14502 4638 14554
rect 4476 14500 4500 14502
rect 4556 14500 4580 14502
rect 4636 14500 4660 14502
rect 4420 14480 4716 14500
rect 9748 14556 10044 14576
rect 9804 14554 9828 14556
rect 9884 14554 9908 14556
rect 9964 14554 9988 14556
rect 9826 14502 9828 14554
rect 9890 14502 9902 14554
rect 9964 14502 9966 14554
rect 9804 14500 9828 14502
rect 9884 14500 9908 14502
rect 9964 14500 9988 14502
rect 9748 14480 10044 14500
rect 15076 14556 15372 14576
rect 15132 14554 15156 14556
rect 15212 14554 15236 14556
rect 15292 14554 15316 14556
rect 15154 14502 15156 14554
rect 15218 14502 15230 14554
rect 15292 14502 15294 14554
rect 15132 14500 15156 14502
rect 15212 14500 15236 14502
rect 15292 14500 15316 14502
rect 15076 14480 15372 14500
rect 20152 14458 20180 14734
rect 20140 14452 20192 14458
rect 20140 14394 20192 14400
rect 2292 14316 2344 14322
rect 2292 14258 2344 14264
rect 2304 13846 2332 14258
rect 7084 14012 7380 14032
rect 7140 14010 7164 14012
rect 7220 14010 7244 14012
rect 7300 14010 7324 14012
rect 7162 13958 7164 14010
rect 7226 13958 7238 14010
rect 7300 13958 7302 14010
rect 7140 13956 7164 13958
rect 7220 13956 7244 13958
rect 7300 13956 7324 13958
rect 7084 13936 7380 13956
rect 12412 14012 12708 14032
rect 12468 14010 12492 14012
rect 12548 14010 12572 14012
rect 12628 14010 12652 14012
rect 12490 13958 12492 14010
rect 12554 13958 12566 14010
rect 12628 13958 12630 14010
rect 12468 13956 12492 13958
rect 12548 13956 12572 13958
rect 12628 13956 12652 13958
rect 12412 13936 12708 13956
rect 17740 14012 18036 14032
rect 17796 14010 17820 14012
rect 17876 14010 17900 14012
rect 17956 14010 17980 14012
rect 17818 13958 17820 14010
rect 17882 13958 17894 14010
rect 17956 13958 17958 14010
rect 17796 13956 17820 13958
rect 17876 13956 17900 13958
rect 17956 13956 17980 13958
rect 17740 13936 18036 13956
rect 2292 13840 2344 13846
rect 2292 13782 2344 13788
rect 2476 13772 2528 13778
rect 2476 13714 2528 13720
rect 2488 13681 2516 13714
rect 19680 13704 19732 13710
rect 2474 13672 2530 13681
rect 19680 13646 19732 13652
rect 2474 13607 2530 13616
rect 2292 13568 2344 13574
rect 2292 13510 2344 13516
rect 2304 9970 2332 13510
rect 4420 13468 4716 13488
rect 4476 13466 4500 13468
rect 4556 13466 4580 13468
rect 4636 13466 4660 13468
rect 4498 13414 4500 13466
rect 4562 13414 4574 13466
rect 4636 13414 4638 13466
rect 4476 13412 4500 13414
rect 4556 13412 4580 13414
rect 4636 13412 4660 13414
rect 4420 13392 4716 13412
rect 9748 13468 10044 13488
rect 9804 13466 9828 13468
rect 9884 13466 9908 13468
rect 9964 13466 9988 13468
rect 9826 13414 9828 13466
rect 9890 13414 9902 13466
rect 9964 13414 9966 13466
rect 9804 13412 9828 13414
rect 9884 13412 9908 13414
rect 9964 13412 9988 13414
rect 9748 13392 10044 13412
rect 15076 13468 15372 13488
rect 15132 13466 15156 13468
rect 15212 13466 15236 13468
rect 15292 13466 15316 13468
rect 15154 13414 15156 13466
rect 15218 13414 15230 13466
rect 15292 13414 15294 13466
rect 15132 13412 15156 13414
rect 15212 13412 15236 13414
rect 15292 13412 15316 13414
rect 15076 13392 15372 13412
rect 19692 13370 19720 13646
rect 19680 13364 19732 13370
rect 19680 13306 19732 13312
rect 3764 13092 3816 13098
rect 3764 13034 3816 13040
rect 3776 12826 3804 13034
rect 7084 12924 7380 12944
rect 7140 12922 7164 12924
rect 7220 12922 7244 12924
rect 7300 12922 7324 12924
rect 7162 12870 7164 12922
rect 7226 12870 7238 12922
rect 7300 12870 7302 12922
rect 7140 12868 7164 12870
rect 7220 12868 7244 12870
rect 7300 12868 7324 12870
rect 7084 12848 7380 12868
rect 12412 12924 12708 12944
rect 12468 12922 12492 12924
rect 12548 12922 12572 12924
rect 12628 12922 12652 12924
rect 12490 12870 12492 12922
rect 12554 12870 12566 12922
rect 12628 12870 12630 12922
rect 12468 12868 12492 12870
rect 12548 12868 12572 12870
rect 12628 12868 12652 12870
rect 12412 12848 12708 12868
rect 17740 12924 18036 12944
rect 17796 12922 17820 12924
rect 17876 12922 17900 12924
rect 17956 12922 17980 12924
rect 17818 12870 17820 12922
rect 17882 12870 17894 12922
rect 17956 12870 17958 12922
rect 17796 12868 17820 12870
rect 17876 12868 17900 12870
rect 17956 12868 17980 12870
rect 17740 12848 18036 12868
rect 3764 12820 3816 12826
rect 3764 12762 3816 12768
rect 20140 12616 20192 12622
rect 20140 12558 20192 12564
rect 4420 12380 4716 12400
rect 4476 12378 4500 12380
rect 4556 12378 4580 12380
rect 4636 12378 4660 12380
rect 4498 12326 4500 12378
rect 4562 12326 4574 12378
rect 4636 12326 4638 12378
rect 4476 12324 4500 12326
rect 4556 12324 4580 12326
rect 4636 12324 4660 12326
rect 4420 12304 4716 12324
rect 9748 12380 10044 12400
rect 9804 12378 9828 12380
rect 9884 12378 9908 12380
rect 9964 12378 9988 12380
rect 9826 12326 9828 12378
rect 9890 12326 9902 12378
rect 9964 12326 9966 12378
rect 9804 12324 9828 12326
rect 9884 12324 9908 12326
rect 9964 12324 9988 12326
rect 9748 12304 10044 12324
rect 15076 12380 15372 12400
rect 15132 12378 15156 12380
rect 15212 12378 15236 12380
rect 15292 12378 15316 12380
rect 15154 12326 15156 12378
rect 15218 12326 15230 12378
rect 15292 12326 15294 12378
rect 15132 12324 15156 12326
rect 15212 12324 15236 12326
rect 15292 12324 15316 12326
rect 15076 12304 15372 12324
rect 20152 12282 20180 12558
rect 20140 12276 20192 12282
rect 20140 12218 20192 12224
rect 3764 12004 3816 12010
rect 3764 11946 3816 11952
rect 3776 11602 3804 11946
rect 7084 11836 7380 11856
rect 7140 11834 7164 11836
rect 7220 11834 7244 11836
rect 7300 11834 7324 11836
rect 7162 11782 7164 11834
rect 7226 11782 7238 11834
rect 7300 11782 7302 11834
rect 7140 11780 7164 11782
rect 7220 11780 7244 11782
rect 7300 11780 7324 11782
rect 7084 11760 7380 11780
rect 12412 11836 12708 11856
rect 12468 11834 12492 11836
rect 12548 11834 12572 11836
rect 12628 11834 12652 11836
rect 12490 11782 12492 11834
rect 12554 11782 12566 11834
rect 12628 11782 12630 11834
rect 12468 11780 12492 11782
rect 12548 11780 12572 11782
rect 12628 11780 12652 11782
rect 12412 11760 12708 11780
rect 17740 11836 18036 11856
rect 17796 11834 17820 11836
rect 17876 11834 17900 11836
rect 17956 11834 17980 11836
rect 17818 11782 17820 11834
rect 17882 11782 17894 11834
rect 17956 11782 17958 11834
rect 17796 11780 17820 11782
rect 17876 11780 17900 11782
rect 17956 11780 17980 11782
rect 17740 11760 18036 11780
rect 3764 11596 3816 11602
rect 3764 11538 3816 11544
rect 19680 11528 19732 11534
rect 19680 11470 19732 11476
rect 4420 11292 4716 11312
rect 4476 11290 4500 11292
rect 4556 11290 4580 11292
rect 4636 11290 4660 11292
rect 4498 11238 4500 11290
rect 4562 11238 4574 11290
rect 4636 11238 4638 11290
rect 4476 11236 4500 11238
rect 4556 11236 4580 11238
rect 4636 11236 4660 11238
rect 4420 11216 4716 11236
rect 9748 11292 10044 11312
rect 9804 11290 9828 11292
rect 9884 11290 9908 11292
rect 9964 11290 9988 11292
rect 9826 11238 9828 11290
rect 9890 11238 9902 11290
rect 9964 11238 9966 11290
rect 9804 11236 9828 11238
rect 9884 11236 9908 11238
rect 9964 11236 9988 11238
rect 9748 11216 10044 11236
rect 15076 11292 15372 11312
rect 15132 11290 15156 11292
rect 15212 11290 15236 11292
rect 15292 11290 15316 11292
rect 15154 11238 15156 11290
rect 15218 11238 15230 11290
rect 15292 11238 15294 11290
rect 15132 11236 15156 11238
rect 15212 11236 15236 11238
rect 15292 11236 15316 11238
rect 15076 11216 15372 11236
rect 19692 11194 19720 11470
rect 19680 11188 19732 11194
rect 19680 11130 19732 11136
rect 3764 10916 3816 10922
rect 3764 10858 3816 10864
rect 3776 10650 3804 10858
rect 7084 10748 7380 10768
rect 7140 10746 7164 10748
rect 7220 10746 7244 10748
rect 7300 10746 7324 10748
rect 7162 10694 7164 10746
rect 7226 10694 7238 10746
rect 7300 10694 7302 10746
rect 7140 10692 7164 10694
rect 7220 10692 7244 10694
rect 7300 10692 7324 10694
rect 7084 10672 7380 10692
rect 12412 10748 12708 10768
rect 12468 10746 12492 10748
rect 12548 10746 12572 10748
rect 12628 10746 12652 10748
rect 12490 10694 12492 10746
rect 12554 10694 12566 10746
rect 12628 10694 12630 10746
rect 12468 10692 12492 10694
rect 12548 10692 12572 10694
rect 12628 10692 12652 10694
rect 12412 10672 12708 10692
rect 17740 10748 18036 10768
rect 17796 10746 17820 10748
rect 17876 10746 17900 10748
rect 17956 10746 17980 10748
rect 17818 10694 17820 10746
rect 17882 10694 17894 10746
rect 17956 10694 17958 10746
rect 17796 10692 17820 10694
rect 17876 10692 17900 10694
rect 17956 10692 17980 10694
rect 17740 10672 18036 10692
rect 3764 10644 3816 10650
rect 3764 10586 3816 10592
rect 20140 10440 20192 10446
rect 20140 10382 20192 10388
rect 4420 10204 4716 10224
rect 4476 10202 4500 10204
rect 4556 10202 4580 10204
rect 4636 10202 4660 10204
rect 4498 10150 4500 10202
rect 4562 10150 4574 10202
rect 4636 10150 4638 10202
rect 4476 10148 4500 10150
rect 4556 10148 4580 10150
rect 4636 10148 4660 10150
rect 4420 10128 4716 10148
rect 9748 10204 10044 10224
rect 9804 10202 9828 10204
rect 9884 10202 9908 10204
rect 9964 10202 9988 10204
rect 9826 10150 9828 10202
rect 9890 10150 9902 10202
rect 9964 10150 9966 10202
rect 9804 10148 9828 10150
rect 9884 10148 9908 10150
rect 9964 10148 9988 10150
rect 9748 10128 10044 10148
rect 15076 10204 15372 10224
rect 15132 10202 15156 10204
rect 15212 10202 15236 10204
rect 15292 10202 15316 10204
rect 15154 10150 15156 10202
rect 15218 10150 15230 10202
rect 15292 10150 15294 10202
rect 15132 10148 15156 10150
rect 15212 10148 15236 10150
rect 15292 10148 15316 10150
rect 15076 10128 15372 10148
rect 20152 10106 20180 10382
rect 20140 10100 20192 10106
rect 20140 10042 20192 10048
rect 2292 9964 2344 9970
rect 2292 9906 2344 9912
rect 2304 9358 2332 9906
rect 7084 9660 7380 9680
rect 7140 9658 7164 9660
rect 7220 9658 7244 9660
rect 7300 9658 7324 9660
rect 7162 9606 7164 9658
rect 7226 9606 7238 9658
rect 7300 9606 7302 9658
rect 7140 9604 7164 9606
rect 7220 9604 7244 9606
rect 7300 9604 7324 9606
rect 7084 9584 7380 9604
rect 12412 9660 12708 9680
rect 12468 9658 12492 9660
rect 12548 9658 12572 9660
rect 12628 9658 12652 9660
rect 12490 9606 12492 9658
rect 12554 9606 12566 9658
rect 12628 9606 12630 9658
rect 12468 9604 12492 9606
rect 12548 9604 12572 9606
rect 12628 9604 12652 9606
rect 12412 9584 12708 9604
rect 17740 9660 18036 9680
rect 17796 9658 17820 9660
rect 17876 9658 17900 9660
rect 17956 9658 17980 9660
rect 17818 9606 17820 9658
rect 17882 9606 17894 9658
rect 17956 9606 17958 9658
rect 17796 9604 17820 9606
rect 17876 9604 17900 9606
rect 17956 9604 17980 9606
rect 17740 9584 18036 9604
rect 2476 9420 2528 9426
rect 2476 9362 2528 9368
rect 2292 9352 2344 9358
rect 2292 9294 2344 9300
rect 2292 9216 2344 9222
rect 2292 9158 2344 9164
rect 2304 1169 2332 9158
rect 2488 8785 2516 9362
rect 19680 9352 19732 9358
rect 19680 9294 19732 9300
rect 4420 9116 4716 9136
rect 4476 9114 4500 9116
rect 4556 9114 4580 9116
rect 4636 9114 4660 9116
rect 4498 9062 4500 9114
rect 4562 9062 4574 9114
rect 4636 9062 4638 9114
rect 4476 9060 4500 9062
rect 4556 9060 4580 9062
rect 4636 9060 4660 9062
rect 4420 9040 4716 9060
rect 9748 9116 10044 9136
rect 9804 9114 9828 9116
rect 9884 9114 9908 9116
rect 9964 9114 9988 9116
rect 9826 9062 9828 9114
rect 9890 9062 9902 9114
rect 9964 9062 9966 9114
rect 9804 9060 9828 9062
rect 9884 9060 9908 9062
rect 9964 9060 9988 9062
rect 9748 9040 10044 9060
rect 15076 9116 15372 9136
rect 15132 9114 15156 9116
rect 15212 9114 15236 9116
rect 15292 9114 15316 9116
rect 15154 9062 15156 9114
rect 15218 9062 15230 9114
rect 15292 9062 15294 9114
rect 15132 9060 15156 9062
rect 15212 9060 15236 9062
rect 15292 9060 15316 9062
rect 15076 9040 15372 9060
rect 19692 9018 19720 9294
rect 19680 9012 19732 9018
rect 19680 8954 19732 8960
rect 2474 8776 2530 8785
rect 2474 8711 2530 8720
rect 3764 8740 3816 8746
rect 3764 8682 3816 8688
rect 3776 8474 3804 8682
rect 7084 8572 7380 8592
rect 7140 8570 7164 8572
rect 7220 8570 7244 8572
rect 7300 8570 7324 8572
rect 7162 8518 7164 8570
rect 7226 8518 7238 8570
rect 7300 8518 7302 8570
rect 7140 8516 7164 8518
rect 7220 8516 7244 8518
rect 7300 8516 7324 8518
rect 7084 8496 7380 8516
rect 12412 8572 12708 8592
rect 12468 8570 12492 8572
rect 12548 8570 12572 8572
rect 12628 8570 12652 8572
rect 12490 8518 12492 8570
rect 12554 8518 12566 8570
rect 12628 8518 12630 8570
rect 12468 8516 12492 8518
rect 12548 8516 12572 8518
rect 12628 8516 12652 8518
rect 12412 8496 12708 8516
rect 17740 8572 18036 8592
rect 17796 8570 17820 8572
rect 17876 8570 17900 8572
rect 17956 8570 17980 8572
rect 17818 8518 17820 8570
rect 17882 8518 17894 8570
rect 17956 8518 17958 8570
rect 17796 8516 17820 8518
rect 17876 8516 17900 8518
rect 17956 8516 17980 8518
rect 17740 8496 18036 8516
rect 3764 8468 3816 8474
rect 3764 8410 3816 8416
rect 20140 8264 20192 8270
rect 20140 8206 20192 8212
rect 4420 8028 4716 8048
rect 4476 8026 4500 8028
rect 4556 8026 4580 8028
rect 4636 8026 4660 8028
rect 4498 7974 4500 8026
rect 4562 7974 4574 8026
rect 4636 7974 4638 8026
rect 4476 7972 4500 7974
rect 4556 7972 4580 7974
rect 4636 7972 4660 7974
rect 4420 7952 4716 7972
rect 9748 8028 10044 8048
rect 9804 8026 9828 8028
rect 9884 8026 9908 8028
rect 9964 8026 9988 8028
rect 9826 7974 9828 8026
rect 9890 7974 9902 8026
rect 9964 7974 9966 8026
rect 9804 7972 9828 7974
rect 9884 7972 9908 7974
rect 9964 7972 9988 7974
rect 9748 7952 10044 7972
rect 15076 8028 15372 8048
rect 15132 8026 15156 8028
rect 15212 8026 15236 8028
rect 15292 8026 15316 8028
rect 15154 7974 15156 8026
rect 15218 7974 15230 8026
rect 15292 7974 15294 8026
rect 15132 7972 15156 7974
rect 15212 7972 15236 7974
rect 15292 7972 15316 7974
rect 15076 7952 15372 7972
rect 20152 7930 20180 8206
rect 20140 7924 20192 7930
rect 20140 7866 20192 7872
rect 3764 7652 3816 7658
rect 3764 7594 3816 7600
rect 3776 7182 3804 7594
rect 7084 7484 7380 7504
rect 7140 7482 7164 7484
rect 7220 7482 7244 7484
rect 7300 7482 7324 7484
rect 7162 7430 7164 7482
rect 7226 7430 7238 7482
rect 7300 7430 7302 7482
rect 7140 7428 7164 7430
rect 7220 7428 7244 7430
rect 7300 7428 7324 7430
rect 7084 7408 7380 7428
rect 12412 7484 12708 7504
rect 12468 7482 12492 7484
rect 12548 7482 12572 7484
rect 12628 7482 12652 7484
rect 12490 7430 12492 7482
rect 12554 7430 12566 7482
rect 12628 7430 12630 7482
rect 12468 7428 12492 7430
rect 12548 7428 12572 7430
rect 12628 7428 12652 7430
rect 12412 7408 12708 7428
rect 17740 7484 18036 7504
rect 17796 7482 17820 7484
rect 17876 7482 17900 7484
rect 17956 7482 17980 7484
rect 17818 7430 17820 7482
rect 17882 7430 17894 7482
rect 17956 7430 17958 7482
rect 17796 7428 17820 7430
rect 17876 7428 17900 7430
rect 17956 7428 17980 7430
rect 17740 7408 18036 7428
rect 3764 7176 3816 7182
rect 3764 7118 3816 7124
rect 19680 7176 19732 7182
rect 19680 7118 19732 7124
rect 4420 6940 4716 6960
rect 4476 6938 4500 6940
rect 4556 6938 4580 6940
rect 4636 6938 4660 6940
rect 4498 6886 4500 6938
rect 4562 6886 4574 6938
rect 4636 6886 4638 6938
rect 4476 6884 4500 6886
rect 4556 6884 4580 6886
rect 4636 6884 4660 6886
rect 4420 6864 4716 6884
rect 9748 6940 10044 6960
rect 9804 6938 9828 6940
rect 9884 6938 9908 6940
rect 9964 6938 9988 6940
rect 9826 6886 9828 6938
rect 9890 6886 9902 6938
rect 9964 6886 9966 6938
rect 9804 6884 9828 6886
rect 9884 6884 9908 6886
rect 9964 6884 9988 6886
rect 9748 6864 10044 6884
rect 15076 6940 15372 6960
rect 15132 6938 15156 6940
rect 15212 6938 15236 6940
rect 15292 6938 15316 6940
rect 15154 6886 15156 6938
rect 15218 6886 15230 6938
rect 15292 6886 15294 6938
rect 15132 6884 15156 6886
rect 15212 6884 15236 6886
rect 15292 6884 15316 6886
rect 15076 6864 15372 6884
rect 19692 6842 19720 7118
rect 19680 6836 19732 6842
rect 19680 6778 19732 6784
rect 3764 6564 3816 6570
rect 3764 6506 3816 6512
rect 3776 6298 3804 6506
rect 7084 6396 7380 6416
rect 7140 6394 7164 6396
rect 7220 6394 7244 6396
rect 7300 6394 7324 6396
rect 7162 6342 7164 6394
rect 7226 6342 7238 6394
rect 7300 6342 7302 6394
rect 7140 6340 7164 6342
rect 7220 6340 7244 6342
rect 7300 6340 7324 6342
rect 7084 6320 7380 6340
rect 12412 6396 12708 6416
rect 12468 6394 12492 6396
rect 12548 6394 12572 6396
rect 12628 6394 12652 6396
rect 12490 6342 12492 6394
rect 12554 6342 12566 6394
rect 12628 6342 12630 6394
rect 12468 6340 12492 6342
rect 12548 6340 12572 6342
rect 12628 6340 12652 6342
rect 12412 6320 12708 6340
rect 17740 6396 18036 6416
rect 17796 6394 17820 6396
rect 17876 6394 17900 6396
rect 17956 6394 17980 6396
rect 17818 6342 17820 6394
rect 17882 6342 17894 6394
rect 17956 6342 17958 6394
rect 17796 6340 17820 6342
rect 17876 6340 17900 6342
rect 17956 6340 17980 6342
rect 17740 6320 18036 6340
rect 3764 6292 3816 6298
rect 3764 6234 3816 6240
rect 20140 6088 20192 6094
rect 20140 6030 20192 6036
rect 4420 5852 4716 5872
rect 4476 5850 4500 5852
rect 4556 5850 4580 5852
rect 4636 5850 4660 5852
rect 4498 5798 4500 5850
rect 4562 5798 4574 5850
rect 4636 5798 4638 5850
rect 4476 5796 4500 5798
rect 4556 5796 4580 5798
rect 4636 5796 4660 5798
rect 4420 5776 4716 5796
rect 9748 5852 10044 5872
rect 9804 5850 9828 5852
rect 9884 5850 9908 5852
rect 9964 5850 9988 5852
rect 9826 5798 9828 5850
rect 9890 5798 9902 5850
rect 9964 5798 9966 5850
rect 9804 5796 9828 5798
rect 9884 5796 9908 5798
rect 9964 5796 9988 5798
rect 9748 5776 10044 5796
rect 15076 5852 15372 5872
rect 15132 5850 15156 5852
rect 15212 5850 15236 5852
rect 15292 5850 15316 5852
rect 15154 5798 15156 5850
rect 15218 5798 15230 5850
rect 15292 5798 15294 5850
rect 15132 5796 15156 5798
rect 15212 5796 15236 5798
rect 15292 5796 15316 5798
rect 15076 5776 15372 5796
rect 20152 5754 20180 6030
rect 20140 5748 20192 5754
rect 20140 5690 20192 5696
rect 3764 5476 3816 5482
rect 3764 5418 3816 5424
rect 3776 5006 3804 5418
rect 7084 5308 7380 5328
rect 7140 5306 7164 5308
rect 7220 5306 7244 5308
rect 7300 5306 7324 5308
rect 7162 5254 7164 5306
rect 7226 5254 7238 5306
rect 7300 5254 7302 5306
rect 7140 5252 7164 5254
rect 7220 5252 7244 5254
rect 7300 5252 7324 5254
rect 7084 5232 7380 5252
rect 12412 5308 12708 5328
rect 12468 5306 12492 5308
rect 12548 5306 12572 5308
rect 12628 5306 12652 5308
rect 12490 5254 12492 5306
rect 12554 5254 12566 5306
rect 12628 5254 12630 5306
rect 12468 5252 12492 5254
rect 12548 5252 12572 5254
rect 12628 5252 12652 5254
rect 12412 5232 12708 5252
rect 17740 5308 18036 5328
rect 17796 5306 17820 5308
rect 17876 5306 17900 5308
rect 17956 5306 17980 5308
rect 17818 5254 17820 5306
rect 17882 5254 17894 5306
rect 17956 5254 17958 5306
rect 17796 5252 17820 5254
rect 17876 5252 17900 5254
rect 17956 5252 17980 5254
rect 17740 5232 18036 5252
rect 3764 5000 3816 5006
rect 3764 4942 3816 4948
rect 19680 5000 19732 5006
rect 19680 4942 19732 4948
rect 4420 4764 4716 4784
rect 4476 4762 4500 4764
rect 4556 4762 4580 4764
rect 4636 4762 4660 4764
rect 4498 4710 4500 4762
rect 4562 4710 4574 4762
rect 4636 4710 4638 4762
rect 4476 4708 4500 4710
rect 4556 4708 4580 4710
rect 4636 4708 4660 4710
rect 4420 4688 4716 4708
rect 9748 4764 10044 4784
rect 9804 4762 9828 4764
rect 9884 4762 9908 4764
rect 9964 4762 9988 4764
rect 9826 4710 9828 4762
rect 9890 4710 9902 4762
rect 9964 4710 9966 4762
rect 9804 4708 9828 4710
rect 9884 4708 9908 4710
rect 9964 4708 9988 4710
rect 9748 4688 10044 4708
rect 15076 4764 15372 4784
rect 15132 4762 15156 4764
rect 15212 4762 15236 4764
rect 15292 4762 15316 4764
rect 15154 4710 15156 4762
rect 15218 4710 15230 4762
rect 15292 4710 15294 4762
rect 15132 4708 15156 4710
rect 15212 4708 15236 4710
rect 15292 4708 15316 4710
rect 15076 4688 15372 4708
rect 19692 4666 19720 4942
rect 19680 4660 19732 4666
rect 19680 4602 19732 4608
rect 3764 4388 3816 4394
rect 3764 4330 3816 4336
rect 3776 4122 3804 4330
rect 7084 4220 7380 4240
rect 7140 4218 7164 4220
rect 7220 4218 7244 4220
rect 7300 4218 7324 4220
rect 7162 4166 7164 4218
rect 7226 4166 7238 4218
rect 7300 4166 7302 4218
rect 7140 4164 7164 4166
rect 7220 4164 7244 4166
rect 7300 4164 7324 4166
rect 7084 4144 7380 4164
rect 12412 4220 12708 4240
rect 12468 4218 12492 4220
rect 12548 4218 12572 4220
rect 12628 4218 12652 4220
rect 12490 4166 12492 4218
rect 12554 4166 12566 4218
rect 12628 4166 12630 4218
rect 12468 4164 12492 4166
rect 12548 4164 12572 4166
rect 12628 4164 12652 4166
rect 12412 4144 12708 4164
rect 17740 4220 18036 4240
rect 17796 4218 17820 4220
rect 17876 4218 17900 4220
rect 17956 4218 17980 4220
rect 17818 4166 17820 4218
rect 17882 4166 17894 4218
rect 17956 4166 17958 4218
rect 17796 4164 17820 4166
rect 17876 4164 17900 4166
rect 17956 4164 17980 4166
rect 17740 4144 18036 4164
rect 3764 4116 3816 4122
rect 3764 4058 3816 4064
rect 20232 3912 20284 3918
rect 20232 3854 20284 3860
rect 4420 3676 4716 3696
rect 4476 3674 4500 3676
rect 4556 3674 4580 3676
rect 4636 3674 4660 3676
rect 4498 3622 4500 3674
rect 4562 3622 4574 3674
rect 4636 3622 4638 3674
rect 4476 3620 4500 3622
rect 4556 3620 4580 3622
rect 4636 3620 4660 3622
rect 4420 3600 4716 3620
rect 9748 3676 10044 3696
rect 9804 3674 9828 3676
rect 9884 3674 9908 3676
rect 9964 3674 9988 3676
rect 9826 3622 9828 3674
rect 9890 3622 9902 3674
rect 9964 3622 9966 3674
rect 9804 3620 9828 3622
rect 9884 3620 9908 3622
rect 9964 3620 9988 3622
rect 9748 3600 10044 3620
rect 15076 3676 15372 3696
rect 15132 3674 15156 3676
rect 15212 3674 15236 3676
rect 15292 3674 15316 3676
rect 15154 3622 15156 3674
rect 15218 3622 15230 3674
rect 15292 3622 15294 3674
rect 15132 3620 15156 3622
rect 15212 3620 15236 3622
rect 15292 3620 15316 3622
rect 15076 3600 15372 3620
rect 20244 3510 20272 3854
rect 20232 3504 20284 3510
rect 20232 3446 20284 3452
rect 3764 3300 3816 3306
rect 3764 3242 3816 3248
rect 3776 3034 3804 3242
rect 7084 3132 7380 3152
rect 7140 3130 7164 3132
rect 7220 3130 7244 3132
rect 7300 3130 7324 3132
rect 7162 3078 7164 3130
rect 7226 3078 7238 3130
rect 7300 3078 7302 3130
rect 7140 3076 7164 3078
rect 7220 3076 7244 3078
rect 7300 3076 7324 3078
rect 7084 3056 7380 3076
rect 12412 3132 12708 3152
rect 12468 3130 12492 3132
rect 12548 3130 12572 3132
rect 12628 3130 12652 3132
rect 12490 3078 12492 3130
rect 12554 3078 12566 3130
rect 12628 3078 12630 3130
rect 12468 3076 12492 3078
rect 12548 3076 12572 3078
rect 12628 3076 12652 3078
rect 12412 3056 12708 3076
rect 17740 3132 18036 3152
rect 17796 3130 17820 3132
rect 17876 3130 17900 3132
rect 17956 3130 17980 3132
rect 17818 3078 17820 3130
rect 17882 3078 17894 3130
rect 17956 3078 17958 3130
rect 17796 3076 17820 3078
rect 17876 3076 17900 3078
rect 17956 3076 17980 3078
rect 17740 3056 18036 3076
rect 3764 3028 3816 3034
rect 3764 2970 3816 2976
rect 14988 2824 15040 2830
rect 14988 2766 15040 2772
rect 20140 2824 20192 2830
rect 20140 2766 20192 2772
rect 15000 2694 15028 2766
rect 14988 2688 15040 2694
rect 14988 2630 15040 2636
rect 4420 2588 4716 2608
rect 4476 2586 4500 2588
rect 4556 2586 4580 2588
rect 4636 2586 4660 2588
rect 4498 2534 4500 2586
rect 4562 2534 4574 2586
rect 4636 2534 4638 2586
rect 4476 2532 4500 2534
rect 4556 2532 4580 2534
rect 4636 2532 4660 2534
rect 4420 2512 4716 2532
rect 9748 2588 10044 2608
rect 9804 2586 9828 2588
rect 9884 2586 9908 2588
rect 9964 2586 9988 2588
rect 9826 2534 9828 2586
rect 9890 2534 9902 2586
rect 9964 2534 9966 2586
rect 9804 2532 9828 2534
rect 9884 2532 9908 2534
rect 9964 2532 9988 2534
rect 9748 2512 10044 2532
rect 15076 2588 15372 2608
rect 15132 2586 15156 2588
rect 15212 2586 15236 2588
rect 15292 2586 15316 2588
rect 15154 2534 15156 2586
rect 15218 2534 15230 2586
rect 15292 2534 15294 2586
rect 15132 2532 15156 2534
rect 15212 2532 15236 2534
rect 15292 2532 15316 2534
rect 15076 2512 15372 2532
rect 20152 2490 20180 2766
rect 20140 2484 20192 2490
rect 20140 2426 20192 2432
rect 3764 2212 3816 2218
rect 3764 2154 3816 2160
rect 3776 1946 3804 2154
rect 7084 2044 7380 2064
rect 7140 2042 7164 2044
rect 7220 2042 7244 2044
rect 7300 2042 7324 2044
rect 7162 1990 7164 2042
rect 7226 1990 7238 2042
rect 7300 1990 7302 2042
rect 7140 1988 7164 1990
rect 7220 1988 7244 1990
rect 7300 1988 7324 1990
rect 7084 1968 7380 1988
rect 12412 2044 12708 2064
rect 12468 2042 12492 2044
rect 12548 2042 12572 2044
rect 12628 2042 12652 2044
rect 12490 1990 12492 2042
rect 12554 1990 12566 2042
rect 12628 1990 12630 2042
rect 12468 1988 12492 1990
rect 12548 1988 12572 1990
rect 12628 1988 12652 1990
rect 12412 1968 12708 1988
rect 17740 2044 18036 2064
rect 17796 2042 17820 2044
rect 17876 2042 17900 2044
rect 17956 2042 17980 2044
rect 17818 1990 17820 2042
rect 17882 1990 17894 2042
rect 17956 1990 17958 2042
rect 17796 1988 17820 1990
rect 17876 1988 17900 1990
rect 17956 1988 17980 1990
rect 17740 1968 18036 1988
rect 3764 1940 3816 1946
rect 3764 1882 3816 1888
rect 20140 1736 20192 1742
rect 20140 1678 20192 1684
rect 4420 1500 4716 1520
rect 4476 1498 4500 1500
rect 4556 1498 4580 1500
rect 4636 1498 4660 1500
rect 4498 1446 4500 1498
rect 4562 1446 4574 1498
rect 4636 1446 4638 1498
rect 4476 1444 4500 1446
rect 4556 1444 4580 1446
rect 4636 1444 4660 1446
rect 4420 1424 4716 1444
rect 9748 1500 10044 1520
rect 9804 1498 9828 1500
rect 9884 1498 9908 1500
rect 9964 1498 9988 1500
rect 9826 1446 9828 1498
rect 9890 1446 9902 1498
rect 9964 1446 9966 1498
rect 9804 1444 9828 1446
rect 9884 1444 9908 1446
rect 9964 1444 9988 1446
rect 9748 1424 10044 1444
rect 15076 1500 15372 1520
rect 15132 1498 15156 1500
rect 15212 1498 15236 1500
rect 15292 1498 15316 1500
rect 15154 1446 15156 1498
rect 15218 1446 15230 1498
rect 15292 1446 15294 1498
rect 15132 1444 15156 1446
rect 15212 1444 15236 1446
rect 15292 1444 15316 1446
rect 15076 1424 15372 1444
rect 20152 1402 20180 1678
rect 20140 1396 20192 1402
rect 20140 1338 20192 1344
rect 2936 1260 2988 1266
rect 2936 1202 2988 1208
rect 2948 1169 2976 1202
rect 2290 1160 2346 1169
rect 2290 1095 2346 1104
rect 2934 1160 2990 1169
rect 2934 1095 2990 1104
rect 7084 956 7380 976
rect 7140 954 7164 956
rect 7220 954 7244 956
rect 7300 954 7324 956
rect 7162 902 7164 954
rect 7226 902 7238 954
rect 7300 902 7302 954
rect 7140 900 7164 902
rect 7220 900 7244 902
rect 7300 900 7324 902
rect 7084 880 7380 900
rect 12412 956 12708 976
rect 12468 954 12492 956
rect 12548 954 12572 956
rect 12628 954 12652 956
rect 12490 902 12492 954
rect 12554 902 12566 954
rect 12628 902 12630 954
rect 12468 900 12492 902
rect 12548 900 12572 902
rect 12628 900 12652 902
rect 12412 880 12708 900
rect 17740 956 18036 976
rect 17796 954 17820 956
rect 17876 954 17900 956
rect 17956 954 17980 956
rect 17818 902 17820 954
rect 17882 902 17894 954
rect 17956 902 17958 954
rect 17796 900 17820 902
rect 17876 900 17900 902
rect 17956 900 17980 902
rect 17740 880 18036 900
<< via2 >>
rect 1922 22320 1978 22376
rect 4420 22170 4476 22172
rect 4500 22170 4556 22172
rect 4580 22170 4636 22172
rect 4660 22170 4716 22172
rect 4420 22118 4446 22170
rect 4446 22118 4476 22170
rect 4500 22118 4510 22170
rect 4510 22118 4556 22170
rect 4580 22118 4626 22170
rect 4626 22118 4636 22170
rect 4660 22118 4690 22170
rect 4690 22118 4716 22170
rect 4420 22116 4476 22118
rect 4500 22116 4556 22118
rect 4580 22116 4636 22118
rect 4660 22116 4716 22118
rect 9748 22170 9804 22172
rect 9828 22170 9884 22172
rect 9908 22170 9964 22172
rect 9988 22170 10044 22172
rect 9748 22118 9774 22170
rect 9774 22118 9804 22170
rect 9828 22118 9838 22170
rect 9838 22118 9884 22170
rect 9908 22118 9954 22170
rect 9954 22118 9964 22170
rect 9988 22118 10018 22170
rect 10018 22118 10044 22170
rect 9748 22116 9804 22118
rect 9828 22116 9884 22118
rect 9908 22116 9964 22118
rect 9988 22116 10044 22118
rect 15076 22170 15132 22172
rect 15156 22170 15212 22172
rect 15236 22170 15292 22172
rect 15316 22170 15372 22172
rect 15076 22118 15102 22170
rect 15102 22118 15132 22170
rect 15156 22118 15166 22170
rect 15166 22118 15212 22170
rect 15236 22118 15282 22170
rect 15282 22118 15292 22170
rect 15316 22118 15346 22170
rect 15346 22118 15372 22170
rect 15076 22116 15132 22118
rect 15156 22116 15212 22118
rect 15236 22116 15292 22118
rect 15316 22116 15372 22118
rect 2474 21812 2476 21832
rect 2476 21812 2528 21832
rect 2528 21812 2530 21832
rect 2474 21776 2530 21812
rect 7084 21626 7140 21628
rect 7164 21626 7220 21628
rect 7244 21626 7300 21628
rect 7324 21626 7380 21628
rect 7084 21574 7110 21626
rect 7110 21574 7140 21626
rect 7164 21574 7174 21626
rect 7174 21574 7220 21626
rect 7244 21574 7290 21626
rect 7290 21574 7300 21626
rect 7324 21574 7354 21626
rect 7354 21574 7380 21626
rect 7084 21572 7140 21574
rect 7164 21572 7220 21574
rect 7244 21572 7300 21574
rect 7324 21572 7380 21574
rect 12412 21626 12468 21628
rect 12492 21626 12548 21628
rect 12572 21626 12628 21628
rect 12652 21626 12708 21628
rect 12412 21574 12438 21626
rect 12438 21574 12468 21626
rect 12492 21574 12502 21626
rect 12502 21574 12548 21626
rect 12572 21574 12618 21626
rect 12618 21574 12628 21626
rect 12652 21574 12682 21626
rect 12682 21574 12708 21626
rect 12412 21572 12468 21574
rect 12492 21572 12548 21574
rect 12572 21572 12628 21574
rect 12652 21572 12708 21574
rect 17740 21626 17796 21628
rect 17820 21626 17876 21628
rect 17900 21626 17956 21628
rect 17980 21626 18036 21628
rect 17740 21574 17766 21626
rect 17766 21574 17796 21626
rect 17820 21574 17830 21626
rect 17830 21574 17876 21626
rect 17900 21574 17946 21626
rect 17946 21574 17956 21626
rect 17980 21574 18010 21626
rect 18010 21574 18036 21626
rect 17740 21572 17796 21574
rect 17820 21572 17876 21574
rect 17900 21572 17956 21574
rect 17980 21572 18036 21574
rect 2474 21232 2530 21288
rect 4420 21082 4476 21084
rect 4500 21082 4556 21084
rect 4580 21082 4636 21084
rect 4660 21082 4716 21084
rect 4420 21030 4446 21082
rect 4446 21030 4476 21082
rect 4500 21030 4510 21082
rect 4510 21030 4556 21082
rect 4580 21030 4626 21082
rect 4626 21030 4636 21082
rect 4660 21030 4690 21082
rect 4690 21030 4716 21082
rect 4420 21028 4476 21030
rect 4500 21028 4556 21030
rect 4580 21028 4636 21030
rect 4660 21028 4716 21030
rect 9748 21082 9804 21084
rect 9828 21082 9884 21084
rect 9908 21082 9964 21084
rect 9988 21082 10044 21084
rect 9748 21030 9774 21082
rect 9774 21030 9804 21082
rect 9828 21030 9838 21082
rect 9838 21030 9884 21082
rect 9908 21030 9954 21082
rect 9954 21030 9964 21082
rect 9988 21030 10018 21082
rect 10018 21030 10044 21082
rect 9748 21028 9804 21030
rect 9828 21028 9884 21030
rect 9908 21028 9964 21030
rect 9988 21028 10044 21030
rect 15076 21082 15132 21084
rect 15156 21082 15212 21084
rect 15236 21082 15292 21084
rect 15316 21082 15372 21084
rect 15076 21030 15102 21082
rect 15102 21030 15132 21082
rect 15156 21030 15166 21082
rect 15166 21030 15212 21082
rect 15236 21030 15282 21082
rect 15282 21030 15292 21082
rect 15316 21030 15346 21082
rect 15346 21030 15372 21082
rect 15076 21028 15132 21030
rect 15156 21028 15212 21030
rect 15236 21028 15292 21030
rect 15316 21028 15372 21030
rect 7084 20538 7140 20540
rect 7164 20538 7220 20540
rect 7244 20538 7300 20540
rect 7324 20538 7380 20540
rect 7084 20486 7110 20538
rect 7110 20486 7140 20538
rect 7164 20486 7174 20538
rect 7174 20486 7220 20538
rect 7244 20486 7290 20538
rect 7290 20486 7300 20538
rect 7324 20486 7354 20538
rect 7354 20486 7380 20538
rect 7084 20484 7140 20486
rect 7164 20484 7220 20486
rect 7244 20484 7300 20486
rect 7324 20484 7380 20486
rect 12412 20538 12468 20540
rect 12492 20538 12548 20540
rect 12572 20538 12628 20540
rect 12652 20538 12708 20540
rect 12412 20486 12438 20538
rect 12438 20486 12468 20538
rect 12492 20486 12502 20538
rect 12502 20486 12548 20538
rect 12572 20486 12618 20538
rect 12618 20486 12628 20538
rect 12652 20486 12682 20538
rect 12682 20486 12708 20538
rect 12412 20484 12468 20486
rect 12492 20484 12548 20486
rect 12572 20484 12628 20486
rect 12652 20484 12708 20486
rect 17740 20538 17796 20540
rect 17820 20538 17876 20540
rect 17900 20538 17956 20540
rect 17980 20538 18036 20540
rect 17740 20486 17766 20538
rect 17766 20486 17796 20538
rect 17820 20486 17830 20538
rect 17830 20486 17876 20538
rect 17900 20486 17946 20538
rect 17946 20486 17956 20538
rect 17980 20486 18010 20538
rect 18010 20486 18036 20538
rect 17740 20484 17796 20486
rect 17820 20484 17876 20486
rect 17900 20484 17956 20486
rect 17980 20484 18036 20486
rect 2474 20144 2530 20200
rect 4420 19994 4476 19996
rect 4500 19994 4556 19996
rect 4580 19994 4636 19996
rect 4660 19994 4716 19996
rect 4420 19942 4446 19994
rect 4446 19942 4476 19994
rect 4500 19942 4510 19994
rect 4510 19942 4556 19994
rect 4580 19942 4626 19994
rect 4626 19942 4636 19994
rect 4660 19942 4690 19994
rect 4690 19942 4716 19994
rect 4420 19940 4476 19942
rect 4500 19940 4556 19942
rect 4580 19940 4636 19942
rect 4660 19940 4716 19942
rect 9748 19994 9804 19996
rect 9828 19994 9884 19996
rect 9908 19994 9964 19996
rect 9988 19994 10044 19996
rect 9748 19942 9774 19994
rect 9774 19942 9804 19994
rect 9828 19942 9838 19994
rect 9838 19942 9884 19994
rect 9908 19942 9954 19994
rect 9954 19942 9964 19994
rect 9988 19942 10018 19994
rect 10018 19942 10044 19994
rect 9748 19940 9804 19942
rect 9828 19940 9884 19942
rect 9908 19940 9964 19942
rect 9988 19940 10044 19942
rect 15076 19994 15132 19996
rect 15156 19994 15212 19996
rect 15236 19994 15292 19996
rect 15316 19994 15372 19996
rect 15076 19942 15102 19994
rect 15102 19942 15132 19994
rect 15156 19942 15166 19994
rect 15166 19942 15212 19994
rect 15236 19942 15282 19994
rect 15282 19942 15292 19994
rect 15316 19942 15346 19994
rect 15346 19942 15372 19994
rect 15076 19940 15132 19942
rect 15156 19940 15212 19942
rect 15236 19940 15292 19942
rect 15316 19940 15372 19942
rect 7084 19450 7140 19452
rect 7164 19450 7220 19452
rect 7244 19450 7300 19452
rect 7324 19450 7380 19452
rect 7084 19398 7110 19450
rect 7110 19398 7140 19450
rect 7164 19398 7174 19450
rect 7174 19398 7220 19450
rect 7244 19398 7290 19450
rect 7290 19398 7300 19450
rect 7324 19398 7354 19450
rect 7354 19398 7380 19450
rect 7084 19396 7140 19398
rect 7164 19396 7220 19398
rect 7244 19396 7300 19398
rect 7324 19396 7380 19398
rect 12412 19450 12468 19452
rect 12492 19450 12548 19452
rect 12572 19450 12628 19452
rect 12652 19450 12708 19452
rect 12412 19398 12438 19450
rect 12438 19398 12468 19450
rect 12492 19398 12502 19450
rect 12502 19398 12548 19450
rect 12572 19398 12618 19450
rect 12618 19398 12628 19450
rect 12652 19398 12682 19450
rect 12682 19398 12708 19450
rect 12412 19396 12468 19398
rect 12492 19396 12548 19398
rect 12572 19396 12628 19398
rect 12652 19396 12708 19398
rect 17740 19450 17796 19452
rect 17820 19450 17876 19452
rect 17900 19450 17956 19452
rect 17980 19450 18036 19452
rect 17740 19398 17766 19450
rect 17766 19398 17796 19450
rect 17820 19398 17830 19450
rect 17830 19398 17876 19450
rect 17900 19398 17946 19450
rect 17946 19398 17956 19450
rect 17980 19398 18010 19450
rect 18010 19398 18036 19450
rect 17740 19396 17796 19398
rect 17820 19396 17876 19398
rect 17900 19396 17956 19398
rect 17980 19396 18036 19398
rect 2474 19056 2530 19112
rect 4420 18906 4476 18908
rect 4500 18906 4556 18908
rect 4580 18906 4636 18908
rect 4660 18906 4716 18908
rect 4420 18854 4446 18906
rect 4446 18854 4476 18906
rect 4500 18854 4510 18906
rect 4510 18854 4556 18906
rect 4580 18854 4626 18906
rect 4626 18854 4636 18906
rect 4660 18854 4690 18906
rect 4690 18854 4716 18906
rect 4420 18852 4476 18854
rect 4500 18852 4556 18854
rect 4580 18852 4636 18854
rect 4660 18852 4716 18854
rect 9748 18906 9804 18908
rect 9828 18906 9884 18908
rect 9908 18906 9964 18908
rect 9988 18906 10044 18908
rect 9748 18854 9774 18906
rect 9774 18854 9804 18906
rect 9828 18854 9838 18906
rect 9838 18854 9884 18906
rect 9908 18854 9954 18906
rect 9954 18854 9964 18906
rect 9988 18854 10018 18906
rect 10018 18854 10044 18906
rect 9748 18852 9804 18854
rect 9828 18852 9884 18854
rect 9908 18852 9964 18854
rect 9988 18852 10044 18854
rect 15076 18906 15132 18908
rect 15156 18906 15212 18908
rect 15236 18906 15292 18908
rect 15316 18906 15372 18908
rect 15076 18854 15102 18906
rect 15102 18854 15132 18906
rect 15156 18854 15166 18906
rect 15166 18854 15212 18906
rect 15236 18854 15282 18906
rect 15282 18854 15292 18906
rect 15316 18854 15346 18906
rect 15346 18854 15372 18906
rect 15076 18852 15132 18854
rect 15156 18852 15212 18854
rect 15236 18852 15292 18854
rect 15316 18852 15372 18854
rect 7084 18362 7140 18364
rect 7164 18362 7220 18364
rect 7244 18362 7300 18364
rect 7324 18362 7380 18364
rect 7084 18310 7110 18362
rect 7110 18310 7140 18362
rect 7164 18310 7174 18362
rect 7174 18310 7220 18362
rect 7244 18310 7290 18362
rect 7290 18310 7300 18362
rect 7324 18310 7354 18362
rect 7354 18310 7380 18362
rect 7084 18308 7140 18310
rect 7164 18308 7220 18310
rect 7244 18308 7300 18310
rect 7324 18308 7380 18310
rect 12412 18362 12468 18364
rect 12492 18362 12548 18364
rect 12572 18362 12628 18364
rect 12652 18362 12708 18364
rect 12412 18310 12438 18362
rect 12438 18310 12468 18362
rect 12492 18310 12502 18362
rect 12502 18310 12548 18362
rect 12572 18310 12618 18362
rect 12618 18310 12628 18362
rect 12652 18310 12682 18362
rect 12682 18310 12708 18362
rect 12412 18308 12468 18310
rect 12492 18308 12548 18310
rect 12572 18308 12628 18310
rect 12652 18308 12708 18310
rect 17740 18362 17796 18364
rect 17820 18362 17876 18364
rect 17900 18362 17956 18364
rect 17980 18362 18036 18364
rect 17740 18310 17766 18362
rect 17766 18310 17796 18362
rect 17820 18310 17830 18362
rect 17830 18310 17876 18362
rect 17900 18310 17946 18362
rect 17946 18310 17956 18362
rect 17980 18310 18010 18362
rect 18010 18310 18036 18362
rect 17740 18308 17796 18310
rect 17820 18308 17876 18310
rect 17900 18308 17956 18310
rect 17980 18308 18036 18310
rect 2474 17968 2530 18024
rect 4420 17818 4476 17820
rect 4500 17818 4556 17820
rect 4580 17818 4636 17820
rect 4660 17818 4716 17820
rect 4420 17766 4446 17818
rect 4446 17766 4476 17818
rect 4500 17766 4510 17818
rect 4510 17766 4556 17818
rect 4580 17766 4626 17818
rect 4626 17766 4636 17818
rect 4660 17766 4690 17818
rect 4690 17766 4716 17818
rect 4420 17764 4476 17766
rect 4500 17764 4556 17766
rect 4580 17764 4636 17766
rect 4660 17764 4716 17766
rect 9748 17818 9804 17820
rect 9828 17818 9884 17820
rect 9908 17818 9964 17820
rect 9988 17818 10044 17820
rect 9748 17766 9774 17818
rect 9774 17766 9804 17818
rect 9828 17766 9838 17818
rect 9838 17766 9884 17818
rect 9908 17766 9954 17818
rect 9954 17766 9964 17818
rect 9988 17766 10018 17818
rect 10018 17766 10044 17818
rect 9748 17764 9804 17766
rect 9828 17764 9884 17766
rect 9908 17764 9964 17766
rect 9988 17764 10044 17766
rect 15076 17818 15132 17820
rect 15156 17818 15212 17820
rect 15236 17818 15292 17820
rect 15316 17818 15372 17820
rect 15076 17766 15102 17818
rect 15102 17766 15132 17818
rect 15156 17766 15166 17818
rect 15166 17766 15212 17818
rect 15236 17766 15282 17818
rect 15282 17766 15292 17818
rect 15316 17766 15346 17818
rect 15346 17766 15372 17818
rect 15076 17764 15132 17766
rect 15156 17764 15212 17766
rect 15236 17764 15292 17766
rect 15316 17764 15372 17766
rect 7084 17274 7140 17276
rect 7164 17274 7220 17276
rect 7244 17274 7300 17276
rect 7324 17274 7380 17276
rect 7084 17222 7110 17274
rect 7110 17222 7140 17274
rect 7164 17222 7174 17274
rect 7174 17222 7220 17274
rect 7244 17222 7290 17274
rect 7290 17222 7300 17274
rect 7324 17222 7354 17274
rect 7354 17222 7380 17274
rect 7084 17220 7140 17222
rect 7164 17220 7220 17222
rect 7244 17220 7300 17222
rect 7324 17220 7380 17222
rect 12412 17274 12468 17276
rect 12492 17274 12548 17276
rect 12572 17274 12628 17276
rect 12652 17274 12708 17276
rect 12412 17222 12438 17274
rect 12438 17222 12468 17274
rect 12492 17222 12502 17274
rect 12502 17222 12548 17274
rect 12572 17222 12618 17274
rect 12618 17222 12628 17274
rect 12652 17222 12682 17274
rect 12682 17222 12708 17274
rect 12412 17220 12468 17222
rect 12492 17220 12548 17222
rect 12572 17220 12628 17222
rect 12652 17220 12708 17222
rect 17740 17274 17796 17276
rect 17820 17274 17876 17276
rect 17900 17274 17956 17276
rect 17980 17274 18036 17276
rect 17740 17222 17766 17274
rect 17766 17222 17796 17274
rect 17820 17222 17830 17274
rect 17830 17222 17876 17274
rect 17900 17222 17946 17274
rect 17946 17222 17956 17274
rect 17980 17222 18010 17274
rect 18010 17222 18036 17274
rect 17740 17220 17796 17222
rect 17820 17220 17876 17222
rect 17900 17220 17956 17222
rect 17980 17220 18036 17222
rect 4420 16730 4476 16732
rect 4500 16730 4556 16732
rect 4580 16730 4636 16732
rect 4660 16730 4716 16732
rect 4420 16678 4446 16730
rect 4446 16678 4476 16730
rect 4500 16678 4510 16730
rect 4510 16678 4556 16730
rect 4580 16678 4626 16730
rect 4626 16678 4636 16730
rect 4660 16678 4690 16730
rect 4690 16678 4716 16730
rect 4420 16676 4476 16678
rect 4500 16676 4556 16678
rect 4580 16676 4636 16678
rect 4660 16676 4716 16678
rect 2474 16608 2530 16664
rect 9748 16730 9804 16732
rect 9828 16730 9884 16732
rect 9908 16730 9964 16732
rect 9988 16730 10044 16732
rect 9748 16678 9774 16730
rect 9774 16678 9804 16730
rect 9828 16678 9838 16730
rect 9838 16678 9884 16730
rect 9908 16678 9954 16730
rect 9954 16678 9964 16730
rect 9988 16678 10018 16730
rect 10018 16678 10044 16730
rect 9748 16676 9804 16678
rect 9828 16676 9884 16678
rect 9908 16676 9964 16678
rect 9988 16676 10044 16678
rect 15076 16730 15132 16732
rect 15156 16730 15212 16732
rect 15236 16730 15292 16732
rect 15316 16730 15372 16732
rect 15076 16678 15102 16730
rect 15102 16678 15132 16730
rect 15156 16678 15166 16730
rect 15166 16678 15212 16730
rect 15236 16678 15282 16730
rect 15282 16678 15292 16730
rect 15316 16678 15346 16730
rect 15346 16678 15372 16730
rect 15076 16676 15132 16678
rect 15156 16676 15212 16678
rect 15236 16676 15292 16678
rect 15316 16676 15372 16678
rect 7084 16186 7140 16188
rect 7164 16186 7220 16188
rect 7244 16186 7300 16188
rect 7324 16186 7380 16188
rect 7084 16134 7110 16186
rect 7110 16134 7140 16186
rect 7164 16134 7174 16186
rect 7174 16134 7220 16186
rect 7244 16134 7290 16186
rect 7290 16134 7300 16186
rect 7324 16134 7354 16186
rect 7354 16134 7380 16186
rect 7084 16132 7140 16134
rect 7164 16132 7220 16134
rect 7244 16132 7300 16134
rect 7324 16132 7380 16134
rect 12412 16186 12468 16188
rect 12492 16186 12548 16188
rect 12572 16186 12628 16188
rect 12652 16186 12708 16188
rect 12412 16134 12438 16186
rect 12438 16134 12468 16186
rect 12492 16134 12502 16186
rect 12502 16134 12548 16186
rect 12572 16134 12618 16186
rect 12618 16134 12628 16186
rect 12652 16134 12682 16186
rect 12682 16134 12708 16186
rect 12412 16132 12468 16134
rect 12492 16132 12548 16134
rect 12572 16132 12628 16134
rect 12652 16132 12708 16134
rect 17740 16186 17796 16188
rect 17820 16186 17876 16188
rect 17900 16186 17956 16188
rect 17980 16186 18036 16188
rect 17740 16134 17766 16186
rect 17766 16134 17796 16186
rect 17820 16134 17830 16186
rect 17830 16134 17876 16186
rect 17900 16134 17946 16186
rect 17946 16134 17956 16186
rect 17980 16134 18010 16186
rect 18010 16134 18036 16186
rect 17740 16132 17796 16134
rect 17820 16132 17876 16134
rect 17900 16132 17956 16134
rect 17980 16132 18036 16134
rect 2474 15792 2530 15848
rect 4420 15642 4476 15644
rect 4500 15642 4556 15644
rect 4580 15642 4636 15644
rect 4660 15642 4716 15644
rect 4420 15590 4446 15642
rect 4446 15590 4476 15642
rect 4500 15590 4510 15642
rect 4510 15590 4556 15642
rect 4580 15590 4626 15642
rect 4626 15590 4636 15642
rect 4660 15590 4690 15642
rect 4690 15590 4716 15642
rect 4420 15588 4476 15590
rect 4500 15588 4556 15590
rect 4580 15588 4636 15590
rect 4660 15588 4716 15590
rect 9748 15642 9804 15644
rect 9828 15642 9884 15644
rect 9908 15642 9964 15644
rect 9988 15642 10044 15644
rect 9748 15590 9774 15642
rect 9774 15590 9804 15642
rect 9828 15590 9838 15642
rect 9838 15590 9884 15642
rect 9908 15590 9954 15642
rect 9954 15590 9964 15642
rect 9988 15590 10018 15642
rect 10018 15590 10044 15642
rect 9748 15588 9804 15590
rect 9828 15588 9884 15590
rect 9908 15588 9964 15590
rect 9988 15588 10044 15590
rect 15076 15642 15132 15644
rect 15156 15642 15212 15644
rect 15236 15642 15292 15644
rect 15316 15642 15372 15644
rect 15076 15590 15102 15642
rect 15102 15590 15132 15642
rect 15156 15590 15166 15642
rect 15166 15590 15212 15642
rect 15236 15590 15282 15642
rect 15282 15590 15292 15642
rect 15316 15590 15346 15642
rect 15346 15590 15372 15642
rect 15076 15588 15132 15590
rect 15156 15588 15212 15590
rect 15236 15588 15292 15590
rect 15316 15588 15372 15590
rect 7084 15098 7140 15100
rect 7164 15098 7220 15100
rect 7244 15098 7300 15100
rect 7324 15098 7380 15100
rect 7084 15046 7110 15098
rect 7110 15046 7140 15098
rect 7164 15046 7174 15098
rect 7174 15046 7220 15098
rect 7244 15046 7290 15098
rect 7290 15046 7300 15098
rect 7324 15046 7354 15098
rect 7354 15046 7380 15098
rect 7084 15044 7140 15046
rect 7164 15044 7220 15046
rect 7244 15044 7300 15046
rect 7324 15044 7380 15046
rect 12412 15098 12468 15100
rect 12492 15098 12548 15100
rect 12572 15098 12628 15100
rect 12652 15098 12708 15100
rect 12412 15046 12438 15098
rect 12438 15046 12468 15098
rect 12492 15046 12502 15098
rect 12502 15046 12548 15098
rect 12572 15046 12618 15098
rect 12618 15046 12628 15098
rect 12652 15046 12682 15098
rect 12682 15046 12708 15098
rect 12412 15044 12468 15046
rect 12492 15044 12548 15046
rect 12572 15044 12628 15046
rect 12652 15044 12708 15046
rect 17740 15098 17796 15100
rect 17820 15098 17876 15100
rect 17900 15098 17956 15100
rect 17980 15098 18036 15100
rect 17740 15046 17766 15098
rect 17766 15046 17796 15098
rect 17820 15046 17830 15098
rect 17830 15046 17876 15098
rect 17900 15046 17946 15098
rect 17946 15046 17956 15098
rect 17980 15046 18010 15098
rect 18010 15046 18036 15098
rect 17740 15044 17796 15046
rect 17820 15044 17876 15046
rect 17900 15044 17956 15046
rect 17980 15044 18036 15046
rect 4420 14554 4476 14556
rect 4500 14554 4556 14556
rect 4580 14554 4636 14556
rect 4660 14554 4716 14556
rect 4420 14502 4446 14554
rect 4446 14502 4476 14554
rect 4500 14502 4510 14554
rect 4510 14502 4556 14554
rect 4580 14502 4626 14554
rect 4626 14502 4636 14554
rect 4660 14502 4690 14554
rect 4690 14502 4716 14554
rect 4420 14500 4476 14502
rect 4500 14500 4556 14502
rect 4580 14500 4636 14502
rect 4660 14500 4716 14502
rect 9748 14554 9804 14556
rect 9828 14554 9884 14556
rect 9908 14554 9964 14556
rect 9988 14554 10044 14556
rect 9748 14502 9774 14554
rect 9774 14502 9804 14554
rect 9828 14502 9838 14554
rect 9838 14502 9884 14554
rect 9908 14502 9954 14554
rect 9954 14502 9964 14554
rect 9988 14502 10018 14554
rect 10018 14502 10044 14554
rect 9748 14500 9804 14502
rect 9828 14500 9884 14502
rect 9908 14500 9964 14502
rect 9988 14500 10044 14502
rect 15076 14554 15132 14556
rect 15156 14554 15212 14556
rect 15236 14554 15292 14556
rect 15316 14554 15372 14556
rect 15076 14502 15102 14554
rect 15102 14502 15132 14554
rect 15156 14502 15166 14554
rect 15166 14502 15212 14554
rect 15236 14502 15282 14554
rect 15282 14502 15292 14554
rect 15316 14502 15346 14554
rect 15346 14502 15372 14554
rect 15076 14500 15132 14502
rect 15156 14500 15212 14502
rect 15236 14500 15292 14502
rect 15316 14500 15372 14502
rect 7084 14010 7140 14012
rect 7164 14010 7220 14012
rect 7244 14010 7300 14012
rect 7324 14010 7380 14012
rect 7084 13958 7110 14010
rect 7110 13958 7140 14010
rect 7164 13958 7174 14010
rect 7174 13958 7220 14010
rect 7244 13958 7290 14010
rect 7290 13958 7300 14010
rect 7324 13958 7354 14010
rect 7354 13958 7380 14010
rect 7084 13956 7140 13958
rect 7164 13956 7220 13958
rect 7244 13956 7300 13958
rect 7324 13956 7380 13958
rect 12412 14010 12468 14012
rect 12492 14010 12548 14012
rect 12572 14010 12628 14012
rect 12652 14010 12708 14012
rect 12412 13958 12438 14010
rect 12438 13958 12468 14010
rect 12492 13958 12502 14010
rect 12502 13958 12548 14010
rect 12572 13958 12618 14010
rect 12618 13958 12628 14010
rect 12652 13958 12682 14010
rect 12682 13958 12708 14010
rect 12412 13956 12468 13958
rect 12492 13956 12548 13958
rect 12572 13956 12628 13958
rect 12652 13956 12708 13958
rect 17740 14010 17796 14012
rect 17820 14010 17876 14012
rect 17900 14010 17956 14012
rect 17980 14010 18036 14012
rect 17740 13958 17766 14010
rect 17766 13958 17796 14010
rect 17820 13958 17830 14010
rect 17830 13958 17876 14010
rect 17900 13958 17946 14010
rect 17946 13958 17956 14010
rect 17980 13958 18010 14010
rect 18010 13958 18036 14010
rect 17740 13956 17796 13958
rect 17820 13956 17876 13958
rect 17900 13956 17956 13958
rect 17980 13956 18036 13958
rect 2474 13616 2530 13672
rect 4420 13466 4476 13468
rect 4500 13466 4556 13468
rect 4580 13466 4636 13468
rect 4660 13466 4716 13468
rect 4420 13414 4446 13466
rect 4446 13414 4476 13466
rect 4500 13414 4510 13466
rect 4510 13414 4556 13466
rect 4580 13414 4626 13466
rect 4626 13414 4636 13466
rect 4660 13414 4690 13466
rect 4690 13414 4716 13466
rect 4420 13412 4476 13414
rect 4500 13412 4556 13414
rect 4580 13412 4636 13414
rect 4660 13412 4716 13414
rect 9748 13466 9804 13468
rect 9828 13466 9884 13468
rect 9908 13466 9964 13468
rect 9988 13466 10044 13468
rect 9748 13414 9774 13466
rect 9774 13414 9804 13466
rect 9828 13414 9838 13466
rect 9838 13414 9884 13466
rect 9908 13414 9954 13466
rect 9954 13414 9964 13466
rect 9988 13414 10018 13466
rect 10018 13414 10044 13466
rect 9748 13412 9804 13414
rect 9828 13412 9884 13414
rect 9908 13412 9964 13414
rect 9988 13412 10044 13414
rect 15076 13466 15132 13468
rect 15156 13466 15212 13468
rect 15236 13466 15292 13468
rect 15316 13466 15372 13468
rect 15076 13414 15102 13466
rect 15102 13414 15132 13466
rect 15156 13414 15166 13466
rect 15166 13414 15212 13466
rect 15236 13414 15282 13466
rect 15282 13414 15292 13466
rect 15316 13414 15346 13466
rect 15346 13414 15372 13466
rect 15076 13412 15132 13414
rect 15156 13412 15212 13414
rect 15236 13412 15292 13414
rect 15316 13412 15372 13414
rect 7084 12922 7140 12924
rect 7164 12922 7220 12924
rect 7244 12922 7300 12924
rect 7324 12922 7380 12924
rect 7084 12870 7110 12922
rect 7110 12870 7140 12922
rect 7164 12870 7174 12922
rect 7174 12870 7220 12922
rect 7244 12870 7290 12922
rect 7290 12870 7300 12922
rect 7324 12870 7354 12922
rect 7354 12870 7380 12922
rect 7084 12868 7140 12870
rect 7164 12868 7220 12870
rect 7244 12868 7300 12870
rect 7324 12868 7380 12870
rect 12412 12922 12468 12924
rect 12492 12922 12548 12924
rect 12572 12922 12628 12924
rect 12652 12922 12708 12924
rect 12412 12870 12438 12922
rect 12438 12870 12468 12922
rect 12492 12870 12502 12922
rect 12502 12870 12548 12922
rect 12572 12870 12618 12922
rect 12618 12870 12628 12922
rect 12652 12870 12682 12922
rect 12682 12870 12708 12922
rect 12412 12868 12468 12870
rect 12492 12868 12548 12870
rect 12572 12868 12628 12870
rect 12652 12868 12708 12870
rect 17740 12922 17796 12924
rect 17820 12922 17876 12924
rect 17900 12922 17956 12924
rect 17980 12922 18036 12924
rect 17740 12870 17766 12922
rect 17766 12870 17796 12922
rect 17820 12870 17830 12922
rect 17830 12870 17876 12922
rect 17900 12870 17946 12922
rect 17946 12870 17956 12922
rect 17980 12870 18010 12922
rect 18010 12870 18036 12922
rect 17740 12868 17796 12870
rect 17820 12868 17876 12870
rect 17900 12868 17956 12870
rect 17980 12868 18036 12870
rect 4420 12378 4476 12380
rect 4500 12378 4556 12380
rect 4580 12378 4636 12380
rect 4660 12378 4716 12380
rect 4420 12326 4446 12378
rect 4446 12326 4476 12378
rect 4500 12326 4510 12378
rect 4510 12326 4556 12378
rect 4580 12326 4626 12378
rect 4626 12326 4636 12378
rect 4660 12326 4690 12378
rect 4690 12326 4716 12378
rect 4420 12324 4476 12326
rect 4500 12324 4556 12326
rect 4580 12324 4636 12326
rect 4660 12324 4716 12326
rect 9748 12378 9804 12380
rect 9828 12378 9884 12380
rect 9908 12378 9964 12380
rect 9988 12378 10044 12380
rect 9748 12326 9774 12378
rect 9774 12326 9804 12378
rect 9828 12326 9838 12378
rect 9838 12326 9884 12378
rect 9908 12326 9954 12378
rect 9954 12326 9964 12378
rect 9988 12326 10018 12378
rect 10018 12326 10044 12378
rect 9748 12324 9804 12326
rect 9828 12324 9884 12326
rect 9908 12324 9964 12326
rect 9988 12324 10044 12326
rect 15076 12378 15132 12380
rect 15156 12378 15212 12380
rect 15236 12378 15292 12380
rect 15316 12378 15372 12380
rect 15076 12326 15102 12378
rect 15102 12326 15132 12378
rect 15156 12326 15166 12378
rect 15166 12326 15212 12378
rect 15236 12326 15282 12378
rect 15282 12326 15292 12378
rect 15316 12326 15346 12378
rect 15346 12326 15372 12378
rect 15076 12324 15132 12326
rect 15156 12324 15212 12326
rect 15236 12324 15292 12326
rect 15316 12324 15372 12326
rect 7084 11834 7140 11836
rect 7164 11834 7220 11836
rect 7244 11834 7300 11836
rect 7324 11834 7380 11836
rect 7084 11782 7110 11834
rect 7110 11782 7140 11834
rect 7164 11782 7174 11834
rect 7174 11782 7220 11834
rect 7244 11782 7290 11834
rect 7290 11782 7300 11834
rect 7324 11782 7354 11834
rect 7354 11782 7380 11834
rect 7084 11780 7140 11782
rect 7164 11780 7220 11782
rect 7244 11780 7300 11782
rect 7324 11780 7380 11782
rect 12412 11834 12468 11836
rect 12492 11834 12548 11836
rect 12572 11834 12628 11836
rect 12652 11834 12708 11836
rect 12412 11782 12438 11834
rect 12438 11782 12468 11834
rect 12492 11782 12502 11834
rect 12502 11782 12548 11834
rect 12572 11782 12618 11834
rect 12618 11782 12628 11834
rect 12652 11782 12682 11834
rect 12682 11782 12708 11834
rect 12412 11780 12468 11782
rect 12492 11780 12548 11782
rect 12572 11780 12628 11782
rect 12652 11780 12708 11782
rect 17740 11834 17796 11836
rect 17820 11834 17876 11836
rect 17900 11834 17956 11836
rect 17980 11834 18036 11836
rect 17740 11782 17766 11834
rect 17766 11782 17796 11834
rect 17820 11782 17830 11834
rect 17830 11782 17876 11834
rect 17900 11782 17946 11834
rect 17946 11782 17956 11834
rect 17980 11782 18010 11834
rect 18010 11782 18036 11834
rect 17740 11780 17796 11782
rect 17820 11780 17876 11782
rect 17900 11780 17956 11782
rect 17980 11780 18036 11782
rect 4420 11290 4476 11292
rect 4500 11290 4556 11292
rect 4580 11290 4636 11292
rect 4660 11290 4716 11292
rect 4420 11238 4446 11290
rect 4446 11238 4476 11290
rect 4500 11238 4510 11290
rect 4510 11238 4556 11290
rect 4580 11238 4626 11290
rect 4626 11238 4636 11290
rect 4660 11238 4690 11290
rect 4690 11238 4716 11290
rect 4420 11236 4476 11238
rect 4500 11236 4556 11238
rect 4580 11236 4636 11238
rect 4660 11236 4716 11238
rect 9748 11290 9804 11292
rect 9828 11290 9884 11292
rect 9908 11290 9964 11292
rect 9988 11290 10044 11292
rect 9748 11238 9774 11290
rect 9774 11238 9804 11290
rect 9828 11238 9838 11290
rect 9838 11238 9884 11290
rect 9908 11238 9954 11290
rect 9954 11238 9964 11290
rect 9988 11238 10018 11290
rect 10018 11238 10044 11290
rect 9748 11236 9804 11238
rect 9828 11236 9884 11238
rect 9908 11236 9964 11238
rect 9988 11236 10044 11238
rect 15076 11290 15132 11292
rect 15156 11290 15212 11292
rect 15236 11290 15292 11292
rect 15316 11290 15372 11292
rect 15076 11238 15102 11290
rect 15102 11238 15132 11290
rect 15156 11238 15166 11290
rect 15166 11238 15212 11290
rect 15236 11238 15282 11290
rect 15282 11238 15292 11290
rect 15316 11238 15346 11290
rect 15346 11238 15372 11290
rect 15076 11236 15132 11238
rect 15156 11236 15212 11238
rect 15236 11236 15292 11238
rect 15316 11236 15372 11238
rect 7084 10746 7140 10748
rect 7164 10746 7220 10748
rect 7244 10746 7300 10748
rect 7324 10746 7380 10748
rect 7084 10694 7110 10746
rect 7110 10694 7140 10746
rect 7164 10694 7174 10746
rect 7174 10694 7220 10746
rect 7244 10694 7290 10746
rect 7290 10694 7300 10746
rect 7324 10694 7354 10746
rect 7354 10694 7380 10746
rect 7084 10692 7140 10694
rect 7164 10692 7220 10694
rect 7244 10692 7300 10694
rect 7324 10692 7380 10694
rect 12412 10746 12468 10748
rect 12492 10746 12548 10748
rect 12572 10746 12628 10748
rect 12652 10746 12708 10748
rect 12412 10694 12438 10746
rect 12438 10694 12468 10746
rect 12492 10694 12502 10746
rect 12502 10694 12548 10746
rect 12572 10694 12618 10746
rect 12618 10694 12628 10746
rect 12652 10694 12682 10746
rect 12682 10694 12708 10746
rect 12412 10692 12468 10694
rect 12492 10692 12548 10694
rect 12572 10692 12628 10694
rect 12652 10692 12708 10694
rect 17740 10746 17796 10748
rect 17820 10746 17876 10748
rect 17900 10746 17956 10748
rect 17980 10746 18036 10748
rect 17740 10694 17766 10746
rect 17766 10694 17796 10746
rect 17820 10694 17830 10746
rect 17830 10694 17876 10746
rect 17900 10694 17946 10746
rect 17946 10694 17956 10746
rect 17980 10694 18010 10746
rect 18010 10694 18036 10746
rect 17740 10692 17796 10694
rect 17820 10692 17876 10694
rect 17900 10692 17956 10694
rect 17980 10692 18036 10694
rect 4420 10202 4476 10204
rect 4500 10202 4556 10204
rect 4580 10202 4636 10204
rect 4660 10202 4716 10204
rect 4420 10150 4446 10202
rect 4446 10150 4476 10202
rect 4500 10150 4510 10202
rect 4510 10150 4556 10202
rect 4580 10150 4626 10202
rect 4626 10150 4636 10202
rect 4660 10150 4690 10202
rect 4690 10150 4716 10202
rect 4420 10148 4476 10150
rect 4500 10148 4556 10150
rect 4580 10148 4636 10150
rect 4660 10148 4716 10150
rect 9748 10202 9804 10204
rect 9828 10202 9884 10204
rect 9908 10202 9964 10204
rect 9988 10202 10044 10204
rect 9748 10150 9774 10202
rect 9774 10150 9804 10202
rect 9828 10150 9838 10202
rect 9838 10150 9884 10202
rect 9908 10150 9954 10202
rect 9954 10150 9964 10202
rect 9988 10150 10018 10202
rect 10018 10150 10044 10202
rect 9748 10148 9804 10150
rect 9828 10148 9884 10150
rect 9908 10148 9964 10150
rect 9988 10148 10044 10150
rect 15076 10202 15132 10204
rect 15156 10202 15212 10204
rect 15236 10202 15292 10204
rect 15316 10202 15372 10204
rect 15076 10150 15102 10202
rect 15102 10150 15132 10202
rect 15156 10150 15166 10202
rect 15166 10150 15212 10202
rect 15236 10150 15282 10202
rect 15282 10150 15292 10202
rect 15316 10150 15346 10202
rect 15346 10150 15372 10202
rect 15076 10148 15132 10150
rect 15156 10148 15212 10150
rect 15236 10148 15292 10150
rect 15316 10148 15372 10150
rect 7084 9658 7140 9660
rect 7164 9658 7220 9660
rect 7244 9658 7300 9660
rect 7324 9658 7380 9660
rect 7084 9606 7110 9658
rect 7110 9606 7140 9658
rect 7164 9606 7174 9658
rect 7174 9606 7220 9658
rect 7244 9606 7290 9658
rect 7290 9606 7300 9658
rect 7324 9606 7354 9658
rect 7354 9606 7380 9658
rect 7084 9604 7140 9606
rect 7164 9604 7220 9606
rect 7244 9604 7300 9606
rect 7324 9604 7380 9606
rect 12412 9658 12468 9660
rect 12492 9658 12548 9660
rect 12572 9658 12628 9660
rect 12652 9658 12708 9660
rect 12412 9606 12438 9658
rect 12438 9606 12468 9658
rect 12492 9606 12502 9658
rect 12502 9606 12548 9658
rect 12572 9606 12618 9658
rect 12618 9606 12628 9658
rect 12652 9606 12682 9658
rect 12682 9606 12708 9658
rect 12412 9604 12468 9606
rect 12492 9604 12548 9606
rect 12572 9604 12628 9606
rect 12652 9604 12708 9606
rect 17740 9658 17796 9660
rect 17820 9658 17876 9660
rect 17900 9658 17956 9660
rect 17980 9658 18036 9660
rect 17740 9606 17766 9658
rect 17766 9606 17796 9658
rect 17820 9606 17830 9658
rect 17830 9606 17876 9658
rect 17900 9606 17946 9658
rect 17946 9606 17956 9658
rect 17980 9606 18010 9658
rect 18010 9606 18036 9658
rect 17740 9604 17796 9606
rect 17820 9604 17876 9606
rect 17900 9604 17956 9606
rect 17980 9604 18036 9606
rect 4420 9114 4476 9116
rect 4500 9114 4556 9116
rect 4580 9114 4636 9116
rect 4660 9114 4716 9116
rect 4420 9062 4446 9114
rect 4446 9062 4476 9114
rect 4500 9062 4510 9114
rect 4510 9062 4556 9114
rect 4580 9062 4626 9114
rect 4626 9062 4636 9114
rect 4660 9062 4690 9114
rect 4690 9062 4716 9114
rect 4420 9060 4476 9062
rect 4500 9060 4556 9062
rect 4580 9060 4636 9062
rect 4660 9060 4716 9062
rect 9748 9114 9804 9116
rect 9828 9114 9884 9116
rect 9908 9114 9964 9116
rect 9988 9114 10044 9116
rect 9748 9062 9774 9114
rect 9774 9062 9804 9114
rect 9828 9062 9838 9114
rect 9838 9062 9884 9114
rect 9908 9062 9954 9114
rect 9954 9062 9964 9114
rect 9988 9062 10018 9114
rect 10018 9062 10044 9114
rect 9748 9060 9804 9062
rect 9828 9060 9884 9062
rect 9908 9060 9964 9062
rect 9988 9060 10044 9062
rect 15076 9114 15132 9116
rect 15156 9114 15212 9116
rect 15236 9114 15292 9116
rect 15316 9114 15372 9116
rect 15076 9062 15102 9114
rect 15102 9062 15132 9114
rect 15156 9062 15166 9114
rect 15166 9062 15212 9114
rect 15236 9062 15282 9114
rect 15282 9062 15292 9114
rect 15316 9062 15346 9114
rect 15346 9062 15372 9114
rect 15076 9060 15132 9062
rect 15156 9060 15212 9062
rect 15236 9060 15292 9062
rect 15316 9060 15372 9062
rect 2474 8720 2530 8776
rect 7084 8570 7140 8572
rect 7164 8570 7220 8572
rect 7244 8570 7300 8572
rect 7324 8570 7380 8572
rect 7084 8518 7110 8570
rect 7110 8518 7140 8570
rect 7164 8518 7174 8570
rect 7174 8518 7220 8570
rect 7244 8518 7290 8570
rect 7290 8518 7300 8570
rect 7324 8518 7354 8570
rect 7354 8518 7380 8570
rect 7084 8516 7140 8518
rect 7164 8516 7220 8518
rect 7244 8516 7300 8518
rect 7324 8516 7380 8518
rect 12412 8570 12468 8572
rect 12492 8570 12548 8572
rect 12572 8570 12628 8572
rect 12652 8570 12708 8572
rect 12412 8518 12438 8570
rect 12438 8518 12468 8570
rect 12492 8518 12502 8570
rect 12502 8518 12548 8570
rect 12572 8518 12618 8570
rect 12618 8518 12628 8570
rect 12652 8518 12682 8570
rect 12682 8518 12708 8570
rect 12412 8516 12468 8518
rect 12492 8516 12548 8518
rect 12572 8516 12628 8518
rect 12652 8516 12708 8518
rect 17740 8570 17796 8572
rect 17820 8570 17876 8572
rect 17900 8570 17956 8572
rect 17980 8570 18036 8572
rect 17740 8518 17766 8570
rect 17766 8518 17796 8570
rect 17820 8518 17830 8570
rect 17830 8518 17876 8570
rect 17900 8518 17946 8570
rect 17946 8518 17956 8570
rect 17980 8518 18010 8570
rect 18010 8518 18036 8570
rect 17740 8516 17796 8518
rect 17820 8516 17876 8518
rect 17900 8516 17956 8518
rect 17980 8516 18036 8518
rect 4420 8026 4476 8028
rect 4500 8026 4556 8028
rect 4580 8026 4636 8028
rect 4660 8026 4716 8028
rect 4420 7974 4446 8026
rect 4446 7974 4476 8026
rect 4500 7974 4510 8026
rect 4510 7974 4556 8026
rect 4580 7974 4626 8026
rect 4626 7974 4636 8026
rect 4660 7974 4690 8026
rect 4690 7974 4716 8026
rect 4420 7972 4476 7974
rect 4500 7972 4556 7974
rect 4580 7972 4636 7974
rect 4660 7972 4716 7974
rect 9748 8026 9804 8028
rect 9828 8026 9884 8028
rect 9908 8026 9964 8028
rect 9988 8026 10044 8028
rect 9748 7974 9774 8026
rect 9774 7974 9804 8026
rect 9828 7974 9838 8026
rect 9838 7974 9884 8026
rect 9908 7974 9954 8026
rect 9954 7974 9964 8026
rect 9988 7974 10018 8026
rect 10018 7974 10044 8026
rect 9748 7972 9804 7974
rect 9828 7972 9884 7974
rect 9908 7972 9964 7974
rect 9988 7972 10044 7974
rect 15076 8026 15132 8028
rect 15156 8026 15212 8028
rect 15236 8026 15292 8028
rect 15316 8026 15372 8028
rect 15076 7974 15102 8026
rect 15102 7974 15132 8026
rect 15156 7974 15166 8026
rect 15166 7974 15212 8026
rect 15236 7974 15282 8026
rect 15282 7974 15292 8026
rect 15316 7974 15346 8026
rect 15346 7974 15372 8026
rect 15076 7972 15132 7974
rect 15156 7972 15212 7974
rect 15236 7972 15292 7974
rect 15316 7972 15372 7974
rect 7084 7482 7140 7484
rect 7164 7482 7220 7484
rect 7244 7482 7300 7484
rect 7324 7482 7380 7484
rect 7084 7430 7110 7482
rect 7110 7430 7140 7482
rect 7164 7430 7174 7482
rect 7174 7430 7220 7482
rect 7244 7430 7290 7482
rect 7290 7430 7300 7482
rect 7324 7430 7354 7482
rect 7354 7430 7380 7482
rect 7084 7428 7140 7430
rect 7164 7428 7220 7430
rect 7244 7428 7300 7430
rect 7324 7428 7380 7430
rect 12412 7482 12468 7484
rect 12492 7482 12548 7484
rect 12572 7482 12628 7484
rect 12652 7482 12708 7484
rect 12412 7430 12438 7482
rect 12438 7430 12468 7482
rect 12492 7430 12502 7482
rect 12502 7430 12548 7482
rect 12572 7430 12618 7482
rect 12618 7430 12628 7482
rect 12652 7430 12682 7482
rect 12682 7430 12708 7482
rect 12412 7428 12468 7430
rect 12492 7428 12548 7430
rect 12572 7428 12628 7430
rect 12652 7428 12708 7430
rect 17740 7482 17796 7484
rect 17820 7482 17876 7484
rect 17900 7482 17956 7484
rect 17980 7482 18036 7484
rect 17740 7430 17766 7482
rect 17766 7430 17796 7482
rect 17820 7430 17830 7482
rect 17830 7430 17876 7482
rect 17900 7430 17946 7482
rect 17946 7430 17956 7482
rect 17980 7430 18010 7482
rect 18010 7430 18036 7482
rect 17740 7428 17796 7430
rect 17820 7428 17876 7430
rect 17900 7428 17956 7430
rect 17980 7428 18036 7430
rect 4420 6938 4476 6940
rect 4500 6938 4556 6940
rect 4580 6938 4636 6940
rect 4660 6938 4716 6940
rect 4420 6886 4446 6938
rect 4446 6886 4476 6938
rect 4500 6886 4510 6938
rect 4510 6886 4556 6938
rect 4580 6886 4626 6938
rect 4626 6886 4636 6938
rect 4660 6886 4690 6938
rect 4690 6886 4716 6938
rect 4420 6884 4476 6886
rect 4500 6884 4556 6886
rect 4580 6884 4636 6886
rect 4660 6884 4716 6886
rect 9748 6938 9804 6940
rect 9828 6938 9884 6940
rect 9908 6938 9964 6940
rect 9988 6938 10044 6940
rect 9748 6886 9774 6938
rect 9774 6886 9804 6938
rect 9828 6886 9838 6938
rect 9838 6886 9884 6938
rect 9908 6886 9954 6938
rect 9954 6886 9964 6938
rect 9988 6886 10018 6938
rect 10018 6886 10044 6938
rect 9748 6884 9804 6886
rect 9828 6884 9884 6886
rect 9908 6884 9964 6886
rect 9988 6884 10044 6886
rect 15076 6938 15132 6940
rect 15156 6938 15212 6940
rect 15236 6938 15292 6940
rect 15316 6938 15372 6940
rect 15076 6886 15102 6938
rect 15102 6886 15132 6938
rect 15156 6886 15166 6938
rect 15166 6886 15212 6938
rect 15236 6886 15282 6938
rect 15282 6886 15292 6938
rect 15316 6886 15346 6938
rect 15346 6886 15372 6938
rect 15076 6884 15132 6886
rect 15156 6884 15212 6886
rect 15236 6884 15292 6886
rect 15316 6884 15372 6886
rect 7084 6394 7140 6396
rect 7164 6394 7220 6396
rect 7244 6394 7300 6396
rect 7324 6394 7380 6396
rect 7084 6342 7110 6394
rect 7110 6342 7140 6394
rect 7164 6342 7174 6394
rect 7174 6342 7220 6394
rect 7244 6342 7290 6394
rect 7290 6342 7300 6394
rect 7324 6342 7354 6394
rect 7354 6342 7380 6394
rect 7084 6340 7140 6342
rect 7164 6340 7220 6342
rect 7244 6340 7300 6342
rect 7324 6340 7380 6342
rect 12412 6394 12468 6396
rect 12492 6394 12548 6396
rect 12572 6394 12628 6396
rect 12652 6394 12708 6396
rect 12412 6342 12438 6394
rect 12438 6342 12468 6394
rect 12492 6342 12502 6394
rect 12502 6342 12548 6394
rect 12572 6342 12618 6394
rect 12618 6342 12628 6394
rect 12652 6342 12682 6394
rect 12682 6342 12708 6394
rect 12412 6340 12468 6342
rect 12492 6340 12548 6342
rect 12572 6340 12628 6342
rect 12652 6340 12708 6342
rect 17740 6394 17796 6396
rect 17820 6394 17876 6396
rect 17900 6394 17956 6396
rect 17980 6394 18036 6396
rect 17740 6342 17766 6394
rect 17766 6342 17796 6394
rect 17820 6342 17830 6394
rect 17830 6342 17876 6394
rect 17900 6342 17946 6394
rect 17946 6342 17956 6394
rect 17980 6342 18010 6394
rect 18010 6342 18036 6394
rect 17740 6340 17796 6342
rect 17820 6340 17876 6342
rect 17900 6340 17956 6342
rect 17980 6340 18036 6342
rect 4420 5850 4476 5852
rect 4500 5850 4556 5852
rect 4580 5850 4636 5852
rect 4660 5850 4716 5852
rect 4420 5798 4446 5850
rect 4446 5798 4476 5850
rect 4500 5798 4510 5850
rect 4510 5798 4556 5850
rect 4580 5798 4626 5850
rect 4626 5798 4636 5850
rect 4660 5798 4690 5850
rect 4690 5798 4716 5850
rect 4420 5796 4476 5798
rect 4500 5796 4556 5798
rect 4580 5796 4636 5798
rect 4660 5796 4716 5798
rect 9748 5850 9804 5852
rect 9828 5850 9884 5852
rect 9908 5850 9964 5852
rect 9988 5850 10044 5852
rect 9748 5798 9774 5850
rect 9774 5798 9804 5850
rect 9828 5798 9838 5850
rect 9838 5798 9884 5850
rect 9908 5798 9954 5850
rect 9954 5798 9964 5850
rect 9988 5798 10018 5850
rect 10018 5798 10044 5850
rect 9748 5796 9804 5798
rect 9828 5796 9884 5798
rect 9908 5796 9964 5798
rect 9988 5796 10044 5798
rect 15076 5850 15132 5852
rect 15156 5850 15212 5852
rect 15236 5850 15292 5852
rect 15316 5850 15372 5852
rect 15076 5798 15102 5850
rect 15102 5798 15132 5850
rect 15156 5798 15166 5850
rect 15166 5798 15212 5850
rect 15236 5798 15282 5850
rect 15282 5798 15292 5850
rect 15316 5798 15346 5850
rect 15346 5798 15372 5850
rect 15076 5796 15132 5798
rect 15156 5796 15212 5798
rect 15236 5796 15292 5798
rect 15316 5796 15372 5798
rect 7084 5306 7140 5308
rect 7164 5306 7220 5308
rect 7244 5306 7300 5308
rect 7324 5306 7380 5308
rect 7084 5254 7110 5306
rect 7110 5254 7140 5306
rect 7164 5254 7174 5306
rect 7174 5254 7220 5306
rect 7244 5254 7290 5306
rect 7290 5254 7300 5306
rect 7324 5254 7354 5306
rect 7354 5254 7380 5306
rect 7084 5252 7140 5254
rect 7164 5252 7220 5254
rect 7244 5252 7300 5254
rect 7324 5252 7380 5254
rect 12412 5306 12468 5308
rect 12492 5306 12548 5308
rect 12572 5306 12628 5308
rect 12652 5306 12708 5308
rect 12412 5254 12438 5306
rect 12438 5254 12468 5306
rect 12492 5254 12502 5306
rect 12502 5254 12548 5306
rect 12572 5254 12618 5306
rect 12618 5254 12628 5306
rect 12652 5254 12682 5306
rect 12682 5254 12708 5306
rect 12412 5252 12468 5254
rect 12492 5252 12548 5254
rect 12572 5252 12628 5254
rect 12652 5252 12708 5254
rect 17740 5306 17796 5308
rect 17820 5306 17876 5308
rect 17900 5306 17956 5308
rect 17980 5306 18036 5308
rect 17740 5254 17766 5306
rect 17766 5254 17796 5306
rect 17820 5254 17830 5306
rect 17830 5254 17876 5306
rect 17900 5254 17946 5306
rect 17946 5254 17956 5306
rect 17980 5254 18010 5306
rect 18010 5254 18036 5306
rect 17740 5252 17796 5254
rect 17820 5252 17876 5254
rect 17900 5252 17956 5254
rect 17980 5252 18036 5254
rect 4420 4762 4476 4764
rect 4500 4762 4556 4764
rect 4580 4762 4636 4764
rect 4660 4762 4716 4764
rect 4420 4710 4446 4762
rect 4446 4710 4476 4762
rect 4500 4710 4510 4762
rect 4510 4710 4556 4762
rect 4580 4710 4626 4762
rect 4626 4710 4636 4762
rect 4660 4710 4690 4762
rect 4690 4710 4716 4762
rect 4420 4708 4476 4710
rect 4500 4708 4556 4710
rect 4580 4708 4636 4710
rect 4660 4708 4716 4710
rect 9748 4762 9804 4764
rect 9828 4762 9884 4764
rect 9908 4762 9964 4764
rect 9988 4762 10044 4764
rect 9748 4710 9774 4762
rect 9774 4710 9804 4762
rect 9828 4710 9838 4762
rect 9838 4710 9884 4762
rect 9908 4710 9954 4762
rect 9954 4710 9964 4762
rect 9988 4710 10018 4762
rect 10018 4710 10044 4762
rect 9748 4708 9804 4710
rect 9828 4708 9884 4710
rect 9908 4708 9964 4710
rect 9988 4708 10044 4710
rect 15076 4762 15132 4764
rect 15156 4762 15212 4764
rect 15236 4762 15292 4764
rect 15316 4762 15372 4764
rect 15076 4710 15102 4762
rect 15102 4710 15132 4762
rect 15156 4710 15166 4762
rect 15166 4710 15212 4762
rect 15236 4710 15282 4762
rect 15282 4710 15292 4762
rect 15316 4710 15346 4762
rect 15346 4710 15372 4762
rect 15076 4708 15132 4710
rect 15156 4708 15212 4710
rect 15236 4708 15292 4710
rect 15316 4708 15372 4710
rect 7084 4218 7140 4220
rect 7164 4218 7220 4220
rect 7244 4218 7300 4220
rect 7324 4218 7380 4220
rect 7084 4166 7110 4218
rect 7110 4166 7140 4218
rect 7164 4166 7174 4218
rect 7174 4166 7220 4218
rect 7244 4166 7290 4218
rect 7290 4166 7300 4218
rect 7324 4166 7354 4218
rect 7354 4166 7380 4218
rect 7084 4164 7140 4166
rect 7164 4164 7220 4166
rect 7244 4164 7300 4166
rect 7324 4164 7380 4166
rect 12412 4218 12468 4220
rect 12492 4218 12548 4220
rect 12572 4218 12628 4220
rect 12652 4218 12708 4220
rect 12412 4166 12438 4218
rect 12438 4166 12468 4218
rect 12492 4166 12502 4218
rect 12502 4166 12548 4218
rect 12572 4166 12618 4218
rect 12618 4166 12628 4218
rect 12652 4166 12682 4218
rect 12682 4166 12708 4218
rect 12412 4164 12468 4166
rect 12492 4164 12548 4166
rect 12572 4164 12628 4166
rect 12652 4164 12708 4166
rect 17740 4218 17796 4220
rect 17820 4218 17876 4220
rect 17900 4218 17956 4220
rect 17980 4218 18036 4220
rect 17740 4166 17766 4218
rect 17766 4166 17796 4218
rect 17820 4166 17830 4218
rect 17830 4166 17876 4218
rect 17900 4166 17946 4218
rect 17946 4166 17956 4218
rect 17980 4166 18010 4218
rect 18010 4166 18036 4218
rect 17740 4164 17796 4166
rect 17820 4164 17876 4166
rect 17900 4164 17956 4166
rect 17980 4164 18036 4166
rect 4420 3674 4476 3676
rect 4500 3674 4556 3676
rect 4580 3674 4636 3676
rect 4660 3674 4716 3676
rect 4420 3622 4446 3674
rect 4446 3622 4476 3674
rect 4500 3622 4510 3674
rect 4510 3622 4556 3674
rect 4580 3622 4626 3674
rect 4626 3622 4636 3674
rect 4660 3622 4690 3674
rect 4690 3622 4716 3674
rect 4420 3620 4476 3622
rect 4500 3620 4556 3622
rect 4580 3620 4636 3622
rect 4660 3620 4716 3622
rect 9748 3674 9804 3676
rect 9828 3674 9884 3676
rect 9908 3674 9964 3676
rect 9988 3674 10044 3676
rect 9748 3622 9774 3674
rect 9774 3622 9804 3674
rect 9828 3622 9838 3674
rect 9838 3622 9884 3674
rect 9908 3622 9954 3674
rect 9954 3622 9964 3674
rect 9988 3622 10018 3674
rect 10018 3622 10044 3674
rect 9748 3620 9804 3622
rect 9828 3620 9884 3622
rect 9908 3620 9964 3622
rect 9988 3620 10044 3622
rect 15076 3674 15132 3676
rect 15156 3674 15212 3676
rect 15236 3674 15292 3676
rect 15316 3674 15372 3676
rect 15076 3622 15102 3674
rect 15102 3622 15132 3674
rect 15156 3622 15166 3674
rect 15166 3622 15212 3674
rect 15236 3622 15282 3674
rect 15282 3622 15292 3674
rect 15316 3622 15346 3674
rect 15346 3622 15372 3674
rect 15076 3620 15132 3622
rect 15156 3620 15212 3622
rect 15236 3620 15292 3622
rect 15316 3620 15372 3622
rect 7084 3130 7140 3132
rect 7164 3130 7220 3132
rect 7244 3130 7300 3132
rect 7324 3130 7380 3132
rect 7084 3078 7110 3130
rect 7110 3078 7140 3130
rect 7164 3078 7174 3130
rect 7174 3078 7220 3130
rect 7244 3078 7290 3130
rect 7290 3078 7300 3130
rect 7324 3078 7354 3130
rect 7354 3078 7380 3130
rect 7084 3076 7140 3078
rect 7164 3076 7220 3078
rect 7244 3076 7300 3078
rect 7324 3076 7380 3078
rect 12412 3130 12468 3132
rect 12492 3130 12548 3132
rect 12572 3130 12628 3132
rect 12652 3130 12708 3132
rect 12412 3078 12438 3130
rect 12438 3078 12468 3130
rect 12492 3078 12502 3130
rect 12502 3078 12548 3130
rect 12572 3078 12618 3130
rect 12618 3078 12628 3130
rect 12652 3078 12682 3130
rect 12682 3078 12708 3130
rect 12412 3076 12468 3078
rect 12492 3076 12548 3078
rect 12572 3076 12628 3078
rect 12652 3076 12708 3078
rect 17740 3130 17796 3132
rect 17820 3130 17876 3132
rect 17900 3130 17956 3132
rect 17980 3130 18036 3132
rect 17740 3078 17766 3130
rect 17766 3078 17796 3130
rect 17820 3078 17830 3130
rect 17830 3078 17876 3130
rect 17900 3078 17946 3130
rect 17946 3078 17956 3130
rect 17980 3078 18010 3130
rect 18010 3078 18036 3130
rect 17740 3076 17796 3078
rect 17820 3076 17876 3078
rect 17900 3076 17956 3078
rect 17980 3076 18036 3078
rect 4420 2586 4476 2588
rect 4500 2586 4556 2588
rect 4580 2586 4636 2588
rect 4660 2586 4716 2588
rect 4420 2534 4446 2586
rect 4446 2534 4476 2586
rect 4500 2534 4510 2586
rect 4510 2534 4556 2586
rect 4580 2534 4626 2586
rect 4626 2534 4636 2586
rect 4660 2534 4690 2586
rect 4690 2534 4716 2586
rect 4420 2532 4476 2534
rect 4500 2532 4556 2534
rect 4580 2532 4636 2534
rect 4660 2532 4716 2534
rect 9748 2586 9804 2588
rect 9828 2586 9884 2588
rect 9908 2586 9964 2588
rect 9988 2586 10044 2588
rect 9748 2534 9774 2586
rect 9774 2534 9804 2586
rect 9828 2534 9838 2586
rect 9838 2534 9884 2586
rect 9908 2534 9954 2586
rect 9954 2534 9964 2586
rect 9988 2534 10018 2586
rect 10018 2534 10044 2586
rect 9748 2532 9804 2534
rect 9828 2532 9884 2534
rect 9908 2532 9964 2534
rect 9988 2532 10044 2534
rect 15076 2586 15132 2588
rect 15156 2586 15212 2588
rect 15236 2586 15292 2588
rect 15316 2586 15372 2588
rect 15076 2534 15102 2586
rect 15102 2534 15132 2586
rect 15156 2534 15166 2586
rect 15166 2534 15212 2586
rect 15236 2534 15282 2586
rect 15282 2534 15292 2586
rect 15316 2534 15346 2586
rect 15346 2534 15372 2586
rect 15076 2532 15132 2534
rect 15156 2532 15212 2534
rect 15236 2532 15292 2534
rect 15316 2532 15372 2534
rect 7084 2042 7140 2044
rect 7164 2042 7220 2044
rect 7244 2042 7300 2044
rect 7324 2042 7380 2044
rect 7084 1990 7110 2042
rect 7110 1990 7140 2042
rect 7164 1990 7174 2042
rect 7174 1990 7220 2042
rect 7244 1990 7290 2042
rect 7290 1990 7300 2042
rect 7324 1990 7354 2042
rect 7354 1990 7380 2042
rect 7084 1988 7140 1990
rect 7164 1988 7220 1990
rect 7244 1988 7300 1990
rect 7324 1988 7380 1990
rect 12412 2042 12468 2044
rect 12492 2042 12548 2044
rect 12572 2042 12628 2044
rect 12652 2042 12708 2044
rect 12412 1990 12438 2042
rect 12438 1990 12468 2042
rect 12492 1990 12502 2042
rect 12502 1990 12548 2042
rect 12572 1990 12618 2042
rect 12618 1990 12628 2042
rect 12652 1990 12682 2042
rect 12682 1990 12708 2042
rect 12412 1988 12468 1990
rect 12492 1988 12548 1990
rect 12572 1988 12628 1990
rect 12652 1988 12708 1990
rect 17740 2042 17796 2044
rect 17820 2042 17876 2044
rect 17900 2042 17956 2044
rect 17980 2042 18036 2044
rect 17740 1990 17766 2042
rect 17766 1990 17796 2042
rect 17820 1990 17830 2042
rect 17830 1990 17876 2042
rect 17900 1990 17946 2042
rect 17946 1990 17956 2042
rect 17980 1990 18010 2042
rect 18010 1990 18036 2042
rect 17740 1988 17796 1990
rect 17820 1988 17876 1990
rect 17900 1988 17956 1990
rect 17980 1988 18036 1990
rect 4420 1498 4476 1500
rect 4500 1498 4556 1500
rect 4580 1498 4636 1500
rect 4660 1498 4716 1500
rect 4420 1446 4446 1498
rect 4446 1446 4476 1498
rect 4500 1446 4510 1498
rect 4510 1446 4556 1498
rect 4580 1446 4626 1498
rect 4626 1446 4636 1498
rect 4660 1446 4690 1498
rect 4690 1446 4716 1498
rect 4420 1444 4476 1446
rect 4500 1444 4556 1446
rect 4580 1444 4636 1446
rect 4660 1444 4716 1446
rect 9748 1498 9804 1500
rect 9828 1498 9884 1500
rect 9908 1498 9964 1500
rect 9988 1498 10044 1500
rect 9748 1446 9774 1498
rect 9774 1446 9804 1498
rect 9828 1446 9838 1498
rect 9838 1446 9884 1498
rect 9908 1446 9954 1498
rect 9954 1446 9964 1498
rect 9988 1446 10018 1498
rect 10018 1446 10044 1498
rect 9748 1444 9804 1446
rect 9828 1444 9884 1446
rect 9908 1444 9964 1446
rect 9988 1444 10044 1446
rect 15076 1498 15132 1500
rect 15156 1498 15212 1500
rect 15236 1498 15292 1500
rect 15316 1498 15372 1500
rect 15076 1446 15102 1498
rect 15102 1446 15132 1498
rect 15156 1446 15166 1498
rect 15166 1446 15212 1498
rect 15236 1446 15282 1498
rect 15282 1446 15292 1498
rect 15316 1446 15346 1498
rect 15346 1446 15372 1498
rect 15076 1444 15132 1446
rect 15156 1444 15212 1446
rect 15236 1444 15292 1446
rect 15316 1444 15372 1446
rect 2290 1104 2346 1160
rect 2934 1104 2990 1160
rect 7084 954 7140 956
rect 7164 954 7220 956
rect 7244 954 7300 956
rect 7324 954 7380 956
rect 7084 902 7110 954
rect 7110 902 7140 954
rect 7164 902 7174 954
rect 7174 902 7220 954
rect 7244 902 7290 954
rect 7290 902 7300 954
rect 7324 902 7354 954
rect 7354 902 7380 954
rect 7084 900 7140 902
rect 7164 900 7220 902
rect 7244 900 7300 902
rect 7324 900 7380 902
rect 12412 954 12468 956
rect 12492 954 12548 956
rect 12572 954 12628 956
rect 12652 954 12708 956
rect 12412 902 12438 954
rect 12438 902 12468 954
rect 12492 902 12502 954
rect 12502 902 12548 954
rect 12572 902 12618 954
rect 12618 902 12628 954
rect 12652 902 12682 954
rect 12682 902 12708 954
rect 12412 900 12468 902
rect 12492 900 12548 902
rect 12572 900 12628 902
rect 12652 900 12708 902
rect 17740 954 17796 956
rect 17820 954 17876 956
rect 17900 954 17956 956
rect 17980 954 18036 956
rect 17740 902 17766 954
rect 17766 902 17796 954
rect 17820 902 17830 954
rect 17830 902 17876 954
rect 17900 902 17946 954
rect 17946 902 17956 954
rect 17980 902 18010 954
rect 18010 902 18036 954
rect 17740 900 17796 902
rect 17820 900 17876 902
rect 17900 900 17956 902
rect 17980 900 18036 902
<< metal3 >>
rect 1917 22378 1983 22381
rect 830 22376 1983 22378
rect 830 22320 1922 22376
rect 1978 22320 1983 22376
rect 830 22318 1983 22320
rect 830 22136 890 22318
rect 1917 22315 1983 22318
rect 4408 22176 4728 22177
rect 800 22016 920 22136
rect 4408 22112 4416 22176
rect 4480 22112 4496 22176
rect 4560 22112 4576 22176
rect 4640 22112 4656 22176
rect 4720 22112 4728 22176
rect 4408 22111 4728 22112
rect 9736 22176 10056 22177
rect 9736 22112 9744 22176
rect 9808 22112 9824 22176
rect 9888 22112 9904 22176
rect 9968 22112 9984 22176
rect 10048 22112 10056 22176
rect 9736 22111 10056 22112
rect 15064 22176 15384 22177
rect 15064 22112 15072 22176
rect 15136 22112 15152 22176
rect 15216 22112 15232 22176
rect 15296 22112 15312 22176
rect 15376 22112 15384 22176
rect 15064 22111 15384 22112
rect 2469 21834 2535 21837
rect 830 21832 2535 21834
rect 830 21776 2474 21832
rect 2530 21776 2535 21832
rect 830 21774 2535 21776
rect 830 21592 890 21774
rect 2469 21771 2535 21774
rect 7072 21632 7392 21633
rect 800 21472 920 21592
rect 7072 21568 7080 21632
rect 7144 21568 7160 21632
rect 7224 21568 7240 21632
rect 7304 21568 7320 21632
rect 7384 21568 7392 21632
rect 7072 21567 7392 21568
rect 12400 21632 12720 21633
rect 12400 21568 12408 21632
rect 12472 21568 12488 21632
rect 12552 21568 12568 21632
rect 12632 21568 12648 21632
rect 12712 21568 12720 21632
rect 12400 21567 12720 21568
rect 17728 21632 18048 21633
rect 17728 21568 17736 21632
rect 17800 21568 17816 21632
rect 17880 21568 17896 21632
rect 17960 21568 17976 21632
rect 18040 21568 18048 21632
rect 17728 21567 18048 21568
rect 2469 21290 2535 21293
rect 830 21288 2535 21290
rect 830 21232 2474 21288
rect 2530 21232 2535 21288
rect 830 21230 2535 21232
rect 830 21048 890 21230
rect 2469 21227 2535 21230
rect 4408 21088 4728 21089
rect 800 20928 920 21048
rect 4408 21024 4416 21088
rect 4480 21024 4496 21088
rect 4560 21024 4576 21088
rect 4640 21024 4656 21088
rect 4720 21024 4728 21088
rect 4408 21023 4728 21024
rect 9736 21088 10056 21089
rect 9736 21024 9744 21088
rect 9808 21024 9824 21088
rect 9888 21024 9904 21088
rect 9968 21024 9984 21088
rect 10048 21024 10056 21088
rect 9736 21023 10056 21024
rect 15064 21088 15384 21089
rect 15064 21024 15072 21088
rect 15136 21024 15152 21088
rect 15216 21024 15232 21088
rect 15296 21024 15312 21088
rect 15376 21024 15384 21088
rect 15064 21023 15384 21024
rect 7072 20544 7392 20545
rect 7072 20480 7080 20544
rect 7144 20480 7160 20544
rect 7224 20480 7240 20544
rect 7304 20480 7320 20544
rect 7384 20480 7392 20544
rect 7072 20479 7392 20480
rect 12400 20544 12720 20545
rect 12400 20480 12408 20544
rect 12472 20480 12488 20544
rect 12552 20480 12568 20544
rect 12632 20480 12648 20544
rect 12712 20480 12720 20544
rect 12400 20479 12720 20480
rect 17728 20544 18048 20545
rect 17728 20480 17736 20544
rect 17800 20480 17816 20544
rect 17880 20480 17896 20544
rect 17960 20480 17976 20544
rect 18040 20480 18048 20544
rect 17728 20479 18048 20480
rect 2469 20202 2535 20205
rect 830 20200 2535 20202
rect 830 20144 2474 20200
rect 2530 20144 2535 20200
rect 830 20142 2535 20144
rect 830 19960 890 20142
rect 2469 20139 2535 20142
rect 4408 20000 4728 20001
rect 800 19840 920 19960
rect 4408 19936 4416 20000
rect 4480 19936 4496 20000
rect 4560 19936 4576 20000
rect 4640 19936 4656 20000
rect 4720 19936 4728 20000
rect 4408 19935 4728 19936
rect 9736 20000 10056 20001
rect 9736 19936 9744 20000
rect 9808 19936 9824 20000
rect 9888 19936 9904 20000
rect 9968 19936 9984 20000
rect 10048 19936 10056 20000
rect 9736 19935 10056 19936
rect 15064 20000 15384 20001
rect 15064 19936 15072 20000
rect 15136 19936 15152 20000
rect 15216 19936 15232 20000
rect 15296 19936 15312 20000
rect 15376 19936 15384 20000
rect 15064 19935 15384 19936
rect 7072 19456 7392 19457
rect 7072 19392 7080 19456
rect 7144 19392 7160 19456
rect 7224 19392 7240 19456
rect 7304 19392 7320 19456
rect 7384 19392 7392 19456
rect 7072 19391 7392 19392
rect 12400 19456 12720 19457
rect 12400 19392 12408 19456
rect 12472 19392 12488 19456
rect 12552 19392 12568 19456
rect 12632 19392 12648 19456
rect 12712 19392 12720 19456
rect 12400 19391 12720 19392
rect 17728 19456 18048 19457
rect 17728 19392 17736 19456
rect 17800 19392 17816 19456
rect 17880 19392 17896 19456
rect 17960 19392 17976 19456
rect 18040 19392 18048 19456
rect 17728 19391 18048 19392
rect 2469 19114 2535 19117
rect 830 19112 2535 19114
rect 830 19056 2474 19112
rect 2530 19056 2535 19112
rect 830 19054 2535 19056
rect 830 18872 890 19054
rect 2469 19051 2535 19054
rect 4408 18912 4728 18913
rect 800 18752 920 18872
rect 4408 18848 4416 18912
rect 4480 18848 4496 18912
rect 4560 18848 4576 18912
rect 4640 18848 4656 18912
rect 4720 18848 4728 18912
rect 4408 18847 4728 18848
rect 9736 18912 10056 18913
rect 9736 18848 9744 18912
rect 9808 18848 9824 18912
rect 9888 18848 9904 18912
rect 9968 18848 9984 18912
rect 10048 18848 10056 18912
rect 9736 18847 10056 18848
rect 15064 18912 15384 18913
rect 15064 18848 15072 18912
rect 15136 18848 15152 18912
rect 15216 18848 15232 18912
rect 15296 18848 15312 18912
rect 15376 18848 15384 18912
rect 15064 18847 15384 18848
rect 7072 18368 7392 18369
rect 7072 18304 7080 18368
rect 7144 18304 7160 18368
rect 7224 18304 7240 18368
rect 7304 18304 7320 18368
rect 7384 18304 7392 18368
rect 7072 18303 7392 18304
rect 12400 18368 12720 18369
rect 12400 18304 12408 18368
rect 12472 18304 12488 18368
rect 12552 18304 12568 18368
rect 12632 18304 12648 18368
rect 12712 18304 12720 18368
rect 12400 18303 12720 18304
rect 17728 18368 18048 18369
rect 17728 18304 17736 18368
rect 17800 18304 17816 18368
rect 17880 18304 17896 18368
rect 17960 18304 17976 18368
rect 18040 18304 18048 18368
rect 17728 18303 18048 18304
rect 2469 18026 2535 18029
rect 830 18024 2535 18026
rect 830 17968 2474 18024
rect 2530 17968 2535 18024
rect 830 17966 2535 17968
rect 830 17784 890 17966
rect 2469 17963 2535 17966
rect 4408 17824 4728 17825
rect 800 17664 920 17784
rect 4408 17760 4416 17824
rect 4480 17760 4496 17824
rect 4560 17760 4576 17824
rect 4640 17760 4656 17824
rect 4720 17760 4728 17824
rect 4408 17759 4728 17760
rect 9736 17824 10056 17825
rect 9736 17760 9744 17824
rect 9808 17760 9824 17824
rect 9888 17760 9904 17824
rect 9968 17760 9984 17824
rect 10048 17760 10056 17824
rect 9736 17759 10056 17760
rect 15064 17824 15384 17825
rect 15064 17760 15072 17824
rect 15136 17760 15152 17824
rect 15216 17760 15232 17824
rect 15296 17760 15312 17824
rect 15376 17760 15384 17824
rect 15064 17759 15384 17760
rect 7072 17280 7392 17281
rect 7072 17216 7080 17280
rect 7144 17216 7160 17280
rect 7224 17216 7240 17280
rect 7304 17216 7320 17280
rect 7384 17216 7392 17280
rect 7072 17215 7392 17216
rect 12400 17280 12720 17281
rect 12400 17216 12408 17280
rect 12472 17216 12488 17280
rect 12552 17216 12568 17280
rect 12632 17216 12648 17280
rect 12712 17216 12720 17280
rect 12400 17215 12720 17216
rect 17728 17280 18048 17281
rect 17728 17216 17736 17280
rect 17800 17216 17816 17280
rect 17880 17216 17896 17280
rect 17960 17216 17976 17280
rect 18040 17216 18048 17280
rect 17728 17215 18048 17216
rect 4408 16736 4728 16737
rect 800 16576 920 16696
rect 4408 16672 4416 16736
rect 4480 16672 4496 16736
rect 4560 16672 4576 16736
rect 4640 16672 4656 16736
rect 4720 16672 4728 16736
rect 4408 16671 4728 16672
rect 9736 16736 10056 16737
rect 9736 16672 9744 16736
rect 9808 16672 9824 16736
rect 9888 16672 9904 16736
rect 9968 16672 9984 16736
rect 10048 16672 10056 16736
rect 9736 16671 10056 16672
rect 15064 16736 15384 16737
rect 15064 16672 15072 16736
rect 15136 16672 15152 16736
rect 15216 16672 15232 16736
rect 15296 16672 15312 16736
rect 15376 16672 15384 16736
rect 15064 16671 15384 16672
rect 2469 16666 2535 16669
rect 1046 16664 2535 16666
rect 1046 16608 2474 16664
rect 2530 16608 2535 16664
rect 1046 16606 2535 16608
rect 830 16394 890 16576
rect 1046 16394 1106 16606
rect 2469 16603 2535 16606
rect 830 16334 1106 16394
rect 7072 16192 7392 16193
rect 7072 16128 7080 16192
rect 7144 16128 7160 16192
rect 7224 16128 7240 16192
rect 7304 16128 7320 16192
rect 7384 16128 7392 16192
rect 7072 16127 7392 16128
rect 12400 16192 12720 16193
rect 12400 16128 12408 16192
rect 12472 16128 12488 16192
rect 12552 16128 12568 16192
rect 12632 16128 12648 16192
rect 12712 16128 12720 16192
rect 12400 16127 12720 16128
rect 17728 16192 18048 16193
rect 17728 16128 17736 16192
rect 17800 16128 17816 16192
rect 17880 16128 17896 16192
rect 17960 16128 17976 16192
rect 18040 16128 18048 16192
rect 17728 16127 18048 16128
rect 2469 15850 2535 15853
rect 830 15848 2535 15850
rect 830 15792 2474 15848
rect 2530 15792 2535 15848
rect 830 15790 2535 15792
rect 830 15608 890 15790
rect 2469 15787 2535 15790
rect 4408 15648 4728 15649
rect 800 15488 920 15608
rect 4408 15584 4416 15648
rect 4480 15584 4496 15648
rect 4560 15584 4576 15648
rect 4640 15584 4656 15648
rect 4720 15584 4728 15648
rect 4408 15583 4728 15584
rect 9736 15648 10056 15649
rect 9736 15584 9744 15648
rect 9808 15584 9824 15648
rect 9888 15584 9904 15648
rect 9968 15584 9984 15648
rect 10048 15584 10056 15648
rect 9736 15583 10056 15584
rect 15064 15648 15384 15649
rect 15064 15584 15072 15648
rect 15136 15584 15152 15648
rect 15216 15584 15232 15648
rect 15296 15584 15312 15648
rect 15376 15584 15384 15648
rect 15064 15583 15384 15584
rect 7072 15104 7392 15105
rect 7072 15040 7080 15104
rect 7144 15040 7160 15104
rect 7224 15040 7240 15104
rect 7304 15040 7320 15104
rect 7384 15040 7392 15104
rect 7072 15039 7392 15040
rect 12400 15104 12720 15105
rect 12400 15040 12408 15104
rect 12472 15040 12488 15104
rect 12552 15040 12568 15104
rect 12632 15040 12648 15104
rect 12712 15040 12720 15104
rect 12400 15039 12720 15040
rect 17728 15104 18048 15105
rect 17728 15040 17736 15104
rect 17800 15040 17816 15104
rect 17880 15040 17896 15104
rect 17960 15040 17976 15104
rect 18040 15040 18048 15104
rect 17728 15039 18048 15040
rect 4408 14560 4728 14561
rect 4408 14496 4416 14560
rect 4480 14496 4496 14560
rect 4560 14496 4576 14560
rect 4640 14496 4656 14560
rect 4720 14496 4728 14560
rect 4408 14495 4728 14496
rect 9736 14560 10056 14561
rect 9736 14496 9744 14560
rect 9808 14496 9824 14560
rect 9888 14496 9904 14560
rect 9968 14496 9984 14560
rect 10048 14496 10056 14560
rect 9736 14495 10056 14496
rect 15064 14560 15384 14561
rect 15064 14496 15072 14560
rect 15136 14496 15152 14560
rect 15216 14496 15232 14560
rect 15296 14496 15312 14560
rect 15376 14496 15384 14560
rect 15064 14495 15384 14496
rect 7072 14016 7392 14017
rect 7072 13952 7080 14016
rect 7144 13952 7160 14016
rect 7224 13952 7240 14016
rect 7304 13952 7320 14016
rect 7384 13952 7392 14016
rect 7072 13951 7392 13952
rect 12400 14016 12720 14017
rect 12400 13952 12408 14016
rect 12472 13952 12488 14016
rect 12552 13952 12568 14016
rect 12632 13952 12648 14016
rect 12712 13952 12720 14016
rect 12400 13951 12720 13952
rect 17728 14016 18048 14017
rect 17728 13952 17736 14016
rect 17800 13952 17816 14016
rect 17880 13952 17896 14016
rect 17960 13952 17976 14016
rect 18040 13952 18048 14016
rect 17728 13951 18048 13952
rect 2469 13674 2535 13677
rect 830 13672 2535 13674
rect 830 13616 2474 13672
rect 2530 13616 2535 13672
rect 830 13614 2535 13616
rect 830 13432 890 13614
rect 2469 13611 2535 13614
rect 4408 13472 4728 13473
rect 800 13312 920 13432
rect 4408 13408 4416 13472
rect 4480 13408 4496 13472
rect 4560 13408 4576 13472
rect 4640 13408 4656 13472
rect 4720 13408 4728 13472
rect 4408 13407 4728 13408
rect 9736 13472 10056 13473
rect 9736 13408 9744 13472
rect 9808 13408 9824 13472
rect 9888 13408 9904 13472
rect 9968 13408 9984 13472
rect 10048 13408 10056 13472
rect 9736 13407 10056 13408
rect 15064 13472 15384 13473
rect 15064 13408 15072 13472
rect 15136 13408 15152 13472
rect 15216 13408 15232 13472
rect 15296 13408 15312 13472
rect 15376 13408 15384 13472
rect 15064 13407 15384 13408
rect 7072 12928 7392 12929
rect 7072 12864 7080 12928
rect 7144 12864 7160 12928
rect 7224 12864 7240 12928
rect 7304 12864 7320 12928
rect 7384 12864 7392 12928
rect 7072 12863 7392 12864
rect 12400 12928 12720 12929
rect 12400 12864 12408 12928
rect 12472 12864 12488 12928
rect 12552 12864 12568 12928
rect 12632 12864 12648 12928
rect 12712 12864 12720 12928
rect 12400 12863 12720 12864
rect 17728 12928 18048 12929
rect 17728 12864 17736 12928
rect 17800 12864 17816 12928
rect 17880 12864 17896 12928
rect 17960 12864 17976 12928
rect 18040 12864 18048 12928
rect 17728 12863 18048 12864
rect 4408 12384 4728 12385
rect 4408 12320 4416 12384
rect 4480 12320 4496 12384
rect 4560 12320 4576 12384
rect 4640 12320 4656 12384
rect 4720 12320 4728 12384
rect 4408 12319 4728 12320
rect 9736 12384 10056 12385
rect 9736 12320 9744 12384
rect 9808 12320 9824 12384
rect 9888 12320 9904 12384
rect 9968 12320 9984 12384
rect 10048 12320 10056 12384
rect 9736 12319 10056 12320
rect 15064 12384 15384 12385
rect 15064 12320 15072 12384
rect 15136 12320 15152 12384
rect 15216 12320 15232 12384
rect 15296 12320 15312 12384
rect 15376 12320 15384 12384
rect 15064 12319 15384 12320
rect 7072 11840 7392 11841
rect 7072 11776 7080 11840
rect 7144 11776 7160 11840
rect 7224 11776 7240 11840
rect 7304 11776 7320 11840
rect 7384 11776 7392 11840
rect 7072 11775 7392 11776
rect 12400 11840 12720 11841
rect 12400 11776 12408 11840
rect 12472 11776 12488 11840
rect 12552 11776 12568 11840
rect 12632 11776 12648 11840
rect 12712 11776 12720 11840
rect 12400 11775 12720 11776
rect 17728 11840 18048 11841
rect 17728 11776 17736 11840
rect 17800 11776 17816 11840
rect 17880 11776 17896 11840
rect 17960 11776 17976 11840
rect 18040 11776 18048 11840
rect 17728 11775 18048 11776
rect 4408 11296 4728 11297
rect 4408 11232 4416 11296
rect 4480 11232 4496 11296
rect 4560 11232 4576 11296
rect 4640 11232 4656 11296
rect 4720 11232 4728 11296
rect 4408 11231 4728 11232
rect 9736 11296 10056 11297
rect 9736 11232 9744 11296
rect 9808 11232 9824 11296
rect 9888 11232 9904 11296
rect 9968 11232 9984 11296
rect 10048 11232 10056 11296
rect 9736 11231 10056 11232
rect 15064 11296 15384 11297
rect 15064 11232 15072 11296
rect 15136 11232 15152 11296
rect 15216 11232 15232 11296
rect 15296 11232 15312 11296
rect 15376 11232 15384 11296
rect 15064 11231 15384 11232
rect 7072 10752 7392 10753
rect 7072 10688 7080 10752
rect 7144 10688 7160 10752
rect 7224 10688 7240 10752
rect 7304 10688 7320 10752
rect 7384 10688 7392 10752
rect 7072 10687 7392 10688
rect 12400 10752 12720 10753
rect 12400 10688 12408 10752
rect 12472 10688 12488 10752
rect 12552 10688 12568 10752
rect 12632 10688 12648 10752
rect 12712 10688 12720 10752
rect 12400 10687 12720 10688
rect 17728 10752 18048 10753
rect 17728 10688 17736 10752
rect 17800 10688 17816 10752
rect 17880 10688 17896 10752
rect 17960 10688 17976 10752
rect 18040 10688 18048 10752
rect 17728 10687 18048 10688
rect 4408 10208 4728 10209
rect 4408 10144 4416 10208
rect 4480 10144 4496 10208
rect 4560 10144 4576 10208
rect 4640 10144 4656 10208
rect 4720 10144 4728 10208
rect 4408 10143 4728 10144
rect 9736 10208 10056 10209
rect 9736 10144 9744 10208
rect 9808 10144 9824 10208
rect 9888 10144 9904 10208
rect 9968 10144 9984 10208
rect 10048 10144 10056 10208
rect 9736 10143 10056 10144
rect 15064 10208 15384 10209
rect 15064 10144 15072 10208
rect 15136 10144 15152 10208
rect 15216 10144 15232 10208
rect 15296 10144 15312 10208
rect 15376 10144 15384 10208
rect 15064 10143 15384 10144
rect 7072 9664 7392 9665
rect 7072 9600 7080 9664
rect 7144 9600 7160 9664
rect 7224 9600 7240 9664
rect 7304 9600 7320 9664
rect 7384 9600 7392 9664
rect 7072 9599 7392 9600
rect 12400 9664 12720 9665
rect 12400 9600 12408 9664
rect 12472 9600 12488 9664
rect 12552 9600 12568 9664
rect 12632 9600 12648 9664
rect 12712 9600 12720 9664
rect 12400 9599 12720 9600
rect 17728 9664 18048 9665
rect 17728 9600 17736 9664
rect 17800 9600 17816 9664
rect 17880 9600 17896 9664
rect 17960 9600 17976 9664
rect 18040 9600 18048 9664
rect 17728 9599 18048 9600
rect 4408 9120 4728 9121
rect 800 8960 920 9080
rect 4408 9056 4416 9120
rect 4480 9056 4496 9120
rect 4560 9056 4576 9120
rect 4640 9056 4656 9120
rect 4720 9056 4728 9120
rect 4408 9055 4728 9056
rect 9736 9120 10056 9121
rect 9736 9056 9744 9120
rect 9808 9056 9824 9120
rect 9888 9056 9904 9120
rect 9968 9056 9984 9120
rect 10048 9056 10056 9120
rect 9736 9055 10056 9056
rect 15064 9120 15384 9121
rect 15064 9056 15072 9120
rect 15136 9056 15152 9120
rect 15216 9056 15232 9120
rect 15296 9056 15312 9120
rect 15376 9056 15384 9120
rect 15064 9055 15384 9056
rect 830 8778 890 8960
rect 2469 8778 2535 8781
rect 830 8776 2535 8778
rect 830 8720 2474 8776
rect 2530 8720 2535 8776
rect 830 8718 2535 8720
rect 2469 8715 2535 8718
rect 7072 8576 7392 8577
rect 7072 8512 7080 8576
rect 7144 8512 7160 8576
rect 7224 8512 7240 8576
rect 7304 8512 7320 8576
rect 7384 8512 7392 8576
rect 7072 8511 7392 8512
rect 12400 8576 12720 8577
rect 12400 8512 12408 8576
rect 12472 8512 12488 8576
rect 12552 8512 12568 8576
rect 12632 8512 12648 8576
rect 12712 8512 12720 8576
rect 12400 8511 12720 8512
rect 17728 8576 18048 8577
rect 17728 8512 17736 8576
rect 17800 8512 17816 8576
rect 17880 8512 17896 8576
rect 17960 8512 17976 8576
rect 18040 8512 18048 8576
rect 17728 8511 18048 8512
rect 4408 8032 4728 8033
rect 4408 7968 4416 8032
rect 4480 7968 4496 8032
rect 4560 7968 4576 8032
rect 4640 7968 4656 8032
rect 4720 7968 4728 8032
rect 4408 7967 4728 7968
rect 9736 8032 10056 8033
rect 9736 7968 9744 8032
rect 9808 7968 9824 8032
rect 9888 7968 9904 8032
rect 9968 7968 9984 8032
rect 10048 7968 10056 8032
rect 9736 7967 10056 7968
rect 15064 8032 15384 8033
rect 15064 7968 15072 8032
rect 15136 7968 15152 8032
rect 15216 7968 15232 8032
rect 15296 7968 15312 8032
rect 15376 7968 15384 8032
rect 15064 7967 15384 7968
rect 7072 7488 7392 7489
rect 7072 7424 7080 7488
rect 7144 7424 7160 7488
rect 7224 7424 7240 7488
rect 7304 7424 7320 7488
rect 7384 7424 7392 7488
rect 7072 7423 7392 7424
rect 12400 7488 12720 7489
rect 12400 7424 12408 7488
rect 12472 7424 12488 7488
rect 12552 7424 12568 7488
rect 12632 7424 12648 7488
rect 12712 7424 12720 7488
rect 12400 7423 12720 7424
rect 17728 7488 18048 7489
rect 17728 7424 17736 7488
rect 17800 7424 17816 7488
rect 17880 7424 17896 7488
rect 17960 7424 17976 7488
rect 18040 7424 18048 7488
rect 17728 7423 18048 7424
rect 4408 6944 4728 6945
rect 4408 6880 4416 6944
rect 4480 6880 4496 6944
rect 4560 6880 4576 6944
rect 4640 6880 4656 6944
rect 4720 6880 4728 6944
rect 4408 6879 4728 6880
rect 9736 6944 10056 6945
rect 9736 6880 9744 6944
rect 9808 6880 9824 6944
rect 9888 6880 9904 6944
rect 9968 6880 9984 6944
rect 10048 6880 10056 6944
rect 9736 6879 10056 6880
rect 15064 6944 15384 6945
rect 15064 6880 15072 6944
rect 15136 6880 15152 6944
rect 15216 6880 15232 6944
rect 15296 6880 15312 6944
rect 15376 6880 15384 6944
rect 15064 6879 15384 6880
rect 7072 6400 7392 6401
rect 7072 6336 7080 6400
rect 7144 6336 7160 6400
rect 7224 6336 7240 6400
rect 7304 6336 7320 6400
rect 7384 6336 7392 6400
rect 7072 6335 7392 6336
rect 12400 6400 12720 6401
rect 12400 6336 12408 6400
rect 12472 6336 12488 6400
rect 12552 6336 12568 6400
rect 12632 6336 12648 6400
rect 12712 6336 12720 6400
rect 12400 6335 12720 6336
rect 17728 6400 18048 6401
rect 17728 6336 17736 6400
rect 17800 6336 17816 6400
rect 17880 6336 17896 6400
rect 17960 6336 17976 6400
rect 18040 6336 18048 6400
rect 17728 6335 18048 6336
rect 4408 5856 4728 5857
rect 4408 5792 4416 5856
rect 4480 5792 4496 5856
rect 4560 5792 4576 5856
rect 4640 5792 4656 5856
rect 4720 5792 4728 5856
rect 4408 5791 4728 5792
rect 9736 5856 10056 5857
rect 9736 5792 9744 5856
rect 9808 5792 9824 5856
rect 9888 5792 9904 5856
rect 9968 5792 9984 5856
rect 10048 5792 10056 5856
rect 9736 5791 10056 5792
rect 15064 5856 15384 5857
rect 15064 5792 15072 5856
rect 15136 5792 15152 5856
rect 15216 5792 15232 5856
rect 15296 5792 15312 5856
rect 15376 5792 15384 5856
rect 15064 5791 15384 5792
rect 7072 5312 7392 5313
rect 7072 5248 7080 5312
rect 7144 5248 7160 5312
rect 7224 5248 7240 5312
rect 7304 5248 7320 5312
rect 7384 5248 7392 5312
rect 7072 5247 7392 5248
rect 12400 5312 12720 5313
rect 12400 5248 12408 5312
rect 12472 5248 12488 5312
rect 12552 5248 12568 5312
rect 12632 5248 12648 5312
rect 12712 5248 12720 5312
rect 12400 5247 12720 5248
rect 17728 5312 18048 5313
rect 17728 5248 17736 5312
rect 17800 5248 17816 5312
rect 17880 5248 17896 5312
rect 17960 5248 17976 5312
rect 18040 5248 18048 5312
rect 17728 5247 18048 5248
rect 4408 4768 4728 4769
rect 4408 4704 4416 4768
rect 4480 4704 4496 4768
rect 4560 4704 4576 4768
rect 4640 4704 4656 4768
rect 4720 4704 4728 4768
rect 4408 4703 4728 4704
rect 9736 4768 10056 4769
rect 9736 4704 9744 4768
rect 9808 4704 9824 4768
rect 9888 4704 9904 4768
rect 9968 4704 9984 4768
rect 10048 4704 10056 4768
rect 9736 4703 10056 4704
rect 15064 4768 15384 4769
rect 15064 4704 15072 4768
rect 15136 4704 15152 4768
rect 15216 4704 15232 4768
rect 15296 4704 15312 4768
rect 15376 4704 15384 4768
rect 15064 4703 15384 4704
rect 7072 4224 7392 4225
rect 7072 4160 7080 4224
rect 7144 4160 7160 4224
rect 7224 4160 7240 4224
rect 7304 4160 7320 4224
rect 7384 4160 7392 4224
rect 7072 4159 7392 4160
rect 12400 4224 12720 4225
rect 12400 4160 12408 4224
rect 12472 4160 12488 4224
rect 12552 4160 12568 4224
rect 12632 4160 12648 4224
rect 12712 4160 12720 4224
rect 12400 4159 12720 4160
rect 17728 4224 18048 4225
rect 17728 4160 17736 4224
rect 17800 4160 17816 4224
rect 17880 4160 17896 4224
rect 17960 4160 17976 4224
rect 18040 4160 18048 4224
rect 17728 4159 18048 4160
rect 4408 3680 4728 3681
rect 4408 3616 4416 3680
rect 4480 3616 4496 3680
rect 4560 3616 4576 3680
rect 4640 3616 4656 3680
rect 4720 3616 4728 3680
rect 4408 3615 4728 3616
rect 9736 3680 10056 3681
rect 9736 3616 9744 3680
rect 9808 3616 9824 3680
rect 9888 3616 9904 3680
rect 9968 3616 9984 3680
rect 10048 3616 10056 3680
rect 9736 3615 10056 3616
rect 15064 3680 15384 3681
rect 15064 3616 15072 3680
rect 15136 3616 15152 3680
rect 15216 3616 15232 3680
rect 15296 3616 15312 3680
rect 15376 3616 15384 3680
rect 15064 3615 15384 3616
rect 7072 3136 7392 3137
rect 7072 3072 7080 3136
rect 7144 3072 7160 3136
rect 7224 3072 7240 3136
rect 7304 3072 7320 3136
rect 7384 3072 7392 3136
rect 7072 3071 7392 3072
rect 12400 3136 12720 3137
rect 12400 3072 12408 3136
rect 12472 3072 12488 3136
rect 12552 3072 12568 3136
rect 12632 3072 12648 3136
rect 12712 3072 12720 3136
rect 12400 3071 12720 3072
rect 17728 3136 18048 3137
rect 17728 3072 17736 3136
rect 17800 3072 17816 3136
rect 17880 3072 17896 3136
rect 17960 3072 17976 3136
rect 18040 3072 18048 3136
rect 17728 3071 18048 3072
rect 4408 2592 4728 2593
rect 4408 2528 4416 2592
rect 4480 2528 4496 2592
rect 4560 2528 4576 2592
rect 4640 2528 4656 2592
rect 4720 2528 4728 2592
rect 4408 2527 4728 2528
rect 9736 2592 10056 2593
rect 9736 2528 9744 2592
rect 9808 2528 9824 2592
rect 9888 2528 9904 2592
rect 9968 2528 9984 2592
rect 10048 2528 10056 2592
rect 9736 2527 10056 2528
rect 15064 2592 15384 2593
rect 15064 2528 15072 2592
rect 15136 2528 15152 2592
rect 15216 2528 15232 2592
rect 15296 2528 15312 2592
rect 15376 2528 15384 2592
rect 15064 2527 15384 2528
rect 7072 2048 7392 2049
rect 7072 1984 7080 2048
rect 7144 1984 7160 2048
rect 7224 1984 7240 2048
rect 7304 1984 7320 2048
rect 7384 1984 7392 2048
rect 7072 1983 7392 1984
rect 12400 2048 12720 2049
rect 12400 1984 12408 2048
rect 12472 1984 12488 2048
rect 12552 1984 12568 2048
rect 12632 1984 12648 2048
rect 12712 1984 12720 2048
rect 12400 1983 12720 1984
rect 17728 2048 18048 2049
rect 17728 1984 17736 2048
rect 17800 1984 17816 2048
rect 17880 1984 17896 2048
rect 17960 1984 17976 2048
rect 18040 1984 18048 2048
rect 17728 1983 18048 1984
rect 4408 1504 4728 1505
rect 4408 1440 4416 1504
rect 4480 1440 4496 1504
rect 4560 1440 4576 1504
rect 4640 1440 4656 1504
rect 4720 1440 4728 1504
rect 4408 1439 4728 1440
rect 9736 1504 10056 1505
rect 9736 1440 9744 1504
rect 9808 1440 9824 1504
rect 9888 1440 9904 1504
rect 9968 1440 9984 1504
rect 10048 1440 10056 1504
rect 9736 1439 10056 1440
rect 15064 1504 15384 1505
rect 15064 1440 15072 1504
rect 15136 1440 15152 1504
rect 15216 1440 15232 1504
rect 15296 1440 15312 1504
rect 15376 1440 15384 1504
rect 15064 1439 15384 1440
rect 2285 1162 2351 1165
rect 2929 1162 2995 1165
rect 830 1160 2995 1162
rect 830 1104 2290 1160
rect 2346 1104 2934 1160
rect 2990 1104 2995 1160
rect 830 1102 2995 1104
rect 830 920 890 1102
rect 2285 1099 2351 1102
rect 2929 1099 2995 1102
rect 7072 960 7392 961
rect 800 800 920 920
rect 7072 896 7080 960
rect 7144 896 7160 960
rect 7224 896 7240 960
rect 7304 896 7320 960
rect 7384 896 7392 960
rect 7072 895 7392 896
rect 12400 960 12720 961
rect 12400 896 12408 960
rect 12472 896 12488 960
rect 12552 896 12568 960
rect 12632 896 12648 960
rect 12712 896 12720 960
rect 12400 895 12720 896
rect 17728 960 18048 961
rect 17728 896 17736 960
rect 17800 896 17816 960
rect 17880 896 17896 960
rect 17960 896 17976 960
rect 18040 896 18048 960
rect 17728 895 18048 896
<< via3 >>
rect 4416 22172 4480 22176
rect 4416 22116 4420 22172
rect 4420 22116 4476 22172
rect 4476 22116 4480 22172
rect 4416 22112 4480 22116
rect 4496 22172 4560 22176
rect 4496 22116 4500 22172
rect 4500 22116 4556 22172
rect 4556 22116 4560 22172
rect 4496 22112 4560 22116
rect 4576 22172 4640 22176
rect 4576 22116 4580 22172
rect 4580 22116 4636 22172
rect 4636 22116 4640 22172
rect 4576 22112 4640 22116
rect 4656 22172 4720 22176
rect 4656 22116 4660 22172
rect 4660 22116 4716 22172
rect 4716 22116 4720 22172
rect 4656 22112 4720 22116
rect 9744 22172 9808 22176
rect 9744 22116 9748 22172
rect 9748 22116 9804 22172
rect 9804 22116 9808 22172
rect 9744 22112 9808 22116
rect 9824 22172 9888 22176
rect 9824 22116 9828 22172
rect 9828 22116 9884 22172
rect 9884 22116 9888 22172
rect 9824 22112 9888 22116
rect 9904 22172 9968 22176
rect 9904 22116 9908 22172
rect 9908 22116 9964 22172
rect 9964 22116 9968 22172
rect 9904 22112 9968 22116
rect 9984 22172 10048 22176
rect 9984 22116 9988 22172
rect 9988 22116 10044 22172
rect 10044 22116 10048 22172
rect 9984 22112 10048 22116
rect 15072 22172 15136 22176
rect 15072 22116 15076 22172
rect 15076 22116 15132 22172
rect 15132 22116 15136 22172
rect 15072 22112 15136 22116
rect 15152 22172 15216 22176
rect 15152 22116 15156 22172
rect 15156 22116 15212 22172
rect 15212 22116 15216 22172
rect 15152 22112 15216 22116
rect 15232 22172 15296 22176
rect 15232 22116 15236 22172
rect 15236 22116 15292 22172
rect 15292 22116 15296 22172
rect 15232 22112 15296 22116
rect 15312 22172 15376 22176
rect 15312 22116 15316 22172
rect 15316 22116 15372 22172
rect 15372 22116 15376 22172
rect 15312 22112 15376 22116
rect 7080 21628 7144 21632
rect 7080 21572 7084 21628
rect 7084 21572 7140 21628
rect 7140 21572 7144 21628
rect 7080 21568 7144 21572
rect 7160 21628 7224 21632
rect 7160 21572 7164 21628
rect 7164 21572 7220 21628
rect 7220 21572 7224 21628
rect 7160 21568 7224 21572
rect 7240 21628 7304 21632
rect 7240 21572 7244 21628
rect 7244 21572 7300 21628
rect 7300 21572 7304 21628
rect 7240 21568 7304 21572
rect 7320 21628 7384 21632
rect 7320 21572 7324 21628
rect 7324 21572 7380 21628
rect 7380 21572 7384 21628
rect 7320 21568 7384 21572
rect 12408 21628 12472 21632
rect 12408 21572 12412 21628
rect 12412 21572 12468 21628
rect 12468 21572 12472 21628
rect 12408 21568 12472 21572
rect 12488 21628 12552 21632
rect 12488 21572 12492 21628
rect 12492 21572 12548 21628
rect 12548 21572 12552 21628
rect 12488 21568 12552 21572
rect 12568 21628 12632 21632
rect 12568 21572 12572 21628
rect 12572 21572 12628 21628
rect 12628 21572 12632 21628
rect 12568 21568 12632 21572
rect 12648 21628 12712 21632
rect 12648 21572 12652 21628
rect 12652 21572 12708 21628
rect 12708 21572 12712 21628
rect 12648 21568 12712 21572
rect 17736 21628 17800 21632
rect 17736 21572 17740 21628
rect 17740 21572 17796 21628
rect 17796 21572 17800 21628
rect 17736 21568 17800 21572
rect 17816 21628 17880 21632
rect 17816 21572 17820 21628
rect 17820 21572 17876 21628
rect 17876 21572 17880 21628
rect 17816 21568 17880 21572
rect 17896 21628 17960 21632
rect 17896 21572 17900 21628
rect 17900 21572 17956 21628
rect 17956 21572 17960 21628
rect 17896 21568 17960 21572
rect 17976 21628 18040 21632
rect 17976 21572 17980 21628
rect 17980 21572 18036 21628
rect 18036 21572 18040 21628
rect 17976 21568 18040 21572
rect 4416 21084 4480 21088
rect 4416 21028 4420 21084
rect 4420 21028 4476 21084
rect 4476 21028 4480 21084
rect 4416 21024 4480 21028
rect 4496 21084 4560 21088
rect 4496 21028 4500 21084
rect 4500 21028 4556 21084
rect 4556 21028 4560 21084
rect 4496 21024 4560 21028
rect 4576 21084 4640 21088
rect 4576 21028 4580 21084
rect 4580 21028 4636 21084
rect 4636 21028 4640 21084
rect 4576 21024 4640 21028
rect 4656 21084 4720 21088
rect 4656 21028 4660 21084
rect 4660 21028 4716 21084
rect 4716 21028 4720 21084
rect 4656 21024 4720 21028
rect 9744 21084 9808 21088
rect 9744 21028 9748 21084
rect 9748 21028 9804 21084
rect 9804 21028 9808 21084
rect 9744 21024 9808 21028
rect 9824 21084 9888 21088
rect 9824 21028 9828 21084
rect 9828 21028 9884 21084
rect 9884 21028 9888 21084
rect 9824 21024 9888 21028
rect 9904 21084 9968 21088
rect 9904 21028 9908 21084
rect 9908 21028 9964 21084
rect 9964 21028 9968 21084
rect 9904 21024 9968 21028
rect 9984 21084 10048 21088
rect 9984 21028 9988 21084
rect 9988 21028 10044 21084
rect 10044 21028 10048 21084
rect 9984 21024 10048 21028
rect 15072 21084 15136 21088
rect 15072 21028 15076 21084
rect 15076 21028 15132 21084
rect 15132 21028 15136 21084
rect 15072 21024 15136 21028
rect 15152 21084 15216 21088
rect 15152 21028 15156 21084
rect 15156 21028 15212 21084
rect 15212 21028 15216 21084
rect 15152 21024 15216 21028
rect 15232 21084 15296 21088
rect 15232 21028 15236 21084
rect 15236 21028 15292 21084
rect 15292 21028 15296 21084
rect 15232 21024 15296 21028
rect 15312 21084 15376 21088
rect 15312 21028 15316 21084
rect 15316 21028 15372 21084
rect 15372 21028 15376 21084
rect 15312 21024 15376 21028
rect 7080 20540 7144 20544
rect 7080 20484 7084 20540
rect 7084 20484 7140 20540
rect 7140 20484 7144 20540
rect 7080 20480 7144 20484
rect 7160 20540 7224 20544
rect 7160 20484 7164 20540
rect 7164 20484 7220 20540
rect 7220 20484 7224 20540
rect 7160 20480 7224 20484
rect 7240 20540 7304 20544
rect 7240 20484 7244 20540
rect 7244 20484 7300 20540
rect 7300 20484 7304 20540
rect 7240 20480 7304 20484
rect 7320 20540 7384 20544
rect 7320 20484 7324 20540
rect 7324 20484 7380 20540
rect 7380 20484 7384 20540
rect 7320 20480 7384 20484
rect 12408 20540 12472 20544
rect 12408 20484 12412 20540
rect 12412 20484 12468 20540
rect 12468 20484 12472 20540
rect 12408 20480 12472 20484
rect 12488 20540 12552 20544
rect 12488 20484 12492 20540
rect 12492 20484 12548 20540
rect 12548 20484 12552 20540
rect 12488 20480 12552 20484
rect 12568 20540 12632 20544
rect 12568 20484 12572 20540
rect 12572 20484 12628 20540
rect 12628 20484 12632 20540
rect 12568 20480 12632 20484
rect 12648 20540 12712 20544
rect 12648 20484 12652 20540
rect 12652 20484 12708 20540
rect 12708 20484 12712 20540
rect 12648 20480 12712 20484
rect 17736 20540 17800 20544
rect 17736 20484 17740 20540
rect 17740 20484 17796 20540
rect 17796 20484 17800 20540
rect 17736 20480 17800 20484
rect 17816 20540 17880 20544
rect 17816 20484 17820 20540
rect 17820 20484 17876 20540
rect 17876 20484 17880 20540
rect 17816 20480 17880 20484
rect 17896 20540 17960 20544
rect 17896 20484 17900 20540
rect 17900 20484 17956 20540
rect 17956 20484 17960 20540
rect 17896 20480 17960 20484
rect 17976 20540 18040 20544
rect 17976 20484 17980 20540
rect 17980 20484 18036 20540
rect 18036 20484 18040 20540
rect 17976 20480 18040 20484
rect 4416 19996 4480 20000
rect 4416 19940 4420 19996
rect 4420 19940 4476 19996
rect 4476 19940 4480 19996
rect 4416 19936 4480 19940
rect 4496 19996 4560 20000
rect 4496 19940 4500 19996
rect 4500 19940 4556 19996
rect 4556 19940 4560 19996
rect 4496 19936 4560 19940
rect 4576 19996 4640 20000
rect 4576 19940 4580 19996
rect 4580 19940 4636 19996
rect 4636 19940 4640 19996
rect 4576 19936 4640 19940
rect 4656 19996 4720 20000
rect 4656 19940 4660 19996
rect 4660 19940 4716 19996
rect 4716 19940 4720 19996
rect 4656 19936 4720 19940
rect 9744 19996 9808 20000
rect 9744 19940 9748 19996
rect 9748 19940 9804 19996
rect 9804 19940 9808 19996
rect 9744 19936 9808 19940
rect 9824 19996 9888 20000
rect 9824 19940 9828 19996
rect 9828 19940 9884 19996
rect 9884 19940 9888 19996
rect 9824 19936 9888 19940
rect 9904 19996 9968 20000
rect 9904 19940 9908 19996
rect 9908 19940 9964 19996
rect 9964 19940 9968 19996
rect 9904 19936 9968 19940
rect 9984 19996 10048 20000
rect 9984 19940 9988 19996
rect 9988 19940 10044 19996
rect 10044 19940 10048 19996
rect 9984 19936 10048 19940
rect 15072 19996 15136 20000
rect 15072 19940 15076 19996
rect 15076 19940 15132 19996
rect 15132 19940 15136 19996
rect 15072 19936 15136 19940
rect 15152 19996 15216 20000
rect 15152 19940 15156 19996
rect 15156 19940 15212 19996
rect 15212 19940 15216 19996
rect 15152 19936 15216 19940
rect 15232 19996 15296 20000
rect 15232 19940 15236 19996
rect 15236 19940 15292 19996
rect 15292 19940 15296 19996
rect 15232 19936 15296 19940
rect 15312 19996 15376 20000
rect 15312 19940 15316 19996
rect 15316 19940 15372 19996
rect 15372 19940 15376 19996
rect 15312 19936 15376 19940
rect 7080 19452 7144 19456
rect 7080 19396 7084 19452
rect 7084 19396 7140 19452
rect 7140 19396 7144 19452
rect 7080 19392 7144 19396
rect 7160 19452 7224 19456
rect 7160 19396 7164 19452
rect 7164 19396 7220 19452
rect 7220 19396 7224 19452
rect 7160 19392 7224 19396
rect 7240 19452 7304 19456
rect 7240 19396 7244 19452
rect 7244 19396 7300 19452
rect 7300 19396 7304 19452
rect 7240 19392 7304 19396
rect 7320 19452 7384 19456
rect 7320 19396 7324 19452
rect 7324 19396 7380 19452
rect 7380 19396 7384 19452
rect 7320 19392 7384 19396
rect 12408 19452 12472 19456
rect 12408 19396 12412 19452
rect 12412 19396 12468 19452
rect 12468 19396 12472 19452
rect 12408 19392 12472 19396
rect 12488 19452 12552 19456
rect 12488 19396 12492 19452
rect 12492 19396 12548 19452
rect 12548 19396 12552 19452
rect 12488 19392 12552 19396
rect 12568 19452 12632 19456
rect 12568 19396 12572 19452
rect 12572 19396 12628 19452
rect 12628 19396 12632 19452
rect 12568 19392 12632 19396
rect 12648 19452 12712 19456
rect 12648 19396 12652 19452
rect 12652 19396 12708 19452
rect 12708 19396 12712 19452
rect 12648 19392 12712 19396
rect 17736 19452 17800 19456
rect 17736 19396 17740 19452
rect 17740 19396 17796 19452
rect 17796 19396 17800 19452
rect 17736 19392 17800 19396
rect 17816 19452 17880 19456
rect 17816 19396 17820 19452
rect 17820 19396 17876 19452
rect 17876 19396 17880 19452
rect 17816 19392 17880 19396
rect 17896 19452 17960 19456
rect 17896 19396 17900 19452
rect 17900 19396 17956 19452
rect 17956 19396 17960 19452
rect 17896 19392 17960 19396
rect 17976 19452 18040 19456
rect 17976 19396 17980 19452
rect 17980 19396 18036 19452
rect 18036 19396 18040 19452
rect 17976 19392 18040 19396
rect 4416 18908 4480 18912
rect 4416 18852 4420 18908
rect 4420 18852 4476 18908
rect 4476 18852 4480 18908
rect 4416 18848 4480 18852
rect 4496 18908 4560 18912
rect 4496 18852 4500 18908
rect 4500 18852 4556 18908
rect 4556 18852 4560 18908
rect 4496 18848 4560 18852
rect 4576 18908 4640 18912
rect 4576 18852 4580 18908
rect 4580 18852 4636 18908
rect 4636 18852 4640 18908
rect 4576 18848 4640 18852
rect 4656 18908 4720 18912
rect 4656 18852 4660 18908
rect 4660 18852 4716 18908
rect 4716 18852 4720 18908
rect 4656 18848 4720 18852
rect 9744 18908 9808 18912
rect 9744 18852 9748 18908
rect 9748 18852 9804 18908
rect 9804 18852 9808 18908
rect 9744 18848 9808 18852
rect 9824 18908 9888 18912
rect 9824 18852 9828 18908
rect 9828 18852 9884 18908
rect 9884 18852 9888 18908
rect 9824 18848 9888 18852
rect 9904 18908 9968 18912
rect 9904 18852 9908 18908
rect 9908 18852 9964 18908
rect 9964 18852 9968 18908
rect 9904 18848 9968 18852
rect 9984 18908 10048 18912
rect 9984 18852 9988 18908
rect 9988 18852 10044 18908
rect 10044 18852 10048 18908
rect 9984 18848 10048 18852
rect 15072 18908 15136 18912
rect 15072 18852 15076 18908
rect 15076 18852 15132 18908
rect 15132 18852 15136 18908
rect 15072 18848 15136 18852
rect 15152 18908 15216 18912
rect 15152 18852 15156 18908
rect 15156 18852 15212 18908
rect 15212 18852 15216 18908
rect 15152 18848 15216 18852
rect 15232 18908 15296 18912
rect 15232 18852 15236 18908
rect 15236 18852 15292 18908
rect 15292 18852 15296 18908
rect 15232 18848 15296 18852
rect 15312 18908 15376 18912
rect 15312 18852 15316 18908
rect 15316 18852 15372 18908
rect 15372 18852 15376 18908
rect 15312 18848 15376 18852
rect 7080 18364 7144 18368
rect 7080 18308 7084 18364
rect 7084 18308 7140 18364
rect 7140 18308 7144 18364
rect 7080 18304 7144 18308
rect 7160 18364 7224 18368
rect 7160 18308 7164 18364
rect 7164 18308 7220 18364
rect 7220 18308 7224 18364
rect 7160 18304 7224 18308
rect 7240 18364 7304 18368
rect 7240 18308 7244 18364
rect 7244 18308 7300 18364
rect 7300 18308 7304 18364
rect 7240 18304 7304 18308
rect 7320 18364 7384 18368
rect 7320 18308 7324 18364
rect 7324 18308 7380 18364
rect 7380 18308 7384 18364
rect 7320 18304 7384 18308
rect 12408 18364 12472 18368
rect 12408 18308 12412 18364
rect 12412 18308 12468 18364
rect 12468 18308 12472 18364
rect 12408 18304 12472 18308
rect 12488 18364 12552 18368
rect 12488 18308 12492 18364
rect 12492 18308 12548 18364
rect 12548 18308 12552 18364
rect 12488 18304 12552 18308
rect 12568 18364 12632 18368
rect 12568 18308 12572 18364
rect 12572 18308 12628 18364
rect 12628 18308 12632 18364
rect 12568 18304 12632 18308
rect 12648 18364 12712 18368
rect 12648 18308 12652 18364
rect 12652 18308 12708 18364
rect 12708 18308 12712 18364
rect 12648 18304 12712 18308
rect 17736 18364 17800 18368
rect 17736 18308 17740 18364
rect 17740 18308 17796 18364
rect 17796 18308 17800 18364
rect 17736 18304 17800 18308
rect 17816 18364 17880 18368
rect 17816 18308 17820 18364
rect 17820 18308 17876 18364
rect 17876 18308 17880 18364
rect 17816 18304 17880 18308
rect 17896 18364 17960 18368
rect 17896 18308 17900 18364
rect 17900 18308 17956 18364
rect 17956 18308 17960 18364
rect 17896 18304 17960 18308
rect 17976 18364 18040 18368
rect 17976 18308 17980 18364
rect 17980 18308 18036 18364
rect 18036 18308 18040 18364
rect 17976 18304 18040 18308
rect 4416 17820 4480 17824
rect 4416 17764 4420 17820
rect 4420 17764 4476 17820
rect 4476 17764 4480 17820
rect 4416 17760 4480 17764
rect 4496 17820 4560 17824
rect 4496 17764 4500 17820
rect 4500 17764 4556 17820
rect 4556 17764 4560 17820
rect 4496 17760 4560 17764
rect 4576 17820 4640 17824
rect 4576 17764 4580 17820
rect 4580 17764 4636 17820
rect 4636 17764 4640 17820
rect 4576 17760 4640 17764
rect 4656 17820 4720 17824
rect 4656 17764 4660 17820
rect 4660 17764 4716 17820
rect 4716 17764 4720 17820
rect 4656 17760 4720 17764
rect 9744 17820 9808 17824
rect 9744 17764 9748 17820
rect 9748 17764 9804 17820
rect 9804 17764 9808 17820
rect 9744 17760 9808 17764
rect 9824 17820 9888 17824
rect 9824 17764 9828 17820
rect 9828 17764 9884 17820
rect 9884 17764 9888 17820
rect 9824 17760 9888 17764
rect 9904 17820 9968 17824
rect 9904 17764 9908 17820
rect 9908 17764 9964 17820
rect 9964 17764 9968 17820
rect 9904 17760 9968 17764
rect 9984 17820 10048 17824
rect 9984 17764 9988 17820
rect 9988 17764 10044 17820
rect 10044 17764 10048 17820
rect 9984 17760 10048 17764
rect 15072 17820 15136 17824
rect 15072 17764 15076 17820
rect 15076 17764 15132 17820
rect 15132 17764 15136 17820
rect 15072 17760 15136 17764
rect 15152 17820 15216 17824
rect 15152 17764 15156 17820
rect 15156 17764 15212 17820
rect 15212 17764 15216 17820
rect 15152 17760 15216 17764
rect 15232 17820 15296 17824
rect 15232 17764 15236 17820
rect 15236 17764 15292 17820
rect 15292 17764 15296 17820
rect 15232 17760 15296 17764
rect 15312 17820 15376 17824
rect 15312 17764 15316 17820
rect 15316 17764 15372 17820
rect 15372 17764 15376 17820
rect 15312 17760 15376 17764
rect 7080 17276 7144 17280
rect 7080 17220 7084 17276
rect 7084 17220 7140 17276
rect 7140 17220 7144 17276
rect 7080 17216 7144 17220
rect 7160 17276 7224 17280
rect 7160 17220 7164 17276
rect 7164 17220 7220 17276
rect 7220 17220 7224 17276
rect 7160 17216 7224 17220
rect 7240 17276 7304 17280
rect 7240 17220 7244 17276
rect 7244 17220 7300 17276
rect 7300 17220 7304 17276
rect 7240 17216 7304 17220
rect 7320 17276 7384 17280
rect 7320 17220 7324 17276
rect 7324 17220 7380 17276
rect 7380 17220 7384 17276
rect 7320 17216 7384 17220
rect 12408 17276 12472 17280
rect 12408 17220 12412 17276
rect 12412 17220 12468 17276
rect 12468 17220 12472 17276
rect 12408 17216 12472 17220
rect 12488 17276 12552 17280
rect 12488 17220 12492 17276
rect 12492 17220 12548 17276
rect 12548 17220 12552 17276
rect 12488 17216 12552 17220
rect 12568 17276 12632 17280
rect 12568 17220 12572 17276
rect 12572 17220 12628 17276
rect 12628 17220 12632 17276
rect 12568 17216 12632 17220
rect 12648 17276 12712 17280
rect 12648 17220 12652 17276
rect 12652 17220 12708 17276
rect 12708 17220 12712 17276
rect 12648 17216 12712 17220
rect 17736 17276 17800 17280
rect 17736 17220 17740 17276
rect 17740 17220 17796 17276
rect 17796 17220 17800 17276
rect 17736 17216 17800 17220
rect 17816 17276 17880 17280
rect 17816 17220 17820 17276
rect 17820 17220 17876 17276
rect 17876 17220 17880 17276
rect 17816 17216 17880 17220
rect 17896 17276 17960 17280
rect 17896 17220 17900 17276
rect 17900 17220 17956 17276
rect 17956 17220 17960 17276
rect 17896 17216 17960 17220
rect 17976 17276 18040 17280
rect 17976 17220 17980 17276
rect 17980 17220 18036 17276
rect 18036 17220 18040 17276
rect 17976 17216 18040 17220
rect 4416 16732 4480 16736
rect 4416 16676 4420 16732
rect 4420 16676 4476 16732
rect 4476 16676 4480 16732
rect 4416 16672 4480 16676
rect 4496 16732 4560 16736
rect 4496 16676 4500 16732
rect 4500 16676 4556 16732
rect 4556 16676 4560 16732
rect 4496 16672 4560 16676
rect 4576 16732 4640 16736
rect 4576 16676 4580 16732
rect 4580 16676 4636 16732
rect 4636 16676 4640 16732
rect 4576 16672 4640 16676
rect 4656 16732 4720 16736
rect 4656 16676 4660 16732
rect 4660 16676 4716 16732
rect 4716 16676 4720 16732
rect 4656 16672 4720 16676
rect 9744 16732 9808 16736
rect 9744 16676 9748 16732
rect 9748 16676 9804 16732
rect 9804 16676 9808 16732
rect 9744 16672 9808 16676
rect 9824 16732 9888 16736
rect 9824 16676 9828 16732
rect 9828 16676 9884 16732
rect 9884 16676 9888 16732
rect 9824 16672 9888 16676
rect 9904 16732 9968 16736
rect 9904 16676 9908 16732
rect 9908 16676 9964 16732
rect 9964 16676 9968 16732
rect 9904 16672 9968 16676
rect 9984 16732 10048 16736
rect 9984 16676 9988 16732
rect 9988 16676 10044 16732
rect 10044 16676 10048 16732
rect 9984 16672 10048 16676
rect 15072 16732 15136 16736
rect 15072 16676 15076 16732
rect 15076 16676 15132 16732
rect 15132 16676 15136 16732
rect 15072 16672 15136 16676
rect 15152 16732 15216 16736
rect 15152 16676 15156 16732
rect 15156 16676 15212 16732
rect 15212 16676 15216 16732
rect 15152 16672 15216 16676
rect 15232 16732 15296 16736
rect 15232 16676 15236 16732
rect 15236 16676 15292 16732
rect 15292 16676 15296 16732
rect 15232 16672 15296 16676
rect 15312 16732 15376 16736
rect 15312 16676 15316 16732
rect 15316 16676 15372 16732
rect 15372 16676 15376 16732
rect 15312 16672 15376 16676
rect 7080 16188 7144 16192
rect 7080 16132 7084 16188
rect 7084 16132 7140 16188
rect 7140 16132 7144 16188
rect 7080 16128 7144 16132
rect 7160 16188 7224 16192
rect 7160 16132 7164 16188
rect 7164 16132 7220 16188
rect 7220 16132 7224 16188
rect 7160 16128 7224 16132
rect 7240 16188 7304 16192
rect 7240 16132 7244 16188
rect 7244 16132 7300 16188
rect 7300 16132 7304 16188
rect 7240 16128 7304 16132
rect 7320 16188 7384 16192
rect 7320 16132 7324 16188
rect 7324 16132 7380 16188
rect 7380 16132 7384 16188
rect 7320 16128 7384 16132
rect 12408 16188 12472 16192
rect 12408 16132 12412 16188
rect 12412 16132 12468 16188
rect 12468 16132 12472 16188
rect 12408 16128 12472 16132
rect 12488 16188 12552 16192
rect 12488 16132 12492 16188
rect 12492 16132 12548 16188
rect 12548 16132 12552 16188
rect 12488 16128 12552 16132
rect 12568 16188 12632 16192
rect 12568 16132 12572 16188
rect 12572 16132 12628 16188
rect 12628 16132 12632 16188
rect 12568 16128 12632 16132
rect 12648 16188 12712 16192
rect 12648 16132 12652 16188
rect 12652 16132 12708 16188
rect 12708 16132 12712 16188
rect 12648 16128 12712 16132
rect 17736 16188 17800 16192
rect 17736 16132 17740 16188
rect 17740 16132 17796 16188
rect 17796 16132 17800 16188
rect 17736 16128 17800 16132
rect 17816 16188 17880 16192
rect 17816 16132 17820 16188
rect 17820 16132 17876 16188
rect 17876 16132 17880 16188
rect 17816 16128 17880 16132
rect 17896 16188 17960 16192
rect 17896 16132 17900 16188
rect 17900 16132 17956 16188
rect 17956 16132 17960 16188
rect 17896 16128 17960 16132
rect 17976 16188 18040 16192
rect 17976 16132 17980 16188
rect 17980 16132 18036 16188
rect 18036 16132 18040 16188
rect 17976 16128 18040 16132
rect 4416 15644 4480 15648
rect 4416 15588 4420 15644
rect 4420 15588 4476 15644
rect 4476 15588 4480 15644
rect 4416 15584 4480 15588
rect 4496 15644 4560 15648
rect 4496 15588 4500 15644
rect 4500 15588 4556 15644
rect 4556 15588 4560 15644
rect 4496 15584 4560 15588
rect 4576 15644 4640 15648
rect 4576 15588 4580 15644
rect 4580 15588 4636 15644
rect 4636 15588 4640 15644
rect 4576 15584 4640 15588
rect 4656 15644 4720 15648
rect 4656 15588 4660 15644
rect 4660 15588 4716 15644
rect 4716 15588 4720 15644
rect 4656 15584 4720 15588
rect 9744 15644 9808 15648
rect 9744 15588 9748 15644
rect 9748 15588 9804 15644
rect 9804 15588 9808 15644
rect 9744 15584 9808 15588
rect 9824 15644 9888 15648
rect 9824 15588 9828 15644
rect 9828 15588 9884 15644
rect 9884 15588 9888 15644
rect 9824 15584 9888 15588
rect 9904 15644 9968 15648
rect 9904 15588 9908 15644
rect 9908 15588 9964 15644
rect 9964 15588 9968 15644
rect 9904 15584 9968 15588
rect 9984 15644 10048 15648
rect 9984 15588 9988 15644
rect 9988 15588 10044 15644
rect 10044 15588 10048 15644
rect 9984 15584 10048 15588
rect 15072 15644 15136 15648
rect 15072 15588 15076 15644
rect 15076 15588 15132 15644
rect 15132 15588 15136 15644
rect 15072 15584 15136 15588
rect 15152 15644 15216 15648
rect 15152 15588 15156 15644
rect 15156 15588 15212 15644
rect 15212 15588 15216 15644
rect 15152 15584 15216 15588
rect 15232 15644 15296 15648
rect 15232 15588 15236 15644
rect 15236 15588 15292 15644
rect 15292 15588 15296 15644
rect 15232 15584 15296 15588
rect 15312 15644 15376 15648
rect 15312 15588 15316 15644
rect 15316 15588 15372 15644
rect 15372 15588 15376 15644
rect 15312 15584 15376 15588
rect 7080 15100 7144 15104
rect 7080 15044 7084 15100
rect 7084 15044 7140 15100
rect 7140 15044 7144 15100
rect 7080 15040 7144 15044
rect 7160 15100 7224 15104
rect 7160 15044 7164 15100
rect 7164 15044 7220 15100
rect 7220 15044 7224 15100
rect 7160 15040 7224 15044
rect 7240 15100 7304 15104
rect 7240 15044 7244 15100
rect 7244 15044 7300 15100
rect 7300 15044 7304 15100
rect 7240 15040 7304 15044
rect 7320 15100 7384 15104
rect 7320 15044 7324 15100
rect 7324 15044 7380 15100
rect 7380 15044 7384 15100
rect 7320 15040 7384 15044
rect 12408 15100 12472 15104
rect 12408 15044 12412 15100
rect 12412 15044 12468 15100
rect 12468 15044 12472 15100
rect 12408 15040 12472 15044
rect 12488 15100 12552 15104
rect 12488 15044 12492 15100
rect 12492 15044 12548 15100
rect 12548 15044 12552 15100
rect 12488 15040 12552 15044
rect 12568 15100 12632 15104
rect 12568 15044 12572 15100
rect 12572 15044 12628 15100
rect 12628 15044 12632 15100
rect 12568 15040 12632 15044
rect 12648 15100 12712 15104
rect 12648 15044 12652 15100
rect 12652 15044 12708 15100
rect 12708 15044 12712 15100
rect 12648 15040 12712 15044
rect 17736 15100 17800 15104
rect 17736 15044 17740 15100
rect 17740 15044 17796 15100
rect 17796 15044 17800 15100
rect 17736 15040 17800 15044
rect 17816 15100 17880 15104
rect 17816 15044 17820 15100
rect 17820 15044 17876 15100
rect 17876 15044 17880 15100
rect 17816 15040 17880 15044
rect 17896 15100 17960 15104
rect 17896 15044 17900 15100
rect 17900 15044 17956 15100
rect 17956 15044 17960 15100
rect 17896 15040 17960 15044
rect 17976 15100 18040 15104
rect 17976 15044 17980 15100
rect 17980 15044 18036 15100
rect 18036 15044 18040 15100
rect 17976 15040 18040 15044
rect 4416 14556 4480 14560
rect 4416 14500 4420 14556
rect 4420 14500 4476 14556
rect 4476 14500 4480 14556
rect 4416 14496 4480 14500
rect 4496 14556 4560 14560
rect 4496 14500 4500 14556
rect 4500 14500 4556 14556
rect 4556 14500 4560 14556
rect 4496 14496 4560 14500
rect 4576 14556 4640 14560
rect 4576 14500 4580 14556
rect 4580 14500 4636 14556
rect 4636 14500 4640 14556
rect 4576 14496 4640 14500
rect 4656 14556 4720 14560
rect 4656 14500 4660 14556
rect 4660 14500 4716 14556
rect 4716 14500 4720 14556
rect 4656 14496 4720 14500
rect 9744 14556 9808 14560
rect 9744 14500 9748 14556
rect 9748 14500 9804 14556
rect 9804 14500 9808 14556
rect 9744 14496 9808 14500
rect 9824 14556 9888 14560
rect 9824 14500 9828 14556
rect 9828 14500 9884 14556
rect 9884 14500 9888 14556
rect 9824 14496 9888 14500
rect 9904 14556 9968 14560
rect 9904 14500 9908 14556
rect 9908 14500 9964 14556
rect 9964 14500 9968 14556
rect 9904 14496 9968 14500
rect 9984 14556 10048 14560
rect 9984 14500 9988 14556
rect 9988 14500 10044 14556
rect 10044 14500 10048 14556
rect 9984 14496 10048 14500
rect 15072 14556 15136 14560
rect 15072 14500 15076 14556
rect 15076 14500 15132 14556
rect 15132 14500 15136 14556
rect 15072 14496 15136 14500
rect 15152 14556 15216 14560
rect 15152 14500 15156 14556
rect 15156 14500 15212 14556
rect 15212 14500 15216 14556
rect 15152 14496 15216 14500
rect 15232 14556 15296 14560
rect 15232 14500 15236 14556
rect 15236 14500 15292 14556
rect 15292 14500 15296 14556
rect 15232 14496 15296 14500
rect 15312 14556 15376 14560
rect 15312 14500 15316 14556
rect 15316 14500 15372 14556
rect 15372 14500 15376 14556
rect 15312 14496 15376 14500
rect 7080 14012 7144 14016
rect 7080 13956 7084 14012
rect 7084 13956 7140 14012
rect 7140 13956 7144 14012
rect 7080 13952 7144 13956
rect 7160 14012 7224 14016
rect 7160 13956 7164 14012
rect 7164 13956 7220 14012
rect 7220 13956 7224 14012
rect 7160 13952 7224 13956
rect 7240 14012 7304 14016
rect 7240 13956 7244 14012
rect 7244 13956 7300 14012
rect 7300 13956 7304 14012
rect 7240 13952 7304 13956
rect 7320 14012 7384 14016
rect 7320 13956 7324 14012
rect 7324 13956 7380 14012
rect 7380 13956 7384 14012
rect 7320 13952 7384 13956
rect 12408 14012 12472 14016
rect 12408 13956 12412 14012
rect 12412 13956 12468 14012
rect 12468 13956 12472 14012
rect 12408 13952 12472 13956
rect 12488 14012 12552 14016
rect 12488 13956 12492 14012
rect 12492 13956 12548 14012
rect 12548 13956 12552 14012
rect 12488 13952 12552 13956
rect 12568 14012 12632 14016
rect 12568 13956 12572 14012
rect 12572 13956 12628 14012
rect 12628 13956 12632 14012
rect 12568 13952 12632 13956
rect 12648 14012 12712 14016
rect 12648 13956 12652 14012
rect 12652 13956 12708 14012
rect 12708 13956 12712 14012
rect 12648 13952 12712 13956
rect 17736 14012 17800 14016
rect 17736 13956 17740 14012
rect 17740 13956 17796 14012
rect 17796 13956 17800 14012
rect 17736 13952 17800 13956
rect 17816 14012 17880 14016
rect 17816 13956 17820 14012
rect 17820 13956 17876 14012
rect 17876 13956 17880 14012
rect 17816 13952 17880 13956
rect 17896 14012 17960 14016
rect 17896 13956 17900 14012
rect 17900 13956 17956 14012
rect 17956 13956 17960 14012
rect 17896 13952 17960 13956
rect 17976 14012 18040 14016
rect 17976 13956 17980 14012
rect 17980 13956 18036 14012
rect 18036 13956 18040 14012
rect 17976 13952 18040 13956
rect 4416 13468 4480 13472
rect 4416 13412 4420 13468
rect 4420 13412 4476 13468
rect 4476 13412 4480 13468
rect 4416 13408 4480 13412
rect 4496 13468 4560 13472
rect 4496 13412 4500 13468
rect 4500 13412 4556 13468
rect 4556 13412 4560 13468
rect 4496 13408 4560 13412
rect 4576 13468 4640 13472
rect 4576 13412 4580 13468
rect 4580 13412 4636 13468
rect 4636 13412 4640 13468
rect 4576 13408 4640 13412
rect 4656 13468 4720 13472
rect 4656 13412 4660 13468
rect 4660 13412 4716 13468
rect 4716 13412 4720 13468
rect 4656 13408 4720 13412
rect 9744 13468 9808 13472
rect 9744 13412 9748 13468
rect 9748 13412 9804 13468
rect 9804 13412 9808 13468
rect 9744 13408 9808 13412
rect 9824 13468 9888 13472
rect 9824 13412 9828 13468
rect 9828 13412 9884 13468
rect 9884 13412 9888 13468
rect 9824 13408 9888 13412
rect 9904 13468 9968 13472
rect 9904 13412 9908 13468
rect 9908 13412 9964 13468
rect 9964 13412 9968 13468
rect 9904 13408 9968 13412
rect 9984 13468 10048 13472
rect 9984 13412 9988 13468
rect 9988 13412 10044 13468
rect 10044 13412 10048 13468
rect 9984 13408 10048 13412
rect 15072 13468 15136 13472
rect 15072 13412 15076 13468
rect 15076 13412 15132 13468
rect 15132 13412 15136 13468
rect 15072 13408 15136 13412
rect 15152 13468 15216 13472
rect 15152 13412 15156 13468
rect 15156 13412 15212 13468
rect 15212 13412 15216 13468
rect 15152 13408 15216 13412
rect 15232 13468 15296 13472
rect 15232 13412 15236 13468
rect 15236 13412 15292 13468
rect 15292 13412 15296 13468
rect 15232 13408 15296 13412
rect 15312 13468 15376 13472
rect 15312 13412 15316 13468
rect 15316 13412 15372 13468
rect 15372 13412 15376 13468
rect 15312 13408 15376 13412
rect 7080 12924 7144 12928
rect 7080 12868 7084 12924
rect 7084 12868 7140 12924
rect 7140 12868 7144 12924
rect 7080 12864 7144 12868
rect 7160 12924 7224 12928
rect 7160 12868 7164 12924
rect 7164 12868 7220 12924
rect 7220 12868 7224 12924
rect 7160 12864 7224 12868
rect 7240 12924 7304 12928
rect 7240 12868 7244 12924
rect 7244 12868 7300 12924
rect 7300 12868 7304 12924
rect 7240 12864 7304 12868
rect 7320 12924 7384 12928
rect 7320 12868 7324 12924
rect 7324 12868 7380 12924
rect 7380 12868 7384 12924
rect 7320 12864 7384 12868
rect 12408 12924 12472 12928
rect 12408 12868 12412 12924
rect 12412 12868 12468 12924
rect 12468 12868 12472 12924
rect 12408 12864 12472 12868
rect 12488 12924 12552 12928
rect 12488 12868 12492 12924
rect 12492 12868 12548 12924
rect 12548 12868 12552 12924
rect 12488 12864 12552 12868
rect 12568 12924 12632 12928
rect 12568 12868 12572 12924
rect 12572 12868 12628 12924
rect 12628 12868 12632 12924
rect 12568 12864 12632 12868
rect 12648 12924 12712 12928
rect 12648 12868 12652 12924
rect 12652 12868 12708 12924
rect 12708 12868 12712 12924
rect 12648 12864 12712 12868
rect 17736 12924 17800 12928
rect 17736 12868 17740 12924
rect 17740 12868 17796 12924
rect 17796 12868 17800 12924
rect 17736 12864 17800 12868
rect 17816 12924 17880 12928
rect 17816 12868 17820 12924
rect 17820 12868 17876 12924
rect 17876 12868 17880 12924
rect 17816 12864 17880 12868
rect 17896 12924 17960 12928
rect 17896 12868 17900 12924
rect 17900 12868 17956 12924
rect 17956 12868 17960 12924
rect 17896 12864 17960 12868
rect 17976 12924 18040 12928
rect 17976 12868 17980 12924
rect 17980 12868 18036 12924
rect 18036 12868 18040 12924
rect 17976 12864 18040 12868
rect 4416 12380 4480 12384
rect 4416 12324 4420 12380
rect 4420 12324 4476 12380
rect 4476 12324 4480 12380
rect 4416 12320 4480 12324
rect 4496 12380 4560 12384
rect 4496 12324 4500 12380
rect 4500 12324 4556 12380
rect 4556 12324 4560 12380
rect 4496 12320 4560 12324
rect 4576 12380 4640 12384
rect 4576 12324 4580 12380
rect 4580 12324 4636 12380
rect 4636 12324 4640 12380
rect 4576 12320 4640 12324
rect 4656 12380 4720 12384
rect 4656 12324 4660 12380
rect 4660 12324 4716 12380
rect 4716 12324 4720 12380
rect 4656 12320 4720 12324
rect 9744 12380 9808 12384
rect 9744 12324 9748 12380
rect 9748 12324 9804 12380
rect 9804 12324 9808 12380
rect 9744 12320 9808 12324
rect 9824 12380 9888 12384
rect 9824 12324 9828 12380
rect 9828 12324 9884 12380
rect 9884 12324 9888 12380
rect 9824 12320 9888 12324
rect 9904 12380 9968 12384
rect 9904 12324 9908 12380
rect 9908 12324 9964 12380
rect 9964 12324 9968 12380
rect 9904 12320 9968 12324
rect 9984 12380 10048 12384
rect 9984 12324 9988 12380
rect 9988 12324 10044 12380
rect 10044 12324 10048 12380
rect 9984 12320 10048 12324
rect 15072 12380 15136 12384
rect 15072 12324 15076 12380
rect 15076 12324 15132 12380
rect 15132 12324 15136 12380
rect 15072 12320 15136 12324
rect 15152 12380 15216 12384
rect 15152 12324 15156 12380
rect 15156 12324 15212 12380
rect 15212 12324 15216 12380
rect 15152 12320 15216 12324
rect 15232 12380 15296 12384
rect 15232 12324 15236 12380
rect 15236 12324 15292 12380
rect 15292 12324 15296 12380
rect 15232 12320 15296 12324
rect 15312 12380 15376 12384
rect 15312 12324 15316 12380
rect 15316 12324 15372 12380
rect 15372 12324 15376 12380
rect 15312 12320 15376 12324
rect 7080 11836 7144 11840
rect 7080 11780 7084 11836
rect 7084 11780 7140 11836
rect 7140 11780 7144 11836
rect 7080 11776 7144 11780
rect 7160 11836 7224 11840
rect 7160 11780 7164 11836
rect 7164 11780 7220 11836
rect 7220 11780 7224 11836
rect 7160 11776 7224 11780
rect 7240 11836 7304 11840
rect 7240 11780 7244 11836
rect 7244 11780 7300 11836
rect 7300 11780 7304 11836
rect 7240 11776 7304 11780
rect 7320 11836 7384 11840
rect 7320 11780 7324 11836
rect 7324 11780 7380 11836
rect 7380 11780 7384 11836
rect 7320 11776 7384 11780
rect 12408 11836 12472 11840
rect 12408 11780 12412 11836
rect 12412 11780 12468 11836
rect 12468 11780 12472 11836
rect 12408 11776 12472 11780
rect 12488 11836 12552 11840
rect 12488 11780 12492 11836
rect 12492 11780 12548 11836
rect 12548 11780 12552 11836
rect 12488 11776 12552 11780
rect 12568 11836 12632 11840
rect 12568 11780 12572 11836
rect 12572 11780 12628 11836
rect 12628 11780 12632 11836
rect 12568 11776 12632 11780
rect 12648 11836 12712 11840
rect 12648 11780 12652 11836
rect 12652 11780 12708 11836
rect 12708 11780 12712 11836
rect 12648 11776 12712 11780
rect 17736 11836 17800 11840
rect 17736 11780 17740 11836
rect 17740 11780 17796 11836
rect 17796 11780 17800 11836
rect 17736 11776 17800 11780
rect 17816 11836 17880 11840
rect 17816 11780 17820 11836
rect 17820 11780 17876 11836
rect 17876 11780 17880 11836
rect 17816 11776 17880 11780
rect 17896 11836 17960 11840
rect 17896 11780 17900 11836
rect 17900 11780 17956 11836
rect 17956 11780 17960 11836
rect 17896 11776 17960 11780
rect 17976 11836 18040 11840
rect 17976 11780 17980 11836
rect 17980 11780 18036 11836
rect 18036 11780 18040 11836
rect 17976 11776 18040 11780
rect 4416 11292 4480 11296
rect 4416 11236 4420 11292
rect 4420 11236 4476 11292
rect 4476 11236 4480 11292
rect 4416 11232 4480 11236
rect 4496 11292 4560 11296
rect 4496 11236 4500 11292
rect 4500 11236 4556 11292
rect 4556 11236 4560 11292
rect 4496 11232 4560 11236
rect 4576 11292 4640 11296
rect 4576 11236 4580 11292
rect 4580 11236 4636 11292
rect 4636 11236 4640 11292
rect 4576 11232 4640 11236
rect 4656 11292 4720 11296
rect 4656 11236 4660 11292
rect 4660 11236 4716 11292
rect 4716 11236 4720 11292
rect 4656 11232 4720 11236
rect 9744 11292 9808 11296
rect 9744 11236 9748 11292
rect 9748 11236 9804 11292
rect 9804 11236 9808 11292
rect 9744 11232 9808 11236
rect 9824 11292 9888 11296
rect 9824 11236 9828 11292
rect 9828 11236 9884 11292
rect 9884 11236 9888 11292
rect 9824 11232 9888 11236
rect 9904 11292 9968 11296
rect 9904 11236 9908 11292
rect 9908 11236 9964 11292
rect 9964 11236 9968 11292
rect 9904 11232 9968 11236
rect 9984 11292 10048 11296
rect 9984 11236 9988 11292
rect 9988 11236 10044 11292
rect 10044 11236 10048 11292
rect 9984 11232 10048 11236
rect 15072 11292 15136 11296
rect 15072 11236 15076 11292
rect 15076 11236 15132 11292
rect 15132 11236 15136 11292
rect 15072 11232 15136 11236
rect 15152 11292 15216 11296
rect 15152 11236 15156 11292
rect 15156 11236 15212 11292
rect 15212 11236 15216 11292
rect 15152 11232 15216 11236
rect 15232 11292 15296 11296
rect 15232 11236 15236 11292
rect 15236 11236 15292 11292
rect 15292 11236 15296 11292
rect 15232 11232 15296 11236
rect 15312 11292 15376 11296
rect 15312 11236 15316 11292
rect 15316 11236 15372 11292
rect 15372 11236 15376 11292
rect 15312 11232 15376 11236
rect 7080 10748 7144 10752
rect 7080 10692 7084 10748
rect 7084 10692 7140 10748
rect 7140 10692 7144 10748
rect 7080 10688 7144 10692
rect 7160 10748 7224 10752
rect 7160 10692 7164 10748
rect 7164 10692 7220 10748
rect 7220 10692 7224 10748
rect 7160 10688 7224 10692
rect 7240 10748 7304 10752
rect 7240 10692 7244 10748
rect 7244 10692 7300 10748
rect 7300 10692 7304 10748
rect 7240 10688 7304 10692
rect 7320 10748 7384 10752
rect 7320 10692 7324 10748
rect 7324 10692 7380 10748
rect 7380 10692 7384 10748
rect 7320 10688 7384 10692
rect 12408 10748 12472 10752
rect 12408 10692 12412 10748
rect 12412 10692 12468 10748
rect 12468 10692 12472 10748
rect 12408 10688 12472 10692
rect 12488 10748 12552 10752
rect 12488 10692 12492 10748
rect 12492 10692 12548 10748
rect 12548 10692 12552 10748
rect 12488 10688 12552 10692
rect 12568 10748 12632 10752
rect 12568 10692 12572 10748
rect 12572 10692 12628 10748
rect 12628 10692 12632 10748
rect 12568 10688 12632 10692
rect 12648 10748 12712 10752
rect 12648 10692 12652 10748
rect 12652 10692 12708 10748
rect 12708 10692 12712 10748
rect 12648 10688 12712 10692
rect 17736 10748 17800 10752
rect 17736 10692 17740 10748
rect 17740 10692 17796 10748
rect 17796 10692 17800 10748
rect 17736 10688 17800 10692
rect 17816 10748 17880 10752
rect 17816 10692 17820 10748
rect 17820 10692 17876 10748
rect 17876 10692 17880 10748
rect 17816 10688 17880 10692
rect 17896 10748 17960 10752
rect 17896 10692 17900 10748
rect 17900 10692 17956 10748
rect 17956 10692 17960 10748
rect 17896 10688 17960 10692
rect 17976 10748 18040 10752
rect 17976 10692 17980 10748
rect 17980 10692 18036 10748
rect 18036 10692 18040 10748
rect 17976 10688 18040 10692
rect 4416 10204 4480 10208
rect 4416 10148 4420 10204
rect 4420 10148 4476 10204
rect 4476 10148 4480 10204
rect 4416 10144 4480 10148
rect 4496 10204 4560 10208
rect 4496 10148 4500 10204
rect 4500 10148 4556 10204
rect 4556 10148 4560 10204
rect 4496 10144 4560 10148
rect 4576 10204 4640 10208
rect 4576 10148 4580 10204
rect 4580 10148 4636 10204
rect 4636 10148 4640 10204
rect 4576 10144 4640 10148
rect 4656 10204 4720 10208
rect 4656 10148 4660 10204
rect 4660 10148 4716 10204
rect 4716 10148 4720 10204
rect 4656 10144 4720 10148
rect 9744 10204 9808 10208
rect 9744 10148 9748 10204
rect 9748 10148 9804 10204
rect 9804 10148 9808 10204
rect 9744 10144 9808 10148
rect 9824 10204 9888 10208
rect 9824 10148 9828 10204
rect 9828 10148 9884 10204
rect 9884 10148 9888 10204
rect 9824 10144 9888 10148
rect 9904 10204 9968 10208
rect 9904 10148 9908 10204
rect 9908 10148 9964 10204
rect 9964 10148 9968 10204
rect 9904 10144 9968 10148
rect 9984 10204 10048 10208
rect 9984 10148 9988 10204
rect 9988 10148 10044 10204
rect 10044 10148 10048 10204
rect 9984 10144 10048 10148
rect 15072 10204 15136 10208
rect 15072 10148 15076 10204
rect 15076 10148 15132 10204
rect 15132 10148 15136 10204
rect 15072 10144 15136 10148
rect 15152 10204 15216 10208
rect 15152 10148 15156 10204
rect 15156 10148 15212 10204
rect 15212 10148 15216 10204
rect 15152 10144 15216 10148
rect 15232 10204 15296 10208
rect 15232 10148 15236 10204
rect 15236 10148 15292 10204
rect 15292 10148 15296 10204
rect 15232 10144 15296 10148
rect 15312 10204 15376 10208
rect 15312 10148 15316 10204
rect 15316 10148 15372 10204
rect 15372 10148 15376 10204
rect 15312 10144 15376 10148
rect 7080 9660 7144 9664
rect 7080 9604 7084 9660
rect 7084 9604 7140 9660
rect 7140 9604 7144 9660
rect 7080 9600 7144 9604
rect 7160 9660 7224 9664
rect 7160 9604 7164 9660
rect 7164 9604 7220 9660
rect 7220 9604 7224 9660
rect 7160 9600 7224 9604
rect 7240 9660 7304 9664
rect 7240 9604 7244 9660
rect 7244 9604 7300 9660
rect 7300 9604 7304 9660
rect 7240 9600 7304 9604
rect 7320 9660 7384 9664
rect 7320 9604 7324 9660
rect 7324 9604 7380 9660
rect 7380 9604 7384 9660
rect 7320 9600 7384 9604
rect 12408 9660 12472 9664
rect 12408 9604 12412 9660
rect 12412 9604 12468 9660
rect 12468 9604 12472 9660
rect 12408 9600 12472 9604
rect 12488 9660 12552 9664
rect 12488 9604 12492 9660
rect 12492 9604 12548 9660
rect 12548 9604 12552 9660
rect 12488 9600 12552 9604
rect 12568 9660 12632 9664
rect 12568 9604 12572 9660
rect 12572 9604 12628 9660
rect 12628 9604 12632 9660
rect 12568 9600 12632 9604
rect 12648 9660 12712 9664
rect 12648 9604 12652 9660
rect 12652 9604 12708 9660
rect 12708 9604 12712 9660
rect 12648 9600 12712 9604
rect 17736 9660 17800 9664
rect 17736 9604 17740 9660
rect 17740 9604 17796 9660
rect 17796 9604 17800 9660
rect 17736 9600 17800 9604
rect 17816 9660 17880 9664
rect 17816 9604 17820 9660
rect 17820 9604 17876 9660
rect 17876 9604 17880 9660
rect 17816 9600 17880 9604
rect 17896 9660 17960 9664
rect 17896 9604 17900 9660
rect 17900 9604 17956 9660
rect 17956 9604 17960 9660
rect 17896 9600 17960 9604
rect 17976 9660 18040 9664
rect 17976 9604 17980 9660
rect 17980 9604 18036 9660
rect 18036 9604 18040 9660
rect 17976 9600 18040 9604
rect 4416 9116 4480 9120
rect 4416 9060 4420 9116
rect 4420 9060 4476 9116
rect 4476 9060 4480 9116
rect 4416 9056 4480 9060
rect 4496 9116 4560 9120
rect 4496 9060 4500 9116
rect 4500 9060 4556 9116
rect 4556 9060 4560 9116
rect 4496 9056 4560 9060
rect 4576 9116 4640 9120
rect 4576 9060 4580 9116
rect 4580 9060 4636 9116
rect 4636 9060 4640 9116
rect 4576 9056 4640 9060
rect 4656 9116 4720 9120
rect 4656 9060 4660 9116
rect 4660 9060 4716 9116
rect 4716 9060 4720 9116
rect 4656 9056 4720 9060
rect 9744 9116 9808 9120
rect 9744 9060 9748 9116
rect 9748 9060 9804 9116
rect 9804 9060 9808 9116
rect 9744 9056 9808 9060
rect 9824 9116 9888 9120
rect 9824 9060 9828 9116
rect 9828 9060 9884 9116
rect 9884 9060 9888 9116
rect 9824 9056 9888 9060
rect 9904 9116 9968 9120
rect 9904 9060 9908 9116
rect 9908 9060 9964 9116
rect 9964 9060 9968 9116
rect 9904 9056 9968 9060
rect 9984 9116 10048 9120
rect 9984 9060 9988 9116
rect 9988 9060 10044 9116
rect 10044 9060 10048 9116
rect 9984 9056 10048 9060
rect 15072 9116 15136 9120
rect 15072 9060 15076 9116
rect 15076 9060 15132 9116
rect 15132 9060 15136 9116
rect 15072 9056 15136 9060
rect 15152 9116 15216 9120
rect 15152 9060 15156 9116
rect 15156 9060 15212 9116
rect 15212 9060 15216 9116
rect 15152 9056 15216 9060
rect 15232 9116 15296 9120
rect 15232 9060 15236 9116
rect 15236 9060 15292 9116
rect 15292 9060 15296 9116
rect 15232 9056 15296 9060
rect 15312 9116 15376 9120
rect 15312 9060 15316 9116
rect 15316 9060 15372 9116
rect 15372 9060 15376 9116
rect 15312 9056 15376 9060
rect 7080 8572 7144 8576
rect 7080 8516 7084 8572
rect 7084 8516 7140 8572
rect 7140 8516 7144 8572
rect 7080 8512 7144 8516
rect 7160 8572 7224 8576
rect 7160 8516 7164 8572
rect 7164 8516 7220 8572
rect 7220 8516 7224 8572
rect 7160 8512 7224 8516
rect 7240 8572 7304 8576
rect 7240 8516 7244 8572
rect 7244 8516 7300 8572
rect 7300 8516 7304 8572
rect 7240 8512 7304 8516
rect 7320 8572 7384 8576
rect 7320 8516 7324 8572
rect 7324 8516 7380 8572
rect 7380 8516 7384 8572
rect 7320 8512 7384 8516
rect 12408 8572 12472 8576
rect 12408 8516 12412 8572
rect 12412 8516 12468 8572
rect 12468 8516 12472 8572
rect 12408 8512 12472 8516
rect 12488 8572 12552 8576
rect 12488 8516 12492 8572
rect 12492 8516 12548 8572
rect 12548 8516 12552 8572
rect 12488 8512 12552 8516
rect 12568 8572 12632 8576
rect 12568 8516 12572 8572
rect 12572 8516 12628 8572
rect 12628 8516 12632 8572
rect 12568 8512 12632 8516
rect 12648 8572 12712 8576
rect 12648 8516 12652 8572
rect 12652 8516 12708 8572
rect 12708 8516 12712 8572
rect 12648 8512 12712 8516
rect 17736 8572 17800 8576
rect 17736 8516 17740 8572
rect 17740 8516 17796 8572
rect 17796 8516 17800 8572
rect 17736 8512 17800 8516
rect 17816 8572 17880 8576
rect 17816 8516 17820 8572
rect 17820 8516 17876 8572
rect 17876 8516 17880 8572
rect 17816 8512 17880 8516
rect 17896 8572 17960 8576
rect 17896 8516 17900 8572
rect 17900 8516 17956 8572
rect 17956 8516 17960 8572
rect 17896 8512 17960 8516
rect 17976 8572 18040 8576
rect 17976 8516 17980 8572
rect 17980 8516 18036 8572
rect 18036 8516 18040 8572
rect 17976 8512 18040 8516
rect 4416 8028 4480 8032
rect 4416 7972 4420 8028
rect 4420 7972 4476 8028
rect 4476 7972 4480 8028
rect 4416 7968 4480 7972
rect 4496 8028 4560 8032
rect 4496 7972 4500 8028
rect 4500 7972 4556 8028
rect 4556 7972 4560 8028
rect 4496 7968 4560 7972
rect 4576 8028 4640 8032
rect 4576 7972 4580 8028
rect 4580 7972 4636 8028
rect 4636 7972 4640 8028
rect 4576 7968 4640 7972
rect 4656 8028 4720 8032
rect 4656 7972 4660 8028
rect 4660 7972 4716 8028
rect 4716 7972 4720 8028
rect 4656 7968 4720 7972
rect 9744 8028 9808 8032
rect 9744 7972 9748 8028
rect 9748 7972 9804 8028
rect 9804 7972 9808 8028
rect 9744 7968 9808 7972
rect 9824 8028 9888 8032
rect 9824 7972 9828 8028
rect 9828 7972 9884 8028
rect 9884 7972 9888 8028
rect 9824 7968 9888 7972
rect 9904 8028 9968 8032
rect 9904 7972 9908 8028
rect 9908 7972 9964 8028
rect 9964 7972 9968 8028
rect 9904 7968 9968 7972
rect 9984 8028 10048 8032
rect 9984 7972 9988 8028
rect 9988 7972 10044 8028
rect 10044 7972 10048 8028
rect 9984 7968 10048 7972
rect 15072 8028 15136 8032
rect 15072 7972 15076 8028
rect 15076 7972 15132 8028
rect 15132 7972 15136 8028
rect 15072 7968 15136 7972
rect 15152 8028 15216 8032
rect 15152 7972 15156 8028
rect 15156 7972 15212 8028
rect 15212 7972 15216 8028
rect 15152 7968 15216 7972
rect 15232 8028 15296 8032
rect 15232 7972 15236 8028
rect 15236 7972 15292 8028
rect 15292 7972 15296 8028
rect 15232 7968 15296 7972
rect 15312 8028 15376 8032
rect 15312 7972 15316 8028
rect 15316 7972 15372 8028
rect 15372 7972 15376 8028
rect 15312 7968 15376 7972
rect 7080 7484 7144 7488
rect 7080 7428 7084 7484
rect 7084 7428 7140 7484
rect 7140 7428 7144 7484
rect 7080 7424 7144 7428
rect 7160 7484 7224 7488
rect 7160 7428 7164 7484
rect 7164 7428 7220 7484
rect 7220 7428 7224 7484
rect 7160 7424 7224 7428
rect 7240 7484 7304 7488
rect 7240 7428 7244 7484
rect 7244 7428 7300 7484
rect 7300 7428 7304 7484
rect 7240 7424 7304 7428
rect 7320 7484 7384 7488
rect 7320 7428 7324 7484
rect 7324 7428 7380 7484
rect 7380 7428 7384 7484
rect 7320 7424 7384 7428
rect 12408 7484 12472 7488
rect 12408 7428 12412 7484
rect 12412 7428 12468 7484
rect 12468 7428 12472 7484
rect 12408 7424 12472 7428
rect 12488 7484 12552 7488
rect 12488 7428 12492 7484
rect 12492 7428 12548 7484
rect 12548 7428 12552 7484
rect 12488 7424 12552 7428
rect 12568 7484 12632 7488
rect 12568 7428 12572 7484
rect 12572 7428 12628 7484
rect 12628 7428 12632 7484
rect 12568 7424 12632 7428
rect 12648 7484 12712 7488
rect 12648 7428 12652 7484
rect 12652 7428 12708 7484
rect 12708 7428 12712 7484
rect 12648 7424 12712 7428
rect 17736 7484 17800 7488
rect 17736 7428 17740 7484
rect 17740 7428 17796 7484
rect 17796 7428 17800 7484
rect 17736 7424 17800 7428
rect 17816 7484 17880 7488
rect 17816 7428 17820 7484
rect 17820 7428 17876 7484
rect 17876 7428 17880 7484
rect 17816 7424 17880 7428
rect 17896 7484 17960 7488
rect 17896 7428 17900 7484
rect 17900 7428 17956 7484
rect 17956 7428 17960 7484
rect 17896 7424 17960 7428
rect 17976 7484 18040 7488
rect 17976 7428 17980 7484
rect 17980 7428 18036 7484
rect 18036 7428 18040 7484
rect 17976 7424 18040 7428
rect 4416 6940 4480 6944
rect 4416 6884 4420 6940
rect 4420 6884 4476 6940
rect 4476 6884 4480 6940
rect 4416 6880 4480 6884
rect 4496 6940 4560 6944
rect 4496 6884 4500 6940
rect 4500 6884 4556 6940
rect 4556 6884 4560 6940
rect 4496 6880 4560 6884
rect 4576 6940 4640 6944
rect 4576 6884 4580 6940
rect 4580 6884 4636 6940
rect 4636 6884 4640 6940
rect 4576 6880 4640 6884
rect 4656 6940 4720 6944
rect 4656 6884 4660 6940
rect 4660 6884 4716 6940
rect 4716 6884 4720 6940
rect 4656 6880 4720 6884
rect 9744 6940 9808 6944
rect 9744 6884 9748 6940
rect 9748 6884 9804 6940
rect 9804 6884 9808 6940
rect 9744 6880 9808 6884
rect 9824 6940 9888 6944
rect 9824 6884 9828 6940
rect 9828 6884 9884 6940
rect 9884 6884 9888 6940
rect 9824 6880 9888 6884
rect 9904 6940 9968 6944
rect 9904 6884 9908 6940
rect 9908 6884 9964 6940
rect 9964 6884 9968 6940
rect 9904 6880 9968 6884
rect 9984 6940 10048 6944
rect 9984 6884 9988 6940
rect 9988 6884 10044 6940
rect 10044 6884 10048 6940
rect 9984 6880 10048 6884
rect 15072 6940 15136 6944
rect 15072 6884 15076 6940
rect 15076 6884 15132 6940
rect 15132 6884 15136 6940
rect 15072 6880 15136 6884
rect 15152 6940 15216 6944
rect 15152 6884 15156 6940
rect 15156 6884 15212 6940
rect 15212 6884 15216 6940
rect 15152 6880 15216 6884
rect 15232 6940 15296 6944
rect 15232 6884 15236 6940
rect 15236 6884 15292 6940
rect 15292 6884 15296 6940
rect 15232 6880 15296 6884
rect 15312 6940 15376 6944
rect 15312 6884 15316 6940
rect 15316 6884 15372 6940
rect 15372 6884 15376 6940
rect 15312 6880 15376 6884
rect 7080 6396 7144 6400
rect 7080 6340 7084 6396
rect 7084 6340 7140 6396
rect 7140 6340 7144 6396
rect 7080 6336 7144 6340
rect 7160 6396 7224 6400
rect 7160 6340 7164 6396
rect 7164 6340 7220 6396
rect 7220 6340 7224 6396
rect 7160 6336 7224 6340
rect 7240 6396 7304 6400
rect 7240 6340 7244 6396
rect 7244 6340 7300 6396
rect 7300 6340 7304 6396
rect 7240 6336 7304 6340
rect 7320 6396 7384 6400
rect 7320 6340 7324 6396
rect 7324 6340 7380 6396
rect 7380 6340 7384 6396
rect 7320 6336 7384 6340
rect 12408 6396 12472 6400
rect 12408 6340 12412 6396
rect 12412 6340 12468 6396
rect 12468 6340 12472 6396
rect 12408 6336 12472 6340
rect 12488 6396 12552 6400
rect 12488 6340 12492 6396
rect 12492 6340 12548 6396
rect 12548 6340 12552 6396
rect 12488 6336 12552 6340
rect 12568 6396 12632 6400
rect 12568 6340 12572 6396
rect 12572 6340 12628 6396
rect 12628 6340 12632 6396
rect 12568 6336 12632 6340
rect 12648 6396 12712 6400
rect 12648 6340 12652 6396
rect 12652 6340 12708 6396
rect 12708 6340 12712 6396
rect 12648 6336 12712 6340
rect 17736 6396 17800 6400
rect 17736 6340 17740 6396
rect 17740 6340 17796 6396
rect 17796 6340 17800 6396
rect 17736 6336 17800 6340
rect 17816 6396 17880 6400
rect 17816 6340 17820 6396
rect 17820 6340 17876 6396
rect 17876 6340 17880 6396
rect 17816 6336 17880 6340
rect 17896 6396 17960 6400
rect 17896 6340 17900 6396
rect 17900 6340 17956 6396
rect 17956 6340 17960 6396
rect 17896 6336 17960 6340
rect 17976 6396 18040 6400
rect 17976 6340 17980 6396
rect 17980 6340 18036 6396
rect 18036 6340 18040 6396
rect 17976 6336 18040 6340
rect 4416 5852 4480 5856
rect 4416 5796 4420 5852
rect 4420 5796 4476 5852
rect 4476 5796 4480 5852
rect 4416 5792 4480 5796
rect 4496 5852 4560 5856
rect 4496 5796 4500 5852
rect 4500 5796 4556 5852
rect 4556 5796 4560 5852
rect 4496 5792 4560 5796
rect 4576 5852 4640 5856
rect 4576 5796 4580 5852
rect 4580 5796 4636 5852
rect 4636 5796 4640 5852
rect 4576 5792 4640 5796
rect 4656 5852 4720 5856
rect 4656 5796 4660 5852
rect 4660 5796 4716 5852
rect 4716 5796 4720 5852
rect 4656 5792 4720 5796
rect 9744 5852 9808 5856
rect 9744 5796 9748 5852
rect 9748 5796 9804 5852
rect 9804 5796 9808 5852
rect 9744 5792 9808 5796
rect 9824 5852 9888 5856
rect 9824 5796 9828 5852
rect 9828 5796 9884 5852
rect 9884 5796 9888 5852
rect 9824 5792 9888 5796
rect 9904 5852 9968 5856
rect 9904 5796 9908 5852
rect 9908 5796 9964 5852
rect 9964 5796 9968 5852
rect 9904 5792 9968 5796
rect 9984 5852 10048 5856
rect 9984 5796 9988 5852
rect 9988 5796 10044 5852
rect 10044 5796 10048 5852
rect 9984 5792 10048 5796
rect 15072 5852 15136 5856
rect 15072 5796 15076 5852
rect 15076 5796 15132 5852
rect 15132 5796 15136 5852
rect 15072 5792 15136 5796
rect 15152 5852 15216 5856
rect 15152 5796 15156 5852
rect 15156 5796 15212 5852
rect 15212 5796 15216 5852
rect 15152 5792 15216 5796
rect 15232 5852 15296 5856
rect 15232 5796 15236 5852
rect 15236 5796 15292 5852
rect 15292 5796 15296 5852
rect 15232 5792 15296 5796
rect 15312 5852 15376 5856
rect 15312 5796 15316 5852
rect 15316 5796 15372 5852
rect 15372 5796 15376 5852
rect 15312 5792 15376 5796
rect 7080 5308 7144 5312
rect 7080 5252 7084 5308
rect 7084 5252 7140 5308
rect 7140 5252 7144 5308
rect 7080 5248 7144 5252
rect 7160 5308 7224 5312
rect 7160 5252 7164 5308
rect 7164 5252 7220 5308
rect 7220 5252 7224 5308
rect 7160 5248 7224 5252
rect 7240 5308 7304 5312
rect 7240 5252 7244 5308
rect 7244 5252 7300 5308
rect 7300 5252 7304 5308
rect 7240 5248 7304 5252
rect 7320 5308 7384 5312
rect 7320 5252 7324 5308
rect 7324 5252 7380 5308
rect 7380 5252 7384 5308
rect 7320 5248 7384 5252
rect 12408 5308 12472 5312
rect 12408 5252 12412 5308
rect 12412 5252 12468 5308
rect 12468 5252 12472 5308
rect 12408 5248 12472 5252
rect 12488 5308 12552 5312
rect 12488 5252 12492 5308
rect 12492 5252 12548 5308
rect 12548 5252 12552 5308
rect 12488 5248 12552 5252
rect 12568 5308 12632 5312
rect 12568 5252 12572 5308
rect 12572 5252 12628 5308
rect 12628 5252 12632 5308
rect 12568 5248 12632 5252
rect 12648 5308 12712 5312
rect 12648 5252 12652 5308
rect 12652 5252 12708 5308
rect 12708 5252 12712 5308
rect 12648 5248 12712 5252
rect 17736 5308 17800 5312
rect 17736 5252 17740 5308
rect 17740 5252 17796 5308
rect 17796 5252 17800 5308
rect 17736 5248 17800 5252
rect 17816 5308 17880 5312
rect 17816 5252 17820 5308
rect 17820 5252 17876 5308
rect 17876 5252 17880 5308
rect 17816 5248 17880 5252
rect 17896 5308 17960 5312
rect 17896 5252 17900 5308
rect 17900 5252 17956 5308
rect 17956 5252 17960 5308
rect 17896 5248 17960 5252
rect 17976 5308 18040 5312
rect 17976 5252 17980 5308
rect 17980 5252 18036 5308
rect 18036 5252 18040 5308
rect 17976 5248 18040 5252
rect 4416 4764 4480 4768
rect 4416 4708 4420 4764
rect 4420 4708 4476 4764
rect 4476 4708 4480 4764
rect 4416 4704 4480 4708
rect 4496 4764 4560 4768
rect 4496 4708 4500 4764
rect 4500 4708 4556 4764
rect 4556 4708 4560 4764
rect 4496 4704 4560 4708
rect 4576 4764 4640 4768
rect 4576 4708 4580 4764
rect 4580 4708 4636 4764
rect 4636 4708 4640 4764
rect 4576 4704 4640 4708
rect 4656 4764 4720 4768
rect 4656 4708 4660 4764
rect 4660 4708 4716 4764
rect 4716 4708 4720 4764
rect 4656 4704 4720 4708
rect 9744 4764 9808 4768
rect 9744 4708 9748 4764
rect 9748 4708 9804 4764
rect 9804 4708 9808 4764
rect 9744 4704 9808 4708
rect 9824 4764 9888 4768
rect 9824 4708 9828 4764
rect 9828 4708 9884 4764
rect 9884 4708 9888 4764
rect 9824 4704 9888 4708
rect 9904 4764 9968 4768
rect 9904 4708 9908 4764
rect 9908 4708 9964 4764
rect 9964 4708 9968 4764
rect 9904 4704 9968 4708
rect 9984 4764 10048 4768
rect 9984 4708 9988 4764
rect 9988 4708 10044 4764
rect 10044 4708 10048 4764
rect 9984 4704 10048 4708
rect 15072 4764 15136 4768
rect 15072 4708 15076 4764
rect 15076 4708 15132 4764
rect 15132 4708 15136 4764
rect 15072 4704 15136 4708
rect 15152 4764 15216 4768
rect 15152 4708 15156 4764
rect 15156 4708 15212 4764
rect 15212 4708 15216 4764
rect 15152 4704 15216 4708
rect 15232 4764 15296 4768
rect 15232 4708 15236 4764
rect 15236 4708 15292 4764
rect 15292 4708 15296 4764
rect 15232 4704 15296 4708
rect 15312 4764 15376 4768
rect 15312 4708 15316 4764
rect 15316 4708 15372 4764
rect 15372 4708 15376 4764
rect 15312 4704 15376 4708
rect 7080 4220 7144 4224
rect 7080 4164 7084 4220
rect 7084 4164 7140 4220
rect 7140 4164 7144 4220
rect 7080 4160 7144 4164
rect 7160 4220 7224 4224
rect 7160 4164 7164 4220
rect 7164 4164 7220 4220
rect 7220 4164 7224 4220
rect 7160 4160 7224 4164
rect 7240 4220 7304 4224
rect 7240 4164 7244 4220
rect 7244 4164 7300 4220
rect 7300 4164 7304 4220
rect 7240 4160 7304 4164
rect 7320 4220 7384 4224
rect 7320 4164 7324 4220
rect 7324 4164 7380 4220
rect 7380 4164 7384 4220
rect 7320 4160 7384 4164
rect 12408 4220 12472 4224
rect 12408 4164 12412 4220
rect 12412 4164 12468 4220
rect 12468 4164 12472 4220
rect 12408 4160 12472 4164
rect 12488 4220 12552 4224
rect 12488 4164 12492 4220
rect 12492 4164 12548 4220
rect 12548 4164 12552 4220
rect 12488 4160 12552 4164
rect 12568 4220 12632 4224
rect 12568 4164 12572 4220
rect 12572 4164 12628 4220
rect 12628 4164 12632 4220
rect 12568 4160 12632 4164
rect 12648 4220 12712 4224
rect 12648 4164 12652 4220
rect 12652 4164 12708 4220
rect 12708 4164 12712 4220
rect 12648 4160 12712 4164
rect 17736 4220 17800 4224
rect 17736 4164 17740 4220
rect 17740 4164 17796 4220
rect 17796 4164 17800 4220
rect 17736 4160 17800 4164
rect 17816 4220 17880 4224
rect 17816 4164 17820 4220
rect 17820 4164 17876 4220
rect 17876 4164 17880 4220
rect 17816 4160 17880 4164
rect 17896 4220 17960 4224
rect 17896 4164 17900 4220
rect 17900 4164 17956 4220
rect 17956 4164 17960 4220
rect 17896 4160 17960 4164
rect 17976 4220 18040 4224
rect 17976 4164 17980 4220
rect 17980 4164 18036 4220
rect 18036 4164 18040 4220
rect 17976 4160 18040 4164
rect 4416 3676 4480 3680
rect 4416 3620 4420 3676
rect 4420 3620 4476 3676
rect 4476 3620 4480 3676
rect 4416 3616 4480 3620
rect 4496 3676 4560 3680
rect 4496 3620 4500 3676
rect 4500 3620 4556 3676
rect 4556 3620 4560 3676
rect 4496 3616 4560 3620
rect 4576 3676 4640 3680
rect 4576 3620 4580 3676
rect 4580 3620 4636 3676
rect 4636 3620 4640 3676
rect 4576 3616 4640 3620
rect 4656 3676 4720 3680
rect 4656 3620 4660 3676
rect 4660 3620 4716 3676
rect 4716 3620 4720 3676
rect 4656 3616 4720 3620
rect 9744 3676 9808 3680
rect 9744 3620 9748 3676
rect 9748 3620 9804 3676
rect 9804 3620 9808 3676
rect 9744 3616 9808 3620
rect 9824 3676 9888 3680
rect 9824 3620 9828 3676
rect 9828 3620 9884 3676
rect 9884 3620 9888 3676
rect 9824 3616 9888 3620
rect 9904 3676 9968 3680
rect 9904 3620 9908 3676
rect 9908 3620 9964 3676
rect 9964 3620 9968 3676
rect 9904 3616 9968 3620
rect 9984 3676 10048 3680
rect 9984 3620 9988 3676
rect 9988 3620 10044 3676
rect 10044 3620 10048 3676
rect 9984 3616 10048 3620
rect 15072 3676 15136 3680
rect 15072 3620 15076 3676
rect 15076 3620 15132 3676
rect 15132 3620 15136 3676
rect 15072 3616 15136 3620
rect 15152 3676 15216 3680
rect 15152 3620 15156 3676
rect 15156 3620 15212 3676
rect 15212 3620 15216 3676
rect 15152 3616 15216 3620
rect 15232 3676 15296 3680
rect 15232 3620 15236 3676
rect 15236 3620 15292 3676
rect 15292 3620 15296 3676
rect 15232 3616 15296 3620
rect 15312 3676 15376 3680
rect 15312 3620 15316 3676
rect 15316 3620 15372 3676
rect 15372 3620 15376 3676
rect 15312 3616 15376 3620
rect 7080 3132 7144 3136
rect 7080 3076 7084 3132
rect 7084 3076 7140 3132
rect 7140 3076 7144 3132
rect 7080 3072 7144 3076
rect 7160 3132 7224 3136
rect 7160 3076 7164 3132
rect 7164 3076 7220 3132
rect 7220 3076 7224 3132
rect 7160 3072 7224 3076
rect 7240 3132 7304 3136
rect 7240 3076 7244 3132
rect 7244 3076 7300 3132
rect 7300 3076 7304 3132
rect 7240 3072 7304 3076
rect 7320 3132 7384 3136
rect 7320 3076 7324 3132
rect 7324 3076 7380 3132
rect 7380 3076 7384 3132
rect 7320 3072 7384 3076
rect 12408 3132 12472 3136
rect 12408 3076 12412 3132
rect 12412 3076 12468 3132
rect 12468 3076 12472 3132
rect 12408 3072 12472 3076
rect 12488 3132 12552 3136
rect 12488 3076 12492 3132
rect 12492 3076 12548 3132
rect 12548 3076 12552 3132
rect 12488 3072 12552 3076
rect 12568 3132 12632 3136
rect 12568 3076 12572 3132
rect 12572 3076 12628 3132
rect 12628 3076 12632 3132
rect 12568 3072 12632 3076
rect 12648 3132 12712 3136
rect 12648 3076 12652 3132
rect 12652 3076 12708 3132
rect 12708 3076 12712 3132
rect 12648 3072 12712 3076
rect 17736 3132 17800 3136
rect 17736 3076 17740 3132
rect 17740 3076 17796 3132
rect 17796 3076 17800 3132
rect 17736 3072 17800 3076
rect 17816 3132 17880 3136
rect 17816 3076 17820 3132
rect 17820 3076 17876 3132
rect 17876 3076 17880 3132
rect 17816 3072 17880 3076
rect 17896 3132 17960 3136
rect 17896 3076 17900 3132
rect 17900 3076 17956 3132
rect 17956 3076 17960 3132
rect 17896 3072 17960 3076
rect 17976 3132 18040 3136
rect 17976 3076 17980 3132
rect 17980 3076 18036 3132
rect 18036 3076 18040 3132
rect 17976 3072 18040 3076
rect 4416 2588 4480 2592
rect 4416 2532 4420 2588
rect 4420 2532 4476 2588
rect 4476 2532 4480 2588
rect 4416 2528 4480 2532
rect 4496 2588 4560 2592
rect 4496 2532 4500 2588
rect 4500 2532 4556 2588
rect 4556 2532 4560 2588
rect 4496 2528 4560 2532
rect 4576 2588 4640 2592
rect 4576 2532 4580 2588
rect 4580 2532 4636 2588
rect 4636 2532 4640 2588
rect 4576 2528 4640 2532
rect 4656 2588 4720 2592
rect 4656 2532 4660 2588
rect 4660 2532 4716 2588
rect 4716 2532 4720 2588
rect 4656 2528 4720 2532
rect 9744 2588 9808 2592
rect 9744 2532 9748 2588
rect 9748 2532 9804 2588
rect 9804 2532 9808 2588
rect 9744 2528 9808 2532
rect 9824 2588 9888 2592
rect 9824 2532 9828 2588
rect 9828 2532 9884 2588
rect 9884 2532 9888 2588
rect 9824 2528 9888 2532
rect 9904 2588 9968 2592
rect 9904 2532 9908 2588
rect 9908 2532 9964 2588
rect 9964 2532 9968 2588
rect 9904 2528 9968 2532
rect 9984 2588 10048 2592
rect 9984 2532 9988 2588
rect 9988 2532 10044 2588
rect 10044 2532 10048 2588
rect 9984 2528 10048 2532
rect 15072 2588 15136 2592
rect 15072 2532 15076 2588
rect 15076 2532 15132 2588
rect 15132 2532 15136 2588
rect 15072 2528 15136 2532
rect 15152 2588 15216 2592
rect 15152 2532 15156 2588
rect 15156 2532 15212 2588
rect 15212 2532 15216 2588
rect 15152 2528 15216 2532
rect 15232 2588 15296 2592
rect 15232 2532 15236 2588
rect 15236 2532 15292 2588
rect 15292 2532 15296 2588
rect 15232 2528 15296 2532
rect 15312 2588 15376 2592
rect 15312 2532 15316 2588
rect 15316 2532 15372 2588
rect 15372 2532 15376 2588
rect 15312 2528 15376 2532
rect 7080 2044 7144 2048
rect 7080 1988 7084 2044
rect 7084 1988 7140 2044
rect 7140 1988 7144 2044
rect 7080 1984 7144 1988
rect 7160 2044 7224 2048
rect 7160 1988 7164 2044
rect 7164 1988 7220 2044
rect 7220 1988 7224 2044
rect 7160 1984 7224 1988
rect 7240 2044 7304 2048
rect 7240 1988 7244 2044
rect 7244 1988 7300 2044
rect 7300 1988 7304 2044
rect 7240 1984 7304 1988
rect 7320 2044 7384 2048
rect 7320 1988 7324 2044
rect 7324 1988 7380 2044
rect 7380 1988 7384 2044
rect 7320 1984 7384 1988
rect 12408 2044 12472 2048
rect 12408 1988 12412 2044
rect 12412 1988 12468 2044
rect 12468 1988 12472 2044
rect 12408 1984 12472 1988
rect 12488 2044 12552 2048
rect 12488 1988 12492 2044
rect 12492 1988 12548 2044
rect 12548 1988 12552 2044
rect 12488 1984 12552 1988
rect 12568 2044 12632 2048
rect 12568 1988 12572 2044
rect 12572 1988 12628 2044
rect 12628 1988 12632 2044
rect 12568 1984 12632 1988
rect 12648 2044 12712 2048
rect 12648 1988 12652 2044
rect 12652 1988 12708 2044
rect 12708 1988 12712 2044
rect 12648 1984 12712 1988
rect 17736 2044 17800 2048
rect 17736 1988 17740 2044
rect 17740 1988 17796 2044
rect 17796 1988 17800 2044
rect 17736 1984 17800 1988
rect 17816 2044 17880 2048
rect 17816 1988 17820 2044
rect 17820 1988 17876 2044
rect 17876 1988 17880 2044
rect 17816 1984 17880 1988
rect 17896 2044 17960 2048
rect 17896 1988 17900 2044
rect 17900 1988 17956 2044
rect 17956 1988 17960 2044
rect 17896 1984 17960 1988
rect 17976 2044 18040 2048
rect 17976 1988 17980 2044
rect 17980 1988 18036 2044
rect 18036 1988 18040 2044
rect 17976 1984 18040 1988
rect 4416 1500 4480 1504
rect 4416 1444 4420 1500
rect 4420 1444 4476 1500
rect 4476 1444 4480 1500
rect 4416 1440 4480 1444
rect 4496 1500 4560 1504
rect 4496 1444 4500 1500
rect 4500 1444 4556 1500
rect 4556 1444 4560 1500
rect 4496 1440 4560 1444
rect 4576 1500 4640 1504
rect 4576 1444 4580 1500
rect 4580 1444 4636 1500
rect 4636 1444 4640 1500
rect 4576 1440 4640 1444
rect 4656 1500 4720 1504
rect 4656 1444 4660 1500
rect 4660 1444 4716 1500
rect 4716 1444 4720 1500
rect 4656 1440 4720 1444
rect 9744 1500 9808 1504
rect 9744 1444 9748 1500
rect 9748 1444 9804 1500
rect 9804 1444 9808 1500
rect 9744 1440 9808 1444
rect 9824 1500 9888 1504
rect 9824 1444 9828 1500
rect 9828 1444 9884 1500
rect 9884 1444 9888 1500
rect 9824 1440 9888 1444
rect 9904 1500 9968 1504
rect 9904 1444 9908 1500
rect 9908 1444 9964 1500
rect 9964 1444 9968 1500
rect 9904 1440 9968 1444
rect 9984 1500 10048 1504
rect 9984 1444 9988 1500
rect 9988 1444 10044 1500
rect 10044 1444 10048 1500
rect 9984 1440 10048 1444
rect 15072 1500 15136 1504
rect 15072 1444 15076 1500
rect 15076 1444 15132 1500
rect 15132 1444 15136 1500
rect 15072 1440 15136 1444
rect 15152 1500 15216 1504
rect 15152 1444 15156 1500
rect 15156 1444 15212 1500
rect 15212 1444 15216 1500
rect 15152 1440 15216 1444
rect 15232 1500 15296 1504
rect 15232 1444 15236 1500
rect 15236 1444 15292 1500
rect 15292 1444 15296 1500
rect 15232 1440 15296 1444
rect 15312 1500 15376 1504
rect 15312 1444 15316 1500
rect 15316 1444 15372 1500
rect 15372 1444 15376 1500
rect 15312 1440 15376 1444
rect 7080 956 7144 960
rect 7080 900 7084 956
rect 7084 900 7140 956
rect 7140 900 7144 956
rect 7080 896 7144 900
rect 7160 956 7224 960
rect 7160 900 7164 956
rect 7164 900 7220 956
rect 7220 900 7224 956
rect 7160 896 7224 900
rect 7240 956 7304 960
rect 7240 900 7244 956
rect 7244 900 7300 956
rect 7300 900 7304 956
rect 7240 896 7304 900
rect 7320 956 7384 960
rect 7320 900 7324 956
rect 7324 900 7380 956
rect 7380 900 7384 956
rect 7320 896 7384 900
rect 12408 956 12472 960
rect 12408 900 12412 956
rect 12412 900 12468 956
rect 12468 900 12472 956
rect 12408 896 12472 900
rect 12488 956 12552 960
rect 12488 900 12492 956
rect 12492 900 12548 956
rect 12548 900 12552 956
rect 12488 896 12552 900
rect 12568 956 12632 960
rect 12568 900 12572 956
rect 12572 900 12628 956
rect 12628 900 12632 956
rect 12568 896 12632 900
rect 12648 956 12712 960
rect 12648 900 12652 956
rect 12652 900 12708 956
rect 12708 900 12712 956
rect 12648 896 12712 900
rect 17736 956 17800 960
rect 17736 900 17740 956
rect 17740 900 17796 956
rect 17796 900 17800 956
rect 17736 896 17800 900
rect 17816 956 17880 960
rect 17816 900 17820 956
rect 17820 900 17876 956
rect 17876 900 17880 956
rect 17816 896 17880 900
rect 17896 956 17960 960
rect 17896 900 17900 956
rect 17900 900 17956 956
rect 17956 900 17960 956
rect 17896 896 17960 900
rect 17976 956 18040 960
rect 17976 900 17980 956
rect 17980 900 18036 956
rect 18036 900 18040 956
rect 17976 896 18040 900
<< metal4 >>
rect 4408 22176 4728 22192
rect 4408 22112 4416 22176
rect 4480 22112 4496 22176
rect 4560 22112 4576 22176
rect 4640 22112 4656 22176
rect 4720 22112 4728 22176
rect 4408 21088 4728 22112
rect 4408 21024 4416 21088
rect 4480 21024 4496 21088
rect 4560 21024 4576 21088
rect 4640 21024 4656 21088
rect 4720 21024 4728 21088
rect 4408 20838 4728 21024
rect 4408 20602 4450 20838
rect 4686 20602 4728 20838
rect 4408 20000 4728 20602
rect 4408 19936 4416 20000
rect 4480 19936 4496 20000
rect 4560 19936 4576 20000
rect 4640 19936 4656 20000
rect 4720 19936 4728 20000
rect 4408 18912 4728 19936
rect 4408 18848 4416 18912
rect 4480 18848 4496 18912
rect 4560 18848 4576 18912
rect 4640 18848 4656 18912
rect 4720 18848 4728 18912
rect 4408 17824 4728 18848
rect 4408 17760 4416 17824
rect 4480 17760 4496 17824
rect 4560 17760 4576 17824
rect 4640 17760 4656 17824
rect 4720 17760 4728 17824
rect 4408 16736 4728 17760
rect 4408 16672 4416 16736
rect 4480 16672 4496 16736
rect 4560 16672 4576 16736
rect 4640 16672 4656 16736
rect 4720 16672 4728 16736
rect 4408 15648 4728 16672
rect 4408 15584 4416 15648
rect 4480 15584 4496 15648
rect 4560 15584 4576 15648
rect 4640 15584 4656 15648
rect 4720 15584 4728 15648
rect 4408 14560 4728 15584
rect 4408 14496 4416 14560
rect 4480 14496 4496 14560
rect 4560 14496 4576 14560
rect 4640 14496 4656 14560
rect 4720 14496 4728 14560
rect 4408 13472 4728 14496
rect 4408 13408 4416 13472
rect 4480 13408 4496 13472
rect 4560 13408 4576 13472
rect 4640 13408 4656 13472
rect 4720 13408 4728 13472
rect 4408 12384 4728 13408
rect 4408 12320 4416 12384
rect 4480 12320 4496 12384
rect 4560 12320 4576 12384
rect 4640 12320 4656 12384
rect 4720 12320 4728 12384
rect 4408 11296 4728 12320
rect 4408 11232 4416 11296
rect 4480 11232 4496 11296
rect 4560 11232 4576 11296
rect 4640 11232 4656 11296
rect 4720 11232 4728 11296
rect 4408 10208 4728 11232
rect 4408 10144 4416 10208
rect 4480 10144 4496 10208
rect 4560 10144 4576 10208
rect 4640 10144 4656 10208
rect 4720 10144 4728 10208
rect 4408 9120 4728 10144
rect 4408 9056 4416 9120
rect 4480 9056 4496 9120
rect 4560 9056 4576 9120
rect 4640 9056 4656 9120
rect 4720 9056 4728 9120
rect 4408 8032 4728 9056
rect 4408 7968 4416 8032
rect 4480 7968 4496 8032
rect 4560 7968 4576 8032
rect 4640 7968 4656 8032
rect 4720 7968 4728 8032
rect 4408 6944 4728 7968
rect 4408 6880 4416 6944
rect 4480 6880 4496 6944
rect 4560 6880 4576 6944
rect 4640 6880 4656 6944
rect 4720 6880 4728 6944
rect 4408 5856 4728 6880
rect 4408 5792 4416 5856
rect 4480 5792 4496 5856
rect 4560 5792 4576 5856
rect 4640 5792 4656 5856
rect 4720 5792 4728 5856
rect 4408 4768 4728 5792
rect 4408 4704 4416 4768
rect 4480 4704 4496 4768
rect 4560 4704 4576 4768
rect 4640 4704 4656 4768
rect 4720 4704 4728 4768
rect 4408 3680 4728 4704
rect 4408 3616 4416 3680
rect 4480 3616 4496 3680
rect 4560 3616 4576 3680
rect 4640 3616 4656 3680
rect 4720 3616 4728 3680
rect 4408 2592 4728 3616
rect 4408 2528 4416 2592
rect 4480 2528 4496 2592
rect 4560 2528 4576 2592
rect 4640 2528 4656 2592
rect 4720 2528 4728 2592
rect 4408 1504 4728 2528
rect 4408 1440 4416 1504
rect 4480 1440 4496 1504
rect 4560 1440 4576 1504
rect 4640 1440 4656 1504
rect 4720 1440 4728 1504
rect 4408 880 4728 1440
rect 7072 21632 7392 22192
rect 7072 21568 7080 21632
rect 7144 21568 7160 21632
rect 7224 21568 7240 21632
rect 7304 21568 7320 21632
rect 7384 21568 7392 21632
rect 7072 20544 7392 21568
rect 7072 20480 7080 20544
rect 7144 20480 7160 20544
rect 7224 20480 7240 20544
rect 7304 20480 7320 20544
rect 7384 20480 7392 20544
rect 7072 19456 7392 20480
rect 7072 19392 7080 19456
rect 7144 19392 7160 19456
rect 7224 19392 7240 19456
rect 7304 19392 7320 19456
rect 7384 19392 7392 19456
rect 7072 18368 7392 19392
rect 7072 18304 7080 18368
rect 7144 18304 7160 18368
rect 7224 18304 7240 18368
rect 7304 18304 7320 18368
rect 7384 18304 7392 18368
rect 7072 17280 7392 18304
rect 7072 17216 7080 17280
rect 7144 17216 7160 17280
rect 7224 17216 7240 17280
rect 7304 17216 7320 17280
rect 7384 17216 7392 17280
rect 7072 16192 7392 17216
rect 7072 16128 7080 16192
rect 7144 16128 7160 16192
rect 7224 16128 7240 16192
rect 7304 16128 7320 16192
rect 7384 16128 7392 16192
rect 7072 15104 7392 16128
rect 7072 15040 7080 15104
rect 7144 15040 7160 15104
rect 7224 15040 7240 15104
rect 7304 15040 7320 15104
rect 7384 15040 7392 15104
rect 7072 14016 7392 15040
rect 7072 13952 7080 14016
rect 7144 13952 7160 14016
rect 7224 13952 7240 14016
rect 7304 13952 7320 14016
rect 7384 13952 7392 14016
rect 7072 12928 7392 13952
rect 7072 12864 7080 12928
rect 7144 12864 7160 12928
rect 7224 12864 7240 12928
rect 7304 12864 7320 12928
rect 7384 12864 7392 12928
rect 7072 11840 7392 12864
rect 7072 11776 7080 11840
rect 7144 11776 7160 11840
rect 7224 11776 7240 11840
rect 7304 11776 7320 11840
rect 7384 11776 7392 11840
rect 7072 10752 7392 11776
rect 7072 10688 7080 10752
rect 7144 10688 7160 10752
rect 7224 10688 7240 10752
rect 7304 10688 7320 10752
rect 7384 10688 7392 10752
rect 7072 9664 7392 10688
rect 7072 9600 7080 9664
rect 7144 9600 7160 9664
rect 7224 9600 7240 9664
rect 7304 9600 7320 9664
rect 7384 9600 7392 9664
rect 7072 8576 7392 9600
rect 7072 8512 7080 8576
rect 7144 8512 7160 8576
rect 7224 8512 7240 8576
rect 7304 8512 7320 8576
rect 7384 8512 7392 8576
rect 7072 7488 7392 8512
rect 7072 7424 7080 7488
rect 7144 7424 7160 7488
rect 7224 7424 7240 7488
rect 7304 7424 7320 7488
rect 7384 7424 7392 7488
rect 7072 6400 7392 7424
rect 7072 6336 7080 6400
rect 7144 6336 7160 6400
rect 7224 6336 7240 6400
rect 7304 6336 7320 6400
rect 7384 6336 7392 6400
rect 7072 5312 7392 6336
rect 7072 5248 7080 5312
rect 7144 5248 7160 5312
rect 7224 5248 7240 5312
rect 7304 5248 7320 5312
rect 7384 5248 7392 5312
rect 7072 4224 7392 5248
rect 7072 4160 7080 4224
rect 7144 4160 7160 4224
rect 7224 4160 7240 4224
rect 7304 4160 7320 4224
rect 7384 4160 7392 4224
rect 7072 3136 7392 4160
rect 7072 3072 7080 3136
rect 7144 3072 7160 3136
rect 7224 3072 7240 3136
rect 7304 3072 7320 3136
rect 7384 3072 7392 3136
rect 7072 2838 7392 3072
rect 7072 2602 7114 2838
rect 7350 2602 7392 2838
rect 7072 2048 7392 2602
rect 7072 1984 7080 2048
rect 7144 1984 7160 2048
rect 7224 1984 7240 2048
rect 7304 1984 7320 2048
rect 7384 1984 7392 2048
rect 7072 960 7392 1984
rect 7072 896 7080 960
rect 7144 896 7160 960
rect 7224 896 7240 960
rect 7304 896 7320 960
rect 7384 896 7392 960
rect 7072 880 7392 896
rect 9736 22176 10056 22192
rect 9736 22112 9744 22176
rect 9808 22112 9824 22176
rect 9888 22112 9904 22176
rect 9968 22112 9984 22176
rect 10048 22112 10056 22176
rect 9736 21088 10056 22112
rect 9736 21024 9744 21088
rect 9808 21024 9824 21088
rect 9888 21024 9904 21088
rect 9968 21024 9984 21088
rect 10048 21024 10056 21088
rect 9736 20838 10056 21024
rect 9736 20602 9778 20838
rect 10014 20602 10056 20838
rect 9736 20000 10056 20602
rect 9736 19936 9744 20000
rect 9808 19936 9824 20000
rect 9888 19936 9904 20000
rect 9968 19936 9984 20000
rect 10048 19936 10056 20000
rect 9736 18912 10056 19936
rect 9736 18848 9744 18912
rect 9808 18848 9824 18912
rect 9888 18848 9904 18912
rect 9968 18848 9984 18912
rect 10048 18848 10056 18912
rect 9736 17824 10056 18848
rect 9736 17760 9744 17824
rect 9808 17760 9824 17824
rect 9888 17760 9904 17824
rect 9968 17760 9984 17824
rect 10048 17760 10056 17824
rect 9736 16736 10056 17760
rect 9736 16672 9744 16736
rect 9808 16672 9824 16736
rect 9888 16672 9904 16736
rect 9968 16672 9984 16736
rect 10048 16672 10056 16736
rect 9736 15648 10056 16672
rect 9736 15584 9744 15648
rect 9808 15584 9824 15648
rect 9888 15584 9904 15648
rect 9968 15584 9984 15648
rect 10048 15584 10056 15648
rect 9736 14560 10056 15584
rect 9736 14496 9744 14560
rect 9808 14496 9824 14560
rect 9888 14496 9904 14560
rect 9968 14496 9984 14560
rect 10048 14496 10056 14560
rect 9736 13472 10056 14496
rect 9736 13408 9744 13472
rect 9808 13408 9824 13472
rect 9888 13408 9904 13472
rect 9968 13408 9984 13472
rect 10048 13408 10056 13472
rect 9736 12384 10056 13408
rect 9736 12320 9744 12384
rect 9808 12320 9824 12384
rect 9888 12320 9904 12384
rect 9968 12320 9984 12384
rect 10048 12320 10056 12384
rect 9736 11296 10056 12320
rect 9736 11232 9744 11296
rect 9808 11232 9824 11296
rect 9888 11232 9904 11296
rect 9968 11232 9984 11296
rect 10048 11232 10056 11296
rect 9736 10208 10056 11232
rect 9736 10144 9744 10208
rect 9808 10144 9824 10208
rect 9888 10144 9904 10208
rect 9968 10144 9984 10208
rect 10048 10144 10056 10208
rect 9736 9120 10056 10144
rect 9736 9056 9744 9120
rect 9808 9056 9824 9120
rect 9888 9056 9904 9120
rect 9968 9056 9984 9120
rect 10048 9056 10056 9120
rect 9736 8032 10056 9056
rect 9736 7968 9744 8032
rect 9808 7968 9824 8032
rect 9888 7968 9904 8032
rect 9968 7968 9984 8032
rect 10048 7968 10056 8032
rect 9736 6944 10056 7968
rect 9736 6880 9744 6944
rect 9808 6880 9824 6944
rect 9888 6880 9904 6944
rect 9968 6880 9984 6944
rect 10048 6880 10056 6944
rect 9736 5856 10056 6880
rect 9736 5792 9744 5856
rect 9808 5792 9824 5856
rect 9888 5792 9904 5856
rect 9968 5792 9984 5856
rect 10048 5792 10056 5856
rect 9736 4768 10056 5792
rect 9736 4704 9744 4768
rect 9808 4704 9824 4768
rect 9888 4704 9904 4768
rect 9968 4704 9984 4768
rect 10048 4704 10056 4768
rect 9736 3680 10056 4704
rect 9736 3616 9744 3680
rect 9808 3616 9824 3680
rect 9888 3616 9904 3680
rect 9968 3616 9984 3680
rect 10048 3616 10056 3680
rect 9736 2592 10056 3616
rect 9736 2528 9744 2592
rect 9808 2528 9824 2592
rect 9888 2528 9904 2592
rect 9968 2528 9984 2592
rect 10048 2528 10056 2592
rect 9736 1504 10056 2528
rect 9736 1440 9744 1504
rect 9808 1440 9824 1504
rect 9888 1440 9904 1504
rect 9968 1440 9984 1504
rect 10048 1440 10056 1504
rect 9736 880 10056 1440
rect 12400 21632 12720 22192
rect 12400 21568 12408 21632
rect 12472 21568 12488 21632
rect 12552 21568 12568 21632
rect 12632 21568 12648 21632
rect 12712 21568 12720 21632
rect 12400 20544 12720 21568
rect 12400 20480 12408 20544
rect 12472 20480 12488 20544
rect 12552 20480 12568 20544
rect 12632 20480 12648 20544
rect 12712 20480 12720 20544
rect 12400 19456 12720 20480
rect 12400 19392 12408 19456
rect 12472 19392 12488 19456
rect 12552 19392 12568 19456
rect 12632 19392 12648 19456
rect 12712 19392 12720 19456
rect 12400 18368 12720 19392
rect 12400 18304 12408 18368
rect 12472 18304 12488 18368
rect 12552 18304 12568 18368
rect 12632 18304 12648 18368
rect 12712 18304 12720 18368
rect 12400 17280 12720 18304
rect 12400 17216 12408 17280
rect 12472 17216 12488 17280
rect 12552 17216 12568 17280
rect 12632 17216 12648 17280
rect 12712 17216 12720 17280
rect 12400 16192 12720 17216
rect 12400 16128 12408 16192
rect 12472 16128 12488 16192
rect 12552 16128 12568 16192
rect 12632 16128 12648 16192
rect 12712 16128 12720 16192
rect 12400 15104 12720 16128
rect 12400 15040 12408 15104
rect 12472 15040 12488 15104
rect 12552 15040 12568 15104
rect 12632 15040 12648 15104
rect 12712 15040 12720 15104
rect 12400 14016 12720 15040
rect 12400 13952 12408 14016
rect 12472 13952 12488 14016
rect 12552 13952 12568 14016
rect 12632 13952 12648 14016
rect 12712 13952 12720 14016
rect 12400 12928 12720 13952
rect 12400 12864 12408 12928
rect 12472 12864 12488 12928
rect 12552 12864 12568 12928
rect 12632 12864 12648 12928
rect 12712 12864 12720 12928
rect 12400 11840 12720 12864
rect 12400 11776 12408 11840
rect 12472 11776 12488 11840
rect 12552 11776 12568 11840
rect 12632 11776 12648 11840
rect 12712 11776 12720 11840
rect 12400 10752 12720 11776
rect 12400 10688 12408 10752
rect 12472 10688 12488 10752
rect 12552 10688 12568 10752
rect 12632 10688 12648 10752
rect 12712 10688 12720 10752
rect 12400 9664 12720 10688
rect 12400 9600 12408 9664
rect 12472 9600 12488 9664
rect 12552 9600 12568 9664
rect 12632 9600 12648 9664
rect 12712 9600 12720 9664
rect 12400 8576 12720 9600
rect 12400 8512 12408 8576
rect 12472 8512 12488 8576
rect 12552 8512 12568 8576
rect 12632 8512 12648 8576
rect 12712 8512 12720 8576
rect 12400 7488 12720 8512
rect 12400 7424 12408 7488
rect 12472 7424 12488 7488
rect 12552 7424 12568 7488
rect 12632 7424 12648 7488
rect 12712 7424 12720 7488
rect 12400 6400 12720 7424
rect 12400 6336 12408 6400
rect 12472 6336 12488 6400
rect 12552 6336 12568 6400
rect 12632 6336 12648 6400
rect 12712 6336 12720 6400
rect 12400 5312 12720 6336
rect 12400 5248 12408 5312
rect 12472 5248 12488 5312
rect 12552 5248 12568 5312
rect 12632 5248 12648 5312
rect 12712 5248 12720 5312
rect 12400 4224 12720 5248
rect 12400 4160 12408 4224
rect 12472 4160 12488 4224
rect 12552 4160 12568 4224
rect 12632 4160 12648 4224
rect 12712 4160 12720 4224
rect 12400 3136 12720 4160
rect 12400 3072 12408 3136
rect 12472 3072 12488 3136
rect 12552 3072 12568 3136
rect 12632 3072 12648 3136
rect 12712 3072 12720 3136
rect 12400 2838 12720 3072
rect 12400 2602 12442 2838
rect 12678 2602 12720 2838
rect 12400 2048 12720 2602
rect 12400 1984 12408 2048
rect 12472 1984 12488 2048
rect 12552 1984 12568 2048
rect 12632 1984 12648 2048
rect 12712 1984 12720 2048
rect 12400 960 12720 1984
rect 12400 896 12408 960
rect 12472 896 12488 960
rect 12552 896 12568 960
rect 12632 896 12648 960
rect 12712 896 12720 960
rect 12400 880 12720 896
rect 15064 22176 15384 22192
rect 15064 22112 15072 22176
rect 15136 22112 15152 22176
rect 15216 22112 15232 22176
rect 15296 22112 15312 22176
rect 15376 22112 15384 22176
rect 15064 21088 15384 22112
rect 15064 21024 15072 21088
rect 15136 21024 15152 21088
rect 15216 21024 15232 21088
rect 15296 21024 15312 21088
rect 15376 21024 15384 21088
rect 15064 20838 15384 21024
rect 15064 20602 15106 20838
rect 15342 20602 15384 20838
rect 15064 20000 15384 20602
rect 15064 19936 15072 20000
rect 15136 19936 15152 20000
rect 15216 19936 15232 20000
rect 15296 19936 15312 20000
rect 15376 19936 15384 20000
rect 15064 18912 15384 19936
rect 15064 18848 15072 18912
rect 15136 18848 15152 18912
rect 15216 18848 15232 18912
rect 15296 18848 15312 18912
rect 15376 18848 15384 18912
rect 15064 17824 15384 18848
rect 15064 17760 15072 17824
rect 15136 17760 15152 17824
rect 15216 17760 15232 17824
rect 15296 17760 15312 17824
rect 15376 17760 15384 17824
rect 15064 16736 15384 17760
rect 15064 16672 15072 16736
rect 15136 16672 15152 16736
rect 15216 16672 15232 16736
rect 15296 16672 15312 16736
rect 15376 16672 15384 16736
rect 15064 15648 15384 16672
rect 15064 15584 15072 15648
rect 15136 15584 15152 15648
rect 15216 15584 15232 15648
rect 15296 15584 15312 15648
rect 15376 15584 15384 15648
rect 15064 14560 15384 15584
rect 15064 14496 15072 14560
rect 15136 14496 15152 14560
rect 15216 14496 15232 14560
rect 15296 14496 15312 14560
rect 15376 14496 15384 14560
rect 15064 13472 15384 14496
rect 15064 13408 15072 13472
rect 15136 13408 15152 13472
rect 15216 13408 15232 13472
rect 15296 13408 15312 13472
rect 15376 13408 15384 13472
rect 15064 12384 15384 13408
rect 15064 12320 15072 12384
rect 15136 12320 15152 12384
rect 15216 12320 15232 12384
rect 15296 12320 15312 12384
rect 15376 12320 15384 12384
rect 15064 11296 15384 12320
rect 15064 11232 15072 11296
rect 15136 11232 15152 11296
rect 15216 11232 15232 11296
rect 15296 11232 15312 11296
rect 15376 11232 15384 11296
rect 15064 10208 15384 11232
rect 15064 10144 15072 10208
rect 15136 10144 15152 10208
rect 15216 10144 15232 10208
rect 15296 10144 15312 10208
rect 15376 10144 15384 10208
rect 15064 9120 15384 10144
rect 15064 9056 15072 9120
rect 15136 9056 15152 9120
rect 15216 9056 15232 9120
rect 15296 9056 15312 9120
rect 15376 9056 15384 9120
rect 15064 8032 15384 9056
rect 15064 7968 15072 8032
rect 15136 7968 15152 8032
rect 15216 7968 15232 8032
rect 15296 7968 15312 8032
rect 15376 7968 15384 8032
rect 15064 6944 15384 7968
rect 15064 6880 15072 6944
rect 15136 6880 15152 6944
rect 15216 6880 15232 6944
rect 15296 6880 15312 6944
rect 15376 6880 15384 6944
rect 15064 5856 15384 6880
rect 15064 5792 15072 5856
rect 15136 5792 15152 5856
rect 15216 5792 15232 5856
rect 15296 5792 15312 5856
rect 15376 5792 15384 5856
rect 15064 4768 15384 5792
rect 15064 4704 15072 4768
rect 15136 4704 15152 4768
rect 15216 4704 15232 4768
rect 15296 4704 15312 4768
rect 15376 4704 15384 4768
rect 15064 3680 15384 4704
rect 15064 3616 15072 3680
rect 15136 3616 15152 3680
rect 15216 3616 15232 3680
rect 15296 3616 15312 3680
rect 15376 3616 15384 3680
rect 15064 2592 15384 3616
rect 15064 2528 15072 2592
rect 15136 2528 15152 2592
rect 15216 2528 15232 2592
rect 15296 2528 15312 2592
rect 15376 2528 15384 2592
rect 15064 1504 15384 2528
rect 15064 1440 15072 1504
rect 15136 1440 15152 1504
rect 15216 1440 15232 1504
rect 15296 1440 15312 1504
rect 15376 1440 15384 1504
rect 15064 880 15384 1440
rect 17728 21632 18048 22192
rect 17728 21568 17736 21632
rect 17800 21568 17816 21632
rect 17880 21568 17896 21632
rect 17960 21568 17976 21632
rect 18040 21568 18048 21632
rect 17728 20544 18048 21568
rect 17728 20480 17736 20544
rect 17800 20480 17816 20544
rect 17880 20480 17896 20544
rect 17960 20480 17976 20544
rect 18040 20480 18048 20544
rect 17728 19456 18048 20480
rect 17728 19392 17736 19456
rect 17800 19392 17816 19456
rect 17880 19392 17896 19456
rect 17960 19392 17976 19456
rect 18040 19392 18048 19456
rect 17728 18368 18048 19392
rect 17728 18304 17736 18368
rect 17800 18304 17816 18368
rect 17880 18304 17896 18368
rect 17960 18304 17976 18368
rect 18040 18304 18048 18368
rect 17728 17280 18048 18304
rect 17728 17216 17736 17280
rect 17800 17216 17816 17280
rect 17880 17216 17896 17280
rect 17960 17216 17976 17280
rect 18040 17216 18048 17280
rect 17728 16192 18048 17216
rect 17728 16128 17736 16192
rect 17800 16128 17816 16192
rect 17880 16128 17896 16192
rect 17960 16128 17976 16192
rect 18040 16128 18048 16192
rect 17728 15104 18048 16128
rect 17728 15040 17736 15104
rect 17800 15040 17816 15104
rect 17880 15040 17896 15104
rect 17960 15040 17976 15104
rect 18040 15040 18048 15104
rect 17728 14016 18048 15040
rect 17728 13952 17736 14016
rect 17800 13952 17816 14016
rect 17880 13952 17896 14016
rect 17960 13952 17976 14016
rect 18040 13952 18048 14016
rect 17728 12928 18048 13952
rect 17728 12864 17736 12928
rect 17800 12864 17816 12928
rect 17880 12864 17896 12928
rect 17960 12864 17976 12928
rect 18040 12864 18048 12928
rect 17728 11840 18048 12864
rect 17728 11776 17736 11840
rect 17800 11776 17816 11840
rect 17880 11776 17896 11840
rect 17960 11776 17976 11840
rect 18040 11776 18048 11840
rect 17728 10752 18048 11776
rect 17728 10688 17736 10752
rect 17800 10688 17816 10752
rect 17880 10688 17896 10752
rect 17960 10688 17976 10752
rect 18040 10688 18048 10752
rect 17728 9664 18048 10688
rect 17728 9600 17736 9664
rect 17800 9600 17816 9664
rect 17880 9600 17896 9664
rect 17960 9600 17976 9664
rect 18040 9600 18048 9664
rect 17728 8576 18048 9600
rect 17728 8512 17736 8576
rect 17800 8512 17816 8576
rect 17880 8512 17896 8576
rect 17960 8512 17976 8576
rect 18040 8512 18048 8576
rect 17728 7488 18048 8512
rect 17728 7424 17736 7488
rect 17800 7424 17816 7488
rect 17880 7424 17896 7488
rect 17960 7424 17976 7488
rect 18040 7424 18048 7488
rect 17728 6400 18048 7424
rect 17728 6336 17736 6400
rect 17800 6336 17816 6400
rect 17880 6336 17896 6400
rect 17960 6336 17976 6400
rect 18040 6336 18048 6400
rect 17728 5312 18048 6336
rect 17728 5248 17736 5312
rect 17800 5248 17816 5312
rect 17880 5248 17896 5312
rect 17960 5248 17976 5312
rect 18040 5248 18048 5312
rect 17728 4224 18048 5248
rect 17728 4160 17736 4224
rect 17800 4160 17816 4224
rect 17880 4160 17896 4224
rect 17960 4160 17976 4224
rect 18040 4160 18048 4224
rect 17728 3136 18048 4160
rect 17728 3072 17736 3136
rect 17800 3072 17816 3136
rect 17880 3072 17896 3136
rect 17960 3072 17976 3136
rect 18040 3072 18048 3136
rect 17728 2838 18048 3072
rect 17728 2602 17770 2838
rect 18006 2602 18048 2838
rect 17728 2048 18048 2602
rect 17728 1984 17736 2048
rect 17800 1984 17816 2048
rect 17880 1984 17896 2048
rect 17960 1984 17976 2048
rect 18040 1984 18048 2048
rect 17728 960 18048 1984
rect 17728 896 17736 960
rect 17800 896 17816 960
rect 17880 896 17896 960
rect 17960 896 17976 960
rect 18040 896 18048 960
rect 17728 880 18048 896
<< via4 >>
rect 4450 20602 4686 20838
rect 7114 2602 7350 2838
rect 9778 20602 10014 20838
rect 12442 2602 12678 2838
rect 15106 20602 15342 20838
rect 17770 2602 18006 2838
<< metal5 >>
rect 1904 20838 20764 20880
rect 1904 20602 4450 20838
rect 4686 20602 9778 20838
rect 10014 20602 15106 20838
rect 15342 20602 20764 20838
rect 1904 20560 20764 20602
rect 1904 2838 20764 2880
rect 1904 2602 7114 2838
rect 7350 2602 12442 2838
rect 12678 2602 17770 2838
rect 18006 2602 20764 2838
rect 1904 2560 20764 2602
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 2732 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 1996 0 1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_2
timestamp 1607194113
transform 1 0 1904 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_0
timestamp 1607194113
transform 1 0 2732 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_1
timestamp 1607194113
transform 1 0 1996 0 -1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_0
timestamp 1607194113
transform 1 0 1904 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_31 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 3100 0 1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 2824 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_0
timestamp 1607194113
transform 1 0 3100 0 -1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap0_0
timestamp 1607194113
transform 1 0 2824 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_30
timestamp 1607194113
transform 1 0 4204 0 1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap1_1
timestamp 1607194113
transform 1 0 3928 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_1
timestamp 1607194113
transform 1 0 3836 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_1
timestamp 1607194113
transform 1 0 4204 0 -1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap0_1
timestamp 1607194113
transform 1 0 3928 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_1
timestamp 1607194113
transform 1 0 3836 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_29
timestamp 1607194113
transform 1 0 5308 0 1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap1_2
timestamp 1607194113
transform 1 0 5032 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_2
timestamp 1607194113
transform 1 0 4940 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_2
timestamp 1607194113
transform 1 0 5308 0 -1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap0_2
timestamp 1607194113
transform 1 0 5032 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_2
timestamp 1607194113
transform 1 0 4940 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_28
timestamp 1607194113
transform 1 0 6412 0 1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap1_3
timestamp 1607194113
transform 1 0 6136 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_3
timestamp 1607194113
transform 1 0 6044 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_3
timestamp 1607194113
transform 1 0 6412 0 -1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap0_3
timestamp 1607194113
transform 1 0 6136 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_3
timestamp 1607194113
transform 1 0 6044 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_4
timestamp 1607194113
transform 1 0 7240 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_4
timestamp 1607194113
transform 1 0 7148 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_4
timestamp 1607194113
transform 1 0 7240 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_4
timestamp 1607194113
transform 1 0 7148 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_27
timestamp 1607194113
transform 1 0 7516 0 1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_4
timestamp 1607194113
transform 1 0 7516 0 -1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_26
timestamp 1607194113
transform 1 0 8620 0 1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap1_5
timestamp 1607194113
transform 1 0 8344 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_5
timestamp 1607194113
transform 1 0 8252 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_5
timestamp 1607194113
transform 1 0 8620 0 -1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap0_5
timestamp 1607194113
transform 1 0 8344 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_5
timestamp 1607194113
transform 1 0 8252 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_25
timestamp 1607194113
transform 1 0 9724 0 1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap1_6
timestamp 1607194113
transform 1 0 9448 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_6
timestamp 1607194113
transform 1 0 9356 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_6
timestamp 1607194113
transform 1 0 9724 0 -1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap0_6
timestamp 1607194113
transform 1 0 9448 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_6
timestamp 1607194113
transform 1 0 9356 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_24
timestamp 1607194113
transform 1 0 10828 0 1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap1_7
timestamp 1607194113
transform 1 0 10552 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_7
timestamp 1607194113
transform 1 0 10460 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_7
timestamp 1607194113
transform 1 0 10828 0 -1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap0_7
timestamp 1607194113
transform 1 0 10552 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_7
timestamp 1607194113
transform 1 0 10460 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_8
timestamp 1607194113
transform 1 0 11656 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_8
timestamp 1607194113
transform 1 0 11564 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_8
timestamp 1607194113
transform 1 0 11656 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_8
timestamp 1607194113
transform 1 0 11564 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_9
timestamp 1607194113
transform 1 0 12760 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_9
timestamp 1607194113
transform 1 0 12668 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_23
timestamp 1607194113
transform 1 0 11932 0 1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap0_9
timestamp 1607194113
transform 1 0 12760 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_9
timestamp 1607194113
transform 1 0 12668 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_8
timestamp 1607194113
transform 1 0 11932 0 -1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_22
timestamp 1607194113
transform 1 0 13036 0 1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_9
timestamp 1607194113
transform 1 0 13036 0 -1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_21
timestamp 1607194113
transform 1 0 14140 0 1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap1_10
timestamp 1607194113
transform 1 0 13864 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_10
timestamp 1607194113
transform 1 0 13772 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_10
timestamp 1607194113
transform 1 0 14140 0 -1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap0_10
timestamp 1607194113
transform 1 0 13864 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_10
timestamp 1607194113
transform 1 0 13772 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_20
timestamp 1607194113
transform 1 0 15244 0 1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap1_11
timestamp 1607194113
transform 1 0 14968 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_11
timestamp 1607194113
transform 1 0 14876 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_11
timestamp 1607194113
transform 1 0 15244 0 -1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap0_11
timestamp 1607194113
transform 1 0 14968 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_11
timestamp 1607194113
transform 1 0 14876 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_19
timestamp 1607194113
transform 1 0 16348 0 1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap1_12
timestamp 1607194113
transform 1 0 16072 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_12
timestamp 1607194113
transform 1 0 15980 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_12
timestamp 1607194113
transform 1 0 16348 0 -1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap0_12
timestamp 1607194113
transform 1 0 16072 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_12
timestamp 1607194113
transform 1 0 15980 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_13
timestamp 1607194113
transform 1 0 17176 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_13
timestamp 1607194113
transform 1 0 17084 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_13
timestamp 1607194113
transform 1 0 17176 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_13
timestamp 1607194113
transform 1 0 17084 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_14
timestamp 1607194113
transform 1 0 18188 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_18
timestamp 1607194113
transform 1 0 17452 0 1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_14
timestamp 1607194113
transform 1 0 18188 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_13
timestamp 1607194113
transform 1 0 17452 0 -1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_17
timestamp 1607194113
transform 1 0 18556 0 1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap1_14
timestamp 1607194113
transform 1 0 18280 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_14
timestamp 1607194113
transform 1 0 18556 0 -1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap0_14
timestamp 1607194113
transform 1 0 18280 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_16
timestamp 1607194113
transform 1 0 19660 0 1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap1_15
timestamp 1607194113
transform 1 0 19384 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_15
timestamp 1607194113
transform 1 0 19292 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_15
timestamp 1607194113
transform 1 0 19660 0 -1 1472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap0_15
timestamp 1607194113
transform 1 0 19384 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_15
timestamp 1607194113
transform 1 0 19292 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_16
timestamp 1607194113
transform 1 0 20488 0 1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_16
timestamp 1607194113
transform 1 0 20396 0 1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_16
timestamp 1607194113
transform 1 0 20488 0 -1 1472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_16
timestamp 1607194113
transform 1 0 20396 0 -1 1472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_0
timestamp 1607194113
transform 1 0 2732 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_5
timestamp 1607194113
transform 1 0 1996 0 -1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_4
timestamp 1607194113
transform 1 0 1904 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_32
timestamp 1607194113
transform 1 0 3100 0 -1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap2_0
timestamp 1607194113
transform 1 0 2824 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_33
timestamp 1607194113
transform 1 0 4204 0 -1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap2_1
timestamp 1607194113
transform 1 0 3928 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_1
timestamp 1607194113
transform 1 0 3836 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_34
timestamp 1607194113
transform 1 0 5308 0 -1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap2_2
timestamp 1607194113
transform 1 0 5032 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_2
timestamp 1607194113
transform 1 0 4940 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_35
timestamp 1607194113
transform 1 0 6412 0 -1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap2_3
timestamp 1607194113
transform 1 0 6136 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_3
timestamp 1607194113
transform 1 0 6044 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_4
timestamp 1607194113
transform 1 0 7240 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_4
timestamp 1607194113
transform 1 0 7148 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_36
timestamp 1607194113
transform 1 0 7516 0 -1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_37
timestamp 1607194113
transform 1 0 8620 0 -1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap2_5
timestamp 1607194113
transform 1 0 8344 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_5
timestamp 1607194113
transform 1 0 8252 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_38
timestamp 1607194113
transform 1 0 9724 0 -1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap2_6
timestamp 1607194113
transform 1 0 9448 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_6
timestamp 1607194113
transform 1 0 9356 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_39
timestamp 1607194113
transform 1 0 10828 0 -1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap2_7
timestamp 1607194113
transform 1 0 10552 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_7
timestamp 1607194113
transform 1 0 10460 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_8
timestamp 1607194113
transform 1 0 11656 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_8
timestamp 1607194113
transform 1 0 11564 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_9
timestamp 1607194113
transform 1 0 12760 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_9
timestamp 1607194113
transform 1 0 12668 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_40
timestamp 1607194113
transform 1 0 11932 0 -1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_41
timestamp 1607194113
transform 1 0 13036 0 -1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_42
timestamp 1607194113
transform 1 0 14140 0 -1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap2_10
timestamp 1607194113
transform 1 0 13864 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_10
timestamp 1607194113
transform 1 0 13772 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_43
timestamp 1607194113
transform 1 0 15244 0 -1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap2_11
timestamp 1607194113
transform 1 0 14968 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_11
timestamp 1607194113
transform 1 0 14876 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_44
timestamp 1607194113
transform 1 0 16348 0 -1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap2_12
timestamp 1607194113
transform 1 0 16072 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_12
timestamp 1607194113
transform 1 0 15980 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_13
timestamp 1607194113
transform 1 0 17176 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_13
timestamp 1607194113
transform 1 0 17084 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_14
timestamp 1607194113
transform 1 0 18188 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_45
timestamp 1607194113
transform 1 0 17452 0 -1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_46
timestamp 1607194113
transform 1 0 18556 0 -1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap2_14
timestamp 1607194113
transform 1 0 18280 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_47
timestamp 1607194113
transform 1 0 19660 0 -1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap2_15
timestamp 1607194113
transform 1 0 19384 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_15
timestamp 1607194113
transform 1 0 19292 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_16
timestamp 1607194113
transform 1 0 20488 0 -1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_16
timestamp 1607194113
transform 1 0 20396 0 -1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_0
timestamp 1607194113
transform 1 0 2732 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_7
timestamp 1607194113
transform 1 0 1996 0 1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_6
timestamp 1607194113
transform 1 0 1904 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_63
timestamp 1607194113
transform 1 0 3100 0 1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap3_0
timestamp 1607194113
transform 1 0 2824 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_62
timestamp 1607194113
transform 1 0 4204 0 1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap3_1
timestamp 1607194113
transform 1 0 3928 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_1
timestamp 1607194113
transform 1 0 3836 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_61
timestamp 1607194113
transform 1 0 5308 0 1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap3_2
timestamp 1607194113
transform 1 0 5032 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_2
timestamp 1607194113
transform 1 0 4940 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_60
timestamp 1607194113
transform 1 0 6412 0 1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap3_3
timestamp 1607194113
transform 1 0 6136 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_3
timestamp 1607194113
transform 1 0 6044 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_4
timestamp 1607194113
transform 1 0 7240 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_4
timestamp 1607194113
transform 1 0 7148 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_59
timestamp 1607194113
transform 1 0 7516 0 1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_58
timestamp 1607194113
transform 1 0 8620 0 1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap3_5
timestamp 1607194113
transform 1 0 8344 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_5
timestamp 1607194113
transform 1 0 8252 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_57
timestamp 1607194113
transform 1 0 9724 0 1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap3_6
timestamp 1607194113
transform 1 0 9448 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_6
timestamp 1607194113
transform 1 0 9356 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_56
timestamp 1607194113
transform 1 0 10828 0 1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap3_7
timestamp 1607194113
transform 1 0 10552 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_7
timestamp 1607194113
transform 1 0 10460 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_8
timestamp 1607194113
transform 1 0 11656 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_8
timestamp 1607194113
transform 1 0 11564 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_9
timestamp 1607194113
transform 1 0 12760 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_9
timestamp 1607194113
transform 1 0 12668 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_55
timestamp 1607194113
transform 1 0 11932 0 1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_54
timestamp 1607194113
transform 1 0 13036 0 1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_53
timestamp 1607194113
transform 1 0 14140 0 1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap3_10
timestamp 1607194113
transform 1 0 13864 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_10
timestamp 1607194113
transform 1 0 13772 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_52
timestamp 1607194113
transform 1 0 15244 0 1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap3_11
timestamp 1607194113
transform 1 0 14968 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_11
timestamp 1607194113
transform 1 0 14876 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_51
timestamp 1607194113
transform 1 0 16348 0 1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap3_12
timestamp 1607194113
transform 1 0 16072 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_12
timestamp 1607194113
transform 1 0 15980 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_13
timestamp 1607194113
transform 1 0 17176 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_13
timestamp 1607194113
transform 1 0 17084 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_14
timestamp 1607194113
transform 1 0 18188 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_50
timestamp 1607194113
transform 1 0 17452 0 1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_49
timestamp 1607194113
transform 1 0 18556 0 1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap3_14
timestamp 1607194113
transform 1 0 18280 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_48
timestamp 1607194113
transform 1 0 19660 0 1 2560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap3_15
timestamp 1607194113
transform 1 0 19384 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_15
timestamp 1607194113
transform 1 0 19292 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_16
timestamp 1607194113
transform 1 0 20488 0 1 2560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_16
timestamp 1607194113
transform 1 0 20396 0 1 2560
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_0
timestamp 1607194113
transform 1 0 2732 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_9
timestamp 1607194113
transform 1 0 1996 0 -1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_8
timestamp 1607194113
transform 1 0 1904 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_64
timestamp 1607194113
transform 1 0 3100 0 -1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap4_0
timestamp 1607194113
transform 1 0 2824 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_65
timestamp 1607194113
transform 1 0 4204 0 -1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap4_1
timestamp 1607194113
transform 1 0 3928 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_1
timestamp 1607194113
transform 1 0 3836 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_66
timestamp 1607194113
transform 1 0 5308 0 -1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap4_2
timestamp 1607194113
transform 1 0 5032 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_2
timestamp 1607194113
transform 1 0 4940 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_67
timestamp 1607194113
transform 1 0 6412 0 -1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap4_3
timestamp 1607194113
transform 1 0 6136 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_3
timestamp 1607194113
transform 1 0 6044 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_4
timestamp 1607194113
transform 1 0 7240 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_4
timestamp 1607194113
transform 1 0 7148 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_68
timestamp 1607194113
transform 1 0 7516 0 -1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_69
timestamp 1607194113
transform 1 0 8620 0 -1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap4_5
timestamp 1607194113
transform 1 0 8344 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_5
timestamp 1607194113
transform 1 0 8252 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_70
timestamp 1607194113
transform 1 0 9724 0 -1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap4_6
timestamp 1607194113
transform 1 0 9448 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_6
timestamp 1607194113
transform 1 0 9356 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_71
timestamp 1607194113
transform 1 0 10828 0 -1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap4_7
timestamp 1607194113
transform 1 0 10552 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_7
timestamp 1607194113
transform 1 0 10460 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_8
timestamp 1607194113
transform 1 0 11656 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_8
timestamp 1607194113
transform 1 0 11564 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_9
timestamp 1607194113
transform 1 0 12760 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_9
timestamp 1607194113
transform 1 0 12668 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_72
timestamp 1607194113
transform 1 0 11932 0 -1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_73
timestamp 1607194113
transform 1 0 13036 0 -1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_74
timestamp 1607194113
transform 1 0 14140 0 -1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap4_10
timestamp 1607194113
transform 1 0 13864 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_10
timestamp 1607194113
transform 1 0 13772 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_75
timestamp 1607194113
transform 1 0 15244 0 -1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap4_11
timestamp 1607194113
transform 1 0 14968 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_11
timestamp 1607194113
transform 1 0 14876 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_76
timestamp 1607194113
transform 1 0 16348 0 -1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap4_12
timestamp 1607194113
transform 1 0 16072 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_12
timestamp 1607194113
transform 1 0 15980 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_13
timestamp 1607194113
transform 1 0 17176 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_13
timestamp 1607194113
transform 1 0 17084 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_14
timestamp 1607194113
transform 1 0 18188 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_77
timestamp 1607194113
transform 1 0 17452 0 -1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_78
timestamp 1607194113
transform 1 0 18556 0 -1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap4_14
timestamp 1607194113
transform 1 0 18280 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_79
timestamp 1607194113
transform 1 0 19660 0 -1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap4_15
timestamp 1607194113
transform 1 0 19384 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_15
timestamp 1607194113
transform 1 0 19292 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_16
timestamp 1607194113
transform 1 0 20488 0 -1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_16
timestamp 1607194113
transform 1 0 20396 0 -1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_0
timestamp 1607194113
transform 1 0 2732 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_11
timestamp 1607194113
transform 1 0 1996 0 1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_10
timestamp 1607194113
transform 1 0 1904 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_95
timestamp 1607194113
transform 1 0 3100 0 1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap5_0
timestamp 1607194113
transform 1 0 2824 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_94
timestamp 1607194113
transform 1 0 4204 0 1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap5_1
timestamp 1607194113
transform 1 0 3928 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_1
timestamp 1607194113
transform 1 0 3836 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_93
timestamp 1607194113
transform 1 0 5308 0 1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap5_2
timestamp 1607194113
transform 1 0 5032 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_2
timestamp 1607194113
transform 1 0 4940 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_92
timestamp 1607194113
transform 1 0 6412 0 1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap5_3
timestamp 1607194113
transform 1 0 6136 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_3
timestamp 1607194113
transform 1 0 6044 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_4
timestamp 1607194113
transform 1 0 7240 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_4
timestamp 1607194113
transform 1 0 7148 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_91
timestamp 1607194113
transform 1 0 7516 0 1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_90
timestamp 1607194113
transform 1 0 8620 0 1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap5_5
timestamp 1607194113
transform 1 0 8344 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_5
timestamp 1607194113
transform 1 0 8252 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_89
timestamp 1607194113
transform 1 0 9724 0 1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap5_6
timestamp 1607194113
transform 1 0 9448 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_6
timestamp 1607194113
transform 1 0 9356 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_88
timestamp 1607194113
transform 1 0 10828 0 1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap5_7
timestamp 1607194113
transform 1 0 10552 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_7
timestamp 1607194113
transform 1 0 10460 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_8
timestamp 1607194113
transform 1 0 11656 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_8
timestamp 1607194113
transform 1 0 11564 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_9
timestamp 1607194113
transform 1 0 12760 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_9
timestamp 1607194113
transform 1 0 12668 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_87
timestamp 1607194113
transform 1 0 11932 0 1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_86
timestamp 1607194113
transform 1 0 13036 0 1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_85
timestamp 1607194113
transform 1 0 14140 0 1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap5_10
timestamp 1607194113
transform 1 0 13864 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_10
timestamp 1607194113
transform 1 0 13772 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_84
timestamp 1607194113
transform 1 0 15244 0 1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap5_11
timestamp 1607194113
transform 1 0 14968 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_11
timestamp 1607194113
transform 1 0 14876 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_83
timestamp 1607194113
transform 1 0 16348 0 1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap5_12
timestamp 1607194113
transform 1 0 16072 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_12
timestamp 1607194113
transform 1 0 15980 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_13
timestamp 1607194113
transform 1 0 17176 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_13
timestamp 1607194113
transform 1 0 17084 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_14
timestamp 1607194113
transform 1 0 18188 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_82
timestamp 1607194113
transform 1 0 17452 0 1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_81
timestamp 1607194113
transform 1 0 18556 0 1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap5_14
timestamp 1607194113
transform 1 0 18280 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_80
timestamp 1607194113
transform 1 0 19660 0 1 3648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap5_15
timestamp 1607194113
transform 1 0 19384 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_15
timestamp 1607194113
transform 1 0 19292 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_16
timestamp 1607194113
transform 1 0 20488 0 1 3648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_16
timestamp 1607194113
transform 1 0 20396 0 1 3648
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_0
timestamp 1607194113
transform 1 0 2732 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_15
timestamp 1607194113
transform 1 0 1996 0 1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_14
timestamp 1607194113
transform 1 0 1904 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_0
timestamp 1607194113
transform 1 0 2732 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_13
timestamp 1607194113
transform 1 0 1996 0 -1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_12
timestamp 1607194113
transform 1 0 1904 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_127
timestamp 1607194113
transform 1 0 3100 0 1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap7_0
timestamp 1607194113
transform 1 0 2824 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_96
timestamp 1607194113
transform 1 0 3100 0 -1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap6_0
timestamp 1607194113
transform 1 0 2824 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_126
timestamp 1607194113
transform 1 0 4204 0 1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap7_1
timestamp 1607194113
transform 1 0 3928 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_1
timestamp 1607194113
transform 1 0 3836 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_97
timestamp 1607194113
transform 1 0 4204 0 -1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap6_1
timestamp 1607194113
transform 1 0 3928 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_1
timestamp 1607194113
transform 1 0 3836 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_125
timestamp 1607194113
transform 1 0 5308 0 1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap7_2
timestamp 1607194113
transform 1 0 5032 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_2
timestamp 1607194113
transform 1 0 4940 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_98
timestamp 1607194113
transform 1 0 5308 0 -1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap6_2
timestamp 1607194113
transform 1 0 5032 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_2
timestamp 1607194113
transform 1 0 4940 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_124
timestamp 1607194113
transform 1 0 6412 0 1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap7_3
timestamp 1607194113
transform 1 0 6136 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_3
timestamp 1607194113
transform 1 0 6044 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_99
timestamp 1607194113
transform 1 0 6412 0 -1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap6_3
timestamp 1607194113
transform 1 0 6136 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_3
timestamp 1607194113
transform 1 0 6044 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_4
timestamp 1607194113
transform 1 0 7240 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_4
timestamp 1607194113
transform 1 0 7148 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_4
timestamp 1607194113
transform 1 0 7240 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_4
timestamp 1607194113
transform 1 0 7148 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_123
timestamp 1607194113
transform 1 0 7516 0 1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_100
timestamp 1607194113
transform 1 0 7516 0 -1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_122
timestamp 1607194113
transform 1 0 8620 0 1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap7_5
timestamp 1607194113
transform 1 0 8344 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_5
timestamp 1607194113
transform 1 0 8252 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_101
timestamp 1607194113
transform 1 0 8620 0 -1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap6_5
timestamp 1607194113
transform 1 0 8344 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_5
timestamp 1607194113
transform 1 0 8252 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_121
timestamp 1607194113
transform 1 0 9724 0 1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap7_6
timestamp 1607194113
transform 1 0 9448 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_6
timestamp 1607194113
transform 1 0 9356 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_102
timestamp 1607194113
transform 1 0 9724 0 -1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap6_6
timestamp 1607194113
transform 1 0 9448 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_6
timestamp 1607194113
transform 1 0 9356 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_120
timestamp 1607194113
transform 1 0 10828 0 1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap7_7
timestamp 1607194113
transform 1 0 10552 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_7
timestamp 1607194113
transform 1 0 10460 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_103
timestamp 1607194113
transform 1 0 10828 0 -1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap6_7
timestamp 1607194113
transform 1 0 10552 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_7
timestamp 1607194113
transform 1 0 10460 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_8
timestamp 1607194113
transform 1 0 11656 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_8
timestamp 1607194113
transform 1 0 11564 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_8
timestamp 1607194113
transform 1 0 11656 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_8
timestamp 1607194113
transform 1 0 11564 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_9
timestamp 1607194113
transform 1 0 12760 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_9
timestamp 1607194113
transform 1 0 12668 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_119
timestamp 1607194113
transform 1 0 11932 0 1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap6_9
timestamp 1607194113
transform 1 0 12760 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_9
timestamp 1607194113
transform 1 0 12668 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_104
timestamp 1607194113
transform 1 0 11932 0 -1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_118
timestamp 1607194113
transform 1 0 13036 0 1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_105
timestamp 1607194113
transform 1 0 13036 0 -1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_117
timestamp 1607194113
transform 1 0 14140 0 1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap7_10
timestamp 1607194113
transform 1 0 13864 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_10
timestamp 1607194113
transform 1 0 13772 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_106
timestamp 1607194113
transform 1 0 14140 0 -1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap6_10
timestamp 1607194113
transform 1 0 13864 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_10
timestamp 1607194113
transform 1 0 13772 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_116
timestamp 1607194113
transform 1 0 15244 0 1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap7_11
timestamp 1607194113
transform 1 0 14968 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_11
timestamp 1607194113
transform 1 0 14876 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_107
timestamp 1607194113
transform 1 0 15244 0 -1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap6_11
timestamp 1607194113
transform 1 0 14968 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_11
timestamp 1607194113
transform 1 0 14876 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_115
timestamp 1607194113
transform 1 0 16348 0 1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap7_12
timestamp 1607194113
transform 1 0 16072 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_12
timestamp 1607194113
transform 1 0 15980 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_108
timestamp 1607194113
transform 1 0 16348 0 -1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap6_12
timestamp 1607194113
transform 1 0 16072 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_12
timestamp 1607194113
transform 1 0 15980 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_13
timestamp 1607194113
transform 1 0 17176 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_13
timestamp 1607194113
transform 1 0 17084 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_13
timestamp 1607194113
transform 1 0 17176 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_13
timestamp 1607194113
transform 1 0 17084 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_14
timestamp 1607194113
transform 1 0 18188 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_114
timestamp 1607194113
transform 1 0 17452 0 1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_14
timestamp 1607194113
transform 1 0 18188 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_109
timestamp 1607194113
transform 1 0 17452 0 -1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_113
timestamp 1607194113
transform 1 0 18556 0 1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap7_14
timestamp 1607194113
transform 1 0 18280 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_110
timestamp 1607194113
transform 1 0 18556 0 -1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap6_14
timestamp 1607194113
transform 1 0 18280 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_112
timestamp 1607194113
transform 1 0 19660 0 1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap7_15
timestamp 1607194113
transform 1 0 19384 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_15
timestamp 1607194113
transform 1 0 19292 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_111
timestamp 1607194113
transform 1 0 19660 0 -1 4736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap6_15
timestamp 1607194113
transform 1 0 19384 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_15
timestamp 1607194113
transform 1 0 19292 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_16
timestamp 1607194113
transform 1 0 20488 0 1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_16
timestamp 1607194113
transform 1 0 20396 0 1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_16
timestamp 1607194113
transform 1 0 20488 0 -1 4736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_16
timestamp 1607194113
transform 1 0 20396 0 -1 4736
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_0
timestamp 1607194113
transform 1 0 2732 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_17
timestamp 1607194113
transform 1 0 1996 0 -1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_16
timestamp 1607194113
transform 1 0 1904 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_128
timestamp 1607194113
transform 1 0 3100 0 -1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap8_0
timestamp 1607194113
transform 1 0 2824 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_129
timestamp 1607194113
transform 1 0 4204 0 -1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap8_1
timestamp 1607194113
transform 1 0 3928 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_1
timestamp 1607194113
transform 1 0 3836 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_130
timestamp 1607194113
transform 1 0 5308 0 -1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap8_2
timestamp 1607194113
transform 1 0 5032 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_2
timestamp 1607194113
transform 1 0 4940 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_131
timestamp 1607194113
transform 1 0 6412 0 -1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap8_3
timestamp 1607194113
transform 1 0 6136 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_3
timestamp 1607194113
transform 1 0 6044 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_4
timestamp 1607194113
transform 1 0 7240 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_4
timestamp 1607194113
transform 1 0 7148 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_132
timestamp 1607194113
transform 1 0 7516 0 -1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_133
timestamp 1607194113
transform 1 0 8620 0 -1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap8_5
timestamp 1607194113
transform 1 0 8344 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_5
timestamp 1607194113
transform 1 0 8252 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_134
timestamp 1607194113
transform 1 0 9724 0 -1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap8_6
timestamp 1607194113
transform 1 0 9448 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_6
timestamp 1607194113
transform 1 0 9356 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_135
timestamp 1607194113
transform 1 0 10828 0 -1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap8_7
timestamp 1607194113
transform 1 0 10552 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_7
timestamp 1607194113
transform 1 0 10460 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_8
timestamp 1607194113
transform 1 0 11656 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_8
timestamp 1607194113
transform 1 0 11564 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_9
timestamp 1607194113
transform 1 0 12760 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_9
timestamp 1607194113
transform 1 0 12668 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_136
timestamp 1607194113
transform 1 0 11932 0 -1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_137
timestamp 1607194113
transform 1 0 13036 0 -1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_138
timestamp 1607194113
transform 1 0 14140 0 -1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap8_10
timestamp 1607194113
transform 1 0 13864 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_10
timestamp 1607194113
transform 1 0 13772 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_139
timestamp 1607194113
transform 1 0 15244 0 -1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap8_11
timestamp 1607194113
transform 1 0 14968 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_11
timestamp 1607194113
transform 1 0 14876 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_140
timestamp 1607194113
transform 1 0 16348 0 -1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap8_12
timestamp 1607194113
transform 1 0 16072 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_12
timestamp 1607194113
transform 1 0 15980 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_13
timestamp 1607194113
transform 1 0 17176 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_13
timestamp 1607194113
transform 1 0 17084 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_14
timestamp 1607194113
transform 1 0 18188 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_141
timestamp 1607194113
transform 1 0 17452 0 -1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_142
timestamp 1607194113
transform 1 0 18556 0 -1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap8_14
timestamp 1607194113
transform 1 0 18280 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_143
timestamp 1607194113
transform 1 0 19660 0 -1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap8_15
timestamp 1607194113
transform 1 0 19384 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_15
timestamp 1607194113
transform 1 0 19292 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_16
timestamp 1607194113
transform 1 0 20488 0 -1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_16
timestamp 1607194113
transform 1 0 20396 0 -1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_0
timestamp 1607194113
transform 1 0 2732 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_19
timestamp 1607194113
transform 1 0 1996 0 1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_18
timestamp 1607194113
transform 1 0 1904 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_159
timestamp 1607194113
transform 1 0 3100 0 1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap9_0
timestamp 1607194113
transform 1 0 2824 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_158
timestamp 1607194113
transform 1 0 4204 0 1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap9_1
timestamp 1607194113
transform 1 0 3928 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_1
timestamp 1607194113
transform 1 0 3836 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_157
timestamp 1607194113
transform 1 0 5308 0 1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap9_2
timestamp 1607194113
transform 1 0 5032 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_2
timestamp 1607194113
transform 1 0 4940 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_156
timestamp 1607194113
transform 1 0 6412 0 1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap9_3
timestamp 1607194113
transform 1 0 6136 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_3
timestamp 1607194113
transform 1 0 6044 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_4
timestamp 1607194113
transform 1 0 7240 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_4
timestamp 1607194113
transform 1 0 7148 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_155
timestamp 1607194113
transform 1 0 7516 0 1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_154
timestamp 1607194113
transform 1 0 8620 0 1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap9_5
timestamp 1607194113
transform 1 0 8344 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_5
timestamp 1607194113
transform 1 0 8252 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_153
timestamp 1607194113
transform 1 0 9724 0 1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap9_6
timestamp 1607194113
transform 1 0 9448 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_6
timestamp 1607194113
transform 1 0 9356 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_152
timestamp 1607194113
transform 1 0 10828 0 1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap9_7
timestamp 1607194113
transform 1 0 10552 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_7
timestamp 1607194113
transform 1 0 10460 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_8
timestamp 1607194113
transform 1 0 11656 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_8
timestamp 1607194113
transform 1 0 11564 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_9
timestamp 1607194113
transform 1 0 12760 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_9
timestamp 1607194113
transform 1 0 12668 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_151
timestamp 1607194113
transform 1 0 11932 0 1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_150
timestamp 1607194113
transform 1 0 13036 0 1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_149
timestamp 1607194113
transform 1 0 14140 0 1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap9_10
timestamp 1607194113
transform 1 0 13864 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_10
timestamp 1607194113
transform 1 0 13772 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_148
timestamp 1607194113
transform 1 0 15244 0 1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap9_11
timestamp 1607194113
transform 1 0 14968 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_11
timestamp 1607194113
transform 1 0 14876 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_147
timestamp 1607194113
transform 1 0 16348 0 1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap9_12
timestamp 1607194113
transform 1 0 16072 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_12
timestamp 1607194113
transform 1 0 15980 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_13
timestamp 1607194113
transform 1 0 17176 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_13
timestamp 1607194113
transform 1 0 17084 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_14
timestamp 1607194113
transform 1 0 18188 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_146
timestamp 1607194113
transform 1 0 17452 0 1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_145
timestamp 1607194113
transform 1 0 18556 0 1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap9_14
timestamp 1607194113
transform 1 0 18280 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_144
timestamp 1607194113
transform 1 0 19660 0 1 5824
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap9_15
timestamp 1607194113
transform 1 0 19384 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_15
timestamp 1607194113
transform 1 0 19292 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_16
timestamp 1607194113
transform 1 0 20488 0 1 5824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_16
timestamp 1607194113
transform 1 0 20396 0 1 5824
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_0
timestamp 1607194113
transform 1 0 2732 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_21
timestamp 1607194113
transform 1 0 1996 0 -1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_20
timestamp 1607194113
transform 1 0 1904 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_160
timestamp 1607194113
transform 1 0 3100 0 -1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap10_0
timestamp 1607194113
transform 1 0 2824 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_161
timestamp 1607194113
transform 1 0 4204 0 -1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap10_1
timestamp 1607194113
transform 1 0 3928 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_1
timestamp 1607194113
transform 1 0 3836 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_162
timestamp 1607194113
transform 1 0 5308 0 -1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap10_2
timestamp 1607194113
transform 1 0 5032 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_2
timestamp 1607194113
transform 1 0 4940 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_163
timestamp 1607194113
transform 1 0 6412 0 -1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap10_3
timestamp 1607194113
transform 1 0 6136 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_3
timestamp 1607194113
transform 1 0 6044 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_4
timestamp 1607194113
transform 1 0 7240 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_4
timestamp 1607194113
transform 1 0 7148 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_164
timestamp 1607194113
transform 1 0 7516 0 -1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_165
timestamp 1607194113
transform 1 0 8620 0 -1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap10_5
timestamp 1607194113
transform 1 0 8344 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_5
timestamp 1607194113
transform 1 0 8252 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_166
timestamp 1607194113
transform 1 0 9724 0 -1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap10_6
timestamp 1607194113
transform 1 0 9448 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_6
timestamp 1607194113
transform 1 0 9356 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_167
timestamp 1607194113
transform 1 0 10828 0 -1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap10_7
timestamp 1607194113
transform 1 0 10552 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_7
timestamp 1607194113
transform 1 0 10460 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_8
timestamp 1607194113
transform 1 0 11656 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_8
timestamp 1607194113
transform 1 0 11564 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_9
timestamp 1607194113
transform 1 0 12760 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_9
timestamp 1607194113
transform 1 0 12668 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_168
timestamp 1607194113
transform 1 0 11932 0 -1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_169
timestamp 1607194113
transform 1 0 13036 0 -1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_170
timestamp 1607194113
transform 1 0 14140 0 -1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap10_10
timestamp 1607194113
transform 1 0 13864 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_10
timestamp 1607194113
transform 1 0 13772 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_171
timestamp 1607194113
transform 1 0 15244 0 -1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap10_11
timestamp 1607194113
transform 1 0 14968 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_11
timestamp 1607194113
transform 1 0 14876 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_172
timestamp 1607194113
transform 1 0 16348 0 -1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap10_12
timestamp 1607194113
transform 1 0 16072 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_12
timestamp 1607194113
transform 1 0 15980 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_13
timestamp 1607194113
transform 1 0 17176 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_13
timestamp 1607194113
transform 1 0 17084 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_14
timestamp 1607194113
transform 1 0 18188 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_173
timestamp 1607194113
transform 1 0 17452 0 -1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_174
timestamp 1607194113
transform 1 0 18556 0 -1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap10_14
timestamp 1607194113
transform 1 0 18280 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_175
timestamp 1607194113
transform 1 0 19660 0 -1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap10_15
timestamp 1607194113
transform 1 0 19384 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_15
timestamp 1607194113
transform 1 0 19292 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_16
timestamp 1607194113
transform 1 0 20488 0 -1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_16
timestamp 1607194113
transform 1 0 20396 0 -1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_0
timestamp 1607194113
transform 1 0 2732 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_23
timestamp 1607194113
transform 1 0 1996 0 1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_22
timestamp 1607194113
transform 1 0 1904 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_191
timestamp 1607194113
transform 1 0 3100 0 1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap11_0
timestamp 1607194113
transform 1 0 2824 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_190
timestamp 1607194113
transform 1 0 4204 0 1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap11_1
timestamp 1607194113
transform 1 0 3928 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_1
timestamp 1607194113
transform 1 0 3836 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_189
timestamp 1607194113
transform 1 0 5308 0 1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap11_2
timestamp 1607194113
transform 1 0 5032 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_2
timestamp 1607194113
transform 1 0 4940 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_188
timestamp 1607194113
transform 1 0 6412 0 1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap11_3
timestamp 1607194113
transform 1 0 6136 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_3
timestamp 1607194113
transform 1 0 6044 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_4
timestamp 1607194113
transform 1 0 7240 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_4
timestamp 1607194113
transform 1 0 7148 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_187
timestamp 1607194113
transform 1 0 7516 0 1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_186
timestamp 1607194113
transform 1 0 8620 0 1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap11_5
timestamp 1607194113
transform 1 0 8344 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_5
timestamp 1607194113
transform 1 0 8252 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_185
timestamp 1607194113
transform 1 0 9724 0 1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap11_6
timestamp 1607194113
transform 1 0 9448 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_6
timestamp 1607194113
transform 1 0 9356 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_184
timestamp 1607194113
transform 1 0 10828 0 1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap11_7
timestamp 1607194113
transform 1 0 10552 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_7
timestamp 1607194113
transform 1 0 10460 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_8
timestamp 1607194113
transform 1 0 11656 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_8
timestamp 1607194113
transform 1 0 11564 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_9
timestamp 1607194113
transform 1 0 12760 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_9
timestamp 1607194113
transform 1 0 12668 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_183
timestamp 1607194113
transform 1 0 11932 0 1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_182
timestamp 1607194113
transform 1 0 13036 0 1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_181
timestamp 1607194113
transform 1 0 14140 0 1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap11_10
timestamp 1607194113
transform 1 0 13864 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_10
timestamp 1607194113
transform 1 0 13772 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_180
timestamp 1607194113
transform 1 0 15244 0 1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap11_11
timestamp 1607194113
transform 1 0 14968 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_11
timestamp 1607194113
transform 1 0 14876 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_179
timestamp 1607194113
transform 1 0 16348 0 1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap11_12
timestamp 1607194113
transform 1 0 16072 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_12
timestamp 1607194113
transform 1 0 15980 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_13
timestamp 1607194113
transform 1 0 17176 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_13
timestamp 1607194113
transform 1 0 17084 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_14
timestamp 1607194113
transform 1 0 18188 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_178
timestamp 1607194113
transform 1 0 17452 0 1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_177
timestamp 1607194113
transform 1 0 18556 0 1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap11_14
timestamp 1607194113
transform 1 0 18280 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_176
timestamp 1607194113
transform 1 0 19660 0 1 6912
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap11_15
timestamp 1607194113
transform 1 0 19384 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_15
timestamp 1607194113
transform 1 0 19292 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_16
timestamp 1607194113
transform 1 0 20488 0 1 6912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_16
timestamp 1607194113
transform 1 0 20396 0 1 6912
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_0
timestamp 1607194113
transform 1 0 2732 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_25
timestamp 1607194113
transform 1 0 1996 0 -1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_24
timestamp 1607194113
transform 1 0 1904 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_192
timestamp 1607194113
transform 1 0 3100 0 -1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap12_0
timestamp 1607194113
transform 1 0 2824 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_193
timestamp 1607194113
transform 1 0 4204 0 -1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap12_1
timestamp 1607194113
transform 1 0 3928 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_1
timestamp 1607194113
transform 1 0 3836 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_194
timestamp 1607194113
transform 1 0 5308 0 -1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap12_2
timestamp 1607194113
transform 1 0 5032 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_2
timestamp 1607194113
transform 1 0 4940 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_195
timestamp 1607194113
transform 1 0 6412 0 -1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap12_3
timestamp 1607194113
transform 1 0 6136 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_3
timestamp 1607194113
transform 1 0 6044 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap12_4
timestamp 1607194113
transform 1 0 7240 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_4
timestamp 1607194113
transform 1 0 7148 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_196
timestamp 1607194113
transform 1 0 7516 0 -1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_197
timestamp 1607194113
transform 1 0 8620 0 -1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap12_5
timestamp 1607194113
transform 1 0 8344 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_5
timestamp 1607194113
transform 1 0 8252 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_198
timestamp 1607194113
transform 1 0 9724 0 -1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap12_6
timestamp 1607194113
transform 1 0 9448 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_6
timestamp 1607194113
transform 1 0 9356 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_199
timestamp 1607194113
transform 1 0 10828 0 -1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap12_7
timestamp 1607194113
transform 1 0 10552 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_7
timestamp 1607194113
transform 1 0 10460 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap12_8
timestamp 1607194113
transform 1 0 11656 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_8
timestamp 1607194113
transform 1 0 11564 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap12_9
timestamp 1607194113
transform 1 0 12760 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_9
timestamp 1607194113
transform 1 0 12668 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_200
timestamp 1607194113
transform 1 0 11932 0 -1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_201
timestamp 1607194113
transform 1 0 13036 0 -1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_202
timestamp 1607194113
transform 1 0 14140 0 -1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap12_10
timestamp 1607194113
transform 1 0 13864 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_10
timestamp 1607194113
transform 1 0 13772 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_203
timestamp 1607194113
transform 1 0 15244 0 -1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap12_11
timestamp 1607194113
transform 1 0 14968 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_11
timestamp 1607194113
transform 1 0 14876 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_204
timestamp 1607194113
transform 1 0 16348 0 -1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap12_12
timestamp 1607194113
transform 1 0 16072 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_12
timestamp 1607194113
transform 1 0 15980 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap12_13
timestamp 1607194113
transform 1 0 17176 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_13
timestamp 1607194113
transform 1 0 17084 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_14
timestamp 1607194113
transform 1 0 18188 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_205
timestamp 1607194113
transform 1 0 17452 0 -1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_206
timestamp 1607194113
transform 1 0 18556 0 -1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap12_14
timestamp 1607194113
transform 1 0 18280 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_207
timestamp 1607194113
transform 1 0 19660 0 -1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap12_15
timestamp 1607194113
transform 1 0 19384 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_15
timestamp 1607194113
transform 1 0 19292 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap12_16
timestamp 1607194113
transform 1 0 20488 0 -1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap12_16
timestamp 1607194113
transform 1 0 20396 0 -1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_0
timestamp 1607194113
transform 1 0 2732 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_29
timestamp 1607194113
transform 1 0 1996 0 -1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_28
timestamp 1607194113
transform 1 0 1904 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_0
timestamp 1607194113
transform 1 0 2732 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_27
timestamp 1607194113
transform 1 0 1996 0 1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_26
timestamp 1607194113
transform 1 0 1904 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_224
timestamp 1607194113
transform 1 0 3100 0 -1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap14_0
timestamp 1607194113
transform 1 0 2824 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_223
timestamp 1607194113
transform 1 0 3100 0 1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap13_0
timestamp 1607194113
transform 1 0 2824 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_225
timestamp 1607194113
transform 1 0 4204 0 -1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap14_1
timestamp 1607194113
transform 1 0 3928 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_1
timestamp 1607194113
transform 1 0 3836 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_222
timestamp 1607194113
transform 1 0 4204 0 1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap13_1
timestamp 1607194113
transform 1 0 3928 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_1
timestamp 1607194113
transform 1 0 3836 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_226
timestamp 1607194113
transform 1 0 5308 0 -1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap14_2
timestamp 1607194113
transform 1 0 5032 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_2
timestamp 1607194113
transform 1 0 4940 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_221
timestamp 1607194113
transform 1 0 5308 0 1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap13_2
timestamp 1607194113
transform 1 0 5032 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_2
timestamp 1607194113
transform 1 0 4940 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_227
timestamp 1607194113
transform 1 0 6412 0 -1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap14_3
timestamp 1607194113
transform 1 0 6136 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_3
timestamp 1607194113
transform 1 0 6044 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_220
timestamp 1607194113
transform 1 0 6412 0 1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap13_3
timestamp 1607194113
transform 1 0 6136 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_3
timestamp 1607194113
transform 1 0 6044 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap14_4
timestamp 1607194113
transform 1 0 7240 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_4
timestamp 1607194113
transform 1 0 7148 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap13_4
timestamp 1607194113
transform 1 0 7240 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_4
timestamp 1607194113
transform 1 0 7148 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_228
timestamp 1607194113
transform 1 0 7516 0 -1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_219
timestamp 1607194113
transform 1 0 7516 0 1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_229
timestamp 1607194113
transform 1 0 8620 0 -1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap14_5
timestamp 1607194113
transform 1 0 8344 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_5
timestamp 1607194113
transform 1 0 8252 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_218
timestamp 1607194113
transform 1 0 8620 0 1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap13_5
timestamp 1607194113
transform 1 0 8344 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_5
timestamp 1607194113
transform 1 0 8252 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_230
timestamp 1607194113
transform 1 0 9724 0 -1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap14_6
timestamp 1607194113
transform 1 0 9448 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_6
timestamp 1607194113
transform 1 0 9356 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_217
timestamp 1607194113
transform 1 0 9724 0 1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap13_6
timestamp 1607194113
transform 1 0 9448 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_6
timestamp 1607194113
transform 1 0 9356 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_231
timestamp 1607194113
transform 1 0 10828 0 -1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap14_7
timestamp 1607194113
transform 1 0 10552 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_7
timestamp 1607194113
transform 1 0 10460 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_216
timestamp 1607194113
transform 1 0 10828 0 1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap13_7
timestamp 1607194113
transform 1 0 10552 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_7
timestamp 1607194113
transform 1 0 10460 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap14_8
timestamp 1607194113
transform 1 0 11656 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_8
timestamp 1607194113
transform 1 0 11564 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap13_8
timestamp 1607194113
transform 1 0 11656 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_8
timestamp 1607194113
transform 1 0 11564 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap14_9
timestamp 1607194113
transform 1 0 12760 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_9
timestamp 1607194113
transform 1 0 12668 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_232
timestamp 1607194113
transform 1 0 11932 0 -1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap13_9
timestamp 1607194113
transform 1 0 12760 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_9
timestamp 1607194113
transform 1 0 12668 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_215
timestamp 1607194113
transform 1 0 11932 0 1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_233
timestamp 1607194113
transform 1 0 13036 0 -1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_214
timestamp 1607194113
transform 1 0 13036 0 1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_234
timestamp 1607194113
transform 1 0 14140 0 -1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap14_10
timestamp 1607194113
transform 1 0 13864 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_10
timestamp 1607194113
transform 1 0 13772 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_213
timestamp 1607194113
transform 1 0 14140 0 1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap13_10
timestamp 1607194113
transform 1 0 13864 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_10
timestamp 1607194113
transform 1 0 13772 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_235
timestamp 1607194113
transform 1 0 15244 0 -1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap14_11
timestamp 1607194113
transform 1 0 14968 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_11
timestamp 1607194113
transform 1 0 14876 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_212
timestamp 1607194113
transform 1 0 15244 0 1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap13_11
timestamp 1607194113
transform 1 0 14968 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_11
timestamp 1607194113
transform 1 0 14876 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_236
timestamp 1607194113
transform 1 0 16348 0 -1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap14_12
timestamp 1607194113
transform 1 0 16072 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_12
timestamp 1607194113
transform 1 0 15980 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_211
timestamp 1607194113
transform 1 0 16348 0 1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap13_12
timestamp 1607194113
transform 1 0 16072 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_12
timestamp 1607194113
transform 1 0 15980 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap14_13
timestamp 1607194113
transform 1 0 17176 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_13
timestamp 1607194113
transform 1 0 17084 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap13_13
timestamp 1607194113
transform 1 0 17176 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_13
timestamp 1607194113
transform 1 0 17084 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_14
timestamp 1607194113
transform 1 0 18188 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_237
timestamp 1607194113
transform 1 0 17452 0 -1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_14
timestamp 1607194113
transform 1 0 18188 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_210
timestamp 1607194113
transform 1 0 17452 0 1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_238
timestamp 1607194113
transform 1 0 18556 0 -1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap14_14
timestamp 1607194113
transform 1 0 18280 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_209
timestamp 1607194113
transform 1 0 18556 0 1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap13_14
timestamp 1607194113
transform 1 0 18280 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_239
timestamp 1607194113
transform 1 0 19660 0 -1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap14_15
timestamp 1607194113
transform 1 0 19384 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_15
timestamp 1607194113
transform 1 0 19292 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_208
timestamp 1607194113
transform 1 0 19660 0 1 8000
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap13_15
timestamp 1607194113
transform 1 0 19384 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_15
timestamp 1607194113
transform 1 0 19292 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap14_16
timestamp 1607194113
transform 1 0 20488 0 -1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap14_16
timestamp 1607194113
transform 1 0 20396 0 -1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap13_16
timestamp 1607194113
transform 1 0 20488 0 1 8000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap13_16
timestamp 1607194113
transform 1 0 20396 0 1 8000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_0
timestamp 1607194113
transform 1 0 2732 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 1904 0 1 9088
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_255
timestamp 1607194113
transform 1 0 3100 0 1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap15_0
timestamp 1607194113
transform 1 0 2824 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_254
timestamp 1607194113
transform 1 0 4204 0 1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap15_1
timestamp 1607194113
transform 1 0 3928 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_1
timestamp 1607194113
transform 1 0 3836 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_253
timestamp 1607194113
transform 1 0 5308 0 1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap15_2
timestamp 1607194113
transform 1 0 5032 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_2
timestamp 1607194113
transform 1 0 4940 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_252
timestamp 1607194113
transform 1 0 6412 0 1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap15_3
timestamp 1607194113
transform 1 0 6136 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_3
timestamp 1607194113
transform 1 0 6044 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap15_4
timestamp 1607194113
transform 1 0 7240 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_4
timestamp 1607194113
transform 1 0 7148 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_251
timestamp 1607194113
transform 1 0 7516 0 1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_250
timestamp 1607194113
transform 1 0 8620 0 1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap15_5
timestamp 1607194113
transform 1 0 8344 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_5
timestamp 1607194113
transform 1 0 8252 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_249
timestamp 1607194113
transform 1 0 9724 0 1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap15_6
timestamp 1607194113
transform 1 0 9448 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_6
timestamp 1607194113
transform 1 0 9356 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_248
timestamp 1607194113
transform 1 0 10828 0 1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap15_7
timestamp 1607194113
transform 1 0 10552 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_7
timestamp 1607194113
transform 1 0 10460 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap15_8
timestamp 1607194113
transform 1 0 11656 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_8
timestamp 1607194113
transform 1 0 11564 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap15_9
timestamp 1607194113
transform 1 0 12760 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_9
timestamp 1607194113
transform 1 0 12668 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_247
timestamp 1607194113
transform 1 0 11932 0 1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_246
timestamp 1607194113
transform 1 0 13036 0 1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_245
timestamp 1607194113
transform 1 0 14140 0 1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap15_10
timestamp 1607194113
transform 1 0 13864 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_10
timestamp 1607194113
transform 1 0 13772 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_244
timestamp 1607194113
transform 1 0 15244 0 1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap15_11
timestamp 1607194113
transform 1 0 14968 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_11
timestamp 1607194113
transform 1 0 14876 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_243
timestamp 1607194113
transform 1 0 16348 0 1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap15_12
timestamp 1607194113
transform 1 0 16072 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_12
timestamp 1607194113
transform 1 0 15980 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap15_13
timestamp 1607194113
transform 1 0 17176 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_13
timestamp 1607194113
transform 1 0 17084 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_14
timestamp 1607194113
transform 1 0 18188 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_242
timestamp 1607194113
transform 1 0 17452 0 1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_241
timestamp 1607194113
transform 1 0 18556 0 1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap15_14
timestamp 1607194113
transform 1 0 18280 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_8_240
timestamp 1607194113
transform 1 0 19660 0 1 9088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap15_15
timestamp 1607194113
transform 1 0 19384 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_15
timestamp 1607194113
transform 1 0 19292 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap15_16
timestamp 1607194113
transform 1 0 20488 0 1 9088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap15_16
timestamp 1607194113
transform 1 0 20396 0 1 9088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_0
timestamp 1607194113
transform 1 0 2732 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_31
timestamp 1607194113
transform 1 0 1996 0 -1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_30
timestamp 1607194113
transform 1 0 1904 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_0
timestamp 1607194113
transform 1 0 3100 0 -1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap16_0
timestamp 1607194113
transform 1 0 2824 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_1
timestamp 1607194113
transform 1 0 4204 0 -1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap16_1
timestamp 1607194113
transform 1 0 3928 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_1
timestamp 1607194113
transform 1 0 3836 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_2
timestamp 1607194113
transform 1 0 5308 0 -1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap16_2
timestamp 1607194113
transform 1 0 5032 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_2
timestamp 1607194113
transform 1 0 4940 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_3
timestamp 1607194113
transform 1 0 6412 0 -1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap16_3
timestamp 1607194113
transform 1 0 6136 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_3
timestamp 1607194113
transform 1 0 6044 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap16_4
timestamp 1607194113
transform 1 0 7240 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_4
timestamp 1607194113
transform 1 0 7148 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_4
timestamp 1607194113
transform 1 0 7516 0 -1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_5
timestamp 1607194113
transform 1 0 8620 0 -1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap16_5
timestamp 1607194113
transform 1 0 8344 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_5
timestamp 1607194113
transform 1 0 8252 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_6
timestamp 1607194113
transform 1 0 9724 0 -1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap16_6
timestamp 1607194113
transform 1 0 9448 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_6
timestamp 1607194113
transform 1 0 9356 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_7
timestamp 1607194113
transform 1 0 10828 0 -1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap16_7
timestamp 1607194113
transform 1 0 10552 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_7
timestamp 1607194113
transform 1 0 10460 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap16_8
timestamp 1607194113
transform 1 0 11656 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_8
timestamp 1607194113
transform 1 0 11564 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap16_9
timestamp 1607194113
transform 1 0 12760 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_9
timestamp 1607194113
transform 1 0 12668 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_8
timestamp 1607194113
transform 1 0 11932 0 -1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_9
timestamp 1607194113
transform 1 0 13036 0 -1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_10
timestamp 1607194113
transform 1 0 14140 0 -1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap16_10
timestamp 1607194113
transform 1 0 13864 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_10
timestamp 1607194113
transform 1 0 13772 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_11
timestamp 1607194113
transform 1 0 15244 0 -1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap16_11
timestamp 1607194113
transform 1 0 14968 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_11
timestamp 1607194113
transform 1 0 14876 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_12
timestamp 1607194113
transform 1 0 16348 0 -1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap16_12
timestamp 1607194113
transform 1 0 16072 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_12
timestamp 1607194113
transform 1 0 15980 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap16_13
timestamp 1607194113
transform 1 0 17176 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_13
timestamp 1607194113
transform 1 0 17084 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_14
timestamp 1607194113
transform 1 0 18188 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_13
timestamp 1607194113
transform 1 0 17452 0 -1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_14
timestamp 1607194113
transform 1 0 18556 0 -1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap16_14
timestamp 1607194113
transform 1 0 18280 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_15
timestamp 1607194113
transform 1 0 19660 0 -1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap16_15
timestamp 1607194113
transform 1 0 19384 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_15
timestamp 1607194113
transform 1 0 19292 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap16_16
timestamp 1607194113
transform 1 0 20488 0 -1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap16_16
timestamp 1607194113
transform 1 0 20396 0 -1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_0
timestamp 1607194113
transform 1 0 2732 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_33
timestamp 1607194113
transform 1 0 1996 0 1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_32
timestamp 1607194113
transform 1 0 1904 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_31
timestamp 1607194113
transform 1 0 3100 0 1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap17_0
timestamp 1607194113
transform 1 0 2824 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_30
timestamp 1607194113
transform 1 0 4204 0 1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap17_1
timestamp 1607194113
transform 1 0 3928 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_1
timestamp 1607194113
transform 1 0 3836 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_29
timestamp 1607194113
transform 1 0 5308 0 1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap17_2
timestamp 1607194113
transform 1 0 5032 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_2
timestamp 1607194113
transform 1 0 4940 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_28
timestamp 1607194113
transform 1 0 6412 0 1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap17_3
timestamp 1607194113
transform 1 0 6136 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_3
timestamp 1607194113
transform 1 0 6044 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap17_4
timestamp 1607194113
transform 1 0 7240 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_4
timestamp 1607194113
transform 1 0 7148 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_27
timestamp 1607194113
transform 1 0 7516 0 1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_26
timestamp 1607194113
transform 1 0 8620 0 1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap17_5
timestamp 1607194113
transform 1 0 8344 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_5
timestamp 1607194113
transform 1 0 8252 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_25
timestamp 1607194113
transform 1 0 9724 0 1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap17_6
timestamp 1607194113
transform 1 0 9448 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_6
timestamp 1607194113
transform 1 0 9356 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_24
timestamp 1607194113
transform 1 0 10828 0 1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap17_7
timestamp 1607194113
transform 1 0 10552 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_7
timestamp 1607194113
transform 1 0 10460 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap17_8
timestamp 1607194113
transform 1 0 11656 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_8
timestamp 1607194113
transform 1 0 11564 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap17_9
timestamp 1607194113
transform 1 0 12760 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_9
timestamp 1607194113
transform 1 0 12668 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_23
timestamp 1607194113
transform 1 0 11932 0 1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_22
timestamp 1607194113
transform 1 0 13036 0 1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_21
timestamp 1607194113
transform 1 0 14140 0 1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap17_10
timestamp 1607194113
transform 1 0 13864 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_10
timestamp 1607194113
transform 1 0 13772 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_20
timestamp 1607194113
transform 1 0 15244 0 1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap17_11
timestamp 1607194113
transform 1 0 14968 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_11
timestamp 1607194113
transform 1 0 14876 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_19
timestamp 1607194113
transform 1 0 16348 0 1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap17_12
timestamp 1607194113
transform 1 0 16072 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_12
timestamp 1607194113
transform 1 0 15980 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap17_13
timestamp 1607194113
transform 1 0 17176 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_13
timestamp 1607194113
transform 1 0 17084 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_14
timestamp 1607194113
transform 1 0 18188 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_18
timestamp 1607194113
transform 1 0 17452 0 1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_17
timestamp 1607194113
transform 1 0 18556 0 1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap17_14
timestamp 1607194113
transform 1 0 18280 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_16
timestamp 1607194113
transform 1 0 19660 0 1 10176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap17_15
timestamp 1607194113
transform 1 0 19384 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_15
timestamp 1607194113
transform 1 0 19292 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap17_16
timestamp 1607194113
transform 1 0 20488 0 1 10176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap17_16
timestamp 1607194113
transform 1 0 20396 0 1 10176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_0
timestamp 1607194113
transform 1 0 2732 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_35
timestamp 1607194113
transform 1 0 1996 0 -1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_34
timestamp 1607194113
transform 1 0 1904 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_32
timestamp 1607194113
transform 1 0 3100 0 -1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap18_0
timestamp 1607194113
transform 1 0 2824 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_33
timestamp 1607194113
transform 1 0 4204 0 -1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap18_1
timestamp 1607194113
transform 1 0 3928 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_1
timestamp 1607194113
transform 1 0 3836 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_34
timestamp 1607194113
transform 1 0 5308 0 -1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap18_2
timestamp 1607194113
transform 1 0 5032 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_2
timestamp 1607194113
transform 1 0 4940 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_35
timestamp 1607194113
transform 1 0 6412 0 -1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap18_3
timestamp 1607194113
transform 1 0 6136 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_3
timestamp 1607194113
transform 1 0 6044 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap18_4
timestamp 1607194113
transform 1 0 7240 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_4
timestamp 1607194113
transform 1 0 7148 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_36
timestamp 1607194113
transform 1 0 7516 0 -1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_37
timestamp 1607194113
transform 1 0 8620 0 -1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap18_5
timestamp 1607194113
transform 1 0 8344 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_5
timestamp 1607194113
transform 1 0 8252 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_38
timestamp 1607194113
transform 1 0 9724 0 -1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap18_6
timestamp 1607194113
transform 1 0 9448 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_6
timestamp 1607194113
transform 1 0 9356 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_39
timestamp 1607194113
transform 1 0 10828 0 -1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap18_7
timestamp 1607194113
transform 1 0 10552 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_7
timestamp 1607194113
transform 1 0 10460 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap18_8
timestamp 1607194113
transform 1 0 11656 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_8
timestamp 1607194113
transform 1 0 11564 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap18_9
timestamp 1607194113
transform 1 0 12760 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_9
timestamp 1607194113
transform 1 0 12668 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_40
timestamp 1607194113
transform 1 0 11932 0 -1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_41
timestamp 1607194113
transform 1 0 13036 0 -1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_42
timestamp 1607194113
transform 1 0 14140 0 -1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap18_10
timestamp 1607194113
transform 1 0 13864 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_10
timestamp 1607194113
transform 1 0 13772 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_43
timestamp 1607194113
transform 1 0 15244 0 -1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap18_11
timestamp 1607194113
transform 1 0 14968 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_11
timestamp 1607194113
transform 1 0 14876 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_44
timestamp 1607194113
transform 1 0 16348 0 -1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap18_12
timestamp 1607194113
transform 1 0 16072 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_12
timestamp 1607194113
transform 1 0 15980 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap18_13
timestamp 1607194113
transform 1 0 17176 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_13
timestamp 1607194113
transform 1 0 17084 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_14
timestamp 1607194113
transform 1 0 18188 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_45
timestamp 1607194113
transform 1 0 17452 0 -1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_46
timestamp 1607194113
transform 1 0 18556 0 -1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap18_14
timestamp 1607194113
transform 1 0 18280 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_47
timestamp 1607194113
transform 1 0 19660 0 -1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap18_15
timestamp 1607194113
transform 1 0 19384 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_15
timestamp 1607194113
transform 1 0 19292 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap18_16
timestamp 1607194113
transform 1 0 20488 0 -1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap18_16
timestamp 1607194113
transform 1 0 20396 0 -1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_0
timestamp 1607194113
transform 1 0 2732 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_39
timestamp 1607194113
transform 1 0 1996 0 -1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_38
timestamp 1607194113
transform 1 0 1904 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_0
timestamp 1607194113
transform 1 0 2732 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_37
timestamp 1607194113
transform 1 0 1996 0 1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_36
timestamp 1607194113
transform 1 0 1904 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_64
timestamp 1607194113
transform 1 0 3100 0 -1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap20_0
timestamp 1607194113
transform 1 0 2824 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_63
timestamp 1607194113
transform 1 0 3100 0 1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap19_0
timestamp 1607194113
transform 1 0 2824 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_65
timestamp 1607194113
transform 1 0 4204 0 -1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap20_1
timestamp 1607194113
transform 1 0 3928 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_1
timestamp 1607194113
transform 1 0 3836 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_62
timestamp 1607194113
transform 1 0 4204 0 1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap19_1
timestamp 1607194113
transform 1 0 3928 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_1
timestamp 1607194113
transform 1 0 3836 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_66
timestamp 1607194113
transform 1 0 5308 0 -1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap20_2
timestamp 1607194113
transform 1 0 5032 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_2
timestamp 1607194113
transform 1 0 4940 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_61
timestamp 1607194113
transform 1 0 5308 0 1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap19_2
timestamp 1607194113
transform 1 0 5032 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_2
timestamp 1607194113
transform 1 0 4940 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_67
timestamp 1607194113
transform 1 0 6412 0 -1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap20_3
timestamp 1607194113
transform 1 0 6136 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_3
timestamp 1607194113
transform 1 0 6044 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_60
timestamp 1607194113
transform 1 0 6412 0 1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap19_3
timestamp 1607194113
transform 1 0 6136 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_3
timestamp 1607194113
transform 1 0 6044 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap20_4
timestamp 1607194113
transform 1 0 7240 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_4
timestamp 1607194113
transform 1 0 7148 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap19_4
timestamp 1607194113
transform 1 0 7240 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_4
timestamp 1607194113
transform 1 0 7148 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_68
timestamp 1607194113
transform 1 0 7516 0 -1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_59
timestamp 1607194113
transform 1 0 7516 0 1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_69
timestamp 1607194113
transform 1 0 8620 0 -1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap20_5
timestamp 1607194113
transform 1 0 8344 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_5
timestamp 1607194113
transform 1 0 8252 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_58
timestamp 1607194113
transform 1 0 8620 0 1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap19_5
timestamp 1607194113
transform 1 0 8344 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_5
timestamp 1607194113
transform 1 0 8252 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_70
timestamp 1607194113
transform 1 0 9724 0 -1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap20_6
timestamp 1607194113
transform 1 0 9448 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_6
timestamp 1607194113
transform 1 0 9356 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_57
timestamp 1607194113
transform 1 0 9724 0 1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap19_6
timestamp 1607194113
transform 1 0 9448 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_6
timestamp 1607194113
transform 1 0 9356 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_71
timestamp 1607194113
transform 1 0 10828 0 -1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap20_7
timestamp 1607194113
transform 1 0 10552 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_7
timestamp 1607194113
transform 1 0 10460 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_56
timestamp 1607194113
transform 1 0 10828 0 1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap19_7
timestamp 1607194113
transform 1 0 10552 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_7
timestamp 1607194113
transform 1 0 10460 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap20_8
timestamp 1607194113
transform 1 0 11656 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_8
timestamp 1607194113
transform 1 0 11564 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap19_8
timestamp 1607194113
transform 1 0 11656 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_8
timestamp 1607194113
transform 1 0 11564 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap20_9
timestamp 1607194113
transform 1 0 12760 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_9
timestamp 1607194113
transform 1 0 12668 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_72
timestamp 1607194113
transform 1 0 11932 0 -1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap19_9
timestamp 1607194113
transform 1 0 12760 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_9
timestamp 1607194113
transform 1 0 12668 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_55
timestamp 1607194113
transform 1 0 11932 0 1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_73
timestamp 1607194113
transform 1 0 13036 0 -1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_54
timestamp 1607194113
transform 1 0 13036 0 1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_74
timestamp 1607194113
transform 1 0 14140 0 -1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap20_10
timestamp 1607194113
transform 1 0 13864 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_10
timestamp 1607194113
transform 1 0 13772 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_53
timestamp 1607194113
transform 1 0 14140 0 1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap19_10
timestamp 1607194113
transform 1 0 13864 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_10
timestamp 1607194113
transform 1 0 13772 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_75
timestamp 1607194113
transform 1 0 15244 0 -1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap20_11
timestamp 1607194113
transform 1 0 14968 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_11
timestamp 1607194113
transform 1 0 14876 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_52
timestamp 1607194113
transform 1 0 15244 0 1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap19_11
timestamp 1607194113
transform 1 0 14968 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_11
timestamp 1607194113
transform 1 0 14876 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_76
timestamp 1607194113
transform 1 0 16348 0 -1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap20_12
timestamp 1607194113
transform 1 0 16072 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_12
timestamp 1607194113
transform 1 0 15980 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_51
timestamp 1607194113
transform 1 0 16348 0 1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap19_12
timestamp 1607194113
transform 1 0 16072 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_12
timestamp 1607194113
transform 1 0 15980 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap20_13
timestamp 1607194113
transform 1 0 17176 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_13
timestamp 1607194113
transform 1 0 17084 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap19_13
timestamp 1607194113
transform 1 0 17176 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_13
timestamp 1607194113
transform 1 0 17084 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_14
timestamp 1607194113
transform 1 0 18188 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_77
timestamp 1607194113
transform 1 0 17452 0 -1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_14
timestamp 1607194113
transform 1 0 18188 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_50
timestamp 1607194113
transform 1 0 17452 0 1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_78
timestamp 1607194113
transform 1 0 18556 0 -1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap20_14
timestamp 1607194113
transform 1 0 18280 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_49
timestamp 1607194113
transform 1 0 18556 0 1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap19_14
timestamp 1607194113
transform 1 0 18280 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_79
timestamp 1607194113
transform 1 0 19660 0 -1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap20_15
timestamp 1607194113
transform 1 0 19384 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_15
timestamp 1607194113
transform 1 0 19292 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_48
timestamp 1607194113
transform 1 0 19660 0 1 11264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap19_15
timestamp 1607194113
transform 1 0 19384 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_15
timestamp 1607194113
transform 1 0 19292 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap20_16
timestamp 1607194113
transform 1 0 20488 0 -1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap20_16
timestamp 1607194113
transform 1 0 20396 0 -1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap19_16
timestamp 1607194113
transform 1 0 20488 0 1 11264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap19_16
timestamp 1607194113
transform 1 0 20396 0 1 11264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_0
timestamp 1607194113
transform 1 0 2732 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_41
timestamp 1607194113
transform 1 0 1996 0 1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_40
timestamp 1607194113
transform 1 0 1904 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_95
timestamp 1607194113
transform 1 0 3100 0 1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap21_0
timestamp 1607194113
transform 1 0 2824 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_94
timestamp 1607194113
transform 1 0 4204 0 1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap21_1
timestamp 1607194113
transform 1 0 3928 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_1
timestamp 1607194113
transform 1 0 3836 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_93
timestamp 1607194113
transform 1 0 5308 0 1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap21_2
timestamp 1607194113
transform 1 0 5032 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_2
timestamp 1607194113
transform 1 0 4940 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_92
timestamp 1607194113
transform 1 0 6412 0 1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap21_3
timestamp 1607194113
transform 1 0 6136 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_3
timestamp 1607194113
transform 1 0 6044 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap21_4
timestamp 1607194113
transform 1 0 7240 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_4
timestamp 1607194113
transform 1 0 7148 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_91
timestamp 1607194113
transform 1 0 7516 0 1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_90
timestamp 1607194113
transform 1 0 8620 0 1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap21_5
timestamp 1607194113
transform 1 0 8344 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_5
timestamp 1607194113
transform 1 0 8252 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_89
timestamp 1607194113
transform 1 0 9724 0 1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap21_6
timestamp 1607194113
transform 1 0 9448 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_6
timestamp 1607194113
transform 1 0 9356 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_88
timestamp 1607194113
transform 1 0 10828 0 1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap21_7
timestamp 1607194113
transform 1 0 10552 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_7
timestamp 1607194113
transform 1 0 10460 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap21_8
timestamp 1607194113
transform 1 0 11656 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_8
timestamp 1607194113
transform 1 0 11564 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap21_9
timestamp 1607194113
transform 1 0 12760 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_9
timestamp 1607194113
transform 1 0 12668 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_87
timestamp 1607194113
transform 1 0 11932 0 1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_86
timestamp 1607194113
transform 1 0 13036 0 1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_85
timestamp 1607194113
transform 1 0 14140 0 1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap21_10
timestamp 1607194113
transform 1 0 13864 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_10
timestamp 1607194113
transform 1 0 13772 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_84
timestamp 1607194113
transform 1 0 15244 0 1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap21_11
timestamp 1607194113
transform 1 0 14968 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_11
timestamp 1607194113
transform 1 0 14876 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_83
timestamp 1607194113
transform 1 0 16348 0 1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap21_12
timestamp 1607194113
transform 1 0 16072 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_12
timestamp 1607194113
transform 1 0 15980 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap21_13
timestamp 1607194113
transform 1 0 17176 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_13
timestamp 1607194113
transform 1 0 17084 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_14
timestamp 1607194113
transform 1 0 18188 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_82
timestamp 1607194113
transform 1 0 17452 0 1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_81
timestamp 1607194113
transform 1 0 18556 0 1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap21_14
timestamp 1607194113
transform 1 0 18280 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_80
timestamp 1607194113
transform 1 0 19660 0 1 12352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap21_15
timestamp 1607194113
transform 1 0 19384 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_15
timestamp 1607194113
transform 1 0 19292 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap21_16
timestamp 1607194113
transform 1 0 20488 0 1 12352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap21_16
timestamp 1607194113
transform 1 0 20396 0 1 12352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_0
timestamp 1607194113
transform 1 0 2732 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_43
timestamp 1607194113
transform 1 0 1996 0 -1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_42
timestamp 1607194113
transform 1 0 1904 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_96
timestamp 1607194113
transform 1 0 3100 0 -1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap22_0
timestamp 1607194113
transform 1 0 2824 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_97
timestamp 1607194113
transform 1 0 4204 0 -1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap22_1
timestamp 1607194113
transform 1 0 3928 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_1
timestamp 1607194113
transform 1 0 3836 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_98
timestamp 1607194113
transform 1 0 5308 0 -1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap22_2
timestamp 1607194113
transform 1 0 5032 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_2
timestamp 1607194113
transform 1 0 4940 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_99
timestamp 1607194113
transform 1 0 6412 0 -1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap22_3
timestamp 1607194113
transform 1 0 6136 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_3
timestamp 1607194113
transform 1 0 6044 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap22_4
timestamp 1607194113
transform 1 0 7240 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_4
timestamp 1607194113
transform 1 0 7148 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_100
timestamp 1607194113
transform 1 0 7516 0 -1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_101
timestamp 1607194113
transform 1 0 8620 0 -1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap22_5
timestamp 1607194113
transform 1 0 8344 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_5
timestamp 1607194113
transform 1 0 8252 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_102
timestamp 1607194113
transform 1 0 9724 0 -1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap22_6
timestamp 1607194113
transform 1 0 9448 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_6
timestamp 1607194113
transform 1 0 9356 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_103
timestamp 1607194113
transform 1 0 10828 0 -1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap22_7
timestamp 1607194113
transform 1 0 10552 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_7
timestamp 1607194113
transform 1 0 10460 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap22_8
timestamp 1607194113
transform 1 0 11656 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_8
timestamp 1607194113
transform 1 0 11564 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap22_9
timestamp 1607194113
transform 1 0 12760 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_9
timestamp 1607194113
transform 1 0 12668 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_104
timestamp 1607194113
transform 1 0 11932 0 -1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_105
timestamp 1607194113
transform 1 0 13036 0 -1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_106
timestamp 1607194113
transform 1 0 14140 0 -1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap22_10
timestamp 1607194113
transform 1 0 13864 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_10
timestamp 1607194113
transform 1 0 13772 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_107
timestamp 1607194113
transform 1 0 15244 0 -1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap22_11
timestamp 1607194113
transform 1 0 14968 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_11
timestamp 1607194113
transform 1 0 14876 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_108
timestamp 1607194113
transform 1 0 16348 0 -1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap22_12
timestamp 1607194113
transform 1 0 16072 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_12
timestamp 1607194113
transform 1 0 15980 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap22_13
timestamp 1607194113
transform 1 0 17176 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_13
timestamp 1607194113
transform 1 0 17084 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_14
timestamp 1607194113
transform 1 0 18188 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_109
timestamp 1607194113
transform 1 0 17452 0 -1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_110
timestamp 1607194113
transform 1 0 18556 0 -1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap22_14
timestamp 1607194113
transform 1 0 18280 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_111
timestamp 1607194113
transform 1 0 19660 0 -1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap22_15
timestamp 1607194113
transform 1 0 19384 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_15
timestamp 1607194113
transform 1 0 19292 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap22_16
timestamp 1607194113
transform 1 0 20488 0 -1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap22_16
timestamp 1607194113
transform 1 0 20396 0 -1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_0
timestamp 1607194113
transform 1 0 2732 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_7
timestamp 1607194113
transform 1 0 1904 0 1 13440
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_127
timestamp 1607194113
transform 1 0 3100 0 1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap23_0
timestamp 1607194113
transform 1 0 2824 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_126
timestamp 1607194113
transform 1 0 4204 0 1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap23_1
timestamp 1607194113
transform 1 0 3928 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_1
timestamp 1607194113
transform 1 0 3836 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_125
timestamp 1607194113
transform 1 0 5308 0 1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap23_2
timestamp 1607194113
transform 1 0 5032 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_2
timestamp 1607194113
transform 1 0 4940 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_124
timestamp 1607194113
transform 1 0 6412 0 1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap23_3
timestamp 1607194113
transform 1 0 6136 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_3
timestamp 1607194113
transform 1 0 6044 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap23_4
timestamp 1607194113
transform 1 0 7240 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_4
timestamp 1607194113
transform 1 0 7148 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_123
timestamp 1607194113
transform 1 0 7516 0 1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_122
timestamp 1607194113
transform 1 0 8620 0 1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap23_5
timestamp 1607194113
transform 1 0 8344 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_5
timestamp 1607194113
transform 1 0 8252 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_121
timestamp 1607194113
transform 1 0 9724 0 1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap23_6
timestamp 1607194113
transform 1 0 9448 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_6
timestamp 1607194113
transform 1 0 9356 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_120
timestamp 1607194113
transform 1 0 10828 0 1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap23_7
timestamp 1607194113
transform 1 0 10552 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_7
timestamp 1607194113
transform 1 0 10460 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap23_8
timestamp 1607194113
transform 1 0 11656 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_8
timestamp 1607194113
transform 1 0 11564 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap23_9
timestamp 1607194113
transform 1 0 12760 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_9
timestamp 1607194113
transform 1 0 12668 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_119
timestamp 1607194113
transform 1 0 11932 0 1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_118
timestamp 1607194113
transform 1 0 13036 0 1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_117
timestamp 1607194113
transform 1 0 14140 0 1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap23_10
timestamp 1607194113
transform 1 0 13864 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_10
timestamp 1607194113
transform 1 0 13772 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_116
timestamp 1607194113
transform 1 0 15244 0 1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap23_11
timestamp 1607194113
transform 1 0 14968 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_11
timestamp 1607194113
transform 1 0 14876 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_115
timestamp 1607194113
transform 1 0 16348 0 1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap23_12
timestamp 1607194113
transform 1 0 16072 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_12
timestamp 1607194113
transform 1 0 15980 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap23_13
timestamp 1607194113
transform 1 0 17176 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_13
timestamp 1607194113
transform 1 0 17084 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_14
timestamp 1607194113
transform 1 0 18188 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_114
timestamp 1607194113
transform 1 0 17452 0 1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_113
timestamp 1607194113
transform 1 0 18556 0 1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap23_14
timestamp 1607194113
transform 1 0 18280 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_7_112
timestamp 1607194113
transform 1 0 19660 0 1 13440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap23_15
timestamp 1607194113
transform 1 0 19384 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_15
timestamp 1607194113
transform 1 0 19292 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap23_16
timestamp 1607194113
transform 1 0 20488 0 1 13440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap23_16
timestamp 1607194113
transform 1 0 20396 0 1 13440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_0
timestamp 1607194113
transform 1 0 2732 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_45
timestamp 1607194113
transform 1 0 1996 0 -1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_44
timestamp 1607194113
transform 1 0 1904 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_0
timestamp 1607194113
transform 1 0 3100 0 -1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap24_0
timestamp 1607194113
transform 1 0 2824 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_1
timestamp 1607194113
transform 1 0 4204 0 -1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap24_1
timestamp 1607194113
transform 1 0 3928 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_1
timestamp 1607194113
transform 1 0 3836 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_2
timestamp 1607194113
transform 1 0 5308 0 -1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap24_2
timestamp 1607194113
transform 1 0 5032 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_2
timestamp 1607194113
transform 1 0 4940 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_3
timestamp 1607194113
transform 1 0 6412 0 -1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap24_3
timestamp 1607194113
transform 1 0 6136 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_3
timestamp 1607194113
transform 1 0 6044 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap24_4
timestamp 1607194113
transform 1 0 7240 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_4
timestamp 1607194113
transform 1 0 7148 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_4
timestamp 1607194113
transform 1 0 7516 0 -1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_5
timestamp 1607194113
transform 1 0 8620 0 -1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap24_5
timestamp 1607194113
transform 1 0 8344 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_5
timestamp 1607194113
transform 1 0 8252 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_6
timestamp 1607194113
transform 1 0 9724 0 -1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap24_6
timestamp 1607194113
transform 1 0 9448 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_6
timestamp 1607194113
transform 1 0 9356 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_7
timestamp 1607194113
transform 1 0 10828 0 -1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap24_7
timestamp 1607194113
transform 1 0 10552 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_7
timestamp 1607194113
transform 1 0 10460 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap24_8
timestamp 1607194113
transform 1 0 11656 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_8
timestamp 1607194113
transform 1 0 11564 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap24_9
timestamp 1607194113
transform 1 0 12760 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_9
timestamp 1607194113
transform 1 0 12668 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_8
timestamp 1607194113
transform 1 0 11932 0 -1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_9
timestamp 1607194113
transform 1 0 13036 0 -1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_10
timestamp 1607194113
transform 1 0 14140 0 -1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap24_10
timestamp 1607194113
transform 1 0 13864 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_10
timestamp 1607194113
transform 1 0 13772 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_11
timestamp 1607194113
transform 1 0 15244 0 -1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap24_11
timestamp 1607194113
transform 1 0 14968 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_11
timestamp 1607194113
transform 1 0 14876 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_12
timestamp 1607194113
transform 1 0 16348 0 -1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap24_12
timestamp 1607194113
transform 1 0 16072 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_12
timestamp 1607194113
transform 1 0 15980 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap24_13
timestamp 1607194113
transform 1 0 17176 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_13
timestamp 1607194113
transform 1 0 17084 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_14
timestamp 1607194113
transform 1 0 18188 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_13
timestamp 1607194113
transform 1 0 17452 0 -1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_14
timestamp 1607194113
transform 1 0 18556 0 -1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap24_14
timestamp 1607194113
transform 1 0 18280 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_15
timestamp 1607194113
transform 1 0 19660 0 -1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap24_15
timestamp 1607194113
transform 1 0 19384 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_15
timestamp 1607194113
transform 1 0 19292 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap24_16
timestamp 1607194113
transform 1 0 20488 0 -1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap24_16
timestamp 1607194113
transform 1 0 20396 0 -1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_0
timestamp 1607194113
transform 1 0 2732 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_47
timestamp 1607194113
transform 1 0 1996 0 1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_46
timestamp 1607194113
transform 1 0 1904 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_31
timestamp 1607194113
transform 1 0 3100 0 1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap25_0
timestamp 1607194113
transform 1 0 2824 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_30
timestamp 1607194113
transform 1 0 4204 0 1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap25_1
timestamp 1607194113
transform 1 0 3928 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_1
timestamp 1607194113
transform 1 0 3836 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_29
timestamp 1607194113
transform 1 0 5308 0 1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap25_2
timestamp 1607194113
transform 1 0 5032 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_2
timestamp 1607194113
transform 1 0 4940 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_28
timestamp 1607194113
transform 1 0 6412 0 1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap25_3
timestamp 1607194113
transform 1 0 6136 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_3
timestamp 1607194113
transform 1 0 6044 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap25_4
timestamp 1607194113
transform 1 0 7240 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_4
timestamp 1607194113
transform 1 0 7148 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_27
timestamp 1607194113
transform 1 0 7516 0 1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_26
timestamp 1607194113
transform 1 0 8620 0 1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap25_5
timestamp 1607194113
transform 1 0 8344 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_5
timestamp 1607194113
transform 1 0 8252 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_25
timestamp 1607194113
transform 1 0 9724 0 1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap25_6
timestamp 1607194113
transform 1 0 9448 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_6
timestamp 1607194113
transform 1 0 9356 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_24
timestamp 1607194113
transform 1 0 10828 0 1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap25_7
timestamp 1607194113
transform 1 0 10552 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_7
timestamp 1607194113
transform 1 0 10460 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap25_8
timestamp 1607194113
transform 1 0 11656 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_8
timestamp 1607194113
transform 1 0 11564 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap25_9
timestamp 1607194113
transform 1 0 12760 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_9
timestamp 1607194113
transform 1 0 12668 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_23
timestamp 1607194113
transform 1 0 11932 0 1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_22
timestamp 1607194113
transform 1 0 13036 0 1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_21
timestamp 1607194113
transform 1 0 14140 0 1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap25_10
timestamp 1607194113
transform 1 0 13864 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_10
timestamp 1607194113
transform 1 0 13772 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_20
timestamp 1607194113
transform 1 0 15244 0 1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap25_11
timestamp 1607194113
transform 1 0 14968 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_11
timestamp 1607194113
transform 1 0 14876 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_19
timestamp 1607194113
transform 1 0 16348 0 1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap25_12
timestamp 1607194113
transform 1 0 16072 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_12
timestamp 1607194113
transform 1 0 15980 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap25_13
timestamp 1607194113
transform 1 0 17176 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_13
timestamp 1607194113
transform 1 0 17084 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_14
timestamp 1607194113
transform 1 0 18188 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_18
timestamp 1607194113
transform 1 0 17452 0 1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_17
timestamp 1607194113
transform 1 0 18556 0 1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap25_14
timestamp 1607194113
transform 1 0 18280 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_16
timestamp 1607194113
transform 1 0 19660 0 1 14528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap25_15
timestamp 1607194113
transform 1 0 19384 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_15
timestamp 1607194113
transform 1 0 19292 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap25_16
timestamp 1607194113
transform 1 0 20488 0 1 14528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap25_16
timestamp 1607194113
transform 1 0 20396 0 1 14528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_0
timestamp 1607194113
transform 1 0 2732 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_6
timestamp 1607194113
transform 1 0 1904 0 1 15616
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_0
timestamp 1607194113
transform 1 0 2732 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_49
timestamp 1607194113
transform 1 0 1996 0 -1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_48
timestamp 1607194113
transform 1 0 1904 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_63
timestamp 1607194113
transform 1 0 3100 0 1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap27_0
timestamp 1607194113
transform 1 0 2824 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_32
timestamp 1607194113
transform 1 0 3100 0 -1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap26_0
timestamp 1607194113
transform 1 0 2824 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_62
timestamp 1607194113
transform 1 0 4204 0 1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap27_1
timestamp 1607194113
transform 1 0 3928 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_1
timestamp 1607194113
transform 1 0 3836 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_33
timestamp 1607194113
transform 1 0 4204 0 -1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap26_1
timestamp 1607194113
transform 1 0 3928 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_1
timestamp 1607194113
transform 1 0 3836 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_61
timestamp 1607194113
transform 1 0 5308 0 1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap27_2
timestamp 1607194113
transform 1 0 5032 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_2
timestamp 1607194113
transform 1 0 4940 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_34
timestamp 1607194113
transform 1 0 5308 0 -1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap26_2
timestamp 1607194113
transform 1 0 5032 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_2
timestamp 1607194113
transform 1 0 4940 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_60
timestamp 1607194113
transform 1 0 6412 0 1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap27_3
timestamp 1607194113
transform 1 0 6136 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_3
timestamp 1607194113
transform 1 0 6044 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_35
timestamp 1607194113
transform 1 0 6412 0 -1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap26_3
timestamp 1607194113
transform 1 0 6136 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_3
timestamp 1607194113
transform 1 0 6044 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap27_4
timestamp 1607194113
transform 1 0 7240 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_4
timestamp 1607194113
transform 1 0 7148 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap26_4
timestamp 1607194113
transform 1 0 7240 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_4
timestamp 1607194113
transform 1 0 7148 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_59
timestamp 1607194113
transform 1 0 7516 0 1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_36
timestamp 1607194113
transform 1 0 7516 0 -1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_58
timestamp 1607194113
transform 1 0 8620 0 1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap27_5
timestamp 1607194113
transform 1 0 8344 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_5
timestamp 1607194113
transform 1 0 8252 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_37
timestamp 1607194113
transform 1 0 8620 0 -1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap26_5
timestamp 1607194113
transform 1 0 8344 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_5
timestamp 1607194113
transform 1 0 8252 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_57
timestamp 1607194113
transform 1 0 9724 0 1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap27_6
timestamp 1607194113
transform 1 0 9448 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_6
timestamp 1607194113
transform 1 0 9356 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_38
timestamp 1607194113
transform 1 0 9724 0 -1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap26_6
timestamp 1607194113
transform 1 0 9448 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_6
timestamp 1607194113
transform 1 0 9356 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_56
timestamp 1607194113
transform 1 0 10828 0 1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap27_7
timestamp 1607194113
transform 1 0 10552 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_7
timestamp 1607194113
transform 1 0 10460 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_39
timestamp 1607194113
transform 1 0 10828 0 -1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap26_7
timestamp 1607194113
transform 1 0 10552 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_7
timestamp 1607194113
transform 1 0 10460 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap27_8
timestamp 1607194113
transform 1 0 11656 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_8
timestamp 1607194113
transform 1 0 11564 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap26_8
timestamp 1607194113
transform 1 0 11656 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_8
timestamp 1607194113
transform 1 0 11564 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap27_9
timestamp 1607194113
transform 1 0 12760 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_9
timestamp 1607194113
transform 1 0 12668 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_55
timestamp 1607194113
transform 1 0 11932 0 1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap26_9
timestamp 1607194113
transform 1 0 12760 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_9
timestamp 1607194113
transform 1 0 12668 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_40
timestamp 1607194113
transform 1 0 11932 0 -1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_54
timestamp 1607194113
transform 1 0 13036 0 1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_41
timestamp 1607194113
transform 1 0 13036 0 -1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_53
timestamp 1607194113
transform 1 0 14140 0 1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap27_10
timestamp 1607194113
transform 1 0 13864 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_10
timestamp 1607194113
transform 1 0 13772 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_42
timestamp 1607194113
transform 1 0 14140 0 -1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap26_10
timestamp 1607194113
transform 1 0 13864 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_10
timestamp 1607194113
transform 1 0 13772 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_52
timestamp 1607194113
transform 1 0 15244 0 1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap27_11
timestamp 1607194113
transform 1 0 14968 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_11
timestamp 1607194113
transform 1 0 14876 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_43
timestamp 1607194113
transform 1 0 15244 0 -1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap26_11
timestamp 1607194113
transform 1 0 14968 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_11
timestamp 1607194113
transform 1 0 14876 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_51
timestamp 1607194113
transform 1 0 16348 0 1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap27_12
timestamp 1607194113
transform 1 0 16072 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_12
timestamp 1607194113
transform 1 0 15980 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_44
timestamp 1607194113
transform 1 0 16348 0 -1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap26_12
timestamp 1607194113
transform 1 0 16072 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_12
timestamp 1607194113
transform 1 0 15980 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap27_13
timestamp 1607194113
transform 1 0 17176 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_13
timestamp 1607194113
transform 1 0 17084 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap26_13
timestamp 1607194113
transform 1 0 17176 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_13
timestamp 1607194113
transform 1 0 17084 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_14
timestamp 1607194113
transform 1 0 18188 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_50
timestamp 1607194113
transform 1 0 17452 0 1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_14
timestamp 1607194113
transform 1 0 18188 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_45
timestamp 1607194113
transform 1 0 17452 0 -1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_49
timestamp 1607194113
transform 1 0 18556 0 1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap27_14
timestamp 1607194113
transform 1 0 18280 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_46
timestamp 1607194113
transform 1 0 18556 0 -1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap26_14
timestamp 1607194113
transform 1 0 18280 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_48
timestamp 1607194113
transform 1 0 19660 0 1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap27_15
timestamp 1607194113
transform 1 0 19384 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_15
timestamp 1607194113
transform 1 0 19292 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_6_47
timestamp 1607194113
transform 1 0 19660 0 -1 15616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap26_15
timestamp 1607194113
transform 1 0 19384 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_15
timestamp 1607194113
transform 1 0 19292 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap27_16
timestamp 1607194113
transform 1 0 20488 0 1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap27_16
timestamp 1607194113
transform 1 0 20396 0 1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap26_16
timestamp 1607194113
transform 1 0 20488 0 -1 15616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap26_16
timestamp 1607194113
transform 1 0 20396 0 -1 15616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_0
timestamp 1607194113
transform 1 0 2732 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_51
timestamp 1607194113
transform 1 0 1996 0 -1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_50
timestamp 1607194113
transform 1 0 1904 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_0
timestamp 1607194113
transform 1 0 3100 0 -1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap28_0
timestamp 1607194113
transform 1 0 2824 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_1
timestamp 1607194113
transform 1 0 4204 0 -1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap28_1
timestamp 1607194113
transform 1 0 3928 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_1
timestamp 1607194113
transform 1 0 3836 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_2
timestamp 1607194113
transform 1 0 5308 0 -1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap28_2
timestamp 1607194113
transform 1 0 5032 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_2
timestamp 1607194113
transform 1 0 4940 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_3
timestamp 1607194113
transform 1 0 6412 0 -1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap28_3
timestamp 1607194113
transform 1 0 6136 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_3
timestamp 1607194113
transform 1 0 6044 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap28_4
timestamp 1607194113
transform 1 0 7240 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_4
timestamp 1607194113
transform 1 0 7148 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_4
timestamp 1607194113
transform 1 0 7516 0 -1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_5
timestamp 1607194113
transform 1 0 8620 0 -1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap28_5
timestamp 1607194113
transform 1 0 8344 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_5
timestamp 1607194113
transform 1 0 8252 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_6
timestamp 1607194113
transform 1 0 9724 0 -1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap28_6
timestamp 1607194113
transform 1 0 9448 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_6
timestamp 1607194113
transform 1 0 9356 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_7
timestamp 1607194113
transform 1 0 10828 0 -1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap28_7
timestamp 1607194113
transform 1 0 10552 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_7
timestamp 1607194113
transform 1 0 10460 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap28_8
timestamp 1607194113
transform 1 0 11656 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_8
timestamp 1607194113
transform 1 0 11564 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap28_9
timestamp 1607194113
transform 1 0 12760 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_9
timestamp 1607194113
transform 1 0 12668 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_8
timestamp 1607194113
transform 1 0 11932 0 -1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_9
timestamp 1607194113
transform 1 0 13036 0 -1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_10
timestamp 1607194113
transform 1 0 14140 0 -1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap28_10
timestamp 1607194113
transform 1 0 13864 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_10
timestamp 1607194113
transform 1 0 13772 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_11
timestamp 1607194113
transform 1 0 15244 0 -1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap28_11
timestamp 1607194113
transform 1 0 14968 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_11
timestamp 1607194113
transform 1 0 14876 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_12
timestamp 1607194113
transform 1 0 16348 0 -1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap28_12
timestamp 1607194113
transform 1 0 16072 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_12
timestamp 1607194113
transform 1 0 15980 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap28_13
timestamp 1607194113
transform 1 0 17176 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_13
timestamp 1607194113
transform 1 0 17084 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_14
timestamp 1607194113
transform 1 0 18188 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_13
timestamp 1607194113
transform 1 0 17452 0 -1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_14
timestamp 1607194113
transform 1 0 18556 0 -1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap28_14
timestamp 1607194113
transform 1 0 18280 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_15
timestamp 1607194113
transform 1 0 19660 0 -1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap28_15
timestamp 1607194113
transform 1 0 19384 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_15
timestamp 1607194113
transform 1 0 19292 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap28_16
timestamp 1607194113
transform 1 0 20488 0 -1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap28_16
timestamp 1607194113
transform 1 0 20396 0 -1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_0
timestamp 1607194113
transform 1 0 2732 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_5
timestamp 1607194113
transform 1 0 1904 0 1 16704
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_31
timestamp 1607194113
transform 1 0 3100 0 1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap29_0
timestamp 1607194113
transform 1 0 2824 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_30
timestamp 1607194113
transform 1 0 4204 0 1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap29_1
timestamp 1607194113
transform 1 0 3928 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_1
timestamp 1607194113
transform 1 0 3836 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_29
timestamp 1607194113
transform 1 0 5308 0 1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap29_2
timestamp 1607194113
transform 1 0 5032 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_2
timestamp 1607194113
transform 1 0 4940 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_28
timestamp 1607194113
transform 1 0 6412 0 1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap29_3
timestamp 1607194113
transform 1 0 6136 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_3
timestamp 1607194113
transform 1 0 6044 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap29_4
timestamp 1607194113
transform 1 0 7240 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_4
timestamp 1607194113
transform 1 0 7148 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_27
timestamp 1607194113
transform 1 0 7516 0 1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_26
timestamp 1607194113
transform 1 0 8620 0 1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap29_5
timestamp 1607194113
transform 1 0 8344 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_5
timestamp 1607194113
transform 1 0 8252 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_25
timestamp 1607194113
transform 1 0 9724 0 1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap29_6
timestamp 1607194113
transform 1 0 9448 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_6
timestamp 1607194113
transform 1 0 9356 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_24
timestamp 1607194113
transform 1 0 10828 0 1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap29_7
timestamp 1607194113
transform 1 0 10552 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_7
timestamp 1607194113
transform 1 0 10460 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap29_8
timestamp 1607194113
transform 1 0 11656 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_8
timestamp 1607194113
transform 1 0 11564 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap29_9
timestamp 1607194113
transform 1 0 12760 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_9
timestamp 1607194113
transform 1 0 12668 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_23
timestamp 1607194113
transform 1 0 11932 0 1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_22
timestamp 1607194113
transform 1 0 13036 0 1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_21
timestamp 1607194113
transform 1 0 14140 0 1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap29_10
timestamp 1607194113
transform 1 0 13864 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_10
timestamp 1607194113
transform 1 0 13772 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_20
timestamp 1607194113
transform 1 0 15244 0 1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap29_11
timestamp 1607194113
transform 1 0 14968 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_11
timestamp 1607194113
transform 1 0 14876 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_19
timestamp 1607194113
transform 1 0 16348 0 1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap29_12
timestamp 1607194113
transform 1 0 16072 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_12
timestamp 1607194113
transform 1 0 15980 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap29_13
timestamp 1607194113
transform 1 0 17176 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_13
timestamp 1607194113
transform 1 0 17084 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_14
timestamp 1607194113
transform 1 0 18188 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_18
timestamp 1607194113
transform 1 0 17452 0 1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_17
timestamp 1607194113
transform 1 0 18556 0 1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap29_14
timestamp 1607194113
transform 1 0 18280 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_5_16
timestamp 1607194113
transform 1 0 19660 0 1 16704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap29_15
timestamp 1607194113
transform 1 0 19384 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_15
timestamp 1607194113
transform 1 0 19292 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap29_16
timestamp 1607194113
transform 1 0 20488 0 1 16704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap29_16
timestamp 1607194113
transform 1 0 20396 0 1 16704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap30_0
timestamp 1607194113
transform 1 0 2732 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_53
timestamp 1607194113
transform 1 0 1996 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_52
timestamp 1607194113
transform 1 0 1904 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_4_0
timestamp 1607194113
transform 1 0 3100 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap30_0
timestamp 1607194113
transform 1 0 2824 0 -1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_4_1
timestamp 1607194113
transform 1 0 4204 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap30_1
timestamp 1607194113
transform 1 0 3928 0 -1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap30_1
timestamp 1607194113
transform 1 0 3836 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_4_2
timestamp 1607194113
transform 1 0 5308 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap30_2
timestamp 1607194113
transform 1 0 5032 0 -1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap30_2
timestamp 1607194113
transform 1 0 4940 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_4_3
timestamp 1607194113
transform 1 0 6412 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap30_3
timestamp 1607194113
transform 1 0 6136 0 -1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap30_3
timestamp 1607194113
transform 1 0 6044 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap30_4
timestamp 1607194113
transform 1 0 7240 0 -1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap30_4
timestamp 1607194113
transform 1 0 7148 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_4_4
timestamp 1607194113
transform 1 0 7516 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_4_5
timestamp 1607194113
transform 1 0 8620 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap30_5
timestamp 1607194113
transform 1 0 8344 0 -1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap30_5
timestamp 1607194113
transform 1 0 8252 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_4_6
timestamp 1607194113
transform 1 0 9724 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap30_6
timestamp 1607194113
transform 1 0 9448 0 -1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap30_6
timestamp 1607194113
transform 1 0 9356 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_4_7
timestamp 1607194113
transform 1 0 10828 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap30_7
timestamp 1607194113
transform 1 0 10552 0 -1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap30_7
timestamp 1607194113
transform 1 0 10460 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap30_8
timestamp 1607194113
transform 1 0 11656 0 -1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap30_8
timestamp 1607194113
transform 1 0 11564 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_62
timestamp 1607194113
transform 1 0 12760 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_61
timestamp 1607194113
transform 1 0 12024 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_60
timestamp 1607194113
transform 1 0 11932 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_64
timestamp 1607194113
transform 1 0 13588 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_63
timestamp 1607194113
transform 1 0 12852 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_67
timestamp 1607194113
transform 1 0 14508 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_66
timestamp 1607194113
transform 1 0 14416 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_65
timestamp 1607194113
transform 1 0 13680 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_69
timestamp 1607194113
transform 1 0 15336 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_68
timestamp 1607194113
transform 1 0 15244 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_71
timestamp 1607194113
transform 1 0 16164 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_70
timestamp 1607194113
transform 1 0 16072 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_73
timestamp 1607194113
transform 1 0 16992 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_72
timestamp 1607194113
transform 1 0 16900 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_75
timestamp 1607194113
transform 1 0 17820 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_74
timestamp 1607194113
transform 1 0 17728 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_77
timestamp 1607194113
transform 1 0 18648 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_76
timestamp 1607194113
transform 1 0 18556 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_79
timestamp 1607194113
transform 1 0 19476 0 -1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_78
timestamp 1607194113
transform 1 0 19384 0 -1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILL_81 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 20580 0 -1 17792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILL_80 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 20212 0 -1 17792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap31_0
timestamp 1607194113
transform 1 0 2732 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_4
timestamp 1607194113
transform 1 0 1904 0 1 17792
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_4_15
timestamp 1607194113
transform 1 0 3100 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap31_0
timestamp 1607194113
transform 1 0 2824 0 1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_4_14
timestamp 1607194113
transform 1 0 4204 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap31_1
timestamp 1607194113
transform 1 0 3928 0 1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap31_1
timestamp 1607194113
transform 1 0 3836 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_4_13
timestamp 1607194113
transform 1 0 5308 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap31_2
timestamp 1607194113
transform 1 0 5032 0 1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap31_2
timestamp 1607194113
transform 1 0 4940 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_4_12
timestamp 1607194113
transform 1 0 6412 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap31_3
timestamp 1607194113
transform 1 0 6136 0 1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap31_3
timestamp 1607194113
transform 1 0 6044 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap31_4
timestamp 1607194113
transform 1 0 7240 0 1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap31_4
timestamp 1607194113
transform 1 0 7148 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_4_11
timestamp 1607194113
transform 1 0 7516 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_4_10
timestamp 1607194113
transform 1 0 8620 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap31_5
timestamp 1607194113
transform 1 0 8344 0 1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap31_5
timestamp 1607194113
transform 1 0 8252 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_4_9
timestamp 1607194113
transform 1 0 9724 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap31_6
timestamp 1607194113
transform 1 0 9448 0 1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap31_6
timestamp 1607194113
transform 1 0 9356 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_4_8
timestamp 1607194113
transform 1 0 10828 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap31_7
timestamp 1607194113
transform 1 0 10552 0 1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap31_7
timestamp 1607194113
transform 1 0 10460 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap31_8
timestamp 1607194113
transform 1 0 11656 0 1 17792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap31_8
timestamp 1607194113
transform 1 0 11564 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_84
timestamp 1607194113
transform 1 0 12760 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_83
timestamp 1607194113
transform 1 0 12024 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_82
timestamp 1607194113
transform 1 0 11932 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_86
timestamp 1607194113
transform 1 0 13588 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_85
timestamp 1607194113
transform 1 0 12852 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_89
timestamp 1607194113
transform 1 0 14508 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_88
timestamp 1607194113
transform 1 0 14416 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_87
timestamp 1607194113
transform 1 0 13680 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_91
timestamp 1607194113
transform 1 0 15336 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_90
timestamp 1607194113
transform 1 0 15244 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_93
timestamp 1607194113
transform 1 0 16164 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_92
timestamp 1607194113
transform 1 0 16072 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_95
timestamp 1607194113
transform 1 0 16992 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_94
timestamp 1607194113
transform 1 0 16900 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_97
timestamp 1607194113
transform 1 0 17820 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_96
timestamp 1607194113
transform 1 0 17728 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_99
timestamp 1607194113
transform 1 0 18648 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_98
timestamp 1607194113
transform 1 0 18556 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_101
timestamp 1607194113
transform 1 0 19476 0 1 17792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_100
timestamp 1607194113
transform 1 0 19384 0 1 17792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILL_103
timestamp 1607194113
transform 1 0 20580 0 1 17792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILL_102
timestamp 1607194113
transform 1 0 20212 0 1 17792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap32_0
timestamp 1607194113
transform 1 0 2732 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_55
timestamp 1607194113
transform 1 0 1996 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_54
timestamp 1607194113
transform 1 0 1904 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_3_0
timestamp 1607194113
transform 1 0 3100 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap32_0
timestamp 1607194113
transform 1 0 2824 0 -1 18880
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_3_1
timestamp 1607194113
transform 1 0 4204 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap32_1
timestamp 1607194113
transform 1 0 3928 0 -1 18880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap32_1
timestamp 1607194113
transform 1 0 3836 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_3_2
timestamp 1607194113
transform 1 0 5308 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap32_2
timestamp 1607194113
transform 1 0 5032 0 -1 18880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap32_2
timestamp 1607194113
transform 1 0 4940 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_3_3
timestamp 1607194113
transform 1 0 6412 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap32_3
timestamp 1607194113
transform 1 0 6136 0 -1 18880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap32_3
timestamp 1607194113
transform 1 0 6044 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap32_4
timestamp 1607194113
transform 1 0 7240 0 -1 18880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap32_4
timestamp 1607194113
transform 1 0 7148 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_105
timestamp 1607194113
transform 1 0 7608 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_104
timestamp 1607194113
transform 1 0 7516 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_107
timestamp 1607194113
transform 1 0 8436 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_106
timestamp 1607194113
transform 1 0 8344 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_110
timestamp 1607194113
transform 1 0 10000 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_109
timestamp 1607194113
transform 1 0 9264 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_108
timestamp 1607194113
transform 1 0 9172 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_113
timestamp 1607194113
transform 1 0 10920 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_112
timestamp 1607194113
transform 1 0 10828 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_111
timestamp 1607194113
transform 1 0 10092 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_115
timestamp 1607194113
transform 1 0 11748 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_114
timestamp 1607194113
transform 1 0 11656 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_117
timestamp 1607194113
transform 1 0 12576 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_116
timestamp 1607194113
transform 1 0 12484 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_119
timestamp 1607194113
transform 1 0 13404 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_118
timestamp 1607194113
transform 1 0 13312 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_121
timestamp 1607194113
transform 1 0 14232 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_120
timestamp 1607194113
transform 1 0 14140 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_123
timestamp 1607194113
transform 1 0 15060 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_122
timestamp 1607194113
transform 1 0 14968 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_125
timestamp 1607194113
transform 1 0 15888 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_124
timestamp 1607194113
transform 1 0 15796 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_127
timestamp 1607194113
transform 1 0 16716 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_126
timestamp 1607194113
transform 1 0 16624 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_129
timestamp 1607194113
transform 1 0 17544 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_128
timestamp 1607194113
transform 1 0 17452 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_131
timestamp 1607194113
transform 1 0 18372 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_130
timestamp 1607194113
transform 1 0 18280 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_134
timestamp 1607194113
transform 1 0 19936 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_133
timestamp 1607194113
transform 1 0 19200 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_132
timestamp 1607194113
transform 1 0 19108 0 -1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_135
timestamp 1607194113
transform 1 0 20028 0 -1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap34_0
timestamp 1607194113
transform 1 0 2732 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_57
timestamp 1607194113
transform 1 0 1996 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_56
timestamp 1607194113
transform 1 0 1904 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap33_0
timestamp 1607194113
transform 1 0 2732 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_3
timestamp 1607194113
transform 1 0 1904 0 1 18880
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_2_0
timestamp 1607194113
transform 1 0 3100 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap34_0
timestamp 1607194113
transform 1 0 2824 0 -1 19968
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_3_7
timestamp 1607194113
transform 1 0 3100 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap33_0
timestamp 1607194113
transform 1 0 2824 0 1 18880
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_2_1
timestamp 1607194113
transform 1 0 4204 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap34_1
timestamp 1607194113
transform 1 0 3928 0 -1 19968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap34_1
timestamp 1607194113
transform 1 0 3836 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_3_6
timestamp 1607194113
transform 1 0 4204 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap33_1
timestamp 1607194113
transform 1 0 3928 0 1 18880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap33_1
timestamp 1607194113
transform 1 0 3836 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_169
timestamp 1607194113
transform 1 0 5400 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_168
timestamp 1607194113
transform 1 0 5308 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap34_2
timestamp 1607194113
transform 1 0 5032 0 -1 19968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap34_2
timestamp 1607194113
transform 1 0 4940 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_3_5
timestamp 1607194113
transform 1 0 5308 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap33_2
timestamp 1607194113
transform 1 0 5032 0 1 18880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap33_2
timestamp 1607194113
transform 1 0 4940 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_171
timestamp 1607194113
transform 1 0 6228 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_170
timestamp 1607194113
transform 1 0 6136 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_3_4
timestamp 1607194113
transform 1 0 6412 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap33_3
timestamp 1607194113
transform 1 0 6136 0 1 18880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap33_3
timestamp 1607194113
transform 1 0 6044 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_173
timestamp 1607194113
transform 1 0 7056 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_172
timestamp 1607194113
transform 1 0 6964 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap33_4
timestamp 1607194113
transform 1 0 7240 0 1 18880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap33_4
timestamp 1607194113
transform 1 0 7148 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_175
timestamp 1607194113
transform 1 0 7884 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_174
timestamp 1607194113
transform 1 0 7792 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_137
timestamp 1607194113
transform 1 0 7608 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_136
timestamp 1607194113
transform 1 0 7516 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_177
timestamp 1607194113
transform 1 0 8712 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_176
timestamp 1607194113
transform 1 0 8620 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_139
timestamp 1607194113
transform 1 0 8436 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_138
timestamp 1607194113
transform 1 0 8344 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_179
timestamp 1607194113
transform 1 0 9540 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_178
timestamp 1607194113
transform 1 0 9448 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_142
timestamp 1607194113
transform 1 0 10000 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_141
timestamp 1607194113
transform 1 0 9264 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_140
timestamp 1607194113
transform 1 0 9172 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_181
timestamp 1607194113
transform 1 0 10368 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_180
timestamp 1607194113
transform 1 0 10276 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_145
timestamp 1607194113
transform 1 0 10920 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_144
timestamp 1607194113
transform 1 0 10828 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_143
timestamp 1607194113
transform 1 0 10092 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_183
timestamp 1607194113
transform 1 0 11196 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_182
timestamp 1607194113
transform 1 0 11104 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_147
timestamp 1607194113
transform 1 0 11748 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_146
timestamp 1607194113
transform 1 0 11656 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_186
timestamp 1607194113
transform 1 0 12760 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_185
timestamp 1607194113
transform 1 0 12024 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_184
timestamp 1607194113
transform 1 0 11932 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_149
timestamp 1607194113
transform 1 0 12576 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_148
timestamp 1607194113
transform 1 0 12484 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_188
timestamp 1607194113
transform 1 0 13588 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_187
timestamp 1607194113
transform 1 0 12852 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_151
timestamp 1607194113
transform 1 0 13404 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_150
timestamp 1607194113
transform 1 0 13312 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_191
timestamp 1607194113
transform 1 0 14508 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_190
timestamp 1607194113
transform 1 0 14416 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_189
timestamp 1607194113
transform 1 0 13680 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_153
timestamp 1607194113
transform 1 0 14232 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_152
timestamp 1607194113
transform 1 0 14140 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_193
timestamp 1607194113
transform 1 0 15336 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_192
timestamp 1607194113
transform 1 0 15244 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_155
timestamp 1607194113
transform 1 0 15060 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_154
timestamp 1607194113
transform 1 0 14968 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_195
timestamp 1607194113
transform 1 0 16164 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_194
timestamp 1607194113
transform 1 0 16072 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_157
timestamp 1607194113
transform 1 0 15888 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_156
timestamp 1607194113
transform 1 0 15796 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_197
timestamp 1607194113
transform 1 0 16992 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_196
timestamp 1607194113
transform 1 0 16900 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_159
timestamp 1607194113
transform 1 0 16716 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_158
timestamp 1607194113
transform 1 0 16624 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_199
timestamp 1607194113
transform 1 0 17820 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_198
timestamp 1607194113
transform 1 0 17728 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_161
timestamp 1607194113
transform 1 0 17544 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_160
timestamp 1607194113
transform 1 0 17452 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_201
timestamp 1607194113
transform 1 0 18648 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_200
timestamp 1607194113
transform 1 0 18556 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_163
timestamp 1607194113
transform 1 0 18372 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_162
timestamp 1607194113
transform 1 0 18280 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_203
timestamp 1607194113
transform 1 0 19476 0 -1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_202
timestamp 1607194113
transform 1 0 19384 0 -1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_166
timestamp 1607194113
transform 1 0 19936 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_165
timestamp 1607194113
transform 1 0 19200 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_164
timestamp 1607194113
transform 1 0 19108 0 1 18880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILL_205
timestamp 1607194113
transform 1 0 20580 0 -1 19968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILL_204
timestamp 1607194113
transform 1 0 20212 0 -1 19968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_8  FILL_167
timestamp 1607194113
transform 1 0 20028 0 1 18880
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap35_0
timestamp 1607194113
transform 1 0 2732 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_2
timestamp 1607194113
transform 1 0 1904 0 1 19968
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_2_3
timestamp 1607194113
transform 1 0 3100 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap35_0
timestamp 1607194113
transform 1 0 2824 0 1 19968
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_2_2
timestamp 1607194113
transform 1 0 4204 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap35_1
timestamp 1607194113
transform 1 0 3928 0 1 19968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap35_1
timestamp 1607194113
transform 1 0 3836 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_207
timestamp 1607194113
transform 1 0 5400 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_206
timestamp 1607194113
transform 1 0 5308 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap35_2
timestamp 1607194113
transform 1 0 5032 0 1 19968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap35_2
timestamp 1607194113
transform 1 0 4940 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_209
timestamp 1607194113
transform 1 0 6228 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_208
timestamp 1607194113
transform 1 0 6136 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_211
timestamp 1607194113
transform 1 0 7056 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_210
timestamp 1607194113
transform 1 0 6964 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_213
timestamp 1607194113
transform 1 0 7884 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_212
timestamp 1607194113
transform 1 0 7792 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_215
timestamp 1607194113
transform 1 0 8712 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_214
timestamp 1607194113
transform 1 0 8620 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_217
timestamp 1607194113
transform 1 0 9540 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_216
timestamp 1607194113
transform 1 0 9448 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_219
timestamp 1607194113
transform 1 0 10368 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_218
timestamp 1607194113
transform 1 0 10276 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_221
timestamp 1607194113
transform 1 0 11196 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_220
timestamp 1607194113
transform 1 0 11104 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_224
timestamp 1607194113
transform 1 0 12760 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_223
timestamp 1607194113
transform 1 0 12024 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_222
timestamp 1607194113
transform 1 0 11932 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_226
timestamp 1607194113
transform 1 0 13588 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_225
timestamp 1607194113
transform 1 0 12852 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_229
timestamp 1607194113
transform 1 0 14508 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_228
timestamp 1607194113
transform 1 0 14416 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_227
timestamp 1607194113
transform 1 0 13680 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_231
timestamp 1607194113
transform 1 0 15336 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_230
timestamp 1607194113
transform 1 0 15244 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_233
timestamp 1607194113
transform 1 0 16164 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_232
timestamp 1607194113
transform 1 0 16072 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_235
timestamp 1607194113
transform 1 0 16992 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_234
timestamp 1607194113
transform 1 0 16900 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_237
timestamp 1607194113
transform 1 0 17820 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_236
timestamp 1607194113
transform 1 0 17728 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_239
timestamp 1607194113
transform 1 0 18648 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_238
timestamp 1607194113
transform 1 0 18556 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_241
timestamp 1607194113
transform 1 0 19476 0 1 19968
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_240
timestamp 1607194113
transform 1 0 19384 0 1 19968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILL_243
timestamp 1607194113
transform 1 0 20580 0 1 19968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_4  FILL_242
timestamp 1607194113
transform 1 0 20212 0 1 19968
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap36_0
timestamp 1607194113
transform 1 0 2732 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_59
timestamp 1607194113
transform 1 0 1996 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_58
timestamp 1607194113
transform 1 0 1904 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_1_0
timestamp 1607194113
transform 1 0 3100 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap36_0
timestamp 1607194113
transform 1 0 2824 0 -1 21056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_8  FILL_245
timestamp 1607194113
transform 1 0 4296 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_244
timestamp 1607194113
transform 1 0 4204 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap36_1
timestamp 1607194113
transform 1 0 3928 0 -1 21056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap36_1
timestamp 1607194113
transform 1 0 3836 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_247
timestamp 1607194113
transform 1 0 5124 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_246
timestamp 1607194113
transform 1 0 5032 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_249
timestamp 1607194113
transform 1 0 5952 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_248
timestamp 1607194113
transform 1 0 5860 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_251
timestamp 1607194113
transform 1 0 6780 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_250
timestamp 1607194113
transform 1 0 6688 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_253
timestamp 1607194113
transform 1 0 7608 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_252
timestamp 1607194113
transform 1 0 7516 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_255
timestamp 1607194113
transform 1 0 8436 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_254
timestamp 1607194113
transform 1 0 8344 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_258
timestamp 1607194113
transform 1 0 10000 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_257
timestamp 1607194113
transform 1 0 9264 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_256
timestamp 1607194113
transform 1 0 9172 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_261
timestamp 1607194113
transform 1 0 10920 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_260
timestamp 1607194113
transform 1 0 10828 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_259
timestamp 1607194113
transform 1 0 10092 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_263
timestamp 1607194113
transform 1 0 11748 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_262
timestamp 1607194113
transform 1 0 11656 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_265
timestamp 1607194113
transform 1 0 12576 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_264
timestamp 1607194113
transform 1 0 12484 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_267
timestamp 1607194113
transform 1 0 13404 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_266
timestamp 1607194113
transform 1 0 13312 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_269
timestamp 1607194113
transform 1 0 14232 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_268
timestamp 1607194113
transform 1 0 14140 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_271
timestamp 1607194113
transform 1 0 15060 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_270
timestamp 1607194113
transform 1 0 14968 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_273
timestamp 1607194113
transform 1 0 15888 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_272
timestamp 1607194113
transform 1 0 15796 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_275
timestamp 1607194113
transform 1 0 16716 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_274
timestamp 1607194113
transform 1 0 16624 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_277
timestamp 1607194113
transform 1 0 17544 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_276
timestamp 1607194113
transform 1 0 17452 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_279
timestamp 1607194113
transform 1 0 18372 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_278
timestamp 1607194113
transform 1 0 18280 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_282
timestamp 1607194113
transform 1 0 19936 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_281
timestamp 1607194113
transform 1 0 19200 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_280
timestamp 1607194113
transform 1 0 19108 0 -1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_283
timestamp 1607194113
transform 1 0 20028 0 -1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap37_0
timestamp 1607194113
transform 1 0 2732 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_1
timestamp 1607194113
transform 1 0 1904 0 1 21056
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_1_1
timestamp 1607194113
transform 1 0 3100 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap37_0
timestamp 1607194113
transform 1 0 2824 0 1 21056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_8  FILL_285
timestamp 1607194113
transform 1 0 4296 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_284
timestamp 1607194113
transform 1 0 4204 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap37_1
timestamp 1607194113
transform 1 0 3928 0 1 21056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap37_1
timestamp 1607194113
transform 1 0 3836 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_287
timestamp 1607194113
transform 1 0 5124 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_286
timestamp 1607194113
transform 1 0 5032 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_289
timestamp 1607194113
transform 1 0 5952 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_288
timestamp 1607194113
transform 1 0 5860 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_291
timestamp 1607194113
transform 1 0 6780 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_290
timestamp 1607194113
transform 1 0 6688 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_293
timestamp 1607194113
transform 1 0 7608 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_292
timestamp 1607194113
transform 1 0 7516 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_295
timestamp 1607194113
transform 1 0 8436 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_294
timestamp 1607194113
transform 1 0 8344 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_298
timestamp 1607194113
transform 1 0 10000 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_297
timestamp 1607194113
transform 1 0 9264 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_296
timestamp 1607194113
transform 1 0 9172 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_301
timestamp 1607194113
transform 1 0 10920 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_300
timestamp 1607194113
transform 1 0 10828 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_299
timestamp 1607194113
transform 1 0 10092 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_303
timestamp 1607194113
transform 1 0 11748 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_302
timestamp 1607194113
transform 1 0 11656 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_305
timestamp 1607194113
transform 1 0 12576 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_304
timestamp 1607194113
transform 1 0 12484 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_307
timestamp 1607194113
transform 1 0 13404 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_306
timestamp 1607194113
transform 1 0 13312 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_309
timestamp 1607194113
transform 1 0 14232 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_308
timestamp 1607194113
transform 1 0 14140 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_311
timestamp 1607194113
transform 1 0 15060 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_310
timestamp 1607194113
transform 1 0 14968 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_313
timestamp 1607194113
transform 1 0 15888 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_312
timestamp 1607194113
transform 1 0 15796 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_315
timestamp 1607194113
transform 1 0 16716 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_314
timestamp 1607194113
transform 1 0 16624 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_317
timestamp 1607194113
transform 1 0 17544 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_316
timestamp 1607194113
transform 1 0 17452 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_319
timestamp 1607194113
transform 1 0 18372 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_318
timestamp 1607194113
transform 1 0 18280 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_322
timestamp 1607194113
transform 1 0 19936 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_321
timestamp 1607194113
transform 1 0 19200 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_320
timestamp 1607194113
transform 1 0 19108 0 1 21056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_323
timestamp 1607194113
transform 1 0 20028 0 1 21056
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap38_0
timestamp 1607194113
transform 1 0 2732 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  mux_0
timestamp 1607194113
transform 1 0 1904 0 -1 22144
box -38 -48 866 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  delay_0_0
timestamp 1607194113
transform 1 0 3100 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  decap38_0
timestamp 1607194113
transform 1 0 2824 0 -1 22144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_8  FILL_325
timestamp 1607194113
transform 1 0 4296 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_324
timestamp 1607194113
transform 1 0 4204 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap38_1
timestamp 1607194113
transform 1 0 3928 0 -1 22144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap38_1
timestamp 1607194113
transform 1 0 3836 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_327
timestamp 1607194113
transform 1 0 5124 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_326
timestamp 1607194113
transform 1 0 5032 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_329
timestamp 1607194113
transform 1 0 5952 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_328
timestamp 1607194113
transform 1 0 5860 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_331
timestamp 1607194113
transform 1 0 6780 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_330
timestamp 1607194113
transform 1 0 6688 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_333
timestamp 1607194113
transform 1 0 7608 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_332
timestamp 1607194113
transform 1 0 7516 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_335
timestamp 1607194113
transform 1 0 8436 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_334
timestamp 1607194113
transform 1 0 8344 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_338
timestamp 1607194113
transform 1 0 10000 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_337
timestamp 1607194113
transform 1 0 9264 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_336
timestamp 1607194113
transform 1 0 9172 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_341
timestamp 1607194113
transform 1 0 10920 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_340
timestamp 1607194113
transform 1 0 10828 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_339
timestamp 1607194113
transform 1 0 10092 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_8  FILL_343
timestamp 1607194113
transform 1 0 11748 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_342
timestamp 1607194113
transform 1 0 11656 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_345
timestamp 1607194113
transform 1 0 12576 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_344
timestamp 1607194113
transform 1 0 12484 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_347
timestamp 1607194113
transform 1 0 13404 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_346
timestamp 1607194113
transform 1 0 13312 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_349
timestamp 1607194113
transform 1 0 14232 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_348
timestamp 1607194113
transform 1 0 14140 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_351
timestamp 1607194113
transform 1 0 15060 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_350
timestamp 1607194113
transform 1 0 14968 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_353
timestamp 1607194113
transform 1 0 15888 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_352
timestamp 1607194113
transform 1 0 15796 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_355
timestamp 1607194113
transform 1 0 16716 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_354
timestamp 1607194113
transform 1 0 16624 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_357
timestamp 1607194113
transform 1 0 17544 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_356
timestamp 1607194113
transform 1 0 17452 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_359
timestamp 1607194113
transform 1 0 18372 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_358
timestamp 1607194113
transform 1 0 18280 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_362
timestamp 1607194113
transform 1 0 19936 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_361
timestamp 1607194113
transform 1 0 19200 0 -1 22144
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_360
timestamp 1607194113
transform 1 0 19108 0 -1 22144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_363
timestamp 1607194113
transform 1 0 20028 0 -1 22144
box -38 -48 774 592
<< labels >>
rlabel metal3 s 800 800 920 920 6 inp_i
port 0 nsew default input
rlabel metal3 s 800 22016 920 22136 6 out_o
port 1 nsew default tristate
rlabel metal3 s 800 8960 920 9080 6 en_i[8]
port 2 nsew default input
rlabel metal3 s 800 13312 920 13432 6 en_i[7]
port 3 nsew default input
rlabel metal3 s 800 15488 920 15608 6 en_i[6]
port 4 nsew default input
rlabel metal3 s 800 16576 920 16696 6 en_i[5]
port 5 nsew default input
rlabel metal3 s 800 17664 920 17784 6 en_i[4]
port 6 nsew default input
rlabel metal3 s 800 18752 920 18872 6 en_i[3]
port 7 nsew default input
rlabel metal3 s 800 19840 920 19960 6 en_i[2]
port 8 nsew default input
rlabel metal3 s 800 20928 920 21048 6 en_i[1]
port 9 nsew default input
rlabel metal3 s 800 21472 920 21592 6 en_i[0]
port 10 nsew default input
rlabel metal5 s 1904 2560 20764 2880 6 VPWR
port 11 nsew default input
rlabel metal5 s 1904 20560 20764 20880 6 VGND
port 12 nsew default input
<< properties >>
string FIXED_BBOX 0 0 21602 23185
<< end >>
