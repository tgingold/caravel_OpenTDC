magic
tech sky130A
magscale 1 2
timestamp 1607276512
<< locali >>
rect 34713 42551 34747 42653
rect 56885 42551 56919 42653
rect 60013 41463 60047 41565
rect 63233 41463 63267 41633
rect 52469 40987 52503 41225
rect 17785 39831 17819 40001
rect 19717 39491 19751 39593
rect 31953 39423 31987 39593
rect 43729 39491 43763 39593
rect 48329 39423 48363 39525
rect 62037 39287 62071 39457
rect 20269 38199 20303 38437
rect 31953 38403 31987 38505
rect 71237 38267 71271 38369
rect 84669 38267 84703 38505
rect 57345 37655 57379 37757
rect 68569 37655 68603 37757
rect 22937 37179 22971 37281
rect 34713 36567 34747 36737
rect 39129 36703 39163 36873
rect 57161 36703 57195 36805
rect 72893 36091 72927 36329
rect 76113 35547 76147 35717
rect 79609 35547 79643 35785
rect 65809 35139 65843 35241
rect 31493 34935 31527 35105
rect 37749 34935 37783 35037
rect 23489 34391 23523 34629
rect 26157 34391 26191 34561
rect 37289 34459 37323 34697
rect 56701 34391 56735 34561
rect 24777 34085 25087 34119
rect 24777 34051 24811 34085
rect 24869 33303 24903 34017
rect 25053 33915 25087 34085
rect 37289 33711 37323 34153
rect 46857 33711 46891 34153
rect 5089 32759 5123 32929
rect 24685 32283 24719 32385
rect 24777 32351 24811 32997
rect 24685 32249 24961 32283
rect 25053 31875 25087 32793
rect 15393 31671 15427 31773
rect 25145 31671 25179 32861
rect 19717 31127 19751 31229
rect 24777 30311 24811 31297
rect 25973 30719 26007 32317
rect 26893 31875 26927 32453
rect 37289 32419 37323 32657
rect 46857 32419 46891 32657
rect 41429 31127 41463 31161
rect 41371 31093 41463 31127
rect 20177 27999 20211 28101
rect 7941 21335 7975 21505
rect 54125 19363 54159 28373
rect 16129 18275 16163 18377
rect 24777 18003 24811 18581
rect 7665 14807 7699 14909
rect 18337 14399 18371 14569
rect 7941 13855 7975 14025
rect 18613 8415 18647 8585
<< viali >>
rect 15945 43809 15979 43843
rect 16497 43809 16531 43843
rect 16681 43809 16715 43843
rect 28273 43809 28307 43843
rect 44649 43809 44683 43843
rect 45109 43809 45143 43843
rect 45201 43809 45235 43843
rect 53665 43809 53699 43843
rect 58541 43809 58575 43843
rect 59553 43809 59587 43843
rect 59737 43809 59771 43843
rect 73813 43809 73847 43843
rect 78505 43809 78539 43843
rect 78781 43809 78815 43843
rect 79333 43809 79367 43843
rect 79793 43809 79827 43843
rect 82277 43809 82311 43843
rect 82369 43809 82403 43843
rect 15669 43741 15703 43775
rect 15761 43741 15795 43775
rect 44281 43741 44315 43775
rect 44465 43741 44499 43775
rect 60105 43741 60139 43775
rect 82829 43741 82863 43775
rect 28365 43673 28399 43707
rect 73905 43673 73939 43707
rect 78873 43673 78907 43707
rect 16957 43605 16991 43639
rect 17325 43605 17359 43639
rect 44189 43605 44223 43639
rect 45661 43605 45695 43639
rect 45937 43605 45971 43639
rect 53849 43605 53883 43639
rect 58633 43605 58667 43639
rect 74089 43605 74123 43639
rect 78689 43605 78723 43639
rect 82093 43605 82127 43639
rect 36829 43401 36863 43435
rect 37013 43401 37047 43435
rect 48329 43401 48363 43435
rect 48421 43401 48455 43435
rect 50169 43401 50203 43435
rect 54585 43401 54619 43435
rect 55045 43401 55079 43435
rect 58725 43401 58759 43435
rect 74641 43401 74675 43435
rect 75561 43401 75595 43435
rect 2421 43265 2455 43299
rect 2789 43265 2823 43299
rect 7573 43265 7607 43299
rect 9321 43265 9355 43299
rect 26985 43265 27019 43299
rect 37197 43265 37231 43299
rect 38485 43265 38519 43299
rect 41337 43265 41371 43299
rect 48605 43265 48639 43299
rect 53481 43265 53515 43299
rect 58817 43265 58851 43299
rect 59093 43265 59127 43299
rect 70317 43265 70351 43299
rect 72065 43265 72099 43299
rect 78413 43265 78447 43299
rect 82369 43265 82403 43299
rect 2513 43197 2547 43231
rect 7849 43197 7883 43231
rect 12449 43197 12483 43231
rect 15485 43197 15519 43231
rect 15761 43197 15795 43231
rect 17141 43197 17175 43231
rect 18061 43197 18095 43231
rect 20453 43197 20487 43231
rect 20637 43197 20671 43231
rect 21189 43197 21223 43231
rect 21373 43197 21407 43231
rect 26709 43197 26743 43231
rect 32597 43197 32631 43231
rect 32781 43197 32815 43231
rect 33241 43197 33275 43231
rect 33333 43197 33367 43231
rect 37381 43197 37415 43231
rect 37841 43197 37875 43231
rect 37933 43197 37967 43231
rect 41061 43197 41095 43231
rect 48789 43197 48823 43231
rect 49249 43197 49283 43231
rect 49341 43197 49375 43231
rect 52193 43197 52227 43231
rect 53205 43197 53239 43231
rect 63693 43197 63727 43231
rect 66913 43197 66947 43231
rect 67189 43197 67223 43231
rect 67373 43197 67407 43231
rect 70593 43197 70627 43231
rect 74181 43197 74215 43231
rect 74457 43197 74491 43231
rect 75745 43197 75779 43231
rect 78689 43197 78723 43231
rect 78873 43197 78907 43231
rect 78965 43197 78999 43231
rect 82001 43197 82035 43231
rect 82553 43197 82587 43231
rect 83565 43197 83599 43231
rect 28365 43129 28399 43163
rect 33885 43129 33919 43163
rect 66361 43129 66395 43163
rect 74365 43129 74399 43163
rect 77861 43129 77895 43163
rect 83657 43129 83691 43163
rect 3893 43061 3927 43095
rect 4353 43061 4387 43095
rect 8953 43061 8987 43095
rect 12541 43061 12575 43095
rect 17233 43061 17267 43095
rect 18153 43061 18187 43095
rect 20269 43061 20303 43095
rect 21649 43061 21683 43095
rect 22017 43061 22051 43095
rect 28457 43061 28491 43095
rect 32045 43061 32079 43095
rect 32229 43061 32263 43095
rect 32413 43061 32447 43095
rect 34161 43061 34195 43095
rect 38761 43061 38795 43095
rect 38853 43061 38887 43095
rect 40969 43061 41003 43095
rect 42625 43061 42659 43095
rect 49801 43061 49835 43095
rect 52285 43061 52319 43095
rect 60197 43061 60231 43095
rect 63785 43061 63819 43095
rect 71881 43061 71915 43095
rect 75929 43061 75963 43095
rect 83841 43061 83875 43095
rect 12357 42857 12391 42891
rect 28273 42857 28307 42891
rect 29285 42857 29319 42891
rect 34253 42857 34287 42891
rect 68477 42857 68511 42891
rect 81449 42857 81483 42891
rect 23949 42789 23983 42823
rect 1961 42721 1995 42755
rect 2513 42721 2547 42755
rect 2697 42721 2731 42755
rect 4169 42721 4203 42755
rect 7573 42721 7607 42755
rect 8125 42721 8159 42755
rect 8309 42721 8343 42755
rect 9689 42721 9723 42755
rect 12541 42721 12575 42755
rect 16773 42721 16807 42755
rect 17049 42721 17083 42755
rect 24409 42721 24443 42755
rect 24961 42721 24995 42755
rect 25145 42721 25179 42755
rect 26985 42721 27019 42755
rect 29193 42721 29227 42755
rect 32229 42721 32263 42755
rect 32413 42721 32447 42755
rect 32873 42721 32907 42755
rect 33425 42721 33459 42755
rect 33609 42721 33643 42755
rect 35265 42721 35299 42755
rect 38301 42721 38335 42755
rect 45017 42721 45051 42755
rect 45477 42721 45511 42755
rect 45569 42721 45603 42755
rect 46397 42721 46431 42755
rect 46581 42721 46615 42755
rect 50905 42721 50939 42755
rect 50997 42721 51031 42755
rect 53481 42721 53515 42755
rect 54585 42721 54619 42755
rect 54769 42721 54803 42755
rect 55229 42721 55263 42755
rect 56977 42721 57011 42755
rect 57161 42721 57195 42755
rect 57345 42721 57379 42755
rect 58541 42721 58575 42755
rect 58817 42721 58851 42755
rect 60381 42721 60415 42755
rect 60473 42721 60507 42755
rect 61761 42721 61795 42755
rect 63417 42721 63451 42755
rect 66177 42721 66211 42755
rect 68569 42721 68603 42755
rect 68937 42721 68971 42755
rect 69213 42721 69247 42755
rect 71605 42721 71639 42755
rect 71973 42721 72007 42755
rect 73905 42721 73939 42755
rect 74089 42721 74123 42755
rect 74365 42721 74399 42755
rect 77033 42721 77067 42755
rect 77309 42721 77343 42755
rect 81173 42721 81207 42755
rect 81357 42721 81391 42755
rect 83013 42721 83047 42755
rect 1869 42653 1903 42687
rect 7389 42653 7423 42687
rect 9781 42653 9815 42687
rect 10793 42653 10827 42687
rect 11069 42653 11103 42687
rect 18521 42653 18555 42687
rect 21281 42653 21315 42687
rect 21557 42653 21591 42687
rect 24225 42653 24259 42687
rect 25513 42653 25547 42687
rect 25789 42653 25823 42687
rect 26709 42653 26743 42687
rect 32505 42653 32539 42687
rect 32689 42653 32723 42687
rect 33977 42653 34011 42687
rect 34713 42653 34747 42687
rect 34989 42653 35023 42687
rect 37841 42653 37875 42687
rect 38032 42653 38066 42687
rect 44465 42653 44499 42687
rect 44649 42653 44683 42687
rect 44833 42653 44867 42687
rect 46029 42653 46063 42687
rect 51273 42653 51307 42687
rect 53573 42653 53607 42687
rect 56885 42653 56919 42687
rect 57713 42653 57747 42687
rect 59001 42653 59035 42687
rect 60933 42653 60967 42687
rect 63049 42653 63083 42687
rect 63141 42653 63175 42687
rect 65901 42653 65935 42687
rect 72433 42653 72467 42687
rect 78597 42653 78631 42687
rect 78873 42653 78907 42687
rect 82461 42653 82495 42687
rect 82737 42653 82771 42687
rect 36553 42585 36587 42619
rect 58633 42585 58667 42619
rect 61853 42585 61887 42619
rect 71513 42585 71547 42619
rect 77125 42585 77159 42619
rect 1685 42517 1719 42551
rect 2973 42517 3007 42551
rect 3341 42517 3375 42551
rect 4261 42517 4295 42551
rect 7205 42517 7239 42551
rect 8585 42517 8619 42551
rect 10057 42517 10091 42551
rect 18337 42517 18371 42551
rect 22661 42517 22695 42551
rect 23121 42517 23155 42551
rect 24041 42517 24075 42551
rect 28457 42517 28491 42551
rect 34713 42517 34747 42551
rect 34805 42517 34839 42551
rect 39589 42517 39623 42551
rect 52377 42517 52411 42551
rect 54861 42517 54895 42551
rect 56885 42517 56919 42551
rect 60197 42517 60231 42551
rect 61025 42517 61059 42551
rect 64521 42517 64555 42551
rect 65533 42517 65567 42551
rect 67281 42517 67315 42551
rect 69581 42517 69615 42551
rect 71237 42517 71271 42551
rect 72709 42517 72743 42551
rect 75469 42517 75503 42551
rect 78413 42517 78447 42551
rect 79977 42517 80011 42551
rect 84301 42517 84335 42551
rect 4169 42313 4203 42347
rect 38761 42313 38795 42347
rect 38945 42313 38979 42347
rect 39497 42313 39531 42347
rect 41981 42313 42015 42347
rect 53757 42313 53791 42347
rect 81081 42313 81115 42347
rect 16681 42245 16715 42279
rect 36829 42245 36863 42279
rect 37013 42245 37047 42279
rect 59093 42245 59127 42279
rect 66729 42245 66763 42279
rect 77861 42245 77895 42279
rect 3065 42177 3099 42211
rect 8585 42177 8619 42211
rect 8861 42177 8895 42211
rect 10241 42177 10275 42211
rect 15485 42177 15519 42211
rect 15669 42177 15703 42211
rect 17141 42177 17175 42211
rect 18429 42177 18463 42211
rect 27169 42177 27203 42211
rect 32137 42177 32171 42211
rect 32229 42177 32263 42211
rect 32597 42177 32631 42211
rect 37197 42177 37231 42211
rect 38485 42177 38519 42211
rect 42073 42177 42107 42211
rect 63877 42177 63911 42211
rect 70593 42177 70627 42211
rect 71145 42177 71179 42211
rect 73261 42177 73295 42211
rect 74549 42177 74583 42211
rect 2789 42109 2823 42143
rect 10333 42109 10367 42143
rect 11069 42109 11103 42143
rect 15761 42109 15795 42143
rect 16221 42109 16255 42143
rect 16313 42109 16347 42143
rect 18337 42109 18371 42143
rect 20085 42109 20119 42143
rect 20269 42109 20303 42143
rect 20821 42109 20855 42143
rect 21005 42109 21039 42143
rect 22569 42109 22603 42143
rect 25789 42109 25823 42143
rect 25973 42109 26007 42143
rect 26157 42109 26191 42143
rect 26617 42109 26651 42143
rect 26709 42109 26743 42143
rect 32781 42109 32815 42143
rect 33333 42109 33367 42143
rect 33517 42109 33551 42143
rect 34345 42109 34379 42143
rect 37381 42109 37415 42143
rect 37841 42109 37875 42143
rect 37933 42109 37967 42143
rect 39405 42109 39439 42143
rect 40509 42109 40543 42143
rect 42349 42109 42383 42143
rect 43729 42109 43763 42143
rect 44557 42109 44591 42143
rect 47593 42109 47627 42143
rect 47961 42109 47995 42143
rect 48145 42109 48179 42143
rect 48605 42109 48639 42143
rect 48697 42109 48731 42143
rect 49617 42109 49651 42143
rect 51733 42109 51767 42143
rect 54309 42109 54343 42143
rect 54401 42109 54435 42143
rect 54677 42109 54711 42143
rect 54861 42109 54895 42143
rect 55689 42109 55723 42143
rect 59645 42109 59679 42143
rect 59737 42109 59771 42143
rect 60013 42109 60047 42143
rect 60197 42109 60231 42143
rect 61025 42109 61059 42143
rect 61209 42109 61243 42143
rect 64521 42109 64555 42143
rect 64613 42109 64647 42143
rect 64889 42109 64923 42143
rect 65073 42109 65107 42143
rect 66637 42109 66671 42143
rect 66913 42109 66947 42143
rect 69489 42109 69523 42143
rect 71283 42109 71317 42143
rect 71421 42109 71455 42143
rect 72893 42109 72927 42143
rect 74181 42109 74215 42143
rect 74733 42109 74767 42143
rect 76573 42109 76607 42143
rect 77677 42109 77711 42143
rect 79885 42109 79919 42143
rect 80903 42109 80937 42143
rect 82829 42109 82863 42143
rect 83105 42109 83139 42143
rect 33885 42041 33919 42075
rect 49249 42041 49283 42075
rect 54953 42041 54987 42075
rect 60289 42041 60323 42075
rect 69857 42041 69891 42075
rect 72709 42041 72743 42075
rect 4629 41973 4663 42007
rect 11253 41973 11287 42007
rect 11437 41973 11471 42007
rect 19993 41973 20027 42007
rect 21281 41973 21315 42007
rect 21649 41973 21683 42007
rect 22661 41973 22695 42007
rect 25697 41973 25731 42007
rect 27537 41973 27571 42007
rect 32413 41973 32447 42007
rect 34161 41973 34195 42007
rect 40601 41973 40635 42007
rect 44649 41973 44683 42007
rect 47869 41973 47903 42007
rect 49525 41973 49559 42007
rect 51825 41973 51859 42007
rect 53481 41973 53515 42007
rect 55781 41973 55815 42007
rect 61301 41973 61335 42007
rect 65257 41973 65291 42007
rect 69673 41973 69707 42007
rect 70409 41973 70443 42007
rect 76757 41973 76791 42007
rect 79977 41973 80011 42007
rect 82737 41973 82771 42007
rect 84209 41973 84243 42007
rect 8033 41769 8067 41803
rect 11529 41769 11563 41803
rect 11897 41769 11931 41803
rect 16773 41769 16807 41803
rect 16957 41769 16991 41803
rect 26617 41769 26651 41803
rect 27905 41769 27939 41803
rect 28089 41769 28123 41803
rect 35541 41769 35575 41803
rect 39405 41769 39439 41803
rect 39589 41769 39623 41803
rect 43729 41769 43763 41803
rect 45477 41769 45511 41803
rect 48513 41769 48547 41803
rect 74733 41769 74767 41803
rect 25789 41701 25823 41735
rect 37473 41701 37507 41735
rect 46121 41701 46155 41735
rect 50537 41701 50571 41735
rect 71881 41701 71915 41735
rect 72709 41701 72743 41735
rect 72893 41701 72927 41735
rect 81725 41701 81759 41735
rect 82829 41701 82863 41735
rect 7021 41633 7055 41667
rect 7481 41633 7515 41667
rect 7573 41633 7607 41667
rect 10517 41633 10551 41667
rect 10977 41633 11011 41667
rect 11069 41633 11103 41667
rect 14197 41633 14231 41667
rect 16037 41633 16071 41667
rect 16405 41633 16439 41667
rect 16589 41633 16623 41667
rect 21189 41633 21223 41667
rect 25053 41633 25087 41667
rect 25421 41633 25455 41667
rect 25605 41633 25639 41667
rect 27169 41633 27203 41667
rect 27537 41633 27571 41667
rect 27721 41633 27755 41667
rect 30941 41633 30975 41667
rect 32321 41633 32355 41667
rect 32781 41633 32815 41667
rect 32873 41633 32907 41667
rect 33977 41633 34011 41667
rect 34161 41633 34195 41667
rect 34345 41633 34379 41667
rect 34529 41633 34563 41667
rect 35081 41633 35115 41667
rect 35265 41633 35299 41667
rect 38025 41633 38059 41667
rect 38485 41633 38519 41667
rect 38577 41633 38611 41667
rect 42257 41633 42291 41667
rect 43913 41633 43947 41667
rect 44097 41633 44131 41667
rect 44557 41633 44591 41667
rect 44649 41633 44683 41667
rect 45569 41633 45603 41667
rect 49157 41633 49191 41667
rect 49709 41633 49743 41667
rect 49893 41633 49927 41667
rect 53113 41633 53147 41667
rect 53297 41633 53331 41667
rect 55045 41633 55079 41667
rect 55149 41633 55183 41667
rect 55249 41633 55283 41667
rect 55781 41633 55815 41667
rect 58725 41633 58759 41667
rect 58909 41633 58943 41667
rect 59001 41633 59035 41667
rect 60197 41633 60231 41667
rect 60473 41633 60507 41667
rect 63233 41633 63267 41667
rect 63325 41633 63359 41667
rect 64337 41633 64371 41667
rect 64521 41633 64555 41667
rect 65809 41633 65843 41667
rect 71789 41633 71823 41667
rect 73040 41633 73074 41667
rect 74457 41633 74491 41667
rect 74641 41633 74675 41667
rect 77953 41633 77987 41667
rect 78413 41633 78447 41667
rect 81173 41633 81207 41667
rect 81357 41633 81391 41667
rect 82645 41633 82679 41667
rect 82921 41633 82955 41667
rect 84209 41633 84243 41667
rect 6929 41565 6963 41599
rect 10241 41565 10275 41599
rect 10333 41565 10367 41599
rect 15393 41565 15427 41599
rect 16129 41565 16163 41599
rect 20913 41565 20947 41599
rect 24409 41565 24443 41599
rect 25145 41565 25179 41599
rect 25973 41565 26007 41599
rect 27261 41565 27295 41599
rect 31861 41565 31895 41599
rect 32137 41565 32171 41599
rect 37933 41565 37967 41599
rect 39037 41565 39071 41599
rect 42349 41565 42383 41599
rect 45201 41565 45235 41599
rect 46489 41565 46523 41599
rect 48697 41565 48731 41599
rect 48973 41565 49007 41599
rect 53665 41565 53699 41599
rect 60013 41565 60047 41599
rect 60289 41565 60323 41599
rect 24225 41497 24259 41531
rect 26249 41497 26283 41531
rect 30757 41497 30791 41531
rect 33241 41497 33275 41531
rect 33701 41497 33735 41531
rect 35909 41497 35943 41531
rect 6653 41429 6687 41463
rect 14289 41429 14323 41463
rect 17141 41429 17175 41463
rect 22293 41429 22327 41463
rect 22753 41429 22787 41463
rect 31585 41429 31619 41463
rect 33885 41429 33919 41463
rect 43545 41429 43579 41463
rect 46259 41429 46293 41463
rect 46397 41429 46431 41463
rect 46581 41429 46615 41463
rect 50169 41429 50203 41463
rect 55413 41429 55447 41463
rect 60013 41429 60047 41463
rect 63417 41565 63451 41599
rect 65533 41565 65567 41599
rect 66177 41565 66211 41599
rect 66361 41565 66395 41599
rect 73261 41565 73295 41599
rect 84301 41565 84335 41599
rect 78137 41497 78171 41531
rect 63233 41429 63267 41463
rect 63601 41429 63635 41463
rect 64613 41429 64647 41463
rect 65947 41429 65981 41463
rect 66085 41429 66119 41463
rect 73169 41429 73203 41463
rect 73537 41429 73571 41463
rect 83105 41429 83139 41463
rect 4629 41225 4663 41259
rect 8769 41225 8803 41259
rect 45017 41225 45051 41259
rect 49893 41225 49927 41259
rect 52469 41225 52503 41259
rect 52745 41225 52779 41259
rect 63785 41225 63819 41259
rect 80253 41225 80287 41259
rect 80897 41225 80931 41259
rect 87153 41225 87187 41259
rect 14105 41157 14139 41191
rect 25329 41157 25363 41191
rect 26157 41157 26191 41191
rect 33977 41157 34011 41191
rect 47961 41157 47995 41191
rect 50077 41157 50111 41191
rect 2789 41089 2823 41123
rect 26801 41089 26835 41123
rect 38301 41089 38335 41123
rect 43913 41089 43947 41123
rect 45293 41089 45327 41123
rect 48421 41089 48455 41123
rect 3065 41021 3099 41055
rect 8401 41021 8435 41055
rect 12725 41021 12759 41055
rect 13001 41021 13035 41055
rect 15209 41021 15243 41055
rect 19717 41021 19751 41055
rect 19993 41021 20027 41055
rect 22293 41021 22327 41055
rect 25145 41021 25179 41055
rect 26893 41021 26927 41055
rect 27261 41021 27295 41055
rect 27445 41021 27479 41055
rect 31585 41021 31619 41055
rect 31769 41021 31803 41055
rect 31953 41021 31987 41055
rect 32413 41021 32447 41055
rect 32505 41021 32539 41055
rect 34161 41021 34195 41055
rect 37013 41021 37047 41055
rect 37197 41021 37231 41055
rect 37657 41021 37691 41055
rect 37749 41021 37783 41055
rect 38485 41021 38519 41055
rect 44005 41021 44039 41055
rect 44465 41021 44499 41055
rect 44557 41021 44591 41055
rect 48513 41021 48547 41055
rect 48973 41021 49007 41055
rect 49065 41021 49099 41055
rect 74457 41157 74491 41191
rect 80786 41157 80820 41191
rect 65165 41089 65199 41123
rect 80989 41089 81023 41123
rect 87337 41089 87371 41123
rect 52653 41021 52687 41055
rect 54769 41021 54803 41055
rect 55045 41021 55079 41055
rect 63693 41021 63727 41055
rect 64889 41021 64923 41055
rect 66269 41021 66303 41055
rect 71697 41021 71731 41055
rect 71789 41021 71823 41055
rect 72893 41021 72927 41055
rect 74365 41021 74399 41055
rect 74641 41021 74675 41055
rect 78413 41021 78447 41055
rect 80621 41021 80655 41055
rect 82645 41021 82679 41055
rect 87613 41021 87647 41055
rect 4445 40953 4479 40987
rect 21373 40953 21407 40987
rect 36829 40953 36863 40987
rect 48145 40953 48179 40987
rect 52469 40953 52503 40987
rect 64705 40953 64739 40987
rect 66085 40953 66119 40987
rect 72709 40953 72743 40987
rect 75193 40953 75227 40987
rect 81357 40953 81391 40987
rect 8493 40885 8527 40919
rect 14473 40885 14507 40919
rect 15393 40885 15427 40919
rect 21465 40885 21499 40919
rect 22385 40885 22419 40919
rect 24961 40885 24995 40919
rect 26341 40885 26375 40919
rect 27629 40885 27663 40919
rect 27813 40885 27847 40919
rect 31401 40885 31435 40919
rect 32965 40885 32999 40919
rect 33333 40885 33367 40919
rect 33517 40885 33551 40919
rect 38761 40885 38795 40919
rect 49525 40885 49559 40919
rect 54585 40885 54619 40919
rect 56149 40885 56183 40919
rect 66361 40885 66395 40919
rect 72065 40885 72099 40919
rect 72985 40885 73019 40919
rect 74825 40885 74859 40919
rect 78597 40885 78631 40919
rect 80529 40885 80563 40919
rect 82829 40885 82863 40919
rect 88717 40885 88751 40919
rect 4169 40681 4203 40715
rect 12541 40681 12575 40715
rect 16681 40681 16715 40715
rect 20729 40681 20763 40715
rect 31953 40681 31987 40715
rect 43177 40681 43211 40715
rect 45109 40681 45143 40715
rect 82921 40681 82955 40715
rect 88993 40681 89027 40715
rect 33701 40613 33735 40647
rect 37565 40613 37599 40647
rect 44649 40613 44683 40647
rect 49433 40613 49467 40647
rect 54677 40613 54711 40647
rect 81357 40613 81391 40647
rect 85681 40613 85715 40647
rect 4353 40545 4387 40579
rect 4629 40545 4663 40579
rect 5641 40545 5675 40579
rect 7573 40545 7607 40579
rect 7757 40545 7791 40579
rect 8125 40545 8159 40579
rect 11529 40545 11563 40579
rect 12081 40545 12115 40579
rect 12265 40545 12299 40579
rect 13553 40545 13587 40579
rect 16405 40545 16439 40579
rect 16497 40545 16531 40579
rect 21557 40545 21591 40579
rect 21925 40545 21959 40579
rect 22109 40545 22143 40579
rect 22477 40545 22511 40579
rect 30481 40545 30515 40579
rect 32137 40545 32171 40579
rect 32321 40545 32355 40579
rect 32781 40545 32815 40579
rect 32873 40545 32907 40579
rect 37933 40545 37967 40579
rect 38393 40545 38427 40579
rect 38485 40545 38519 40579
rect 39405 40545 39439 40579
rect 43545 40545 43579 40579
rect 44005 40545 44039 40579
rect 44097 40545 44131 40579
rect 54861 40545 54895 40579
rect 57805 40545 57839 40579
rect 58817 40545 58851 40579
rect 62773 40545 62807 40579
rect 62957 40545 62991 40579
rect 64337 40545 64371 40579
rect 64429 40545 64463 40579
rect 65809 40545 65843 40579
rect 66177 40545 66211 40579
rect 66361 40545 66395 40579
rect 67373 40545 67407 40579
rect 67557 40545 67591 40579
rect 67925 40545 67959 40579
rect 71421 40545 71455 40579
rect 73077 40545 73111 40579
rect 73445 40545 73479 40579
rect 74733 40545 74767 40579
rect 74917 40545 74951 40579
rect 75377 40545 75411 40579
rect 80805 40545 80839 40579
rect 80989 40545 81023 40579
rect 82645 40545 82679 40579
rect 82829 40545 82863 40579
rect 83289 40545 83323 40579
rect 86509 40545 86543 40579
rect 89177 40545 89211 40579
rect 8033 40477 8067 40511
rect 11345 40477 11379 40511
rect 12909 40477 12943 40511
rect 20913 40477 20947 40511
rect 21649 40477 21683 40511
rect 26525 40477 26559 40511
rect 26801 40477 26835 40511
rect 33425 40477 33459 40511
rect 37841 40477 37875 40511
rect 39037 40477 39071 40511
rect 43361 40477 43395 40511
rect 44925 40477 44959 40511
rect 49801 40477 49835 40511
rect 55137 40477 55171 40511
rect 63325 40477 63359 40511
rect 64889 40477 64923 40511
rect 71513 40477 71547 40511
rect 73169 40477 73203 40511
rect 73537 40477 73571 40511
rect 75193 40477 75227 40511
rect 86233 40477 86267 40511
rect 86693 40477 86727 40511
rect 86785 40477 86819 40511
rect 89453 40477 89487 40511
rect 4997 40409 5031 40443
rect 5733 40341 5767 40375
rect 7389 40341 7423 40375
rect 11161 40341 11195 40375
rect 13737 40341 13771 40375
rect 22293 40341 22327 40375
rect 27905 40341 27939 40375
rect 28273 40341 28307 40375
rect 30297 40341 30331 40375
rect 33885 40341 33919 40375
rect 39313 40341 39347 40375
rect 42901 40341 42935 40375
rect 49571 40341 49605 40375
rect 49709 40341 49743 40375
rect 50077 40341 50111 40375
rect 57897 40341 57931 40375
rect 58909 40341 58943 40375
rect 64153 40341 64187 40375
rect 64981 40341 65015 40375
rect 65533 40341 65567 40375
rect 67189 40341 67223 40375
rect 72525 40341 72559 40375
rect 73721 40341 73755 40375
rect 80713 40341 80747 40375
rect 81449 40341 81483 40375
rect 90557 40341 90591 40375
rect 26433 40137 26467 40171
rect 27537 40137 27571 40171
rect 38853 40137 38887 40171
rect 40785 40137 40819 40171
rect 66729 40137 66763 40171
rect 3801 40069 3835 40103
rect 4261 40069 4295 40103
rect 9137 40069 9171 40103
rect 33517 40069 33551 40103
rect 38945 40069 38979 40103
rect 42257 40069 42291 40103
rect 49479 40069 49513 40103
rect 49617 40069 49651 40103
rect 52929 40069 52963 40103
rect 67557 40069 67591 40103
rect 72157 40069 72191 40103
rect 85681 40069 85715 40103
rect 2605 40001 2639 40035
rect 8309 40001 8343 40035
rect 9229 40001 9263 40035
rect 13001 40001 13035 40035
rect 17785 40001 17819 40035
rect 21741 40001 21775 40035
rect 25145 40001 25179 40035
rect 31769 40001 31803 40035
rect 40656 40001 40690 40035
rect 40877 40001 40911 40035
rect 43545 40001 43579 40035
rect 44833 40001 44867 40035
rect 49709 40001 49743 40035
rect 74181 40001 74215 40035
rect 79425 40001 79459 40035
rect 82369 40001 82403 40035
rect 83105 40001 83139 40035
rect 84577 40001 84611 40035
rect 85221 40001 85255 40035
rect 88625 40001 88659 40035
rect 90741 40001 90775 40035
rect 91017 40001 91051 40035
rect 2881 39933 2915 39967
rect 2973 39933 3007 39967
rect 3433 39933 3467 39967
rect 3617 39933 3651 39967
rect 4905 39933 4939 39967
rect 5457 39933 5491 39967
rect 8391 39933 8425 39967
rect 8769 39933 8803 39967
rect 8861 39933 8895 39967
rect 13185 39933 13219 39967
rect 13737 39933 13771 39967
rect 13912 39933 13946 39967
rect 14473 39933 14507 39967
rect 15209 39933 15243 39967
rect 14289 39865 14323 39899
rect 19993 39933 20027 39967
rect 20269 39933 20303 39967
rect 25421 39933 25455 39967
rect 25513 39933 25547 39967
rect 25973 39933 26007 39967
rect 26157 39933 26191 39967
rect 26801 39933 26835 39967
rect 27445 39933 27479 39967
rect 31953 39933 31987 39967
rect 32413 39933 32447 39967
rect 32505 39933 32539 39967
rect 33333 39933 33367 39967
rect 37289 39933 37323 39967
rect 37473 39933 37507 39967
rect 37933 39933 37967 39967
rect 38025 39933 38059 39967
rect 40509 39933 40543 39967
rect 42441 39933 42475 39967
rect 43729 39933 43763 39967
rect 44189 39933 44223 39967
rect 44281 39933 44315 39967
rect 45109 39933 45143 39967
rect 50077 39933 50111 39967
rect 52009 39933 52043 39967
rect 52101 39933 52135 39967
rect 52469 39933 52503 39967
rect 52561 39933 52595 39967
rect 54309 39933 54343 39967
rect 57069 39933 57103 39967
rect 57345 39933 57379 39967
rect 57621 39933 57655 39967
rect 63233 39933 63267 39967
rect 64245 39933 64279 39967
rect 64521 39933 64555 39967
rect 67005 39933 67039 39967
rect 70685 39933 70719 39967
rect 70777 39933 70811 39967
rect 71053 39933 71087 39967
rect 73997 39933 74031 39967
rect 74457 39933 74491 39967
rect 77493 39933 77527 39967
rect 77769 39933 77803 39967
rect 80437 39933 80471 39967
rect 80529 39933 80563 39967
rect 80805 39933 80839 39967
rect 80897 39933 80931 39967
rect 82645 39933 82679 39967
rect 84209 39933 84243 39967
rect 85405 39933 85439 39967
rect 85957 39933 85991 39967
rect 86233 39933 86267 39967
rect 88533 39933 88567 39967
rect 91293 39933 91327 39967
rect 31585 39865 31619 39899
rect 33057 39865 33091 39899
rect 38577 39865 38611 39899
rect 49341 39865 49375 39899
rect 51549 39865 51583 39899
rect 59001 39865 59035 39899
rect 63325 39865 63359 39899
rect 66913 39865 66947 39899
rect 67465 39865 67499 39899
rect 74365 39865 74399 39899
rect 74917 39865 74951 39899
rect 79793 39865 79827 39899
rect 82565 39865 82599 39899
rect 4997 39797 5031 39831
rect 7849 39797 7883 39831
rect 12817 39797 12851 39831
rect 15393 39797 15427 39831
rect 17785 39797 17819 39831
rect 21557 39797 21591 39831
rect 37105 39797 37139 39831
rect 41153 39797 41187 39831
rect 42625 39797 42659 39831
rect 53389 39797 53423 39831
rect 53573 39797 53607 39831
rect 54125 39797 54159 39831
rect 56793 39797 56827 39831
rect 64153 39797 64187 39831
rect 65625 39797 65659 39831
rect 73813 39797 73847 39831
rect 77585 39797 77619 39831
rect 79241 39797 79275 39831
rect 81081 39797 81115 39831
rect 84393 39797 84427 39831
rect 86601 39797 86635 39831
rect 92397 39797 92431 39831
rect 4169 39593 4203 39627
rect 15485 39593 15519 39627
rect 19717 39593 19751 39627
rect 20177 39593 20211 39627
rect 31953 39593 31987 39627
rect 3341 39525 3375 39559
rect 4997 39525 5031 39559
rect 2605 39457 2639 39491
rect 2973 39457 3007 39491
rect 4353 39457 4387 39491
rect 4537 39457 4571 39491
rect 7297 39457 7331 39491
rect 7619 39457 7653 39491
rect 7849 39457 7883 39491
rect 9689 39457 9723 39491
rect 9965 39457 9999 39491
rect 11805 39457 11839 39491
rect 13093 39457 13127 39491
rect 13645 39457 13679 39491
rect 13829 39457 13863 39491
rect 15301 39457 15335 39491
rect 19717 39457 19751 39491
rect 19809 39457 19843 39491
rect 20913 39457 20947 39491
rect 27537 39457 27571 39491
rect 27629 39457 27663 39491
rect 43729 39593 43763 39627
rect 50169 39593 50203 39627
rect 50721 39593 50755 39627
rect 51365 39593 51399 39627
rect 71605 39593 71639 39627
rect 72617 39593 72651 39627
rect 78781 39593 78815 39627
rect 81357 39593 81391 39627
rect 85957 39593 85991 39627
rect 88809 39593 88843 39627
rect 91109 39593 91143 39627
rect 48329 39525 48363 39559
rect 48697 39525 48731 39559
rect 54677 39525 54711 39559
rect 56425 39525 56459 39559
rect 59553 39525 59587 39559
rect 83749 39525 83783 39559
rect 32321 39457 32355 39491
rect 32873 39457 32907 39491
rect 33057 39457 33091 39491
rect 34345 39457 34379 39491
rect 35081 39457 35115 39491
rect 39405 39457 39439 39491
rect 39497 39457 39531 39491
rect 39865 39457 39899 39491
rect 39957 39457 39991 39491
rect 40785 39457 40819 39491
rect 43729 39457 43763 39491
rect 44189 39457 44223 39491
rect 44373 39457 44407 39491
rect 44833 39457 44867 39491
rect 44925 39457 44959 39491
rect 46397 39457 46431 39491
rect 49157 39457 49191 39491
rect 49617 39457 49651 39491
rect 49709 39457 49743 39491
rect 51549 39457 51583 39491
rect 51825 39457 51859 39491
rect 52101 39457 52135 39491
rect 52653 39457 52687 39491
rect 52837 39457 52871 39491
rect 55045 39457 55079 39491
rect 58081 39457 58115 39491
rect 58541 39457 58575 39491
rect 58633 39457 58667 39491
rect 60197 39457 60231 39491
rect 60841 39457 60875 39491
rect 61209 39457 61243 39491
rect 62037 39457 62071 39491
rect 62497 39457 62531 39491
rect 66269 39457 66303 39491
rect 71513 39457 71547 39491
rect 72525 39457 72559 39491
rect 73813 39457 73847 39491
rect 75377 39457 75411 39491
rect 77309 39457 77343 39491
rect 77401 39457 77435 39491
rect 79885 39457 79919 39491
rect 81265 39457 81299 39491
rect 82737 39457 82771 39491
rect 82829 39457 82863 39491
rect 84393 39457 84427 39491
rect 84761 39457 84795 39491
rect 85037 39457 85071 39491
rect 85773 39457 85807 39491
rect 86141 39457 86175 39491
rect 86877 39457 86911 39491
rect 87153 39457 87187 39491
rect 88717 39457 88751 39491
rect 89913 39457 89947 39491
rect 91017 39457 91051 39491
rect 3157 39389 3191 39423
rect 6653 39389 6687 39423
rect 7389 39389 7423 39423
rect 12173 39389 12207 39423
rect 12909 39389 12943 39423
rect 31861 39389 31895 39423
rect 31953 39389 31987 39423
rect 32137 39389 32171 39423
rect 33701 39389 33735 39423
rect 34713 39389 34747 39423
rect 40969 39389 41003 39423
rect 46544 39389 46578 39423
rect 46765 39389 46799 39423
rect 48329 39389 48363 39423
rect 48513 39389 48547 39423
rect 48973 39389 49007 39423
rect 50537 39389 50571 39423
rect 51917 39389 51951 39423
rect 54769 39389 54803 39423
rect 57989 39389 58023 39423
rect 59185 39389 59219 39423
rect 60749 39389 60783 39423
rect 61301 39389 61335 39423
rect 6377 39321 6411 39355
rect 45385 39321 45419 39355
rect 46673 39321 46707 39355
rect 53021 39321 53055 39355
rect 53665 39321 53699 39355
rect 65993 39389 66027 39423
rect 73537 39389 73571 39423
rect 77677 39389 77711 39423
rect 79977 39389 80011 39423
rect 84485 39389 84519 39423
rect 84853 39389 84887 39423
rect 62313 39321 62347 39355
rect 83657 39321 83691 39355
rect 6561 39253 6595 39287
rect 9781 39253 9815 39287
rect 11989 39253 12023 39287
rect 12725 39253 12759 39287
rect 14105 39253 14139 39287
rect 14473 39253 14507 39287
rect 19901 39253 19935 39287
rect 21005 39253 21039 39287
rect 27813 39253 27847 39287
rect 31677 39253 31711 39287
rect 33333 39253 33367 39287
rect 33885 39253 33919 39287
rect 34483 39253 34517 39287
rect 34621 39253 34655 39287
rect 40417 39253 40451 39287
rect 43821 39253 43855 39287
rect 44005 39253 44039 39287
rect 45753 39253 45787 39287
rect 45937 39253 45971 39287
rect 47041 39253 47075 39287
rect 51641 39253 51675 39287
rect 53481 39253 53515 39287
rect 54309 39253 54343 39287
rect 59369 39253 59403 39287
rect 62037 39253 62071 39287
rect 62129 39253 62163 39287
rect 65809 39253 65843 39287
rect 67373 39253 67407 39287
rect 74917 39253 74951 39287
rect 86969 39253 87003 39287
rect 90005 39253 90039 39287
rect 8953 39049 8987 39083
rect 20729 39049 20763 39083
rect 51871 39049 51905 39083
rect 84025 39049 84059 39083
rect 84577 39049 84611 39083
rect 85681 39049 85715 39083
rect 9137 38981 9171 39015
rect 15301 38981 15335 39015
rect 31861 38981 31895 39015
rect 33149 38981 33183 39015
rect 39018 38981 39052 39015
rect 39129 38981 39163 39015
rect 39773 38981 39807 39015
rect 46397 38981 46431 39015
rect 49893 38981 49927 39015
rect 50445 38981 50479 39015
rect 50629 38981 50663 39015
rect 52009 38981 52043 39015
rect 60749 38981 60783 39015
rect 83565 38981 83599 39015
rect 84209 38981 84243 39015
rect 2789 38913 2823 38947
rect 11437 38913 11471 38947
rect 13001 38913 13035 38947
rect 14381 38913 14415 38947
rect 15117 38913 15151 38947
rect 31585 38913 31619 38947
rect 31953 38913 31987 38947
rect 33701 38913 33735 38947
rect 39221 38913 39255 38947
rect 45109 38913 45143 38947
rect 45385 38913 45419 38947
rect 45569 38913 45603 38947
rect 46489 38913 46523 38947
rect 52101 38913 52135 38947
rect 52469 38913 52503 38947
rect 71605 38913 71639 38947
rect 72525 38913 72559 38947
rect 74641 38913 74675 38947
rect 82553 38913 82587 38947
rect 83896 38913 83930 38947
rect 84117 38913 84151 38947
rect 2513 38845 2547 38879
rect 8033 38845 8067 38879
rect 8217 38845 8251 38879
rect 8585 38845 8619 38879
rect 8769 38845 8803 38879
rect 10149 38845 10183 38879
rect 10333 38845 10367 38879
rect 10793 38845 10827 38879
rect 10885 38845 10919 38879
rect 12725 38845 12759 38879
rect 14473 38845 14507 38879
rect 15209 38845 15243 38879
rect 19165 38845 19199 38879
rect 19441 38845 19475 38879
rect 21649 38845 21683 38879
rect 26157 38845 26191 38879
rect 26433 38845 26467 38879
rect 27813 38845 27847 38879
rect 29285 38845 29319 38879
rect 32137 38845 32171 38879
rect 32689 38845 32723 38879
rect 32873 38845 32907 38879
rect 38853 38845 38887 38879
rect 43821 38845 43855 38879
rect 44005 38845 44039 38879
rect 44465 38845 44499 38879
rect 44557 38845 44591 38879
rect 46121 38845 46155 38879
rect 46268 38845 46302 38879
rect 48513 38845 48547 38879
rect 48697 38845 48731 38879
rect 48881 38845 48915 38879
rect 49433 38845 49467 38879
rect 49617 38845 49651 38879
rect 54317 38845 54351 38879
rect 58265 38845 58299 38879
rect 58449 38845 58483 38879
rect 58633 38845 58667 38879
rect 59093 38845 59127 38879
rect 59185 38845 59219 38879
rect 60013 38845 60047 38879
rect 61223 38845 61257 38879
rect 61393 38845 61427 38879
rect 61669 38845 61703 38879
rect 61853 38845 61887 38879
rect 65533 38845 65567 38879
rect 65809 38845 65843 38879
rect 69673 38845 69707 38879
rect 71145 38845 71179 38879
rect 71329 38845 71363 38879
rect 71697 38845 71731 38879
rect 72893 38845 72927 38879
rect 74181 38845 74215 38879
rect 74365 38845 74399 38879
rect 77033 38845 77067 38879
rect 77309 38845 77343 38879
rect 82461 38845 82495 38879
rect 82921 38845 82955 38879
rect 85589 38845 85623 38879
rect 86049 38845 86083 38879
rect 86877 38845 86911 38879
rect 86969 38845 87003 38879
rect 87153 38845 87187 38879
rect 91569 38845 91603 38879
rect 92857 38845 92891 38879
rect 7573 38777 7607 38811
rect 33517 38777 33551 38811
rect 39589 38777 39623 38811
rect 51733 38777 51767 38811
rect 59737 38777 59771 38811
rect 83381 38777 83415 38811
rect 83749 38777 83783 38811
rect 85405 38777 85439 38811
rect 91661 38777 91695 38811
rect 92673 38777 92707 38811
rect 93225 38777 93259 38811
rect 3893 38709 3927 38743
rect 4353 38709 4387 38743
rect 9965 38709 9999 38743
rect 20913 38709 20947 38743
rect 21741 38709 21775 38743
rect 27905 38709 27939 38743
rect 29377 38709 29411 38743
rect 43453 38709 43487 38743
rect 43637 38709 43671 38743
rect 46765 38709 46799 38743
rect 50169 38709 50203 38743
rect 51457 38709 51491 38743
rect 54125 38709 54159 38743
rect 65625 38709 65659 38743
rect 69765 38709 69799 38743
rect 70501 38709 70535 38743
rect 70961 38709 70995 38743
rect 72709 38709 72743 38743
rect 76941 38709 76975 38743
rect 78413 38709 78447 38743
rect 82001 38709 82035 38743
rect 87337 38709 87371 38743
rect 93409 38709 93443 38743
rect 4169 38505 4203 38539
rect 4997 38505 5031 38539
rect 8677 38505 8711 38539
rect 22109 38505 22143 38539
rect 31953 38505 31987 38539
rect 18521 38437 18555 38471
rect 19901 38437 19935 38471
rect 20177 38437 20211 38471
rect 20269 38437 20303 38471
rect 4353 38369 4387 38403
rect 4629 38369 4663 38403
rect 7389 38369 7423 38403
rect 8493 38369 8527 38403
rect 11437 38369 11471 38403
rect 11989 38369 12023 38403
rect 12173 38369 12207 38403
rect 13461 38369 13495 38403
rect 18797 38369 18831 38403
rect 18889 38369 18923 38403
rect 19395 38369 19429 38403
rect 19533 38369 19567 38403
rect 11253 38301 11287 38335
rect 13553 38301 13587 38335
rect 84669 38505 84703 38539
rect 84761 38505 84795 38539
rect 85957 38505 85991 38539
rect 89085 38505 89119 38539
rect 90097 38505 90131 38539
rect 95709 38505 95743 38539
rect 52929 38437 52963 38471
rect 69305 38437 69339 38471
rect 70133 38437 70167 38471
rect 71145 38437 71179 38471
rect 21097 38369 21131 38403
rect 21649 38369 21683 38403
rect 21833 38369 21867 38403
rect 27905 38369 27939 38403
rect 28457 38369 28491 38403
rect 28641 38369 28675 38403
rect 29285 38369 29319 38403
rect 31953 38369 31987 38403
rect 32873 38369 32907 38403
rect 39037 38369 39071 38403
rect 39497 38369 39531 38403
rect 39589 38369 39623 38403
rect 40325 38369 40359 38403
rect 44465 38369 44499 38403
rect 44925 38369 44959 38403
rect 45017 38369 45051 38403
rect 45845 38369 45879 38403
rect 50353 38369 50387 38403
rect 50813 38369 50847 38403
rect 50905 38369 50939 38403
rect 53076 38369 53110 38403
rect 56609 38369 56643 38403
rect 62865 38369 62899 38403
rect 63417 38369 63451 38403
rect 63601 38369 63635 38403
rect 70317 38369 70351 38403
rect 70961 38369 70995 38403
rect 71237 38369 71271 38403
rect 71881 38369 71915 38403
rect 72065 38369 72099 38403
rect 72433 38369 72467 38403
rect 72525 38369 72559 38403
rect 74365 38369 74399 38403
rect 77401 38369 77435 38403
rect 77677 38369 77711 38403
rect 81541 38369 81575 38403
rect 81817 38369 81851 38403
rect 82829 38369 82863 38403
rect 82921 38369 82955 38403
rect 20729 38301 20763 38335
rect 20913 38301 20947 38335
rect 27721 38301 27755 38335
rect 33241 38301 33275 38335
rect 38945 38301 38979 38335
rect 40141 38301 40175 38335
rect 44281 38301 44315 38335
rect 45477 38301 45511 38335
rect 50261 38301 50295 38335
rect 51733 38301 51767 38335
rect 53297 38301 53331 38335
rect 57621 38301 57655 38335
rect 57897 38301 57931 38335
rect 59093 38301 59127 38335
rect 62681 38301 62715 38335
rect 67649 38301 67683 38335
rect 67925 38301 67959 38335
rect 71421 38301 71455 38335
rect 85865 38437 85899 38471
rect 88441 38437 88475 38471
rect 90465 38437 90499 38471
rect 85129 38369 85163 38403
rect 85276 38369 85310 38403
rect 89269 38369 89303 38403
rect 91109 38369 91143 38403
rect 91477 38369 91511 38403
rect 85497 38301 85531 38335
rect 88588 38301 88622 38335
rect 88809 38301 88843 38335
rect 91017 38301 91051 38335
rect 91569 38301 91603 38335
rect 94329 38301 94363 38335
rect 94605 38301 94639 38335
rect 33038 38233 33072 38267
rect 33517 38233 33551 38267
rect 49801 38233 49835 38267
rect 53849 38233 53883 38267
rect 70409 38233 70443 38267
rect 71237 38233 71271 38267
rect 81633 38233 81667 38267
rect 84669 38233 84703 38267
rect 85405 38233 85439 38267
rect 89453 38233 89487 38267
rect 7573 38165 7607 38199
rect 11069 38165 11103 38199
rect 12449 38165 12483 38199
rect 13829 38165 13863 38199
rect 20269 38165 20303 38199
rect 20453 38165 20487 38199
rect 27537 38165 27571 38199
rect 28917 38165 28951 38199
rect 33149 38165 33183 38199
rect 40509 38165 40543 38199
rect 46029 38165 46063 38199
rect 49985 38165 50019 38199
rect 51365 38165 51399 38199
rect 53205 38165 53239 38199
rect 53389 38165 53423 38199
rect 56701 38165 56735 38199
rect 57437 38165 57471 38199
rect 62129 38165 62163 38199
rect 62313 38165 62347 38199
rect 62589 38165 62623 38199
rect 63877 38165 63911 38199
rect 67281 38165 67315 38199
rect 67465 38165 67499 38199
rect 74181 38165 74215 38199
rect 77493 38165 77527 38199
rect 82461 38165 82495 38199
rect 82645 38165 82679 38199
rect 83105 38165 83139 38199
rect 84945 38165 84979 38199
rect 88717 38165 88751 38199
rect 89637 38165 89671 38199
rect 90281 38165 90315 38199
rect 94237 38165 94271 38199
rect 5181 37961 5215 37995
rect 59001 37961 59035 37995
rect 60270 37961 60304 37995
rect 84117 37961 84151 37995
rect 26617 37893 26651 37927
rect 27077 37893 27111 37927
rect 31493 37893 31527 37927
rect 31677 37893 31711 37927
rect 40785 37893 40819 37927
rect 45385 37893 45419 37927
rect 56333 37893 56367 37927
rect 85865 37893 85899 37927
rect 89177 37893 89211 37927
rect 89453 37893 89487 37927
rect 90189 37893 90223 37927
rect 2789 37825 2823 37859
rect 8309 37825 8343 37859
rect 12725 37825 12759 37859
rect 18521 37825 18555 37859
rect 19257 37825 19291 37859
rect 21097 37825 21131 37859
rect 32229 37825 32263 37859
rect 38117 37825 38151 37859
rect 39497 37825 39531 37859
rect 40656 37825 40690 37859
rect 40877 37825 40911 37859
rect 41245 37825 41279 37859
rect 45569 37825 45603 37859
rect 51273 37825 51307 37859
rect 51733 37825 51767 37859
rect 59921 37825 59955 37859
rect 60473 37825 60507 37859
rect 64429 37825 64463 37859
rect 64705 37825 64739 37859
rect 68753 37825 68787 37859
rect 70225 37825 70259 37859
rect 71605 37825 71639 37859
rect 72709 37825 72743 37859
rect 76757 37825 76791 37859
rect 81633 37825 81667 37859
rect 89913 37825 89947 37859
rect 91569 37825 91603 37859
rect 94053 37825 94087 37859
rect 2513 37757 2547 37791
rect 4997 37757 5031 37791
rect 8217 37757 8251 37791
rect 8585 37757 8619 37791
rect 8769 37757 8803 37791
rect 12449 37757 12483 37791
rect 18153 37757 18187 37791
rect 19533 37757 19567 37791
rect 20913 37757 20947 37791
rect 21741 37757 21775 37791
rect 25651 37757 25685 37791
rect 25789 37757 25823 37791
rect 26157 37757 26191 37791
rect 26249 37757 26283 37791
rect 31861 37757 31895 37791
rect 31953 37757 31987 37791
rect 33609 37757 33643 37791
rect 37841 37757 37875 37791
rect 40509 37757 40543 37791
rect 43821 37757 43855 37791
rect 44005 37757 44039 37791
rect 44465 37757 44499 37791
rect 44557 37757 44591 37791
rect 51457 37757 51491 37791
rect 51917 37757 51951 37791
rect 52377 37757 52411 37791
rect 52469 37757 52503 37791
rect 56241 37757 56275 37791
rect 57345 37757 57379 37791
rect 57621 37757 57655 37791
rect 57897 37757 57931 37791
rect 60335 37757 60369 37791
rect 60841 37757 60875 37791
rect 68569 37757 68603 37791
rect 68661 37757 68695 37791
rect 68937 37757 68971 37791
rect 70685 37757 70719 37791
rect 70869 37757 70903 37791
rect 71237 37757 71271 37791
rect 71329 37757 71363 37791
rect 72249 37757 72283 37791
rect 72341 37757 72375 37791
rect 72525 37757 72559 37791
rect 76849 37757 76883 37791
rect 77493 37757 77527 37791
rect 77677 37757 77711 37791
rect 81265 37757 81299 37791
rect 81357 37757 81391 37791
rect 83841 37757 83875 37791
rect 84025 37757 84059 37791
rect 85681 37757 85715 37791
rect 89361 37757 89395 37791
rect 89607 37757 89641 37791
rect 91201 37757 91235 37791
rect 91661 37757 91695 37791
rect 93317 37757 93351 37791
rect 93501 37757 93535 37791
rect 93593 37757 93627 37791
rect 94973 37757 95007 37791
rect 95249 37757 95283 37791
rect 96629 37757 96663 37791
rect 7573 37689 7607 37723
rect 14105 37689 14139 37723
rect 25421 37689 25455 37723
rect 59737 37689 59771 37723
rect 60105 37689 60139 37723
rect 66085 37689 66119 37723
rect 91017 37689 91051 37723
rect 95157 37689 95191 37723
rect 95709 37689 95743 37723
rect 3893 37621 3927 37655
rect 4261 37621 4295 37655
rect 14197 37621 14231 37655
rect 18337 37621 18371 37655
rect 21833 37621 21867 37655
rect 37657 37621 37691 37655
rect 40233 37621 40267 37655
rect 45017 37621 45051 37655
rect 52929 37621 52963 37655
rect 53297 37621 53331 37655
rect 57345 37621 57379 37655
rect 57437 37621 57471 37655
rect 64245 37621 64279 37655
rect 68569 37621 68603 37655
rect 69121 37621 69155 37655
rect 71789 37621 71823 37655
rect 76941 37621 76975 37655
rect 82737 37621 82771 37655
rect 83657 37621 83691 37655
rect 93133 37621 93167 37655
rect 94789 37621 94823 37655
rect 96721 37621 96755 37655
rect 8953 37417 8987 37451
rect 19441 37417 19475 37451
rect 19809 37417 19843 37451
rect 22109 37417 22143 37451
rect 23397 37417 23431 37451
rect 24501 37417 24535 37451
rect 25789 37417 25823 37451
rect 29009 37417 29043 37451
rect 34437 37417 34471 37451
rect 40049 37417 40083 37451
rect 40877 37417 40911 37451
rect 47961 37417 47995 37451
rect 57989 37417 58023 37451
rect 69581 37417 69615 37451
rect 70685 37417 70719 37451
rect 70869 37417 70903 37451
rect 71697 37417 71731 37451
rect 72801 37417 72835 37451
rect 75377 37417 75411 37451
rect 83197 37417 83231 37451
rect 8217 37349 8251 37383
rect 39405 37349 39439 37383
rect 40233 37349 40267 37383
rect 44649 37349 44683 37383
rect 54585 37349 54619 37383
rect 55321 37349 55355 37383
rect 82921 37349 82955 37383
rect 90189 37349 90223 37383
rect 91293 37349 91327 37383
rect 91477 37349 91511 37383
rect 95249 37349 95283 37383
rect 4353 37281 4387 37315
rect 8401 37281 8435 37315
rect 12449 37281 12483 37315
rect 12541 37281 12575 37315
rect 13185 37281 13219 37315
rect 13921 37281 13955 37315
rect 14565 37281 14599 37315
rect 18153 37281 18187 37315
rect 18245 37281 18279 37315
rect 18429 37281 18463 37315
rect 18981 37281 19015 37315
rect 19165 37281 19199 37315
rect 21097 37281 21131 37315
rect 21649 37281 21683 37315
rect 21833 37281 21867 37315
rect 22937 37281 22971 37315
rect 23213 37281 23247 37315
rect 25053 37281 25087 37315
rect 25421 37281 25455 37315
rect 25605 37281 25639 37315
rect 27353 37281 27387 37315
rect 27537 37281 27571 37315
rect 27721 37281 27755 37315
rect 28273 37281 28307 37315
rect 28457 37281 28491 37315
rect 32505 37281 32539 37315
rect 32689 37281 32723 37315
rect 34621 37281 34655 37315
rect 35173 37281 35207 37315
rect 35633 37281 35667 37315
rect 36185 37281 36219 37315
rect 36369 37281 36403 37315
rect 38025 37281 38059 37315
rect 43821 37281 43855 37315
rect 44833 37281 44867 37315
rect 45109 37281 45143 37315
rect 46489 37281 46523 37315
rect 47869 37281 47903 37315
rect 49065 37281 49099 37315
rect 50077 37281 50111 37315
rect 50261 37281 50295 37315
rect 50445 37281 50479 37315
rect 50905 37281 50939 37315
rect 50997 37281 51031 37315
rect 52009 37281 52043 37315
rect 56977 37281 57011 37315
rect 57437 37281 57471 37315
rect 57529 37281 57563 37315
rect 62221 37281 62255 37315
rect 62405 37281 62439 37315
rect 62957 37281 62991 37315
rect 63509 37281 63543 37315
rect 63693 37281 63727 37315
rect 69949 37281 69983 37315
rect 70317 37281 70351 37315
rect 71881 37281 71915 37315
rect 72065 37281 72099 37315
rect 72433 37281 72467 37315
rect 75193 37281 75227 37315
rect 82829 37281 82863 37315
rect 83105 37281 83139 37315
rect 85037 37281 85071 37315
rect 85313 37281 85347 37315
rect 89453 37281 89487 37315
rect 89729 37281 89763 37315
rect 91661 37281 91695 37315
rect 94053 37281 94087 37315
rect 94237 37281 94271 37315
rect 95433 37281 95467 37315
rect 95709 37281 95743 37315
rect 4077 37213 4111 37247
rect 5825 37213 5859 37247
rect 13829 37213 13863 37247
rect 20913 37213 20947 37247
rect 22477 37213 22511 37247
rect 25145 37213 25179 37247
rect 25973 37213 26007 37247
rect 35265 37213 35299 37247
rect 35449 37213 35483 37247
rect 36737 37213 36771 37247
rect 37565 37213 37599 37247
rect 37749 37213 37783 37247
rect 40601 37213 40635 37247
rect 43913 37213 43947 37247
rect 54732 37213 54766 37247
rect 54953 37213 54987 37247
rect 56241 37213 56275 37247
rect 56425 37213 56459 37247
rect 56793 37213 56827 37247
rect 62773 37213 62807 37247
rect 69765 37213 69799 37247
rect 70225 37213 70259 37247
rect 72341 37213 72375 37247
rect 77033 37213 77067 37247
rect 77309 37213 77343 37247
rect 84485 37213 84519 37247
rect 85497 37213 85531 37247
rect 89545 37213 89579 37247
rect 92029 37213 92063 37247
rect 94605 37213 94639 37247
rect 22937 37145 22971 37179
rect 23029 37145 23063 37179
rect 28733 37145 28767 37179
rect 5457 37077 5491 37111
rect 8493 37077 8527 37111
rect 12725 37077 12759 37111
rect 14105 37077 14139 37111
rect 20637 37077 20671 37111
rect 32873 37077 32907 37111
rect 40371 37077 40405 37111
rect 40509 37077 40543 37111
rect 49157 37077 49191 37111
rect 49341 37077 49375 37111
rect 51457 37077 51491 37111
rect 51733 37077 51767 37111
rect 54861 37077 54895 37111
rect 56609 37077 56643 37111
rect 62589 37077 62623 37111
rect 63969 37077 64003 37111
rect 72985 37077 73019 37111
rect 76757 37077 76791 37111
rect 78413 37077 78447 37111
rect 84301 37077 84335 37111
rect 90373 37077 90407 37111
rect 96997 37077 97031 37111
rect 3893 36873 3927 36907
rect 12725 36873 12759 36907
rect 35633 36873 35667 36907
rect 37013 36873 37047 36907
rect 39129 36873 39163 36907
rect 39405 36873 39439 36907
rect 53757 36873 53791 36907
rect 91109 36873 91143 36907
rect 91385 36873 91419 36907
rect 93869 36873 93903 36907
rect 96905 36873 96939 36907
rect 10057 36805 10091 36839
rect 14197 36805 14231 36839
rect 17049 36805 17083 36839
rect 22661 36805 22695 36839
rect 32045 36805 32079 36839
rect 2513 36737 2547 36771
rect 9413 36737 9447 36771
rect 9873 36737 9907 36771
rect 12817 36737 12851 36771
rect 13185 36737 13219 36771
rect 20821 36737 20855 36771
rect 24133 36737 24167 36771
rect 24961 36737 24995 36771
rect 27813 36737 27847 36771
rect 30297 36737 30331 36771
rect 31953 36737 31987 36771
rect 34713 36737 34747 36771
rect 35817 36737 35851 36771
rect 2789 36669 2823 36703
rect 4261 36669 4295 36703
rect 6929 36669 6963 36703
rect 7665 36669 7699 36703
rect 7941 36669 7975 36703
rect 8861 36669 8895 36703
rect 9689 36669 9723 36703
rect 10149 36669 10183 36703
rect 12596 36669 12630 36703
rect 14013 36669 14047 36703
rect 16681 36669 16715 36703
rect 16865 36669 16899 36703
rect 19073 36669 19107 36703
rect 19349 36669 19383 36703
rect 22385 36669 22419 36703
rect 22477 36669 22511 36703
rect 24317 36669 24351 36703
rect 25053 36669 25087 36703
rect 25421 36669 25455 36703
rect 25513 36669 25547 36703
rect 26893 36669 26927 36703
rect 27077 36669 27111 36703
rect 27445 36669 27479 36703
rect 27629 36669 27663 36703
rect 27997 36669 28031 36703
rect 30573 36669 30607 36703
rect 32965 36669 32999 36703
rect 12449 36601 12483 36635
rect 26433 36601 26467 36635
rect 44189 36805 44223 36839
rect 50721 36805 50755 36839
rect 54861 36805 54895 36839
rect 56609 36805 56643 36839
rect 57161 36805 57195 36839
rect 58449 36805 58483 36839
rect 64429 36805 64463 36839
rect 71697 36805 71731 36839
rect 71881 36805 71915 36839
rect 85129 36805 85163 36839
rect 85589 36805 85623 36839
rect 48697 36737 48731 36771
rect 50261 36737 50295 36771
rect 50592 36737 50626 36771
rect 50813 36737 50847 36771
rect 51181 36737 51215 36771
rect 54309 36737 54343 36771
rect 55321 36737 55355 36771
rect 55965 36737 55999 36771
rect 64521 36737 64555 36771
rect 64797 36737 64831 36771
rect 70317 36737 70351 36771
rect 71053 36737 71087 36771
rect 77309 36737 77343 36771
rect 77769 36737 77803 36771
rect 78689 36737 78723 36771
rect 86233 36737 86267 36771
rect 90097 36737 90131 36771
rect 35541 36669 35575 36703
rect 36001 36669 36035 36703
rect 36553 36669 36587 36703
rect 36737 36669 36771 36703
rect 39129 36669 39163 36703
rect 39313 36669 39347 36703
rect 44097 36669 44131 36703
rect 46949 36669 46983 36703
rect 47041 36669 47075 36703
rect 47317 36669 47351 36703
rect 48973 36669 49007 36703
rect 49157 36669 49191 36703
rect 49617 36669 49651 36703
rect 49709 36669 49743 36703
rect 50445 36669 50479 36703
rect 52745 36669 52779 36703
rect 52837 36669 52871 36703
rect 53205 36669 53239 36703
rect 53297 36669 53331 36703
rect 55873 36669 55907 36703
rect 56241 36669 56275 36703
rect 56333 36669 56367 36703
rect 56793 36669 56827 36703
rect 56977 36669 57011 36703
rect 57161 36669 57195 36703
rect 57345 36669 57379 36703
rect 57529 36669 57563 36703
rect 57989 36669 58023 36703
rect 58081 36669 58115 36703
rect 69305 36669 69339 36703
rect 70961 36669 70995 36703
rect 71329 36669 71363 36703
rect 71421 36669 71455 36703
rect 76757 36669 76791 36703
rect 77585 36669 77619 36703
rect 78597 36669 78631 36703
rect 79977 36669 80011 36703
rect 80437 36669 80471 36703
rect 81541 36669 81575 36703
rect 85405 36669 85439 36703
rect 85957 36669 85991 36703
rect 89729 36669 89763 36703
rect 91017 36669 91051 36703
rect 92949 36669 92983 36703
rect 93041 36669 93075 36703
rect 94605 36669 94639 36703
rect 94697 36669 94731 36703
rect 94973 36669 95007 36703
rect 95065 36669 95099 36703
rect 96813 36669 96847 36703
rect 97273 36669 97307 36703
rect 51273 36601 51307 36635
rect 52469 36601 52503 36635
rect 69397 36601 69431 36635
rect 79793 36601 79827 36635
rect 89545 36601 89579 36635
rect 90189 36601 90223 36635
rect 93961 36601 93995 36635
rect 96629 36601 96663 36635
rect 4537 36533 4571 36567
rect 7021 36533 7055 36567
rect 14473 36533 14507 36567
rect 20637 36533 20671 36567
rect 24501 36533 24535 36567
rect 32781 36533 32815 36567
rect 34713 36533 34747 36567
rect 48789 36533 48823 36567
rect 51549 36533 51583 36567
rect 54125 36533 54159 36567
rect 55045 36533 55079 36567
rect 66085 36533 66119 36567
rect 78413 36533 78447 36567
rect 80069 36533 80103 36567
rect 81725 36533 81759 36567
rect 84853 36533 84887 36567
rect 93593 36533 93627 36567
rect 8953 36329 8987 36363
rect 11805 36329 11839 36363
rect 26801 36329 26835 36363
rect 27169 36329 27203 36363
rect 36645 36329 36679 36363
rect 50997 36329 51031 36363
rect 57529 36329 57563 36363
rect 59185 36329 59219 36363
rect 62313 36329 62347 36363
rect 71513 36329 71547 36363
rect 72893 36329 72927 36363
rect 88809 36329 88843 36363
rect 97273 36329 97307 36363
rect 12449 36261 12483 36295
rect 24317 36261 24351 36295
rect 31125 36261 31159 36295
rect 45017 36261 45051 36295
rect 50721 36261 50755 36295
rect 8585 36193 8619 36227
rect 8769 36193 8803 36227
rect 11345 36193 11379 36227
rect 12788 36193 12822 36227
rect 14013 36193 14047 36227
rect 17877 36193 17911 36227
rect 18429 36193 18463 36227
rect 18613 36193 18647 36227
rect 19165 36193 19199 36227
rect 20913 36193 20947 36227
rect 24133 36193 24167 36227
rect 24961 36193 24995 36227
rect 25329 36193 25363 36227
rect 25513 36193 25547 36227
rect 26985 36193 27019 36227
rect 29009 36193 29043 36227
rect 29561 36193 29595 36227
rect 29745 36193 29779 36227
rect 31033 36193 31067 36227
rect 32137 36193 32171 36227
rect 35633 36193 35667 36227
rect 36185 36193 36219 36227
rect 36369 36193 36403 36227
rect 36921 36193 36955 36227
rect 39037 36193 39071 36227
rect 43177 36193 43211 36227
rect 43361 36193 43395 36227
rect 49617 36193 49651 36227
rect 50169 36193 50203 36227
rect 50353 36193 50387 36227
rect 56517 36193 56551 36227
rect 56977 36193 57011 36227
rect 57069 36193 57103 36227
rect 58541 36193 58575 36227
rect 62497 36193 62531 36227
rect 63325 36193 63359 36227
rect 63693 36193 63727 36227
rect 63877 36193 63911 36227
rect 69857 36193 69891 36227
rect 71421 36193 71455 36227
rect 7757 36125 7791 36159
rect 8309 36125 8343 36159
rect 13185 36125 13219 36159
rect 17693 36125 17727 36159
rect 24041 36125 24075 36159
rect 24869 36125 24903 36159
rect 28825 36125 28859 36159
rect 35449 36125 35483 36159
rect 39129 36125 39163 36159
rect 43637 36125 43671 36159
rect 49433 36125 49467 36159
rect 56333 36125 56367 36159
rect 57805 36125 57839 36159
rect 58909 36125 58943 36159
rect 62681 36125 62715 36159
rect 63141 36125 63175 36159
rect 69949 36125 69983 36159
rect 79333 36261 79367 36295
rect 89177 36261 89211 36295
rect 73077 36193 73111 36227
rect 73629 36193 73663 36227
rect 77585 36193 77619 36227
rect 78229 36193 78263 36227
rect 78505 36193 78539 36227
rect 79241 36193 79275 36227
rect 79425 36193 79459 36227
rect 84485 36193 84519 36227
rect 85865 36193 85899 36227
rect 86693 36193 86727 36227
rect 88993 36193 89027 36227
rect 89269 36193 89303 36227
rect 90557 36193 90591 36227
rect 92765 36193 92799 36227
rect 92857 36193 92891 36227
rect 94881 36193 94915 36227
rect 97089 36193 97123 36227
rect 72985 36125 73019 36159
rect 73813 36125 73847 36159
rect 77953 36125 77987 36159
rect 84209 36125 84243 36159
rect 94605 36125 94639 36159
rect 11529 36057 11563 36091
rect 12587 36057 12621 36091
rect 12725 36057 12759 36091
rect 14197 36057 14231 36091
rect 18797 36057 18831 36091
rect 32229 36057 32263 36091
rect 58081 36057 58115 36091
rect 72893 36057 72927 36091
rect 9045 35989 9079 36023
rect 13921 35989 13955 36023
rect 17509 35989 17543 36023
rect 21005 35989 21039 36023
rect 28641 35989 28675 36023
rect 30021 35989 30055 36023
rect 35357 35989 35391 36023
rect 49065 35989 49099 36023
rect 49341 35989 49375 36023
rect 51181 35989 51215 36023
rect 55965 35989 55999 36023
rect 56241 35989 56275 36023
rect 58679 35989 58713 36023
rect 58817 35989 58851 36023
rect 73261 35989 73295 36023
rect 79609 35989 79643 36023
rect 84025 35989 84059 36023
rect 86785 35989 86819 36023
rect 89453 35989 89487 36023
rect 90649 35989 90683 36023
rect 94421 35989 94455 36023
rect 96169 35989 96203 36023
rect 9781 35785 9815 35819
rect 19625 35785 19659 35819
rect 25237 35785 25271 35819
rect 71421 35785 71455 35819
rect 74273 35785 74307 35819
rect 77934 35785 77968 35819
rect 78045 35785 78079 35819
rect 79609 35785 79643 35819
rect 80069 35785 80103 35819
rect 86049 35785 86083 35819
rect 94145 35785 94179 35819
rect 96721 35785 96755 35819
rect 7205 35717 7239 35751
rect 20729 35717 20763 35751
rect 32137 35717 32171 35751
rect 42809 35717 42843 35751
rect 44465 35717 44499 35751
rect 52009 35717 52043 35751
rect 56149 35717 56183 35751
rect 63325 35717 63359 35751
rect 63693 35717 63727 35751
rect 67465 35717 67499 35751
rect 76113 35717 76147 35751
rect 78413 35717 78447 35751
rect 2789 35649 2823 35683
rect 7941 35649 7975 35683
rect 9505 35649 9539 35683
rect 12817 35649 12851 35683
rect 15301 35649 15335 35683
rect 16037 35649 16071 35683
rect 18337 35649 18371 35683
rect 26893 35649 26927 35683
rect 30573 35649 30607 35683
rect 35357 35649 35391 35683
rect 36645 35649 36679 35683
rect 43177 35649 43211 35683
rect 50445 35649 50479 35683
rect 51880 35649 51914 35683
rect 52101 35649 52135 35683
rect 55045 35649 55079 35683
rect 56701 35649 56735 35683
rect 56977 35649 57011 35683
rect 58633 35649 58667 35683
rect 64153 35649 64187 35683
rect 66269 35649 66303 35683
rect 2513 35581 2547 35615
rect 5457 35581 5491 35615
rect 5733 35581 5767 35615
rect 7113 35581 7147 35615
rect 7849 35581 7883 35615
rect 9229 35581 9263 35615
rect 10977 35581 11011 35615
rect 13001 35581 13035 35615
rect 13185 35581 13219 35615
rect 13553 35581 13587 35615
rect 13645 35581 13679 35615
rect 15209 35581 15243 35615
rect 15577 35581 15611 35615
rect 15761 35581 15795 35615
rect 15853 35581 15887 35615
rect 18061 35581 18095 35615
rect 20637 35581 20671 35615
rect 25053 35581 25087 35615
rect 26801 35581 26835 35615
rect 27169 35581 27203 35615
rect 27353 35581 27387 35615
rect 30297 35581 30331 35615
rect 35541 35581 35575 35615
rect 36093 35581 36127 35615
rect 36277 35581 36311 35615
rect 42901 35581 42935 35615
rect 49157 35581 49191 35615
rect 49341 35581 49375 35615
rect 49801 35581 49835 35615
rect 49893 35581 49927 35615
rect 55229 35581 55263 35615
rect 55689 35581 55723 35615
rect 55781 35581 55815 35615
rect 57345 35581 57379 35615
rect 57529 35581 57563 35615
rect 57989 35581 58023 35615
rect 58081 35581 58115 35615
rect 59093 35581 59127 35615
rect 63141 35581 63175 35615
rect 64061 35581 64095 35615
rect 64429 35581 64463 35615
rect 64613 35581 64647 35615
rect 66453 35581 66487 35615
rect 67005 35581 67039 35615
rect 67189 35581 67223 35615
rect 68845 35581 68879 35615
rect 69115 35581 69149 35615
rect 70501 35581 70535 35615
rect 71329 35581 71363 35615
rect 74181 35581 74215 35615
rect 74457 35581 74491 35615
rect 76205 35581 76239 35615
rect 76481 35581 76515 35615
rect 77769 35581 77803 35615
rect 78108 35581 78142 35615
rect 85681 35717 85715 35751
rect 93869 35717 93903 35751
rect 85552 35649 85586 35683
rect 85773 35649 85807 35683
rect 86417 35649 86451 35683
rect 88441 35649 88475 35683
rect 89729 35649 89763 35683
rect 90741 35649 90775 35683
rect 91017 35649 91051 35683
rect 95249 35649 95283 35683
rect 79977 35581 80011 35615
rect 80437 35581 80471 35615
rect 83749 35581 83783 35615
rect 84117 35581 84151 35615
rect 86233 35581 86267 35615
rect 88165 35581 88199 35615
rect 89545 35581 89579 35615
rect 89913 35581 89947 35615
rect 91293 35581 91327 35615
rect 93685 35581 93719 35615
rect 94973 35581 95007 35615
rect 96629 35581 96663 35615
rect 9045 35513 9079 35547
rect 14565 35513 14599 35547
rect 24869 35513 24903 35547
rect 36921 35513 36955 35547
rect 50905 35513 50939 35547
rect 51732 35513 51766 35547
rect 54861 35513 54895 35547
rect 76113 35513 76147 35547
rect 76389 35513 76423 35547
rect 76941 35513 76975 35547
rect 77677 35513 77711 35547
rect 78689 35513 78723 35547
rect 79609 35513 79643 35547
rect 79793 35513 79827 35547
rect 85405 35513 85439 35547
rect 87981 35513 88015 35547
rect 91201 35513 91235 35547
rect 91753 35513 91787 35547
rect 94789 35513 94823 35547
rect 3893 35445 3927 35479
rect 4353 35445 4387 35479
rect 5273 35445 5307 35479
rect 10885 35445 10919 35479
rect 11161 35445 11195 35479
rect 13829 35445 13863 35479
rect 14013 35445 14047 35479
rect 19901 35445 19935 35479
rect 26433 35445 26467 35479
rect 31861 35445 31895 35479
rect 35173 35445 35207 35479
rect 48789 35445 48823 35479
rect 48973 35445 49007 35479
rect 50721 35445 50755 35479
rect 52377 35445 52411 35479
rect 54677 35445 54711 35479
rect 56517 35445 56551 35479
rect 58909 35445 58943 35479
rect 65717 35445 65751 35479
rect 65901 35445 65935 35479
rect 66085 35445 66119 35479
rect 70593 35445 70627 35479
rect 83933 35445 83967 35479
rect 89177 35445 89211 35479
rect 94605 35445 94639 35479
rect 5825 35241 5859 35275
rect 7389 35241 7423 35275
rect 19441 35241 19475 35275
rect 19809 35241 19843 35275
rect 25145 35241 25179 35275
rect 28273 35241 28307 35275
rect 30389 35241 30423 35275
rect 34345 35241 34379 35275
rect 34713 35241 34747 35275
rect 39037 35241 39071 35275
rect 42257 35241 42291 35275
rect 48145 35241 48179 35275
rect 51641 35241 51675 35275
rect 56333 35241 56367 35275
rect 63325 35241 63359 35275
rect 65809 35241 65843 35275
rect 65901 35241 65935 35275
rect 66085 35241 66119 35275
rect 90649 35241 90683 35275
rect 12909 35173 12943 35207
rect 14381 35173 14415 35207
rect 24409 35173 24443 35207
rect 43085 35173 43119 35207
rect 58081 35173 58115 35207
rect 70501 35173 70535 35207
rect 75929 35173 75963 35207
rect 84761 35173 84795 35207
rect 86049 35173 86083 35207
rect 5733 35105 5767 35139
rect 6285 35105 6319 35139
rect 7297 35105 7331 35139
rect 7849 35105 7883 35139
rect 13553 35105 13587 35139
rect 13921 35105 13955 35139
rect 14105 35105 14139 35139
rect 18429 35105 18463 35139
rect 18981 35105 19015 35139
rect 19165 35105 19199 35139
rect 21833 35105 21867 35139
rect 24317 35105 24351 35139
rect 25329 35105 25363 35139
rect 28089 35105 28123 35139
rect 29193 35105 29227 35139
rect 29377 35105 29411 35139
rect 29929 35105 29963 35139
rect 30113 35105 30147 35139
rect 31493 35105 31527 35139
rect 32306 35105 32340 35139
rect 32781 35105 32815 35139
rect 32873 35105 32907 35139
rect 34529 35105 34563 35139
rect 35541 35105 35575 35139
rect 36277 35105 36311 35139
rect 36616 35105 36650 35139
rect 36737 35105 36771 35139
rect 37841 35105 37875 35139
rect 38025 35105 38059 35139
rect 38485 35105 38519 35139
rect 38577 35105 38611 35139
rect 39405 35105 39439 35139
rect 39589 35105 39623 35139
rect 40601 35105 40635 35139
rect 40785 35105 40819 35139
rect 41245 35105 41279 35139
rect 41797 35105 41831 35139
rect 41981 35105 42015 35139
rect 44005 35105 44039 35139
rect 44373 35105 44407 35139
rect 44465 35105 44499 35139
rect 47133 35105 47167 35139
rect 47593 35105 47627 35139
rect 47685 35105 47719 35139
rect 48513 35105 48547 35139
rect 50077 35105 50111 35139
rect 50261 35105 50295 35139
rect 50721 35105 50755 35139
rect 50813 35105 50847 35139
rect 53297 35105 53331 35139
rect 54585 35105 54619 35139
rect 56701 35105 56735 35139
rect 56977 35105 57011 35139
rect 57437 35105 57471 35139
rect 57529 35105 57563 35139
rect 58357 35105 58391 35139
rect 58541 35105 58575 35139
rect 62313 35105 62347 35139
rect 62773 35105 62807 35139
rect 62865 35105 62899 35139
rect 64705 35105 64739 35139
rect 65809 35105 65843 35139
rect 66637 35105 66671 35139
rect 66729 35105 66763 35139
rect 67097 35105 67131 35139
rect 67189 35105 67223 35139
rect 69121 35105 69155 35139
rect 73169 35105 73203 35139
rect 74641 35105 74675 35139
rect 75377 35105 75411 35139
rect 75561 35105 75595 35139
rect 77033 35105 77067 35139
rect 78505 35105 78539 35139
rect 83289 35105 83323 35139
rect 84025 35105 84059 35139
rect 84393 35105 84427 35139
rect 84577 35105 84611 35139
rect 85405 35105 85439 35139
rect 85589 35105 85623 35139
rect 85957 35105 85991 35139
rect 88257 35105 88291 35139
rect 89085 35105 89119 35139
rect 89545 35105 89579 35139
rect 91753 35105 91787 35139
rect 94145 35105 94179 35139
rect 13645 35037 13679 35071
rect 14657 35037 14691 35071
rect 18245 35037 18279 35071
rect 22109 35037 22143 35071
rect 14197 34969 14231 35003
rect 25513 34969 25547 35003
rect 31769 35037 31803 35071
rect 32137 35037 32171 35071
rect 33425 35037 33459 35071
rect 33885 35037 33919 35071
rect 35633 35037 35667 35071
rect 36369 35037 36403 35071
rect 37013 35037 37047 35071
rect 37749 35037 37783 35071
rect 40969 35037 41003 35071
rect 41153 35037 41187 35071
rect 43453 35037 43487 35071
rect 44097 35037 44131 35071
rect 46949 35037 46983 35071
rect 49893 35037 49927 35071
rect 51365 35037 51399 35071
rect 51825 35037 51859 35071
rect 56793 35037 56827 35071
rect 62129 35037 62163 35071
rect 64797 35037 64831 35071
rect 68845 35037 68879 35071
rect 70593 35037 70627 35071
rect 72893 35037 72927 35071
rect 74273 35037 74307 35071
rect 75193 35037 75227 35071
rect 76021 35037 76055 35071
rect 78229 35037 78263 35071
rect 82093 35037 82127 35071
rect 83933 35037 83967 35071
rect 88349 35037 88383 35071
rect 89269 35037 89303 35071
rect 93593 35037 93627 35071
rect 93869 35037 93903 35071
rect 95249 35037 95283 35071
rect 42901 34969 42935 35003
rect 48697 34969 48731 35003
rect 63693 34969 63727 35003
rect 67649 34969 67683 35003
rect 77217 34969 77251 35003
rect 83473 34969 83507 35003
rect 18061 34901 18095 34935
rect 23397 34901 23431 34935
rect 23673 34901 23707 34935
rect 27905 34901 27939 34935
rect 29009 34901 29043 34935
rect 31493 34901 31527 34935
rect 31585 34901 31619 34935
rect 33701 34901 33735 34935
rect 37289 34901 37323 34935
rect 37473 34901 37507 34935
rect 37749 34901 37783 34935
rect 46581 34901 46615 34935
rect 46765 34901 46799 34935
rect 49709 34901 49743 34935
rect 53389 34901 53423 34935
rect 54033 34901 54067 34935
rect 54217 34901 54251 34935
rect 54769 34901 54803 34935
rect 54953 34901 54987 34935
rect 56425 34901 56459 34935
rect 61761 34901 61795 34935
rect 61945 34901 61979 34935
rect 63877 34901 63911 34935
rect 66269 34901 66303 34935
rect 78045 34901 78079 34935
rect 79609 34901 79643 34935
rect 81817 34901 81851 34935
rect 82185 34901 82219 34935
rect 91937 34901 91971 34935
rect 4353 34697 4387 34731
rect 11437 34697 11471 34731
rect 14473 34697 14507 34731
rect 18797 34697 18831 34731
rect 21741 34697 21775 34731
rect 22293 34697 22327 34731
rect 24869 34697 24903 34731
rect 36001 34697 36035 34731
rect 37289 34697 37323 34731
rect 39037 34697 39071 34731
rect 39405 34697 39439 34731
rect 39589 34697 39623 34731
rect 41245 34697 41279 34731
rect 42993 34697 43027 34731
rect 89269 34697 89303 34731
rect 91293 34697 91327 34731
rect 23489 34629 23523 34663
rect 35633 34629 35667 34663
rect 2513 34561 2547 34595
rect 2789 34561 2823 34595
rect 5457 34493 5491 34527
rect 5733 34493 5767 34527
rect 6837 34493 6871 34527
rect 7297 34493 7331 34527
rect 11345 34493 11379 34527
rect 13093 34493 13127 34527
rect 13369 34493 13403 34527
rect 14841 34493 14875 34527
rect 18613 34493 18647 34527
rect 20545 34493 20579 34527
rect 20729 34493 20763 34527
rect 21189 34493 21223 34527
rect 21281 34493 21315 34527
rect 26157 34561 26191 34595
rect 32229 34561 32263 34595
rect 32689 34561 32723 34595
rect 23673 34493 23707 34527
rect 24777 34493 24811 34527
rect 24041 34425 24075 34459
rect 26433 34493 26467 34527
rect 30757 34493 30791 34527
rect 30941 34493 30975 34527
rect 31125 34493 31159 34527
rect 31585 34493 31619 34527
rect 31677 34493 31711 34527
rect 32505 34493 32539 34527
rect 35817 34493 35851 34527
rect 49893 34629 49927 34663
rect 52285 34629 52319 34663
rect 52469 34629 52503 34663
rect 65809 34629 65843 34663
rect 77769 34629 77803 34663
rect 79885 34629 79919 34663
rect 82185 34629 82219 34663
rect 82553 34629 82587 34663
rect 85773 34629 85807 34663
rect 86601 34629 86635 34663
rect 88257 34629 88291 34663
rect 53021 34561 53055 34595
rect 55045 34561 55079 34595
rect 56701 34561 56735 34595
rect 56977 34561 57011 34595
rect 59001 34561 59035 34595
rect 66269 34561 66303 34595
rect 76481 34561 76515 34595
rect 78965 34561 78999 34595
rect 81265 34561 81299 34595
rect 81633 34561 81667 34595
rect 81817 34561 81851 34595
rect 83013 34561 83047 34595
rect 84393 34561 84427 34595
rect 88073 34561 88107 34595
rect 88809 34561 88843 34595
rect 37473 34493 37507 34527
rect 37657 34493 37691 34527
rect 37841 34493 37875 34527
rect 38025 34493 38059 34527
rect 38485 34493 38519 34527
rect 38577 34493 38611 34527
rect 41613 34493 41647 34527
rect 41797 34493 41831 34527
rect 41981 34493 42015 34527
rect 42533 34493 42567 34527
rect 42717 34493 42751 34527
rect 52653 34493 52687 34527
rect 52745 34493 52779 34527
rect 54493 34493 54527 34527
rect 54677 34493 54711 34527
rect 54861 34493 54895 34527
rect 55413 34493 55447 34527
rect 26249 34425 26283 34459
rect 37289 34425 37323 34459
rect 41521 34425 41555 34459
rect 48513 34425 48547 34459
rect 48605 34425 48639 34459
rect 54401 34425 54435 34459
rect 55229 34425 55263 34459
rect 57345 34493 57379 34527
rect 57529 34493 57563 34527
rect 57989 34493 58023 34527
rect 58081 34493 58115 34527
rect 58909 34493 58943 34527
rect 62957 34493 62991 34527
rect 63141 34493 63175 34527
rect 63601 34493 63635 34527
rect 63693 34493 63727 34527
rect 65993 34493 66027 34527
rect 76205 34493 76239 34527
rect 78689 34493 78723 34527
rect 79793 34493 79827 34527
rect 80989 34493 81023 34527
rect 81449 34493 81483 34527
rect 81733 34493 81767 34527
rect 82369 34493 82403 34527
rect 82737 34493 82771 34527
rect 85405 34493 85439 34527
rect 86509 34493 86543 34527
rect 87981 34493 88015 34527
rect 88993 34493 89027 34527
rect 89177 34493 89211 34527
rect 91201 34493 91235 34527
rect 56793 34425 56827 34459
rect 62497 34425 62531 34459
rect 62681 34425 62715 34459
rect 76021 34425 76055 34459
rect 78781 34425 78815 34459
rect 82001 34425 82035 34459
rect 91017 34425 91051 34459
rect 3893 34357 3927 34391
rect 5273 34357 5307 34391
rect 6929 34357 6963 34391
rect 20177 34357 20211 34391
rect 20361 34357 20395 34391
rect 22109 34357 22143 34391
rect 23489 34357 23523 34391
rect 23857 34357 23891 34391
rect 26157 34357 26191 34391
rect 26617 34357 26651 34391
rect 56701 34357 56735 34391
rect 58541 34357 58575 34391
rect 64153 34357 64187 34391
rect 64521 34357 64555 34391
rect 64705 34357 64739 34391
rect 67373 34357 67407 34391
rect 85589 34357 85623 34391
rect 5089 34153 5123 34187
rect 6101 34153 6135 34187
rect 9873 34153 9907 34187
rect 10149 34153 10183 34187
rect 11529 34153 11563 34187
rect 37289 34153 37323 34187
rect 13737 34085 13771 34119
rect 22753 34085 22787 34119
rect 4905 34017 4939 34051
rect 6285 34017 6319 34051
rect 6561 34017 6595 34051
rect 10057 34017 10091 34051
rect 11345 34017 11379 34051
rect 12633 34017 12667 34051
rect 13185 34017 13219 34051
rect 13369 34017 13403 34051
rect 15301 34017 15335 34051
rect 19625 34017 19659 34051
rect 19717 34017 19751 34051
rect 24777 34017 24811 34051
rect 24869 34017 24903 34051
rect 12357 33949 12391 33983
rect 12449 33949 12483 33983
rect 21097 33949 21131 33983
rect 21373 33949 21407 33983
rect 22937 33949 22971 33983
rect 13921 33813 13955 33847
rect 15393 33813 15427 33847
rect 19901 33813 19935 33847
rect 4813 33609 4847 33643
rect 22201 33609 22235 33643
rect 11253 33541 11287 33575
rect 20453 33473 20487 33507
rect 4629 33405 4663 33439
rect 11069 33405 11103 33439
rect 12265 33405 12299 33439
rect 12449 33405 12483 33439
rect 12725 33405 12759 33439
rect 20637 33405 20671 33439
rect 21097 33405 21131 33439
rect 21277 33405 21311 33439
rect 20361 33337 20395 33371
rect 25053 33881 25087 33915
rect 37289 33677 37323 33711
rect 46857 34153 46891 34187
rect 46857 33677 46891 33711
rect 11529 33269 11563 33303
rect 13829 33269 13863 33303
rect 21649 33269 21683 33303
rect 22017 33269 22051 33303
rect 24869 33269 24903 33303
rect 6561 33065 6595 33099
rect 12909 32997 12943 33031
rect 23581 32997 23615 33031
rect 24777 32997 24811 33031
rect 4077 32929 4111 32963
rect 4353 32929 4387 32963
rect 5089 32929 5123 32963
rect 5181 32929 5215 32963
rect 5457 32929 5491 32963
rect 11805 32929 11839 32963
rect 12265 32929 12299 32963
rect 12357 32929 12391 32963
rect 13829 32929 13863 32963
rect 15301 32929 15335 32963
rect 17417 32929 17451 32963
rect 17969 32929 18003 32963
rect 18153 32929 18187 32963
rect 18705 32929 18739 32963
rect 19625 32929 19659 32963
rect 11529 32861 11563 32895
rect 11713 32861 11747 32895
rect 17233 32861 17267 32895
rect 19717 32861 19751 32895
rect 21925 32861 21959 32895
rect 22201 32861 22235 32895
rect 14013 32793 14047 32827
rect 4169 32725 4203 32759
rect 5089 32725 5123 32759
rect 7021 32725 7055 32759
rect 15485 32725 15519 32759
rect 17141 32725 17175 32759
rect 18429 32725 18463 32759
rect 21741 32725 21775 32759
rect 9781 32453 9815 32487
rect 10609 32453 10643 32487
rect 20453 32453 20487 32487
rect 20821 32453 20855 32487
rect 2973 32385 3007 32419
rect 14105 32385 14139 32419
rect 19625 32385 19659 32419
rect 22661 32385 22695 32419
rect 24685 32385 24719 32419
rect 2697 32317 2731 32351
rect 5181 32317 5215 32351
rect 5641 32317 5675 32351
rect 9689 32317 9723 32351
rect 9965 32317 9999 32351
rect 12449 32317 12483 32351
rect 14381 32317 14415 32351
rect 14473 32317 14507 32351
rect 14933 32317 14967 32351
rect 15117 32317 15151 32351
rect 15761 32317 15795 32351
rect 18153 32317 18187 32351
rect 18423 32317 18457 32351
rect 20637 32317 20671 32351
rect 22569 32317 22603 32351
rect 25145 32861 25179 32895
rect 24777 32317 24811 32351
rect 25053 32793 25087 32827
rect 4537 32249 4571 32283
rect 6101 32249 6135 32283
rect 24961 32249 24995 32283
rect 4077 32181 4111 32215
rect 5457 32181 5491 32215
rect 10149 32181 10183 32215
rect 12633 32181 12667 32215
rect 15393 32181 15427 32215
rect 19993 32181 20027 32215
rect 5825 31977 5859 32011
rect 10885 31977 10919 32011
rect 13737 31977 13771 32011
rect 14013 31977 14047 32011
rect 15669 31977 15703 32011
rect 16497 31977 16531 32011
rect 17785 31977 17819 32011
rect 21741 31977 21775 32011
rect 3341 31909 3375 31943
rect 9689 31909 9723 31943
rect 2697 31841 2731 31875
rect 2973 31841 3007 31875
rect 4077 31841 4111 31875
rect 4629 31841 4663 31875
rect 4813 31841 4847 31875
rect 5641 31841 5675 31875
rect 8585 31841 8619 31875
rect 10241 31841 10275 31875
rect 10517 31841 10551 31875
rect 13553 31841 13587 31875
rect 15485 31841 15519 31875
rect 16589 31841 16623 31875
rect 17693 31841 17727 31875
rect 21925 31841 21959 31875
rect 22201 31841 22235 31875
rect 25053 31841 25087 31875
rect 3157 31773 3191 31807
rect 4905 31773 4939 31807
rect 10701 31773 10735 31807
rect 15393 31773 15427 31807
rect 18061 31773 18095 31807
rect 37289 32657 37323 32691
rect 26893 32453 26927 32487
rect 8677 31637 8711 31671
rect 15393 31637 15427 31671
rect 16773 31637 16807 31671
rect 23489 31637 23523 31671
rect 25145 31637 25179 31671
rect 25973 32317 26007 32351
rect 4445 31433 4479 31467
rect 6009 31433 6043 31467
rect 11713 31433 11747 31467
rect 16957 31365 16991 31399
rect 21557 31365 21591 31399
rect 22661 31365 22695 31399
rect 22937 31365 22971 31399
rect 8769 31297 8803 31331
rect 14657 31297 14691 31331
rect 24777 31297 24811 31331
rect 2421 31229 2455 31263
rect 3801 31229 3835 31263
rect 4077 31229 4111 31263
rect 5089 31229 5123 31263
rect 5641 31229 5675 31263
rect 8493 31229 8527 31263
rect 10241 31229 10275 31263
rect 11161 31229 11195 31263
rect 14381 31229 14415 31263
rect 16865 31229 16899 31263
rect 19717 31229 19751 31263
rect 19993 31229 20027 31263
rect 20177 31229 20211 31263
rect 20637 31229 20671 31263
rect 20729 31229 20763 31263
rect 22569 31229 22603 31263
rect 10149 31161 10183 31195
rect 10977 31161 11011 31195
rect 11529 31161 11563 31195
rect 21281 31161 21315 31195
rect 2605 31093 2639 31127
rect 3801 31093 3835 31127
rect 5181 31093 5215 31127
rect 15761 31093 15795 31127
rect 16221 31093 16255 31127
rect 19717 31093 19751 31127
rect 19901 31093 19935 31127
rect 4169 30889 4203 30923
rect 4997 30889 5031 30923
rect 14289 30889 14323 30923
rect 22385 30889 22419 30923
rect 22661 30889 22695 30923
rect 12081 30821 12115 30855
rect 4077 30753 4111 30787
rect 4629 30753 4663 30787
rect 9689 30753 9723 30787
rect 9781 30753 9815 30787
rect 11713 30753 11747 30787
rect 14197 30753 14231 30787
rect 21373 30753 21407 30787
rect 21925 30753 21959 30787
rect 22109 30753 22143 30787
rect 9965 30685 9999 30719
rect 10885 30685 10919 30719
rect 11437 30685 11471 30719
rect 11897 30685 11931 30719
rect 16221 30685 16255 30719
rect 16497 30685 16531 30719
rect 21189 30685 21223 30719
rect 16037 30549 16071 30583
rect 17601 30549 17635 30583
rect 21005 30549 21039 30583
rect 12541 30345 12575 30379
rect 16497 30345 16531 30379
rect 37289 32385 37323 32419
rect 46857 32657 46891 32691
rect 46857 32385 46891 32419
rect 26893 31841 26927 31875
rect 41429 31161 41463 31195
rect 41337 31093 41371 31127
rect 25973 30685 26007 30719
rect 6009 30277 6043 30311
rect 9321 30277 9355 30311
rect 10885 30277 10919 30311
rect 11713 30277 11747 30311
rect 16865 30277 16899 30311
rect 22569 30277 22603 30311
rect 24777 30277 24811 30311
rect 21373 30209 21407 30243
rect 22293 30209 22327 30243
rect 3801 30141 3835 30175
rect 4077 30141 4111 30175
rect 5089 30141 5123 30175
rect 5641 30141 5675 30175
rect 9229 30141 9263 30175
rect 10793 30141 10827 30175
rect 11069 30141 11103 30175
rect 12449 30141 12483 30175
rect 12725 30141 12759 30175
rect 15301 30141 15335 30175
rect 15485 30141 15519 30175
rect 16037 30141 16071 30175
rect 16221 30141 16255 30175
rect 19993 30141 20027 30175
rect 20269 30141 20303 30175
rect 22477 30141 22511 30175
rect 4445 30073 4479 30107
rect 3617 30005 3651 30039
rect 5181 30005 5215 30039
rect 9505 30005 9539 30039
rect 11253 30005 11287 30039
rect 15209 30005 15243 30039
rect 19901 30005 19935 30039
rect 3341 29801 3375 29835
rect 8953 29801 8987 29835
rect 16497 29801 16531 29835
rect 22109 29801 22143 29835
rect 22477 29801 22511 29835
rect 2697 29665 2731 29699
rect 2881 29665 2915 29699
rect 4077 29665 4111 29699
rect 5825 29665 5859 29699
rect 7573 29665 7607 29699
rect 8125 29665 8159 29699
rect 8309 29665 8343 29699
rect 11621 29665 11655 29699
rect 14933 29665 14967 29699
rect 15301 29665 15335 29699
rect 15485 29665 15519 29699
rect 16037 29665 16071 29699
rect 16221 29665 16255 29699
rect 16773 29665 16807 29699
rect 21097 29665 21131 29699
rect 21649 29665 21683 29699
rect 21833 29665 21867 29699
rect 2973 29597 3007 29631
rect 4353 29597 4387 29631
rect 7481 29597 7515 29631
rect 9873 29597 9907 29631
rect 10149 29597 10183 29631
rect 20913 29597 20947 29631
rect 8493 29529 8527 29563
rect 5457 29461 5491 29495
rect 7297 29461 7331 29495
rect 11437 29461 11471 29495
rect 14749 29461 14783 29495
rect 15025 29461 15059 29495
rect 20729 29461 20763 29495
rect 10793 29257 10827 29291
rect 15117 29257 15151 29291
rect 2513 29121 2547 29155
rect 4261 29121 4295 29155
rect 8217 29121 8251 29155
rect 8493 29121 8527 29155
rect 9597 29121 9631 29155
rect 19441 29121 19475 29155
rect 21649 29121 21683 29155
rect 2789 29053 2823 29087
rect 9965 29053 9999 29087
rect 10701 29053 10735 29087
rect 13461 29053 13495 29087
rect 13553 29053 13587 29087
rect 13737 29053 13771 29087
rect 14289 29053 14323 29087
rect 14473 29053 14507 29087
rect 19165 29053 19199 29087
rect 19533 29053 19567 29087
rect 20085 29053 20119 29087
rect 20269 29053 20303 29087
rect 21557 29053 21591 29087
rect 22569 29053 22603 29087
rect 20637 28985 20671 29019
rect 3893 28917 3927 28951
rect 14749 28917 14783 28951
rect 22661 28917 22695 28951
rect 4169 28713 4203 28747
rect 4997 28713 5031 28747
rect 15393 28713 15427 28747
rect 19809 28713 19843 28747
rect 4353 28577 4387 28611
rect 4629 28577 4663 28611
rect 12909 28577 12943 28611
rect 14197 28577 14231 28611
rect 15301 28577 15335 28611
rect 16589 28577 16623 28611
rect 18797 28577 18831 28611
rect 19349 28577 19383 28611
rect 19533 28577 19567 28611
rect 21281 28577 21315 28611
rect 12817 28509 12851 28543
rect 18613 28509 18647 28543
rect 21005 28509 21039 28543
rect 22569 28509 22603 28543
rect 14013 28441 14047 28475
rect 13093 28373 13127 28407
rect 14289 28373 14323 28407
rect 16405 28373 16439 28407
rect 18429 28373 18463 28407
rect 20637 28373 20671 28407
rect 54125 28373 54159 28407
rect 21833 28169 21867 28203
rect 18797 28101 18831 28135
rect 20177 28101 20211 28135
rect 2513 28033 2547 28067
rect 8401 28033 8435 28067
rect 13829 28033 13863 28067
rect 20729 28033 20763 28067
rect 2789 27965 2823 27999
rect 7941 27965 7975 27999
rect 8033 27965 8067 27999
rect 8309 27965 8343 27999
rect 11253 27965 11287 27999
rect 13553 27965 13587 27999
rect 15301 27965 15335 27999
rect 18981 27965 19015 27999
rect 20177 27965 20211 27999
rect 20453 27965 20487 27999
rect 7297 27897 7331 27931
rect 3893 27829 3927 27863
rect 4353 27829 4387 27863
rect 11437 27829 11471 27863
rect 14933 27829 14967 27863
rect 20361 27829 20395 27863
rect 12541 27557 12575 27591
rect 15669 27557 15703 27591
rect 7113 27489 7147 27523
rect 7665 27489 7699 27523
rect 7840 27489 7874 27523
rect 8493 27489 8527 27523
rect 9689 27489 9723 27523
rect 9781 27489 9815 27523
rect 14381 27489 14415 27523
rect 15301 27489 15335 27523
rect 16313 27489 16347 27523
rect 16497 27489 16531 27523
rect 16681 27489 16715 27523
rect 17233 27489 17267 27523
rect 17417 27489 17451 27523
rect 6929 27421 6963 27455
rect 12725 27421 12759 27455
rect 13001 27421 13035 27455
rect 21649 27421 21683 27455
rect 21925 27421 21959 27455
rect 8033 27353 8067 27387
rect 6745 27285 6779 27319
rect 15393 27285 15427 27319
rect 17693 27285 17727 27319
rect 21465 27285 21499 27319
rect 23213 27285 23247 27319
rect 4353 27013 4387 27047
rect 13553 27013 13587 27047
rect 18337 27013 18371 27047
rect 2513 26945 2547 26979
rect 2789 26945 2823 26979
rect 7113 26945 7147 26979
rect 12265 26945 12299 26979
rect 12449 26945 12483 26979
rect 21189 26945 21223 26979
rect 5733 26877 5767 26911
rect 6837 26877 6871 26911
rect 12587 26877 12621 26911
rect 13093 26877 13127 26911
rect 13185 26877 13219 26911
rect 18245 26877 18279 26911
rect 19901 26877 19935 26911
rect 20085 26877 20119 26911
rect 20637 26877 20671 26911
rect 20821 26877 20855 26911
rect 3893 26741 3927 26775
rect 5825 26741 5859 26775
rect 8401 26741 8435 26775
rect 8585 26741 8619 26775
rect 19809 26741 19843 26775
rect 21465 26741 21499 26775
rect 10793 26537 10827 26571
rect 11713 26537 11747 26571
rect 8309 26469 8343 26503
rect 12817 26469 12851 26503
rect 15393 26469 15427 26503
rect 19257 26469 19291 26503
rect 6745 26401 6779 26435
rect 10609 26401 10643 26435
rect 11897 26401 11931 26435
rect 13001 26401 13035 26435
rect 13185 26401 13219 26435
rect 13737 26401 13771 26435
rect 13921 26401 13955 26435
rect 15301 26401 15335 26435
rect 17877 26401 17911 26435
rect 20913 26401 20947 26435
rect 23213 26401 23247 26435
rect 23305 26401 23339 26435
rect 6469 26333 6503 26367
rect 17601 26333 17635 26367
rect 19441 26333 19475 26367
rect 10425 26265 10459 26299
rect 14105 26265 14139 26299
rect 8033 26197 8067 26231
rect 21097 26197 21131 26231
rect 13369 25993 13403 26027
rect 15117 25993 15151 26027
rect 4353 25925 4387 25959
rect 12633 25925 12667 25959
rect 2789 25857 2823 25891
rect 13553 25857 13587 25891
rect 13829 25857 13863 25891
rect 2513 25789 2547 25823
rect 7941 25789 7975 25823
rect 8125 25789 8159 25823
rect 12449 25789 12483 25823
rect 19625 25789 19659 25823
rect 19901 25789 19935 25823
rect 3893 25653 3927 25687
rect 7941 25653 7975 25687
rect 8585 25653 8619 25687
rect 19533 25653 19567 25687
rect 21005 25653 21039 25687
rect 7389 25381 7423 25415
rect 12817 25381 12851 25415
rect 13553 25381 13587 25415
rect 19625 25381 19659 25415
rect 11713 25313 11747 25347
rect 11897 25313 11931 25347
rect 13001 25313 13035 25347
rect 13185 25313 13219 25347
rect 14565 25313 14599 25347
rect 18521 25313 18555 25347
rect 19073 25313 19107 25347
rect 19257 25313 19291 25347
rect 21097 25313 21131 25347
rect 21649 25313 21683 25347
rect 21833 25313 21867 25347
rect 5733 25245 5767 25279
rect 6009 25245 6043 25279
rect 11989 25245 12023 25279
rect 18245 25245 18279 25279
rect 18337 25245 18371 25279
rect 20913 25245 20947 25279
rect 12265 25177 12299 25211
rect 14381 25177 14415 25211
rect 7573 25109 7607 25143
rect 20729 25109 20763 25143
rect 22109 25109 22143 25143
rect 2789 24769 2823 24803
rect 4353 24769 4387 24803
rect 6837 24769 6871 24803
rect 8493 24769 8527 24803
rect 21373 24769 21407 24803
rect 2513 24701 2547 24735
rect 4537 24701 4571 24735
rect 7113 24701 7147 24735
rect 11437 24701 11471 24735
rect 12449 24701 12483 24735
rect 13553 24701 13587 24735
rect 15301 24701 15335 24735
rect 15669 24701 15703 24735
rect 19349 24701 19383 24735
rect 21097 24701 21131 24735
rect 13461 24633 13495 24667
rect 22753 24633 22787 24667
rect 3893 24565 3927 24599
rect 8677 24565 8711 24599
rect 11253 24565 11287 24599
rect 12541 24565 12575 24599
rect 12725 24565 12759 24599
rect 13737 24565 13771 24599
rect 15393 24565 15427 24599
rect 19257 24565 19291 24599
rect 19533 24565 19567 24599
rect 20913 24565 20947 24599
rect 6469 24361 6503 24395
rect 7389 24361 7423 24395
rect 19533 24361 19567 24395
rect 21005 24361 21039 24395
rect 22017 24361 22051 24395
rect 7573 24293 7607 24327
rect 5457 24225 5491 24259
rect 6009 24225 6043 24259
rect 6193 24225 6227 24259
rect 7481 24225 7515 24259
rect 10885 24225 10919 24259
rect 17785 24225 17819 24259
rect 18061 24225 18095 24259
rect 18797 24225 18831 24259
rect 19165 24225 19199 24259
rect 19349 24225 19383 24259
rect 20913 24225 20947 24259
rect 21925 24225 21959 24259
rect 23121 24225 23155 24259
rect 23397 24225 23431 24259
rect 5181 24157 5215 24191
rect 5365 24157 5399 24191
rect 11161 24157 11195 24191
rect 15301 24157 15335 24191
rect 15577 24157 15611 24191
rect 16681 24157 16715 24191
rect 18153 24157 18187 24191
rect 18889 24157 18923 24191
rect 22937 24089 22971 24123
rect 12449 24021 12483 24055
rect 12725 24021 12759 24055
rect 15025 24021 15059 24055
rect 23489 24021 23523 24055
rect 7665 23817 7699 23851
rect 12633 23817 12667 23851
rect 14933 23817 14967 23851
rect 21189 23817 21223 23851
rect 10057 23749 10091 23783
rect 2789 23681 2823 23715
rect 10241 23681 10275 23715
rect 11345 23681 11379 23715
rect 13553 23681 13587 23715
rect 13737 23681 13771 23715
rect 18061 23681 18095 23715
rect 21373 23681 21407 23715
rect 2513 23613 2547 23647
rect 7297 23613 7331 23647
rect 10333 23613 10367 23647
rect 10885 23613 10919 23647
rect 11069 23613 11103 23647
rect 12449 23613 12483 23647
rect 13921 23613 13955 23647
rect 14473 23613 14507 23647
rect 14657 23613 14691 23647
rect 18245 23613 18279 23647
rect 18797 23613 18831 23647
rect 18981 23613 19015 23647
rect 20269 23613 20303 23647
rect 21557 23613 21591 23647
rect 22109 23613 22143 23647
rect 22293 23613 22327 23647
rect 20361 23545 20395 23579
rect 3893 23477 3927 23511
rect 4353 23477 4387 23511
rect 7389 23477 7423 23511
rect 17785 23477 17819 23511
rect 19257 23477 19291 23511
rect 20177 23477 20211 23511
rect 22569 23477 22603 23511
rect 6745 23205 6779 23239
rect 11713 23205 11747 23239
rect 19717 23205 19751 23239
rect 5641 23137 5675 23171
rect 6193 23137 6227 23171
rect 6377 23137 6411 23171
rect 7665 23137 7699 23171
rect 9689 23137 9723 23171
rect 12449 23137 12483 23171
rect 12817 23137 12851 23171
rect 13001 23137 13035 23171
rect 18337 23137 18371 23171
rect 22201 23137 22235 23171
rect 5365 23069 5399 23103
rect 5549 23069 5583 23103
rect 12541 23069 12575 23103
rect 18061 23069 18095 23103
rect 19901 23069 19935 23103
rect 21741 23069 21775 23103
rect 21925 23069 21959 23103
rect 7849 22933 7883 22967
rect 9781 22933 9815 22967
rect 12081 22933 12115 22967
rect 23489 22933 23523 22967
rect 3893 22729 3927 22763
rect 4537 22729 4571 22763
rect 9045 22729 9079 22763
rect 9689 22729 9723 22763
rect 13829 22729 13863 22763
rect 7297 22593 7331 22627
rect 13185 22593 13219 22627
rect 19533 22593 19567 22627
rect 19625 22593 19659 22627
rect 2513 22525 2547 22559
rect 2789 22525 2823 22559
rect 7573 22525 7607 22559
rect 8953 22525 8987 22559
rect 9781 22525 9815 22559
rect 13093 22525 13127 22559
rect 13461 22525 13495 22559
rect 13645 22525 13679 22559
rect 19901 22525 19935 22559
rect 4353 22457 4387 22491
rect 12449 22457 12483 22491
rect 21281 22457 21315 22491
rect 9873 22389 9907 22423
rect 12265 22389 12299 22423
rect 7941 22185 7975 22219
rect 12449 22185 12483 22219
rect 18337 22185 18371 22219
rect 19993 22185 20027 22219
rect 21281 22117 21315 22151
rect 4077 22049 4111 22083
rect 4353 22049 4387 22083
rect 5825 22049 5859 22083
rect 6929 22049 6963 22083
rect 7481 22049 7515 22083
rect 7665 22049 7699 22083
rect 9689 22049 9723 22083
rect 11529 22049 11563 22083
rect 13001 22049 13035 22083
rect 13185 22049 13219 22083
rect 13461 22049 13495 22083
rect 14013 22049 14047 22083
rect 17325 22049 17359 22083
rect 18521 22049 18555 22083
rect 19257 22049 19291 22083
rect 19625 22049 19659 22083
rect 19809 22049 19843 22083
rect 20913 22049 20947 22083
rect 24041 22049 24075 22083
rect 24317 22049 24351 22083
rect 6745 21981 6779 22015
rect 12541 21981 12575 22015
rect 13737 21981 13771 22015
rect 18613 21981 18647 22015
rect 19165 21981 19199 22015
rect 21005 21981 21039 22015
rect 9873 21913 9907 21947
rect 5457 21845 5491 21879
rect 6653 21845 6687 21879
rect 11621 21845 11655 21879
rect 12265 21845 12299 21879
rect 14197 21845 14231 21879
rect 17509 21845 17543 21879
rect 24133 21845 24167 21879
rect 4353 21641 4387 21675
rect 9321 21641 9355 21675
rect 19625 21641 19659 21675
rect 4537 21573 4571 21607
rect 12265 21573 12299 21607
rect 14013 21573 14047 21607
rect 2789 21505 2823 21539
rect 7941 21505 7975 21539
rect 12449 21505 12483 21539
rect 12725 21505 12759 21539
rect 2513 21437 2547 21471
rect 6837 21437 6871 21471
rect 8033 21437 8067 21471
rect 9137 21437 9171 21471
rect 18429 21437 18463 21471
rect 18613 21437 18647 21471
rect 19073 21437 19107 21471
rect 19165 21437 19199 21471
rect 22201 21437 22235 21471
rect 3893 21301 3927 21335
rect 7021 21301 7055 21335
rect 7941 21301 7975 21335
rect 8217 21301 8251 21335
rect 18337 21301 18371 21335
rect 22293 21301 22327 21335
rect 22569 21301 22603 21335
rect 7389 21097 7423 21131
rect 23029 21097 23063 21131
rect 7021 21029 7055 21063
rect 7481 21029 7515 21063
rect 7849 21029 7883 21063
rect 7297 20961 7331 20995
rect 15301 20961 15335 20995
rect 21557 20961 21591 20995
rect 21649 20961 21683 20995
rect 7113 20893 7147 20927
rect 12725 20893 12759 20927
rect 13001 20893 13035 20927
rect 14381 20893 14415 20927
rect 21925 20893 21959 20927
rect 15485 20825 15519 20859
rect 12633 20757 12667 20791
rect 4353 20553 4387 20587
rect 8217 20553 8251 20587
rect 15393 20553 15427 20587
rect 19717 20553 19751 20587
rect 19901 20553 19935 20587
rect 22753 20553 22787 20587
rect 2513 20417 2547 20451
rect 2789 20417 2823 20451
rect 13737 20417 13771 20451
rect 13829 20417 13863 20451
rect 20177 20417 20211 20451
rect 6929 20349 6963 20383
rect 7481 20349 7515 20383
rect 7849 20349 7883 20383
rect 14105 20349 14139 20383
rect 20361 20349 20395 20383
rect 20821 20349 20855 20383
rect 20913 20349 20947 20383
rect 22385 20349 22419 20383
rect 8033 20281 8067 20315
rect 22477 20281 22511 20315
rect 3893 20213 3927 20247
rect 8401 20213 8435 20247
rect 19993 20213 20027 20247
rect 21373 20213 21407 20247
rect 6193 20009 6227 20043
rect 8125 20009 8159 20043
rect 14565 20009 14599 20043
rect 22569 20009 22603 20043
rect 5641 19941 5675 19975
rect 6009 19941 6043 19975
rect 12909 19941 12943 19975
rect 5457 19873 5491 19907
rect 5549 19873 5583 19907
rect 7021 19873 7055 19907
rect 7389 19873 7423 19907
rect 7757 19873 7791 19907
rect 13369 19873 13403 19907
rect 13645 19873 13679 19907
rect 13829 19873 13863 19907
rect 14105 19873 14139 19907
rect 14381 19873 14415 19907
rect 15301 19873 15335 19907
rect 21281 19873 21315 19907
rect 5273 19805 5307 19839
rect 7849 19805 7883 19839
rect 12633 19805 12667 19839
rect 20729 19805 20763 19839
rect 21005 19805 21039 19839
rect 8217 19669 8251 19703
rect 12725 19669 12759 19703
rect 15485 19669 15519 19703
rect 15209 19465 15243 19499
rect 19993 19465 20027 19499
rect 20085 19465 20119 19499
rect 21649 19465 21683 19499
rect 15669 19397 15703 19431
rect 9321 19329 9355 19363
rect 10885 19329 10919 19363
rect 14933 19329 14967 19363
rect 20453 19329 20487 19363
rect 54125 19329 54159 19363
rect 8769 19261 8803 19295
rect 8937 19261 8971 19295
rect 9413 19261 9447 19295
rect 12449 19261 12483 19295
rect 12817 19261 12851 19295
rect 13553 19261 13587 19295
rect 14105 19261 14139 19295
rect 14197 19261 14231 19295
rect 14381 19261 14415 19295
rect 14841 19261 14875 19295
rect 15853 19261 15887 19295
rect 15945 19261 15979 19295
rect 18061 19261 18095 19295
rect 20637 19261 20671 19295
rect 21189 19261 21223 19295
rect 21373 19261 21407 19295
rect 7021 19193 7055 19227
rect 7297 19193 7331 19227
rect 7389 19193 7423 19227
rect 7757 19193 7791 19227
rect 8585 19193 8619 19227
rect 10149 19193 10183 19227
rect 10425 19193 10459 19227
rect 10517 19193 10551 19227
rect 13277 19193 13311 19227
rect 16405 19193 16439 19227
rect 20269 19193 20303 19227
rect 7205 19125 7239 19159
rect 8861 19125 8895 19159
rect 10333 19125 10367 19159
rect 12633 19125 12667 19159
rect 13461 19125 13495 19159
rect 18153 19125 18187 19159
rect 5733 18853 5767 18887
rect 6101 18853 6135 18887
rect 8953 18853 8987 18887
rect 18613 18853 18647 18887
rect 5917 18785 5951 18819
rect 6009 18785 6043 18819
rect 7665 18785 7699 18819
rect 7849 18785 7883 18819
rect 8125 18785 8159 18819
rect 8309 18785 8343 18819
rect 13461 18785 13495 18819
rect 13645 18785 13679 18819
rect 13829 18785 13863 18819
rect 14013 18785 14047 18819
rect 14381 18785 14415 18819
rect 15393 18785 15427 18819
rect 17969 18785 18003 18819
rect 18061 18785 18095 18819
rect 6469 18717 6503 18751
rect 7297 18717 7331 18751
rect 12909 18717 12943 18751
rect 15301 18717 15335 18751
rect 15945 18717 15979 18751
rect 21833 18717 21867 18751
rect 21925 18717 21959 18751
rect 22201 18717 22235 18751
rect 8677 18581 8711 18615
rect 9137 18581 9171 18615
rect 14473 18581 14507 18615
rect 15577 18581 15611 18615
rect 18245 18581 18279 18615
rect 23489 18581 23523 18615
rect 24777 18581 24811 18615
rect 4353 18377 4387 18411
rect 5825 18377 5859 18411
rect 9045 18377 9079 18411
rect 10977 18377 11011 18411
rect 16129 18377 16163 18411
rect 16221 18377 16255 18411
rect 18705 18377 18739 18411
rect 22201 18377 22235 18411
rect 18797 18309 18831 18343
rect 2513 18241 2547 18275
rect 7481 18241 7515 18275
rect 13277 18241 13311 18275
rect 16129 18241 16163 18275
rect 16405 18241 16439 18275
rect 19717 18241 19751 18275
rect 2789 18173 2823 18207
rect 5641 18173 5675 18207
rect 7849 18173 7883 18207
rect 8033 18173 8067 18207
rect 8217 18173 8251 18207
rect 8493 18173 8527 18207
rect 10793 18173 10827 18207
rect 13829 18173 13863 18207
rect 13921 18173 13955 18207
rect 14105 18173 14139 18207
rect 14565 18173 14599 18207
rect 14749 18173 14783 18207
rect 16497 18173 16531 18207
rect 19625 18173 19659 18207
rect 19947 18173 19981 18207
rect 20177 18173 20211 18207
rect 21005 18173 21039 18207
rect 21189 18173 21223 18207
rect 21649 18173 21683 18207
rect 21741 18173 21775 18207
rect 8953 18105 8987 18139
rect 16957 18105 16991 18139
rect 3893 18037 3927 18071
rect 4537 18037 4571 18071
rect 9321 18037 9355 18071
rect 14933 18037 14967 18071
rect 19257 18037 19291 18071
rect 20821 18037 20855 18071
rect 24777 17969 24811 18003
rect 22845 17833 22879 17867
rect 23121 17833 23155 17867
rect 4353 17697 4387 17731
rect 5457 17697 5491 17731
rect 6561 17697 6595 17731
rect 6837 17697 6871 17731
rect 8217 17697 8251 17731
rect 13093 17697 13127 17731
rect 18245 17697 18279 17731
rect 19533 17697 19567 17731
rect 22753 17697 22787 17731
rect 7297 17629 7331 17663
rect 8125 17629 8159 17663
rect 18153 17629 18187 17663
rect 18797 17629 18831 17663
rect 4537 17561 4571 17595
rect 6653 17561 6687 17595
rect 19625 17561 19659 17595
rect 5641 17493 5675 17527
rect 8401 17493 8435 17527
rect 13185 17493 13219 17527
rect 18429 17493 18463 17527
rect 4077 17289 4111 17323
rect 19441 17289 19475 17323
rect 19993 17289 20027 17323
rect 20177 17289 20211 17323
rect 15853 17221 15887 17255
rect 19901 17221 19935 17255
rect 23305 17221 23339 17255
rect 5733 17153 5767 17187
rect 7941 17153 7975 17187
rect 14197 17153 14231 17187
rect 18061 17153 18095 17187
rect 20821 17153 20855 17187
rect 2881 17085 2915 17119
rect 3893 17085 3927 17119
rect 4997 17085 5031 17119
rect 5089 17085 5123 17119
rect 5273 17085 5307 17119
rect 7297 17085 7331 17119
rect 7481 17085 7515 17119
rect 7665 17085 7699 17119
rect 8309 17085 8343 17119
rect 9137 17085 9171 17119
rect 10977 17085 11011 17119
rect 11110 17085 11144 17119
rect 14565 17085 14599 17119
rect 14749 17085 14783 17119
rect 15025 17085 15059 17119
rect 15209 17085 15243 17119
rect 16957 17085 16991 17119
rect 18245 17085 18279 17119
rect 18613 17085 18647 17119
rect 18889 17085 18923 17119
rect 19073 17085 19107 17119
rect 20361 17085 20395 17119
rect 21005 17085 21039 17119
rect 21373 17085 21407 17119
rect 21557 17085 21591 17119
rect 23489 17085 23523 17119
rect 2973 17017 3007 17051
rect 6837 17017 6871 17051
rect 11529 17017 11563 17051
rect 2789 16949 2823 16983
rect 4813 16949 4847 16983
rect 9321 16949 9355 16983
rect 10885 16949 10919 16983
rect 15577 16949 15611 16983
rect 17049 16949 17083 16983
rect 19625 16949 19659 16983
rect 3065 16745 3099 16779
rect 22661 16745 22695 16779
rect 7205 16677 7239 16711
rect 10333 16677 10367 16711
rect 2881 16609 2915 16643
rect 2973 16609 3007 16643
rect 4537 16609 4571 16643
rect 4905 16609 4939 16643
rect 4997 16609 5031 16643
rect 5181 16609 5215 16643
rect 6469 16609 6503 16643
rect 6561 16609 6595 16643
rect 6745 16609 6779 16643
rect 7849 16609 7883 16643
rect 8033 16609 8067 16643
rect 10149 16609 10183 16643
rect 10241 16609 10275 16643
rect 11437 16609 11471 16643
rect 11584 16609 11618 16643
rect 13093 16609 13127 16643
rect 16681 16609 16715 16643
rect 16957 16609 16991 16643
rect 17233 16609 17267 16643
rect 17417 16609 17451 16643
rect 17601 16609 17635 16643
rect 18521 16609 18555 16643
rect 18981 16609 19015 16643
rect 22569 16609 22603 16643
rect 22845 16609 22879 16643
rect 5549 16541 5583 16575
rect 11805 16541 11839 16575
rect 11897 16541 11931 16575
rect 13001 16541 13035 16575
rect 13553 16541 13587 16575
rect 17969 16541 18003 16575
rect 8217 16473 8251 16507
rect 11713 16473 11747 16507
rect 4813 16405 4847 16439
rect 18245 16405 18279 16439
rect 19165 16405 19199 16439
rect 5181 16201 5215 16235
rect 20729 16201 20763 16235
rect 7113 16133 7147 16167
rect 9781 16065 9815 16099
rect 10793 16065 10827 16099
rect 18061 16065 18095 16099
rect 20913 16065 20947 16099
rect 2513 15997 2547 16031
rect 2789 15997 2823 16031
rect 4261 15997 4295 16031
rect 4997 15997 5031 16031
rect 7021 15997 7055 16031
rect 7297 15997 7331 16031
rect 10149 15997 10183 16031
rect 10425 15997 10459 16031
rect 12449 15997 12483 16031
rect 12541 15997 12575 16031
rect 18429 15997 18463 16031
rect 18613 15997 18647 16031
rect 18797 15997 18831 16031
rect 18981 15997 19015 16031
rect 21097 15997 21131 16031
rect 21557 15997 21591 16031
rect 21649 15997 21683 16031
rect 4905 15929 4939 15963
rect 7757 15929 7791 15963
rect 10701 15929 10735 15963
rect 13001 15929 13035 15963
rect 19717 15929 19751 15963
rect 22201 15929 22235 15963
rect 3893 15861 3927 15895
rect 4537 15861 4571 15895
rect 13185 15861 13219 15895
rect 19441 15861 19475 15895
rect 5457 15657 5491 15691
rect 8677 15657 8711 15691
rect 13921 15657 13955 15691
rect 15117 15657 15151 15691
rect 21741 15657 21775 15691
rect 3801 15589 3835 15623
rect 7941 15589 7975 15623
rect 13001 15589 13035 15623
rect 18061 15589 18095 15623
rect 23581 15589 23615 15623
rect 4353 15521 4387 15555
rect 6377 15521 6411 15555
rect 6561 15521 6595 15555
rect 8125 15521 8159 15555
rect 9965 15521 9999 15555
rect 10057 15521 10091 15555
rect 11621 15521 11655 15555
rect 11989 15521 12023 15555
rect 16037 15521 16071 15555
rect 16129 15521 16163 15555
rect 16405 15521 16439 15555
rect 16589 15521 16623 15555
rect 16681 15521 16715 15555
rect 17969 15521 18003 15555
rect 19533 15521 19567 15555
rect 21925 15521 21959 15555
rect 22201 15521 22235 15555
rect 4077 15453 4111 15487
rect 8401 15453 8435 15487
rect 11529 15453 11563 15487
rect 12081 15453 12115 15487
rect 13148 15453 13182 15487
rect 13369 15453 13403 15487
rect 15393 15453 15427 15487
rect 11069 15385 11103 15419
rect 13461 15385 13495 15419
rect 5825 15317 5859 15351
rect 6745 15317 6779 15351
rect 13277 15317 13311 15351
rect 19625 15317 19659 15351
rect 19901 15317 19935 15351
rect 5365 15113 5399 15147
rect 8401 15113 8435 15147
rect 11161 15113 11195 15147
rect 21925 15113 21959 15147
rect 4353 15045 4387 15079
rect 13277 15045 13311 15079
rect 2513 14977 2547 15011
rect 2789 14977 2823 15011
rect 4537 14977 4571 15011
rect 14749 14977 14783 15011
rect 14933 14977 14967 15011
rect 20269 14977 20303 15011
rect 20361 14977 20395 15011
rect 5181 14909 5215 14943
rect 7665 14909 7699 14943
rect 7941 14909 7975 14943
rect 8217 14909 8251 14943
rect 10425 14909 10459 14943
rect 10609 14909 10643 14943
rect 13461 14909 13495 14943
rect 13553 14909 13587 14943
rect 15117 14909 15151 14943
rect 15577 14909 15611 14943
rect 15669 14909 15703 14943
rect 20637 14909 20671 14943
rect 8125 14841 8159 14875
rect 3893 14773 3927 14807
rect 4997 14773 5031 14807
rect 7665 14773 7699 14807
rect 7757 14773 7791 14807
rect 10701 14773 10735 14807
rect 13737 14773 13771 14807
rect 16129 14773 16163 14807
rect 5549 14569 5583 14603
rect 10241 14569 10275 14603
rect 14289 14569 14323 14603
rect 15761 14569 15795 14603
rect 17233 14569 17267 14603
rect 18337 14569 18371 14603
rect 18429 14569 18463 14603
rect 10609 14501 10643 14535
rect 13001 14501 13035 14535
rect 14565 14501 14599 14535
rect 5457 14433 5491 14467
rect 8585 14433 8619 14467
rect 10425 14433 10459 14467
rect 10701 14433 10735 14467
rect 12541 14433 12575 14467
rect 14197 14433 14231 14467
rect 16129 14433 16163 14467
rect 19901 14501 19935 14535
rect 18797 14433 18831 14467
rect 19349 14433 19383 14467
rect 19533 14433 19567 14467
rect 22753 14433 22787 14467
rect 12449 14365 12483 14399
rect 15853 14365 15887 14399
rect 18337 14365 18371 14399
rect 18613 14365 18647 14399
rect 5365 14229 5399 14263
rect 8677 14229 8711 14263
rect 8953 14229 8987 14263
rect 10885 14229 10919 14263
rect 22845 14229 22879 14263
rect 4353 14025 4387 14059
rect 7941 14025 7975 14059
rect 9597 14025 9631 14059
rect 15117 14025 15151 14059
rect 18429 14025 18463 14059
rect 19441 14025 19475 14059
rect 20729 14025 20763 14059
rect 2789 13889 2823 13923
rect 6101 13889 6135 13923
rect 9873 13957 9907 13991
rect 10701 13957 10735 13991
rect 19809 13957 19843 13991
rect 15025 13889 15059 13923
rect 15485 13889 15519 13923
rect 18153 13889 18187 13923
rect 20913 13889 20947 13923
rect 2513 13821 2547 13855
rect 4445 13821 4479 13855
rect 5733 13821 5767 13855
rect 7941 13821 7975 13855
rect 8033 13821 8067 13855
rect 8309 13821 8343 13855
rect 10517 13821 10551 13855
rect 15301 13821 15335 13855
rect 15577 13821 15611 13855
rect 16129 13821 16163 13855
rect 16313 13821 16347 13855
rect 18061 13821 18095 13855
rect 19625 13821 19659 13855
rect 21097 13821 21131 13855
rect 21649 13821 21683 13855
rect 21833 13821 21867 13855
rect 16681 13753 16715 13787
rect 22201 13753 22235 13787
rect 3893 13685 3927 13719
rect 5825 13685 5859 13719
rect 6101 13481 6135 13515
rect 7297 13481 7331 13515
rect 8585 13481 8619 13515
rect 14105 13481 14139 13515
rect 21741 13481 21775 13515
rect 23489 13481 23523 13515
rect 11345 13413 11379 13447
rect 13829 13413 13863 13447
rect 18245 13413 18279 13447
rect 7573 13345 7607 13379
rect 8125 13345 8159 13379
rect 8309 13345 8343 13379
rect 9689 13345 9723 13379
rect 11529 13345 11563 13379
rect 11713 13345 11747 13379
rect 12265 13345 12299 13379
rect 12449 13345 12483 13379
rect 13737 13345 13771 13379
rect 14933 13345 14967 13379
rect 16865 13345 16899 13379
rect 21925 13345 21959 13379
rect 22201 13345 22235 13379
rect 4537 13277 4571 13311
rect 4813 13277 4847 13311
rect 7389 13277 7423 13311
rect 16589 13277 16623 13311
rect 9873 13209 9907 13243
rect 6285 13141 6319 13175
rect 12725 13141 12759 13175
rect 14749 13141 14783 13175
rect 16405 13141 16439 13175
rect 4445 12937 4479 12971
rect 5733 12937 5767 12971
rect 7941 12937 7975 12971
rect 10517 12937 10551 12971
rect 20545 12937 20579 12971
rect 14013 12869 14047 12903
rect 4629 12801 4663 12835
rect 12725 12801 12759 12835
rect 14197 12801 14231 12835
rect 20637 12801 20671 12835
rect 4721 12733 4755 12767
rect 5273 12733 5307 12767
rect 5457 12733 5491 12767
rect 7573 12733 7607 12767
rect 10333 12733 10367 12767
rect 12449 12733 12483 12767
rect 15025 12733 15059 12767
rect 15209 12733 15243 12767
rect 15761 12733 15795 12767
rect 15945 12733 15979 12767
rect 20821 12733 20855 12767
rect 21373 12733 21407 12767
rect 21557 12733 21591 12767
rect 7665 12597 7699 12631
rect 14841 12597 14875 12631
rect 16221 12597 16255 12631
rect 21833 12597 21867 12631
rect 5089 12393 5123 12427
rect 8493 12393 8527 12427
rect 21373 12393 21407 12427
rect 17325 12325 17359 12359
rect 23121 12325 23155 12359
rect 4905 12257 4939 12291
rect 6193 12257 6227 12291
rect 6745 12257 6779 12291
rect 6929 12257 6963 12291
rect 8217 12257 8251 12291
rect 15945 12257 15979 12291
rect 18337 12257 18371 12291
rect 21465 12257 21499 12291
rect 21741 12257 21775 12291
rect 6009 12189 6043 12223
rect 15669 12189 15703 12223
rect 17417 12189 17451 12223
rect 5825 12053 5859 12087
rect 7205 12053 7239 12087
rect 8309 12053 8343 12087
rect 18153 12053 18187 12087
rect 4353 11849 4387 11883
rect 8401 11849 8435 11883
rect 16589 11849 16623 11883
rect 16865 11849 16899 11883
rect 21373 11849 21407 11883
rect 22293 11849 22327 11883
rect 4537 11781 4571 11815
rect 2789 11713 2823 11747
rect 7021 11713 7055 11747
rect 7297 11713 7331 11747
rect 19533 11713 19567 11747
rect 19809 11713 19843 11747
rect 2513 11645 2547 11679
rect 8769 11645 8803 11679
rect 16497 11645 16531 11679
rect 22201 11645 22235 11679
rect 3893 11509 3927 11543
rect 20913 11509 20947 11543
rect 8493 11305 8527 11339
rect 8861 11305 8895 11339
rect 19073 11305 19107 11339
rect 7113 11169 7147 11203
rect 13277 11169 13311 11203
rect 13645 11169 13679 11203
rect 16405 11169 16439 11203
rect 19901 11169 19935 11203
rect 7389 11101 7423 11135
rect 12725 11101 12759 11135
rect 13369 11101 13403 11135
rect 13553 11101 13587 11135
rect 17233 11101 17267 11135
rect 17509 11101 17543 11135
rect 13921 11033 13955 11067
rect 16221 11033 16255 11067
rect 19257 11033 19291 11067
rect 19717 11033 19751 11067
rect 18613 10965 18647 10999
rect 4353 10761 4387 10795
rect 8033 10761 8067 10795
rect 13829 10761 13863 10795
rect 19441 10761 19475 10795
rect 20361 10761 20395 10795
rect 14289 10693 14323 10727
rect 2513 10625 2547 10659
rect 12725 10625 12759 10659
rect 18337 10625 18371 10659
rect 20545 10625 20579 10659
rect 20821 10625 20855 10659
rect 2789 10557 2823 10591
rect 6837 10557 6871 10591
rect 7021 10557 7055 10591
rect 7573 10557 7607 10591
rect 7757 10557 7791 10591
rect 12449 10557 12483 10591
rect 18061 10557 18095 10591
rect 3893 10421 3927 10455
rect 6561 10421 6595 10455
rect 17785 10421 17819 10455
rect 21925 10421 21959 10455
rect 13829 10217 13863 10251
rect 20913 10217 20947 10251
rect 8217 10149 8251 10183
rect 6561 10081 6595 10115
rect 7757 10081 7791 10115
rect 15301 10081 15335 10115
rect 21097 10081 21131 10115
rect 21373 10081 21407 10115
rect 7665 10013 7699 10047
rect 12265 10013 12299 10047
rect 12541 10013 12575 10047
rect 6745 9945 6779 9979
rect 15393 9945 15427 9979
rect 7021 9877 7055 9911
rect 14013 9877 14047 9911
rect 22477 9877 22511 9911
rect 20729 9673 20763 9707
rect 7757 9605 7791 9639
rect 2789 9537 2823 9571
rect 4261 9537 4295 9571
rect 8493 9537 8527 9571
rect 9321 9537 9355 9571
rect 12909 9537 12943 9571
rect 13829 9537 13863 9571
rect 20361 9537 20395 9571
rect 2513 9469 2547 9503
rect 8033 9469 8067 9503
rect 9413 9469 9447 9503
rect 13369 9469 13403 9503
rect 13553 9469 13587 9503
rect 13921 9469 13955 9503
rect 18981 9469 19015 9503
rect 19257 9469 19291 9503
rect 7941 9401 7975 9435
rect 9873 9401 9907 9435
rect 3893 9333 3927 9367
rect 8677 9333 8711 9367
rect 14289 9333 14323 9367
rect 9965 9129 9999 9163
rect 14105 9129 14139 9163
rect 19441 9129 19475 9163
rect 21373 9129 21407 9163
rect 8677 9061 8711 9095
rect 15393 9061 15427 9095
rect 6469 8993 6503 9027
rect 7757 8993 7791 9027
rect 7941 8993 7975 9027
rect 8033 8993 8067 9027
rect 9689 8993 9723 9027
rect 9873 8993 9907 9027
rect 14473 8993 14507 9027
rect 15301 8993 15335 9027
rect 18613 8993 18647 9027
rect 21557 8993 21591 9027
rect 21833 8993 21867 9027
rect 6377 8925 6411 8959
rect 12725 8925 12759 8959
rect 13001 8925 13035 8959
rect 15669 8857 15703 8891
rect 6653 8789 6687 8823
rect 8217 8789 8251 8823
rect 19257 8789 19291 8823
rect 22937 8789 22971 8823
rect 8401 8585 8435 8619
rect 10149 8585 10183 8619
rect 18613 8585 18647 8619
rect 20085 8585 20119 8619
rect 20545 8585 20579 8619
rect 15761 8517 15795 8551
rect 2789 8449 2823 8483
rect 13553 8449 13587 8483
rect 14473 8449 14507 8483
rect 2513 8381 2547 8415
rect 6837 8381 6871 8415
rect 7113 8381 7147 8415
rect 9689 8381 9723 8415
rect 14013 8381 14047 8415
rect 14197 8381 14231 8415
rect 14565 8381 14599 8415
rect 15577 8381 15611 8415
rect 18613 8381 18647 8415
rect 18705 8381 18739 8415
rect 18981 8381 19015 8415
rect 4353 8313 4387 8347
rect 3893 8245 3927 8279
rect 8585 8245 8619 8279
rect 9873 8245 9907 8279
rect 9965 8041 9999 8075
rect 14105 8041 14139 8075
rect 7389 7973 7423 8007
rect 9689 7973 9723 8007
rect 11805 7973 11839 8007
rect 8033 7905 8067 7939
rect 8401 7905 8435 7939
rect 8493 7905 8527 7939
rect 8769 7905 8803 7939
rect 9873 7905 9907 7939
rect 11989 7905 12023 7939
rect 12357 7905 12391 7939
rect 13369 7905 13403 7939
rect 13461 7905 13495 7939
rect 15485 7905 15519 7939
rect 15577 7905 15611 7939
rect 7849 7837 7883 7871
rect 16037 7837 16071 7871
rect 13093 7769 13127 7803
rect 13185 7769 13219 7803
rect 13645 7701 13679 7735
rect 15117 7701 15151 7735
rect 15301 7701 15335 7735
rect 8585 7497 8619 7531
rect 15301 7497 15335 7531
rect 15485 7497 15519 7531
rect 20729 7497 20763 7531
rect 22293 7497 22327 7531
rect 2789 7361 2823 7395
rect 13737 7361 13771 7395
rect 19349 7361 19383 7395
rect 20913 7361 20947 7395
rect 2513 7293 2547 7327
rect 7021 7293 7055 7327
rect 7297 7293 7331 7327
rect 14013 7293 14047 7327
rect 21189 7293 21223 7327
rect 3893 7157 3927 7191
rect 4353 7157 4387 7191
rect 8769 7157 8803 7191
rect 19993 7157 20027 7191
rect 15117 6953 15151 6987
rect 20729 6953 20763 6987
rect 22293 6953 22327 6987
rect 7113 6885 7147 6919
rect 15301 6885 15335 6919
rect 11161 6817 11195 6851
rect 13829 6817 13863 6851
rect 14013 6817 14047 6851
rect 14381 6817 14415 6851
rect 15945 6817 15979 6851
rect 16313 6817 16347 6851
rect 19257 6817 19291 6851
rect 21189 6817 21223 6851
rect 5457 6749 5491 6783
rect 5733 6749 5767 6783
rect 11437 6749 11471 6783
rect 12541 6749 12575 6783
rect 15761 6749 15795 6783
rect 16221 6749 16255 6783
rect 20913 6749 20947 6783
rect 7297 6613 7331 6647
rect 13001 6613 13035 6647
rect 19901 6613 19935 6647
rect 4353 6409 4387 6443
rect 21649 6409 21683 6443
rect 7849 6273 7883 6307
rect 8401 6273 8435 6307
rect 20177 6273 20211 6307
rect 20269 6273 20303 6307
rect 2513 6205 2547 6239
rect 2789 6205 2823 6239
rect 8493 6205 8527 6239
rect 8861 6205 8895 6239
rect 9045 6205 9079 6239
rect 15393 6205 15427 6239
rect 15577 6205 15611 6239
rect 15945 6205 15979 6239
rect 16129 6205 16163 6239
rect 20545 6205 20579 6239
rect 3893 6069 3927 6103
rect 4537 6069 4571 6103
rect 15209 6069 15243 6103
rect 5917 5865 5951 5899
rect 15025 5865 15059 5899
rect 16681 5865 16715 5899
rect 21557 5865 21591 5899
rect 21741 5865 21775 5899
rect 5733 5797 5767 5831
rect 11529 5797 11563 5831
rect 11989 5729 12023 5763
rect 12173 5729 12207 5763
rect 12541 5729 12575 5763
rect 12725 5729 12759 5763
rect 15577 5729 15611 5763
rect 19165 5729 19199 5763
rect 22201 5729 22235 5763
rect 4077 5661 4111 5695
rect 4353 5661 4387 5695
rect 15301 5661 15335 5695
rect 21925 5661 21959 5695
rect 19809 5525 19843 5559
rect 23489 5525 23523 5559
rect 4261 5321 4295 5355
rect 5641 5321 5675 5355
rect 8493 5321 8527 5355
rect 15301 5321 15335 5355
rect 16865 5321 16899 5355
rect 20913 5321 20947 5355
rect 21373 5321 21407 5355
rect 2789 5185 2823 5219
rect 15485 5185 15519 5219
rect 19809 5185 19843 5219
rect 2513 5117 2547 5151
rect 4997 5117 5031 5151
rect 6929 5117 6963 5151
rect 7205 5117 7239 5151
rect 15761 5117 15795 5151
rect 19533 5117 19567 5151
rect 3893 4981 3927 5015
rect 8769 4981 8803 5015
rect 7297 4777 7331 4811
rect 16681 4777 16715 4811
rect 7205 4709 7239 4743
rect 12449 4709 12483 4743
rect 5549 4641 5583 4675
rect 10793 4641 10827 4675
rect 13277 4641 13311 4675
rect 15577 4641 15611 4675
rect 5825 4573 5859 4607
rect 11069 4573 11103 4607
rect 15301 4573 15335 4607
rect 12633 4505 12667 4539
rect 13921 4437 13955 4471
rect 17049 4437 17083 4471
rect 4261 4233 4295 4267
rect 11161 4233 11195 4267
rect 2513 4097 2547 4131
rect 6837 4097 6871 4131
rect 9873 4097 9907 4131
rect 2789 4029 2823 4063
rect 7481 4029 7515 4063
rect 9597 4029 9631 4063
rect 11345 4029 11379 4063
rect 3893 3893 3927 3927
rect 5273 3145 5307 3179
rect 10517 3145 10551 3179
rect 3249 3009 3283 3043
rect 8677 3009 8711 3043
rect 8953 3009 8987 3043
rect 3525 2941 3559 2975
rect 5089 2941 5123 2975
rect 4629 2805 4663 2839
rect 10057 2805 10091 2839
<< metal1 >>
rect 4062 44140 4068 44192
rect 4120 44180 4126 44192
rect 75546 44180 75552 44192
rect 4120 44152 75552 44180
rect 4120 44140 4126 44152
rect 75546 44140 75552 44152
rect 75604 44140 75610 44192
rect 1104 44090 105616 44112
rect 1104 44038 19606 44090
rect 19658 44038 19670 44090
rect 19722 44038 19734 44090
rect 19786 44038 19798 44090
rect 19850 44038 50326 44090
rect 50378 44038 50390 44090
rect 50442 44038 50454 44090
rect 50506 44038 50518 44090
rect 50570 44038 81046 44090
rect 81098 44038 81110 44090
rect 81162 44038 81174 44090
rect 81226 44038 81238 44090
rect 81290 44038 105616 44090
rect 1104 44016 105616 44038
rect 17862 43908 17868 43920
rect 16500 43880 17868 43908
rect 16500 43849 16528 43880
rect 17862 43868 17868 43880
rect 17920 43868 17926 43920
rect 45922 43908 45928 43920
rect 44652 43880 45928 43908
rect 15933 43843 15991 43849
rect 15933 43809 15945 43843
rect 15979 43840 15991 43843
rect 16485 43843 16543 43849
rect 16485 43840 16497 43843
rect 15979 43812 16497 43840
rect 15979 43809 15991 43812
rect 15933 43803 15991 43809
rect 16485 43809 16497 43812
rect 16531 43809 16543 43843
rect 16485 43803 16543 43809
rect 16669 43843 16727 43849
rect 16669 43809 16681 43843
rect 16715 43840 16727 43843
rect 28258 43840 28264 43852
rect 16715 43812 17356 43840
rect 28219 43812 28264 43840
rect 16715 43809 16727 43812
rect 16669 43803 16727 43809
rect 15654 43772 15660 43784
rect 15567 43744 15660 43772
rect 15654 43732 15660 43744
rect 15712 43772 15718 43784
rect 15749 43775 15807 43781
rect 15749 43772 15761 43775
rect 15712 43744 15761 43772
rect 15712 43732 15718 43744
rect 15749 43741 15761 43744
rect 15795 43741 15807 43775
rect 15749 43735 15807 43741
rect 16945 43639 17003 43645
rect 16945 43605 16957 43639
rect 16991 43636 17003 43639
rect 17034 43636 17040 43648
rect 16991 43608 17040 43636
rect 16991 43605 17003 43608
rect 16945 43599 17003 43605
rect 17034 43596 17040 43608
rect 17092 43596 17098 43648
rect 17328 43645 17356 43812
rect 28258 43800 28264 43812
rect 28316 43800 28322 43852
rect 44652 43849 44680 43880
rect 45922 43868 45928 43880
rect 45980 43868 45986 43920
rect 44637 43843 44695 43849
rect 44284 43812 44588 43840
rect 43622 43732 43628 43784
rect 43680 43772 43686 43784
rect 44284 43781 44312 43812
rect 44269 43775 44327 43781
rect 44269 43772 44281 43775
rect 43680 43744 44281 43772
rect 43680 43732 43686 43744
rect 44269 43741 44281 43744
rect 44315 43741 44327 43775
rect 44450 43772 44456 43784
rect 44411 43744 44456 43772
rect 44269 43735 44327 43741
rect 44450 43732 44456 43744
rect 44508 43732 44514 43784
rect 44560 43772 44588 43812
rect 44637 43809 44649 43843
rect 44683 43809 44695 43843
rect 45097 43843 45155 43849
rect 45097 43840 45109 43843
rect 44637 43803 44695 43809
rect 44744 43812 45109 43840
rect 44744 43772 44772 43812
rect 45097 43809 45109 43812
rect 45143 43809 45155 43843
rect 45097 43803 45155 43809
rect 45189 43843 45247 43849
rect 45189 43809 45201 43843
rect 45235 43840 45247 43843
rect 45235 43812 48728 43840
rect 45235 43809 45247 43812
rect 45189 43803 45247 43809
rect 44560 43744 44772 43772
rect 48700 43772 48728 43812
rect 48774 43800 48780 43852
rect 48832 43840 48838 43852
rect 53653 43843 53711 43849
rect 53653 43840 53665 43843
rect 48832 43812 53665 43840
rect 48832 43800 48838 43812
rect 53653 43809 53665 43812
rect 53699 43840 53711 43843
rect 54570 43840 54576 43852
rect 53699 43812 54576 43840
rect 53699 43809 53711 43812
rect 53653 43803 53711 43809
rect 54570 43800 54576 43812
rect 54628 43800 54634 43852
rect 58526 43840 58532 43852
rect 58487 43812 58532 43840
rect 58526 43800 58532 43812
rect 58584 43800 58590 43852
rect 59538 43840 59544 43852
rect 59499 43812 59544 43840
rect 59538 43800 59544 43812
rect 59596 43800 59602 43852
rect 59725 43843 59783 43849
rect 59725 43809 59737 43843
rect 59771 43840 59783 43843
rect 59998 43840 60004 43852
rect 59771 43812 60004 43840
rect 59771 43809 59783 43812
rect 59725 43803 59783 43809
rect 59998 43800 60004 43812
rect 60056 43800 60062 43852
rect 73801 43843 73859 43849
rect 73801 43809 73813 43843
rect 73847 43840 73859 43843
rect 74074 43840 74080 43852
rect 73847 43812 74080 43840
rect 73847 43809 73859 43812
rect 73801 43803 73859 43809
rect 74074 43800 74080 43812
rect 74132 43800 74138 43852
rect 78493 43843 78551 43849
rect 78493 43809 78505 43843
rect 78539 43840 78551 43843
rect 78582 43840 78588 43852
rect 78539 43812 78588 43840
rect 78539 43809 78551 43812
rect 78493 43803 78551 43809
rect 78582 43800 78588 43812
rect 78640 43840 78646 43852
rect 78769 43843 78827 43849
rect 78769 43840 78781 43843
rect 78640 43812 78781 43840
rect 78640 43800 78646 43812
rect 78769 43809 78781 43812
rect 78815 43809 78827 43843
rect 78769 43803 78827 43809
rect 78858 43800 78864 43852
rect 78916 43840 78922 43852
rect 79321 43843 79379 43849
rect 79321 43840 79333 43843
rect 78916 43812 79333 43840
rect 78916 43800 78922 43812
rect 79321 43809 79333 43812
rect 79367 43809 79379 43843
rect 79321 43803 79379 43809
rect 79781 43843 79839 43849
rect 79781 43809 79793 43843
rect 79827 43840 79839 43843
rect 81434 43840 81440 43852
rect 79827 43812 81440 43840
rect 79827 43809 79839 43812
rect 79781 43803 79839 43809
rect 49602 43772 49608 43784
rect 48700 43744 49608 43772
rect 49602 43732 49608 43744
rect 49660 43732 49666 43784
rect 60093 43775 60151 43781
rect 60093 43741 60105 43775
rect 60139 43772 60151 43775
rect 61010 43772 61016 43784
rect 60139 43744 61016 43772
rect 60139 43741 60151 43744
rect 60093 43735 60151 43741
rect 61010 43732 61016 43744
rect 61068 43732 61074 43784
rect 78674 43732 78680 43784
rect 78732 43772 78738 43784
rect 79796 43772 79824 43803
rect 81434 43800 81440 43812
rect 81492 43840 81498 43852
rect 82265 43843 82323 43849
rect 82265 43840 82277 43843
rect 81492 43812 82277 43840
rect 81492 43800 81498 43812
rect 82265 43809 82277 43812
rect 82311 43809 82323 43843
rect 82265 43803 82323 43809
rect 82354 43800 82360 43852
rect 82412 43840 82418 43852
rect 82412 43812 82457 43840
rect 82412 43800 82418 43812
rect 82814 43772 82820 43784
rect 78732 43744 79824 43772
rect 82775 43744 82820 43772
rect 78732 43732 78738 43744
rect 82814 43732 82820 43744
rect 82872 43732 82878 43784
rect 26234 43664 26240 43716
rect 26292 43704 26298 43716
rect 28353 43707 28411 43713
rect 28353 43704 28365 43707
rect 26292 43676 28365 43704
rect 26292 43664 26298 43676
rect 28353 43673 28365 43676
rect 28399 43704 28411 43707
rect 48314 43704 48320 43716
rect 28399 43676 48320 43704
rect 28399 43673 28411 43676
rect 28353 43667 28411 43673
rect 48314 43664 48320 43676
rect 48372 43664 48378 43716
rect 73893 43707 73951 43713
rect 73893 43673 73905 43707
rect 73939 43704 73951 43707
rect 74258 43704 74264 43716
rect 73939 43676 74264 43704
rect 73939 43673 73951 43676
rect 73893 43667 73951 43673
rect 74258 43664 74264 43676
rect 74316 43664 74322 43716
rect 78490 43664 78496 43716
rect 78548 43704 78554 43716
rect 78861 43707 78919 43713
rect 78861 43704 78873 43707
rect 78548 43676 78873 43704
rect 78548 43664 78554 43676
rect 78861 43673 78873 43676
rect 78907 43673 78919 43707
rect 78861 43667 78919 43673
rect 17313 43639 17371 43645
rect 17313 43605 17325 43639
rect 17359 43636 17371 43639
rect 18414 43636 18420 43648
rect 17359 43608 18420 43636
rect 17359 43605 17371 43608
rect 17313 43599 17371 43605
rect 18414 43596 18420 43608
rect 18472 43596 18478 43648
rect 44177 43639 44235 43645
rect 44177 43605 44189 43639
rect 44223 43636 44235 43639
rect 44542 43636 44548 43648
rect 44223 43608 44548 43636
rect 44223 43605 44235 43608
rect 44177 43599 44235 43605
rect 44542 43596 44548 43608
rect 44600 43596 44606 43648
rect 45646 43636 45652 43648
rect 45607 43608 45652 43636
rect 45646 43596 45652 43608
rect 45704 43596 45710 43648
rect 45922 43636 45928 43648
rect 45883 43608 45928 43636
rect 45922 43596 45928 43608
rect 45980 43596 45986 43648
rect 53834 43636 53840 43648
rect 53795 43608 53840 43636
rect 53834 43596 53840 43608
rect 53892 43596 53898 43648
rect 58621 43639 58679 43645
rect 58621 43605 58633 43639
rect 58667 43636 58679 43639
rect 59078 43636 59084 43648
rect 58667 43608 59084 43636
rect 58667 43605 58679 43608
rect 58621 43599 58679 43605
rect 59078 43596 59084 43608
rect 59136 43596 59142 43648
rect 74074 43636 74080 43648
rect 74035 43608 74080 43636
rect 74074 43596 74080 43608
rect 74132 43596 74138 43648
rect 78677 43639 78735 43645
rect 78677 43605 78689 43639
rect 78723 43636 78735 43639
rect 78766 43636 78772 43648
rect 78723 43608 78772 43636
rect 78723 43605 78735 43608
rect 78677 43599 78735 43605
rect 78766 43596 78772 43608
rect 78824 43596 78830 43648
rect 82078 43636 82084 43648
rect 82039 43608 82084 43636
rect 82078 43596 82084 43608
rect 82136 43596 82142 43648
rect 1104 43546 105616 43568
rect 1104 43494 4246 43546
rect 4298 43494 4310 43546
rect 4362 43494 4374 43546
rect 4426 43494 4438 43546
rect 4490 43494 34966 43546
rect 35018 43494 35030 43546
rect 35082 43494 35094 43546
rect 35146 43494 35158 43546
rect 35210 43494 65686 43546
rect 65738 43494 65750 43546
rect 65802 43494 65814 43546
rect 65866 43494 65878 43546
rect 65930 43494 96406 43546
rect 96458 43494 96470 43546
rect 96522 43494 96534 43546
rect 96586 43494 96598 43546
rect 96650 43494 105616 43546
rect 1104 43472 105616 43494
rect 18414 43392 18420 43444
rect 18472 43432 18478 43444
rect 36817 43435 36875 43441
rect 36817 43432 36829 43435
rect 18472 43404 36829 43432
rect 18472 43392 18478 43404
rect 36817 43401 36829 43404
rect 36863 43432 36875 43435
rect 37001 43435 37059 43441
rect 37001 43432 37013 43435
rect 36863 43404 37013 43432
rect 36863 43401 36875 43404
rect 36817 43395 36875 43401
rect 37001 43401 37013 43404
rect 37047 43401 37059 43435
rect 48314 43432 48320 43444
rect 48275 43404 48320 43432
rect 37001 43395 37059 43401
rect 2409 43299 2467 43305
rect 2409 43265 2421 43299
rect 2455 43296 2467 43299
rect 2774 43296 2780 43308
rect 2455 43268 2780 43296
rect 2455 43265 2467 43268
rect 2409 43259 2467 43265
rect 2774 43256 2780 43268
rect 2832 43296 2838 43308
rect 3142 43296 3148 43308
rect 2832 43268 3148 43296
rect 2832 43256 2838 43268
rect 3142 43256 3148 43268
rect 3200 43256 3206 43308
rect 7561 43299 7619 43305
rect 7561 43265 7573 43299
rect 7607 43296 7619 43299
rect 8570 43296 8576 43308
rect 7607 43268 8576 43296
rect 7607 43265 7619 43268
rect 7561 43259 7619 43265
rect 8570 43256 8576 43268
rect 8628 43296 8634 43308
rect 9309 43299 9367 43305
rect 9309 43296 9321 43299
rect 8628 43268 9321 43296
rect 8628 43256 8634 43268
rect 9309 43265 9321 43268
rect 9355 43265 9367 43299
rect 9309 43259 9367 43265
rect 26973 43299 27031 43305
rect 26973 43265 26985 43299
rect 27019 43296 27031 43299
rect 27154 43296 27160 43308
rect 27019 43268 27160 43296
rect 27019 43265 27031 43268
rect 26973 43259 27031 43265
rect 27154 43256 27160 43268
rect 27212 43256 27218 43308
rect 37016 43296 37044 43395
rect 48314 43392 48320 43404
rect 48372 43432 48378 43444
rect 48409 43435 48467 43441
rect 48409 43432 48421 43435
rect 48372 43404 48421 43432
rect 48372 43392 48378 43404
rect 48409 43401 48421 43404
rect 48455 43401 48467 43435
rect 48409 43395 48467 43401
rect 50157 43435 50215 43441
rect 50157 43401 50169 43435
rect 50203 43432 50215 43435
rect 53834 43432 53840 43444
rect 50203 43404 53840 43432
rect 50203 43401 50215 43404
rect 50157 43395 50215 43401
rect 37185 43299 37243 43305
rect 37185 43296 37197 43299
rect 32232 43268 32812 43296
rect 37016 43268 37197 43296
rect 2501 43231 2559 43237
rect 2501 43197 2513 43231
rect 2547 43197 2559 43231
rect 7834 43228 7840 43240
rect 7795 43200 7840 43228
rect 2501 43191 2559 43197
rect 2516 43092 2544 43191
rect 7834 43188 7840 43200
rect 7892 43188 7898 43240
rect 12342 43188 12348 43240
rect 12400 43228 12406 43240
rect 12437 43231 12495 43237
rect 12437 43228 12449 43231
rect 12400 43200 12449 43228
rect 12400 43188 12406 43200
rect 12437 43197 12449 43200
rect 12483 43197 12495 43231
rect 15470 43228 15476 43240
rect 15431 43200 15476 43228
rect 12437 43191 12495 43197
rect 15470 43188 15476 43200
rect 15528 43188 15534 43240
rect 15749 43231 15807 43237
rect 15749 43197 15761 43231
rect 15795 43228 15807 43231
rect 16666 43228 16672 43240
rect 15795 43200 16672 43228
rect 15795 43197 15807 43200
rect 15749 43191 15807 43197
rect 16666 43188 16672 43200
rect 16724 43188 16730 43240
rect 17129 43231 17187 43237
rect 17129 43197 17141 43231
rect 17175 43228 17187 43231
rect 18049 43231 18107 43237
rect 18049 43228 18061 43231
rect 17175 43200 18061 43228
rect 17175 43197 17187 43200
rect 17129 43191 17187 43197
rect 18049 43197 18061 43200
rect 18095 43197 18107 43231
rect 20441 43231 20499 43237
rect 20441 43228 20453 43231
rect 18049 43191 18107 43197
rect 20272 43200 20453 43228
rect 3712 43132 4384 43160
rect 3712 43092 3740 43132
rect 3878 43092 3884 43104
rect 2516 43064 3740 43092
rect 3839 43064 3884 43092
rect 3878 43052 3884 43064
rect 3936 43052 3942 43104
rect 4356 43101 4384 43132
rect 4341 43095 4399 43101
rect 4341 43061 4353 43095
rect 4387 43092 4399 43095
rect 4798 43092 4804 43104
rect 4387 43064 4804 43092
rect 4387 43061 4399 43064
rect 4341 43055 4399 43061
rect 4798 43052 4804 43064
rect 4856 43052 4862 43104
rect 8938 43092 8944 43104
rect 8899 43064 8944 43092
rect 8938 43052 8944 43064
rect 8996 43052 9002 43104
rect 12526 43092 12532 43104
rect 12487 43064 12532 43092
rect 12526 43052 12532 43064
rect 12584 43052 12590 43104
rect 16482 43052 16488 43104
rect 16540 43092 16546 43104
rect 17221 43095 17279 43101
rect 17221 43092 17233 43095
rect 16540 43064 17233 43092
rect 16540 43052 16546 43064
rect 17221 43061 17233 43064
rect 17267 43061 17279 43095
rect 18138 43092 18144 43104
rect 18099 43064 18144 43092
rect 17221 43055 17279 43061
rect 18138 43052 18144 43064
rect 18196 43052 18202 43104
rect 20162 43052 20168 43104
rect 20220 43092 20226 43104
rect 20272 43101 20300 43200
rect 20441 43197 20453 43200
rect 20487 43197 20499 43231
rect 20441 43191 20499 43197
rect 20625 43231 20683 43237
rect 20625 43197 20637 43231
rect 20671 43228 20683 43231
rect 21174 43228 21180 43240
rect 20671 43200 21180 43228
rect 20671 43197 20683 43200
rect 20625 43191 20683 43197
rect 21174 43188 21180 43200
rect 21232 43188 21238 43240
rect 21361 43231 21419 43237
rect 21361 43197 21373 43231
rect 21407 43228 21419 43231
rect 26697 43231 26755 43237
rect 21407 43200 22048 43228
rect 21407 43197 21419 43200
rect 21361 43191 21419 43197
rect 20257 43095 20315 43101
rect 20257 43092 20269 43095
rect 20220 43064 20269 43092
rect 20220 43052 20226 43064
rect 20257 43061 20269 43064
rect 20303 43061 20315 43095
rect 20257 43055 20315 43061
rect 21450 43052 21456 43104
rect 21508 43092 21514 43104
rect 22020 43101 22048 43200
rect 26697 43197 26709 43231
rect 26743 43197 26755 43231
rect 26697 43191 26755 43197
rect 26712 43104 26740 43191
rect 28353 43163 28411 43169
rect 28353 43129 28365 43163
rect 28399 43160 28411 43163
rect 29178 43160 29184 43172
rect 28399 43132 29184 43160
rect 28399 43129 28411 43132
rect 28353 43123 28411 43129
rect 29178 43120 29184 43132
rect 29236 43120 29242 43172
rect 21637 43095 21695 43101
rect 21637 43092 21649 43095
rect 21508 43064 21649 43092
rect 21508 43052 21514 43064
rect 21637 43061 21649 43064
rect 21683 43061 21695 43095
rect 21637 43055 21695 43061
rect 22005 43095 22063 43101
rect 22005 43061 22017 43095
rect 22051 43092 22063 43095
rect 22094 43092 22100 43104
rect 22051 43064 22100 43092
rect 22051 43061 22063 43064
rect 22005 43055 22063 43061
rect 22094 43052 22100 43064
rect 22152 43052 22158 43104
rect 26694 43092 26700 43104
rect 26607 43064 26700 43092
rect 26694 43052 26700 43064
rect 26752 43092 26758 43104
rect 28442 43092 28448 43104
rect 26752 43064 28448 43092
rect 26752 43052 26758 43064
rect 28442 43052 28448 43064
rect 28500 43052 28506 43104
rect 31938 43052 31944 43104
rect 31996 43092 32002 43104
rect 32232 43101 32260 43268
rect 32784 43237 32812 43268
rect 37185 43265 37197 43268
rect 37231 43296 37243 43299
rect 38473 43299 38531 43305
rect 37231 43268 37504 43296
rect 37231 43265 37243 43268
rect 37185 43259 37243 43265
rect 32585 43231 32643 43237
rect 32585 43228 32597 43231
rect 32416 43200 32597 43228
rect 32033 43095 32091 43101
rect 32033 43092 32045 43095
rect 31996 43064 32045 43092
rect 31996 43052 32002 43064
rect 32033 43061 32045 43064
rect 32079 43092 32091 43095
rect 32217 43095 32275 43101
rect 32217 43092 32229 43095
rect 32079 43064 32229 43092
rect 32079 43061 32091 43064
rect 32033 43055 32091 43061
rect 32217 43061 32229 43064
rect 32263 43061 32275 43095
rect 32217 43055 32275 43061
rect 32306 43052 32312 43104
rect 32364 43092 32370 43104
rect 32416 43101 32444 43200
rect 32585 43197 32597 43200
rect 32631 43197 32643 43231
rect 32585 43191 32643 43197
rect 32769 43231 32827 43237
rect 32769 43197 32781 43231
rect 32815 43197 32827 43231
rect 33226 43228 33232 43240
rect 33187 43200 33232 43228
rect 32769 43191 32827 43197
rect 32784 43160 32812 43191
rect 33226 43188 33232 43200
rect 33284 43188 33290 43240
rect 33321 43231 33379 43237
rect 33321 43197 33333 43231
rect 33367 43228 33379 43231
rect 33962 43228 33968 43240
rect 33367 43200 33968 43228
rect 33367 43197 33379 43200
rect 33321 43191 33379 43197
rect 33336 43160 33364 43191
rect 33962 43188 33968 43200
rect 34020 43188 34026 43240
rect 37369 43231 37427 43237
rect 37369 43197 37381 43231
rect 37415 43197 37427 43231
rect 37476 43228 37504 43268
rect 38473 43265 38485 43299
rect 38519 43296 38531 43299
rect 38838 43296 38844 43308
rect 38519 43268 38844 43296
rect 38519 43265 38531 43268
rect 38473 43259 38531 43265
rect 38838 43256 38844 43268
rect 38896 43256 38902 43308
rect 40034 43256 40040 43308
rect 40092 43296 40098 43308
rect 41325 43299 41383 43305
rect 41325 43296 41337 43299
rect 40092 43268 41337 43296
rect 40092 43256 40098 43268
rect 41325 43265 41337 43268
rect 41371 43265 41383 43299
rect 48424 43296 48452 43395
rect 48593 43299 48651 43305
rect 48593 43296 48605 43299
rect 48424 43268 48605 43296
rect 41325 43259 41383 43265
rect 48593 43265 48605 43268
rect 48639 43296 48651 43299
rect 48639 43268 48912 43296
rect 48639 43265 48651 43268
rect 48593 43259 48651 43265
rect 37829 43231 37887 43237
rect 37829 43228 37841 43231
rect 37476 43200 37841 43228
rect 37369 43191 37427 43197
rect 37829 43197 37841 43200
rect 37875 43197 37887 43231
rect 37829 43191 37887 43197
rect 37921 43231 37979 43237
rect 37921 43197 37933 43231
rect 37967 43228 37979 43231
rect 41049 43231 41107 43237
rect 41049 43228 41061 43231
rect 37967 43200 38792 43228
rect 37967 43197 37979 43200
rect 37921 43191 37979 43197
rect 32784 43132 33364 43160
rect 33873 43163 33931 43169
rect 33873 43129 33885 43163
rect 33919 43160 33931 43163
rect 35250 43160 35256 43172
rect 33919 43132 35256 43160
rect 33919 43129 33931 43132
rect 33873 43123 33931 43129
rect 35250 43120 35256 43132
rect 35308 43120 35314 43172
rect 37384 43160 37412 43191
rect 37936 43160 37964 43191
rect 37384 43132 37964 43160
rect 32401 43095 32459 43101
rect 32401 43092 32413 43095
rect 32364 43064 32413 43092
rect 32364 43052 32370 43064
rect 32401 43061 32413 43064
rect 32447 43061 32459 43095
rect 32401 43055 32459 43061
rect 33226 43052 33232 43104
rect 33284 43092 33290 43104
rect 34146 43092 34152 43104
rect 33284 43064 34152 43092
rect 33284 43052 33290 43064
rect 34146 43052 34152 43064
rect 34204 43052 34210 43104
rect 38764 43101 38792 43200
rect 40972 43200 41061 43228
rect 40972 43104 41000 43200
rect 41049 43197 41061 43200
rect 41095 43197 41107 43231
rect 48774 43228 48780 43240
rect 48735 43200 48780 43228
rect 41049 43191 41107 43197
rect 48774 43188 48780 43200
rect 48832 43188 48838 43240
rect 48884 43228 48912 43268
rect 49237 43231 49295 43237
rect 49237 43228 49249 43231
rect 48884 43200 49249 43228
rect 49237 43197 49249 43200
rect 49283 43197 49295 43231
rect 49237 43191 49295 43197
rect 49329 43231 49387 43237
rect 49329 43197 49341 43231
rect 49375 43228 49387 43231
rect 50172 43228 50200 43395
rect 53834 43392 53840 43404
rect 53892 43392 53898 43444
rect 54570 43432 54576 43444
rect 54531 43404 54576 43432
rect 54570 43392 54576 43404
rect 54628 43392 54634 43444
rect 54662 43392 54668 43444
rect 54720 43432 54726 43444
rect 55033 43435 55091 43441
rect 55033 43432 55045 43435
rect 54720 43404 55045 43432
rect 54720 43392 54726 43404
rect 55033 43401 55045 43404
rect 55079 43432 55091 43435
rect 58713 43435 58771 43441
rect 58713 43432 58725 43435
rect 55079 43404 58725 43432
rect 55079 43401 55091 43404
rect 55033 43395 55091 43401
rect 58713 43401 58725 43404
rect 58759 43432 58771 43435
rect 61102 43432 61108 43444
rect 58759 43404 61108 43432
rect 58759 43401 58771 43404
rect 58713 43395 58771 43401
rect 53374 43296 53380 43308
rect 52196 43268 53380 43296
rect 52196 43237 52224 43268
rect 53374 43256 53380 43268
rect 53432 43256 53438 43308
rect 58820 43305 58848 43404
rect 61102 43392 61108 43404
rect 61160 43392 61166 43444
rect 74626 43432 74632 43444
rect 74587 43404 74632 43432
rect 74626 43392 74632 43404
rect 74684 43392 74690 43444
rect 75546 43432 75552 43444
rect 75507 43404 75552 43432
rect 75546 43392 75552 43404
rect 75604 43392 75610 43444
rect 53469 43299 53527 43305
rect 53469 43265 53481 43299
rect 53515 43296 53527 43299
rect 58805 43299 58863 43305
rect 53515 43268 57100 43296
rect 53515 43265 53527 43268
rect 53469 43259 53527 43265
rect 49375 43200 50200 43228
rect 52181 43231 52239 43237
rect 49375 43197 49387 43200
rect 49329 43191 49387 43197
rect 52181 43197 52193 43231
rect 52227 43197 52239 43231
rect 52181 43191 52239 43197
rect 53193 43231 53251 43237
rect 53193 43197 53205 43231
rect 53239 43228 53251 43231
rect 54662 43228 54668 43240
rect 53239 43200 54668 43228
rect 53239 43197 53251 43200
rect 53193 43191 53251 43197
rect 46566 43120 46572 43172
rect 46624 43160 46630 43172
rect 49344 43160 49372 43191
rect 54662 43188 54668 43200
rect 54720 43188 54726 43240
rect 57072 43228 57100 43268
rect 58805 43265 58817 43299
rect 58851 43265 58863 43299
rect 59078 43296 59084 43308
rect 59039 43268 59084 43296
rect 58805 43259 58863 43265
rect 59078 43256 59084 43268
rect 59136 43256 59142 43308
rect 70305 43299 70363 43305
rect 70305 43265 70317 43299
rect 70351 43296 70363 43299
rect 72053 43299 72111 43305
rect 72053 43296 72065 43299
rect 70351 43268 72065 43296
rect 70351 43265 70363 43268
rect 70305 43259 70363 43265
rect 72053 43265 72065 43268
rect 72099 43296 72111 43299
rect 73890 43296 73896 43308
rect 72099 43268 73896 43296
rect 72099 43265 72111 43268
rect 72053 43259 72111 43265
rect 73890 43256 73896 43268
rect 73948 43256 73954 43308
rect 78401 43299 78459 43305
rect 78401 43265 78413 43299
rect 78447 43296 78459 43299
rect 78490 43296 78496 43308
rect 78447 43268 78496 43296
rect 78447 43265 78459 43268
rect 78401 43259 78459 43265
rect 78490 43256 78496 43268
rect 78548 43256 78554 43308
rect 82354 43296 82360 43308
rect 82315 43268 82360 43296
rect 82354 43256 82360 43268
rect 82412 43256 82418 43308
rect 59354 43228 59360 43240
rect 57072 43200 59360 43228
rect 59354 43188 59360 43200
rect 59412 43188 59418 43240
rect 63681 43231 63739 43237
rect 63681 43197 63693 43231
rect 63727 43228 63739 43231
rect 63862 43228 63868 43240
rect 63727 43200 63868 43228
rect 63727 43197 63739 43200
rect 63681 43191 63739 43197
rect 63862 43188 63868 43200
rect 63920 43188 63926 43240
rect 66898 43228 66904 43240
rect 66859 43200 66904 43228
rect 66898 43188 66904 43200
rect 66956 43188 66962 43240
rect 67177 43231 67235 43237
rect 67177 43197 67189 43231
rect 67223 43197 67235 43231
rect 67358 43228 67364 43240
rect 67319 43200 67364 43228
rect 67177 43191 67235 43197
rect 46624 43132 49372 43160
rect 46624 43120 46630 43132
rect 66254 43120 66260 43172
rect 66312 43160 66318 43172
rect 66349 43163 66407 43169
rect 66349 43160 66361 43163
rect 66312 43132 66361 43160
rect 66312 43120 66318 43132
rect 66349 43129 66361 43132
rect 66395 43129 66407 43163
rect 67192 43160 67220 43191
rect 67358 43188 67364 43200
rect 67416 43188 67422 43240
rect 70578 43228 70584 43240
rect 70539 43200 70584 43228
rect 70578 43188 70584 43200
rect 70636 43188 70642 43240
rect 74166 43228 74172 43240
rect 74127 43200 74172 43228
rect 74166 43188 74172 43200
rect 74224 43188 74230 43240
rect 74445 43231 74503 43237
rect 74445 43197 74457 43231
rect 74491 43228 74503 43231
rect 74534 43228 74540 43240
rect 74491 43200 74540 43228
rect 74491 43197 74503 43200
rect 74445 43191 74503 43197
rect 74534 43188 74540 43200
rect 74592 43188 74598 43240
rect 75546 43188 75552 43240
rect 75604 43228 75610 43240
rect 75733 43231 75791 43237
rect 75733 43228 75745 43231
rect 75604 43200 75745 43228
rect 75604 43188 75610 43200
rect 75733 43197 75745 43200
rect 75779 43197 75791 43231
rect 78674 43228 78680 43240
rect 78635 43200 78680 43228
rect 75733 43191 75791 43197
rect 78674 43188 78680 43200
rect 78732 43188 78738 43240
rect 78858 43228 78864 43240
rect 78819 43200 78864 43228
rect 78858 43188 78864 43200
rect 78916 43228 78922 43240
rect 78953 43231 79011 43237
rect 78953 43228 78965 43231
rect 78916 43200 78965 43228
rect 78916 43188 78922 43200
rect 78953 43197 78965 43200
rect 78999 43197 79011 43231
rect 81986 43228 81992 43240
rect 81947 43200 81992 43228
rect 78953 43191 79011 43197
rect 81986 43188 81992 43200
rect 82044 43188 82050 43240
rect 82541 43231 82599 43237
rect 82541 43197 82553 43231
rect 82587 43197 82599 43231
rect 82541 43191 82599 43197
rect 83553 43231 83611 43237
rect 83553 43197 83565 43231
rect 83599 43228 83611 43231
rect 83599 43200 83872 43228
rect 83599 43197 83611 43200
rect 83553 43191 83611 43197
rect 67910 43160 67916 43172
rect 67192 43132 67916 43160
rect 66349 43123 66407 43129
rect 67910 43120 67916 43132
rect 67968 43160 67974 43172
rect 69198 43160 69204 43172
rect 67968 43132 69204 43160
rect 67968 43120 67974 43132
rect 69198 43120 69204 43132
rect 69256 43120 69262 43172
rect 73246 43120 73252 43172
rect 73304 43160 73310 43172
rect 74353 43163 74411 43169
rect 74353 43160 74365 43163
rect 73304 43132 74365 43160
rect 73304 43120 73310 43132
rect 74353 43129 74365 43132
rect 74399 43129 74411 43163
rect 74353 43123 74411 43129
rect 77849 43163 77907 43169
rect 77849 43129 77861 43163
rect 77895 43160 77907 43163
rect 78766 43160 78772 43172
rect 77895 43132 78772 43160
rect 77895 43129 77907 43132
rect 77849 43123 77907 43129
rect 78766 43120 78772 43132
rect 78824 43120 78830 43172
rect 81526 43120 81532 43172
rect 81584 43160 81590 43172
rect 82556 43160 82584 43191
rect 83645 43163 83703 43169
rect 83645 43160 83657 43163
rect 81584 43132 83657 43160
rect 81584 43120 81590 43132
rect 83645 43129 83657 43132
rect 83691 43129 83703 43163
rect 83645 43123 83703 43129
rect 83844 43104 83872 43200
rect 38749 43095 38807 43101
rect 38749 43061 38761 43095
rect 38795 43092 38807 43095
rect 38841 43095 38899 43101
rect 38841 43092 38853 43095
rect 38795 43064 38853 43092
rect 38795 43061 38807 43064
rect 38749 43055 38807 43061
rect 38841 43061 38853 43064
rect 38887 43092 38899 43095
rect 39022 43092 39028 43104
rect 38887 43064 39028 43092
rect 38887 43061 38899 43064
rect 38841 43055 38899 43061
rect 39022 43052 39028 43064
rect 39080 43052 39086 43104
rect 40954 43092 40960 43104
rect 40915 43064 40960 43092
rect 40954 43052 40960 43064
rect 41012 43052 41018 43104
rect 42610 43092 42616 43104
rect 42571 43064 42616 43092
rect 42610 43052 42616 43064
rect 42668 43052 42674 43104
rect 49786 43092 49792 43104
rect 49747 43064 49792 43092
rect 49786 43052 49792 43064
rect 49844 43052 49850 43104
rect 52270 43092 52276 43104
rect 52231 43064 52276 43092
rect 52270 43052 52276 43064
rect 52328 43052 52334 43104
rect 58434 43052 58440 43104
rect 58492 43092 58498 43104
rect 59906 43092 59912 43104
rect 58492 43064 59912 43092
rect 58492 43052 58498 43064
rect 59906 43052 59912 43064
rect 59964 43092 59970 43104
rect 60185 43095 60243 43101
rect 60185 43092 60197 43095
rect 59964 43064 60197 43092
rect 59964 43052 59970 43064
rect 60185 43061 60197 43064
rect 60231 43061 60243 43095
rect 63770 43092 63776 43104
rect 63731 43064 63776 43092
rect 60185 43055 60243 43061
rect 63770 43052 63776 43064
rect 63828 43052 63834 43104
rect 71774 43052 71780 43104
rect 71832 43092 71838 43104
rect 71869 43095 71927 43101
rect 71869 43092 71881 43095
rect 71832 43064 71881 43092
rect 71832 43052 71838 43064
rect 71869 43061 71881 43064
rect 71915 43061 71927 43095
rect 75914 43092 75920 43104
rect 75875 43064 75920 43092
rect 71869 43055 71927 43061
rect 75914 43052 75920 43064
rect 75972 43052 75978 43104
rect 83826 43092 83832 43104
rect 83787 43064 83832 43092
rect 83826 43052 83832 43064
rect 83884 43052 83890 43104
rect 1104 43002 105616 43024
rect 1104 42950 19606 43002
rect 19658 42950 19670 43002
rect 19722 42950 19734 43002
rect 19786 42950 19798 43002
rect 19850 42950 50326 43002
rect 50378 42950 50390 43002
rect 50442 42950 50454 43002
rect 50506 42950 50518 43002
rect 50570 42950 81046 43002
rect 81098 42950 81110 43002
rect 81162 42950 81174 43002
rect 81226 42950 81238 43002
rect 81290 42950 105616 43002
rect 1104 42928 105616 42950
rect 3510 42848 3516 42900
rect 3568 42888 3574 42900
rect 7558 42888 7564 42900
rect 3568 42860 7564 42888
rect 3568 42848 3574 42860
rect 7558 42848 7564 42860
rect 7616 42848 7622 42900
rect 12342 42888 12348 42900
rect 12303 42860 12348 42888
rect 12342 42848 12348 42860
rect 12400 42848 12406 42900
rect 21174 42848 21180 42900
rect 21232 42888 21238 42900
rect 26050 42888 26056 42900
rect 21232 42860 26056 42888
rect 21232 42848 21238 42860
rect 26050 42848 26056 42860
rect 26108 42848 26114 42900
rect 28258 42888 28264 42900
rect 28219 42860 28264 42888
rect 28258 42848 28264 42860
rect 28316 42848 28322 42900
rect 29273 42891 29331 42897
rect 29273 42857 29285 42891
rect 29319 42888 29331 42891
rect 29362 42888 29368 42900
rect 29319 42860 29368 42888
rect 29319 42857 29331 42860
rect 29273 42851 29331 42857
rect 29362 42848 29368 42860
rect 29420 42848 29426 42900
rect 34241 42891 34299 42897
rect 34241 42857 34253 42891
rect 34287 42888 34299 42891
rect 34287 42860 38976 42888
rect 34287 42857 34299 42860
rect 34241 42851 34299 42857
rect 2608 42792 2912 42820
rect 1949 42755 2007 42761
rect 1949 42721 1961 42755
rect 1995 42752 2007 42755
rect 2501 42755 2559 42761
rect 2501 42752 2513 42755
rect 1995 42724 2513 42752
rect 1995 42721 2007 42724
rect 1949 42715 2007 42721
rect 2501 42721 2513 42724
rect 2547 42752 2559 42755
rect 2608 42752 2636 42792
rect 2547 42724 2636 42752
rect 2547 42721 2559 42724
rect 2501 42715 2559 42721
rect 2682 42712 2688 42764
rect 2740 42752 2746 42764
rect 2740 42724 2785 42752
rect 2740 42712 2746 42724
rect 1857 42687 1915 42693
rect 1857 42653 1869 42687
rect 1903 42653 1915 42687
rect 2884 42684 2912 42792
rect 23842 42780 23848 42832
rect 23900 42820 23906 42832
rect 23937 42823 23995 42829
rect 23937 42820 23949 42823
rect 23900 42792 23949 42820
rect 23900 42780 23906 42792
rect 23937 42789 23949 42792
rect 23983 42820 23995 42823
rect 33226 42820 33232 42832
rect 23983 42792 24532 42820
rect 23983 42789 23995 42792
rect 23937 42783 23995 42789
rect 4062 42712 4068 42764
rect 4120 42752 4126 42764
rect 4157 42755 4215 42761
rect 4157 42752 4169 42755
rect 4120 42724 4169 42752
rect 4120 42712 4126 42724
rect 4157 42721 4169 42724
rect 4203 42721 4215 42755
rect 7561 42755 7619 42761
rect 7561 42752 7573 42755
rect 4157 42715 4215 42721
rect 7116 42724 7573 42752
rect 7116 42684 7144 42724
rect 7561 42721 7573 42724
rect 7607 42752 7619 42755
rect 8110 42752 8116 42764
rect 7607 42724 8116 42752
rect 7607 42721 7619 42724
rect 7561 42715 7619 42721
rect 8110 42712 8116 42724
rect 8168 42712 8174 42764
rect 8297 42755 8355 42761
rect 8297 42721 8309 42755
rect 8343 42752 8355 42755
rect 9677 42755 9735 42761
rect 8343 42724 8800 42752
rect 8343 42721 8355 42724
rect 8297 42715 8355 42721
rect 7377 42687 7435 42693
rect 7377 42684 7389 42687
rect 2884 42656 7144 42684
rect 7208 42656 7389 42684
rect 1857 42647 1915 42653
rect 1673 42551 1731 42557
rect 1673 42517 1685 42551
rect 1719 42548 1731 42551
rect 1872 42548 1900 42647
rect 2682 42576 2688 42628
rect 2740 42616 2746 42628
rect 2740 42588 3372 42616
rect 2740 42576 2746 42588
rect 2774 42548 2780 42560
rect 1719 42520 2780 42548
rect 1719 42517 1731 42520
rect 1673 42511 1731 42517
rect 2774 42508 2780 42520
rect 2832 42508 2838 42560
rect 2961 42551 3019 42557
rect 2961 42517 2973 42551
rect 3007 42548 3019 42551
rect 3050 42548 3056 42560
rect 3007 42520 3056 42548
rect 3007 42517 3019 42520
rect 2961 42511 3019 42517
rect 3050 42508 3056 42520
rect 3108 42508 3114 42560
rect 3344 42557 3372 42588
rect 3329 42551 3387 42557
rect 3329 42517 3341 42551
rect 3375 42548 3387 42551
rect 4249 42551 4307 42557
rect 4249 42548 4261 42551
rect 3375 42520 4261 42548
rect 3375 42517 3387 42520
rect 3329 42511 3387 42517
rect 4249 42517 4261 42520
rect 4295 42548 4307 42551
rect 6546 42548 6552 42560
rect 4295 42520 6552 42548
rect 4295 42517 4307 42520
rect 4249 42511 4307 42517
rect 6546 42508 6552 42520
rect 6604 42508 6610 42560
rect 6914 42508 6920 42560
rect 6972 42548 6978 42560
rect 7208 42557 7236 42656
rect 7377 42653 7389 42656
rect 7423 42653 7435 42687
rect 7377 42647 7435 42653
rect 8018 42576 8024 42628
rect 8076 42616 8082 42628
rect 8496 42616 8524 42724
rect 8772 42684 8800 42724
rect 9677 42721 9689 42755
rect 9723 42752 9735 42755
rect 12529 42755 12587 42761
rect 12529 42752 12541 42755
rect 9723 42724 10088 42752
rect 9723 42721 9735 42724
rect 9677 42715 9735 42721
rect 9769 42687 9827 42693
rect 9769 42684 9781 42687
rect 8772 42656 9781 42684
rect 9769 42653 9781 42656
rect 9815 42653 9827 42687
rect 9769 42647 9827 42653
rect 8076 42588 8524 42616
rect 8076 42576 8082 42588
rect 10060 42560 10088 42724
rect 10796 42724 12541 42752
rect 10796 42696 10824 42724
rect 12529 42721 12541 42724
rect 12575 42752 12587 42755
rect 15470 42752 15476 42764
rect 12575 42724 15476 42752
rect 12575 42721 12587 42724
rect 12529 42715 12587 42721
rect 15470 42712 15476 42724
rect 15528 42752 15534 42764
rect 16482 42752 16488 42764
rect 15528 42724 16488 42752
rect 15528 42712 15534 42724
rect 16482 42712 16488 42724
rect 16540 42752 16546 42764
rect 16761 42755 16819 42761
rect 16761 42752 16773 42755
rect 16540 42724 16773 42752
rect 16540 42712 16546 42724
rect 16761 42721 16773 42724
rect 16807 42721 16819 42755
rect 17034 42752 17040 42764
rect 16995 42724 17040 42752
rect 16761 42715 16819 42721
rect 10778 42684 10784 42696
rect 10739 42656 10784 42684
rect 10778 42644 10784 42656
rect 10836 42644 10842 42696
rect 11057 42687 11115 42693
rect 11057 42653 11069 42687
rect 11103 42684 11115 42687
rect 11514 42684 11520 42696
rect 11103 42656 11520 42684
rect 11103 42653 11115 42656
rect 11057 42647 11115 42653
rect 11514 42644 11520 42656
rect 11572 42644 11578 42696
rect 16776 42684 16804 42715
rect 17034 42712 17040 42724
rect 17092 42712 17098 42764
rect 21376 42724 21680 42752
rect 18509 42687 18567 42693
rect 18509 42684 18521 42687
rect 16776 42656 18521 42684
rect 18509 42653 18521 42656
rect 18555 42684 18567 42687
rect 20898 42684 20904 42696
rect 18555 42656 20904 42684
rect 18555 42653 18567 42656
rect 18509 42647 18567 42653
rect 20898 42644 20904 42656
rect 20956 42684 20962 42696
rect 21269 42687 21327 42693
rect 21269 42684 21281 42687
rect 20956 42656 21281 42684
rect 20956 42644 20962 42656
rect 21269 42653 21281 42656
rect 21315 42684 21327 42687
rect 21376 42684 21404 42724
rect 21315 42656 21404 42684
rect 21315 42653 21327 42656
rect 21269 42647 21327 42653
rect 21450 42644 21456 42696
rect 21508 42684 21514 42696
rect 21545 42687 21603 42693
rect 21545 42684 21557 42687
rect 21508 42656 21557 42684
rect 21508 42644 21514 42656
rect 21545 42653 21557 42656
rect 21591 42653 21603 42687
rect 21652 42684 21680 42724
rect 22002 42712 22008 42764
rect 22060 42752 22066 42764
rect 24397 42755 24455 42761
rect 24397 42752 24409 42755
rect 22060 42724 24409 42752
rect 22060 42712 22066 42724
rect 24397 42721 24409 42724
rect 24443 42721 24455 42755
rect 24504 42752 24532 42792
rect 32048 42792 33232 42820
rect 24762 42752 24768 42764
rect 24504 42724 24768 42752
rect 24397 42715 24455 42721
rect 24762 42712 24768 42724
rect 24820 42752 24826 42764
rect 24949 42755 25007 42761
rect 24949 42752 24961 42755
rect 24820 42724 24961 42752
rect 24820 42712 24826 42724
rect 24949 42721 24961 42724
rect 24995 42721 25007 42755
rect 24949 42715 25007 42721
rect 25133 42755 25191 42761
rect 25133 42721 25145 42755
rect 25179 42752 25191 42755
rect 26973 42755 27031 42761
rect 26973 42752 26985 42755
rect 25179 42724 25452 42752
rect 25179 42721 25191 42724
rect 25133 42715 25191 42721
rect 24213 42687 24271 42693
rect 21652 42656 23152 42684
rect 21545 42647 21603 42653
rect 17696 42588 18644 42616
rect 7193 42551 7251 42557
rect 7193 42548 7205 42551
rect 6972 42520 7205 42548
rect 6972 42508 6978 42520
rect 7193 42517 7205 42520
rect 7239 42517 7251 42551
rect 7193 42511 7251 42517
rect 8573 42551 8631 42557
rect 8573 42517 8585 42551
rect 8619 42548 8631 42551
rect 8846 42548 8852 42560
rect 8619 42520 8852 42548
rect 8619 42517 8631 42520
rect 8573 42511 8631 42517
rect 8846 42508 8852 42520
rect 8904 42508 8910 42560
rect 10042 42548 10048 42560
rect 10003 42520 10048 42548
rect 10042 42508 10048 42520
rect 10100 42508 10106 42560
rect 13722 42508 13728 42560
rect 13780 42548 13786 42560
rect 17696 42548 17724 42588
rect 18322 42548 18328 42560
rect 13780 42520 17724 42548
rect 18283 42520 18328 42548
rect 13780 42508 13786 42520
rect 18322 42508 18328 42520
rect 18380 42508 18386 42560
rect 18616 42548 18644 42588
rect 23124 42560 23152 42656
rect 24213 42653 24225 42687
rect 24259 42653 24271 42687
rect 24213 42647 24271 42653
rect 21910 42548 21916 42560
rect 18616 42520 21916 42548
rect 21910 42508 21916 42520
rect 21968 42508 21974 42560
rect 22554 42508 22560 42560
rect 22612 42548 22618 42560
rect 22649 42551 22707 42557
rect 22649 42548 22661 42551
rect 22612 42520 22661 42548
rect 22612 42508 22618 42520
rect 22649 42517 22661 42520
rect 22695 42517 22707 42551
rect 23106 42548 23112 42560
rect 23067 42520 23112 42548
rect 22649 42511 22707 42517
rect 23106 42508 23112 42520
rect 23164 42508 23170 42560
rect 24026 42548 24032 42560
rect 23987 42520 24032 42548
rect 24026 42508 24032 42520
rect 24084 42548 24090 42560
rect 24228 42548 24256 42647
rect 25424 42616 25452 42724
rect 25516 42724 26985 42752
rect 25516 42693 25544 42724
rect 26973 42721 26985 42724
rect 27019 42721 27031 42755
rect 29178 42752 29184 42764
rect 26973 42715 27031 42721
rect 27632 42724 28580 42752
rect 29139 42724 29184 42752
rect 25501 42687 25559 42693
rect 25501 42653 25513 42687
rect 25547 42653 25559 42687
rect 25501 42647 25559 42653
rect 25777 42687 25835 42693
rect 25777 42653 25789 42687
rect 25823 42684 25835 42687
rect 26234 42684 26240 42696
rect 25823 42656 26240 42684
rect 25823 42653 25835 42656
rect 25777 42647 25835 42653
rect 25792 42616 25820 42647
rect 26234 42644 26240 42656
rect 26292 42644 26298 42696
rect 26694 42684 26700 42696
rect 26655 42656 26700 42684
rect 26694 42644 26700 42656
rect 26752 42644 26758 42696
rect 25424 42588 25820 42616
rect 24084 42520 24256 42548
rect 24084 42508 24090 42520
rect 24762 42508 24768 42560
rect 24820 42548 24826 42560
rect 27632 42548 27660 42724
rect 28552 42684 28580 42724
rect 29178 42712 29184 42724
rect 29236 42712 29242 42764
rect 29270 42712 29276 42764
rect 29328 42752 29334 42764
rect 32048 42752 32076 42792
rect 33226 42780 33232 42792
rect 33284 42780 33290 42832
rect 34256 42820 34284 42851
rect 33612 42792 34284 42820
rect 32214 42752 32220 42764
rect 29328 42724 32076 42752
rect 32127 42724 32220 42752
rect 29328 42712 29334 42724
rect 32214 42712 32220 42724
rect 32272 42752 32278 42764
rect 33612 42761 33640 42792
rect 32401 42755 32459 42761
rect 32401 42752 32413 42755
rect 32272 42724 32413 42752
rect 32272 42712 32278 42724
rect 32401 42721 32413 42724
rect 32447 42752 32459 42755
rect 32861 42755 32919 42761
rect 32861 42752 32873 42755
rect 32447 42724 32873 42752
rect 32447 42721 32459 42724
rect 32401 42715 32459 42721
rect 32861 42721 32873 42724
rect 32907 42752 32919 42755
rect 33413 42755 33471 42761
rect 33413 42752 33425 42755
rect 32907 42724 33425 42752
rect 32907 42721 32919 42724
rect 32861 42715 32919 42721
rect 33413 42721 33425 42724
rect 33459 42721 33471 42755
rect 33413 42715 33471 42721
rect 33597 42755 33655 42761
rect 33597 42721 33609 42755
rect 33643 42752 33655 42755
rect 35250 42752 35256 42764
rect 33643 42724 33824 42752
rect 33643 42721 33655 42724
rect 33597 42715 33655 42721
rect 31938 42684 31944 42696
rect 28552 42656 31944 42684
rect 31938 42644 31944 42656
rect 31996 42644 32002 42696
rect 32306 42644 32312 42696
rect 32364 42684 32370 42696
rect 32493 42687 32551 42693
rect 32493 42684 32505 42687
rect 32364 42656 32505 42684
rect 32364 42644 32370 42656
rect 32493 42653 32505 42656
rect 32539 42684 32551 42687
rect 32677 42687 32735 42693
rect 32677 42684 32689 42687
rect 32539 42656 32689 42684
rect 32539 42653 32551 42656
rect 32493 42647 32551 42653
rect 32677 42653 32689 42656
rect 32723 42653 32735 42687
rect 32677 42647 32735 42653
rect 27890 42576 27896 42628
rect 27948 42616 27954 42628
rect 33796 42616 33824 42724
rect 33980 42724 35112 42752
rect 35211 42724 35256 42752
rect 33980 42693 34008 42724
rect 33965 42687 34023 42693
rect 33965 42653 33977 42687
rect 34011 42653 34023 42687
rect 33965 42647 34023 42653
rect 34701 42687 34759 42693
rect 34701 42653 34713 42687
rect 34747 42684 34759 42687
rect 34974 42684 34980 42696
rect 34747 42656 34980 42684
rect 34747 42653 34759 42656
rect 34701 42647 34759 42653
rect 34974 42644 34980 42656
rect 35032 42644 35038 42696
rect 35084 42684 35112 42724
rect 35250 42712 35256 42724
rect 35308 42712 35314 42764
rect 38289 42755 38347 42761
rect 38289 42752 38301 42755
rect 37660 42724 38301 42752
rect 37660 42684 37688 42724
rect 38289 42721 38301 42724
rect 38335 42721 38347 42755
rect 38948 42752 38976 42860
rect 66898 42848 66904 42900
rect 66956 42888 66962 42900
rect 68465 42891 68523 42897
rect 68465 42888 68477 42891
rect 66956 42860 68477 42888
rect 66956 42848 66962 42860
rect 68465 42857 68477 42860
rect 68511 42857 68523 42891
rect 68465 42851 68523 42857
rect 78582 42848 78588 42900
rect 78640 42888 78646 42900
rect 81434 42888 81440 42900
rect 78640 42860 81296 42888
rect 81395 42860 81440 42888
rect 78640 42848 78646 42860
rect 45020 42792 45600 42820
rect 40126 42752 40132 42764
rect 38948 42724 40132 42752
rect 38289 42715 38347 42721
rect 40126 42712 40132 42724
rect 40184 42712 40190 42764
rect 40494 42712 40500 42764
rect 40552 42752 40558 42764
rect 44910 42752 44916 42764
rect 40552 42724 44916 42752
rect 40552 42712 40558 42724
rect 44910 42712 44916 42724
rect 44968 42712 44974 42764
rect 45020 42761 45048 42792
rect 45572 42761 45600 42792
rect 53834 42780 53840 42832
rect 53892 42820 53898 42832
rect 59998 42820 60004 42832
rect 53892 42792 55352 42820
rect 53892 42780 53898 42792
rect 45005 42755 45063 42761
rect 45005 42721 45017 42755
rect 45051 42721 45063 42755
rect 45465 42755 45523 42761
rect 45465 42752 45477 42755
rect 45005 42715 45063 42721
rect 45112 42724 45477 42752
rect 35084 42656 37688 42684
rect 37734 42644 37740 42696
rect 37792 42684 37798 42696
rect 37829 42687 37887 42693
rect 37829 42684 37841 42687
rect 37792 42656 37841 42684
rect 37792 42644 37798 42656
rect 37829 42653 37841 42656
rect 37875 42684 37887 42687
rect 38020 42687 38078 42693
rect 38020 42684 38032 42687
rect 37875 42656 38032 42684
rect 37875 42653 37887 42656
rect 37829 42647 37887 42653
rect 38020 42653 38032 42656
rect 38066 42653 38078 42687
rect 38020 42647 38078 42653
rect 38194 42644 38200 42696
rect 38252 42684 38258 42696
rect 44453 42687 44511 42693
rect 44453 42684 44465 42687
rect 38252 42656 44465 42684
rect 38252 42644 38258 42656
rect 44453 42653 44465 42656
rect 44499 42684 44511 42687
rect 44637 42687 44695 42693
rect 44637 42684 44649 42687
rect 44499 42656 44649 42684
rect 44499 42653 44511 42656
rect 44453 42647 44511 42653
rect 44637 42653 44649 42656
rect 44683 42684 44695 42687
rect 44821 42687 44879 42693
rect 44821 42684 44833 42687
rect 44683 42656 44833 42684
rect 44683 42653 44695 42656
rect 44637 42647 44695 42653
rect 44821 42653 44833 42656
rect 44867 42684 44879 42687
rect 45112 42684 45140 42724
rect 45465 42721 45477 42724
rect 45511 42721 45523 42755
rect 45465 42715 45523 42721
rect 45557 42755 45615 42761
rect 45557 42721 45569 42755
rect 45603 42752 45615 42755
rect 46385 42755 46443 42761
rect 46385 42752 46397 42755
rect 45603 42724 46397 42752
rect 45603 42721 45615 42724
rect 45557 42715 45615 42721
rect 46385 42721 46397 42724
rect 46431 42752 46443 42755
rect 46566 42752 46572 42764
rect 46431 42724 46572 42752
rect 46431 42721 46443 42724
rect 46385 42715 46443 42721
rect 46566 42712 46572 42724
rect 46624 42712 46630 42764
rect 50893 42755 50951 42761
rect 50893 42721 50905 42755
rect 50939 42752 50951 42755
rect 50985 42755 51043 42761
rect 50985 42752 50997 42755
rect 50939 42724 50997 42752
rect 50939 42721 50951 42724
rect 50893 42715 50951 42721
rect 50985 42721 50997 42724
rect 51031 42721 51043 42755
rect 51350 42752 51356 42764
rect 50985 42715 51043 42721
rect 51184 42724 51356 42752
rect 46014 42684 46020 42696
rect 44867 42656 45140 42684
rect 45975 42656 46020 42684
rect 44867 42653 44879 42656
rect 44821 42647 44879 42653
rect 46014 42644 46020 42656
rect 46072 42644 46078 42696
rect 46106 42644 46112 42696
rect 46164 42684 46170 42696
rect 50908 42684 50936 42715
rect 51184 42684 51212 42724
rect 51350 42712 51356 42724
rect 51408 42712 51414 42764
rect 53469 42755 53527 42761
rect 53469 42721 53481 42755
rect 53515 42752 53527 42755
rect 53742 42752 53748 42764
rect 53515 42724 53748 42752
rect 53515 42721 53527 42724
rect 53469 42715 53527 42721
rect 53742 42712 53748 42724
rect 53800 42712 53806 42764
rect 54573 42755 54631 42761
rect 54573 42721 54585 42755
rect 54619 42721 54631 42755
rect 54573 42715 54631 42721
rect 46164 42656 50936 42684
rect 51000 42656 51212 42684
rect 51261 42687 51319 42693
rect 46164 42644 46170 42656
rect 27948 42588 33824 42616
rect 36541 42619 36599 42625
rect 27948 42576 27954 42588
rect 36541 42585 36553 42619
rect 36587 42616 36599 42619
rect 36587 42588 38056 42616
rect 36587 42585 36599 42588
rect 36541 42579 36599 42585
rect 28442 42548 28448 42560
rect 24820 42520 27660 42548
rect 28403 42520 28448 42548
rect 24820 42508 24826 42520
rect 28442 42508 28448 42520
rect 28500 42508 28506 42560
rect 33870 42508 33876 42560
rect 33928 42548 33934 42560
rect 34701 42551 34759 42557
rect 34701 42548 34713 42551
rect 33928 42520 34713 42548
rect 33928 42508 33934 42520
rect 34701 42517 34713 42520
rect 34747 42548 34759 42551
rect 34793 42551 34851 42557
rect 34793 42548 34805 42551
rect 34747 42520 34805 42548
rect 34747 42517 34759 42520
rect 34701 42511 34759 42517
rect 34793 42517 34805 42520
rect 34839 42517 34851 42551
rect 38028 42548 38056 42588
rect 39022 42576 39028 42628
rect 39080 42616 39086 42628
rect 43530 42616 43536 42628
rect 39080 42588 43536 42616
rect 39080 42576 39086 42588
rect 43530 42576 43536 42588
rect 43588 42576 43594 42628
rect 50798 42616 50804 42628
rect 43640 42588 50804 42616
rect 39298 42548 39304 42560
rect 38028 42520 39304 42548
rect 34793 42511 34851 42517
rect 39298 42508 39304 42520
rect 39356 42508 39362 42560
rect 39574 42548 39580 42560
rect 39535 42520 39580 42548
rect 39574 42508 39580 42520
rect 39632 42508 39638 42560
rect 39666 42508 39672 42560
rect 39724 42548 39730 42560
rect 43640 42548 43668 42588
rect 50798 42576 50804 42588
rect 50856 42576 50862 42628
rect 51000 42616 51028 42656
rect 51261 42653 51273 42687
rect 51307 42684 51319 42687
rect 53561 42687 53619 42693
rect 53561 42684 53573 42687
rect 51307 42656 53573 42684
rect 51307 42653 51319 42656
rect 51261 42647 51319 42653
rect 53561 42653 53573 42656
rect 53607 42653 53619 42687
rect 54588 42684 54616 42715
rect 54662 42712 54668 42764
rect 54720 42752 54726 42764
rect 54757 42755 54815 42761
rect 54757 42752 54769 42755
rect 54720 42724 54769 42752
rect 54720 42712 54726 42724
rect 54757 42721 54769 42724
rect 54803 42752 54815 42755
rect 55217 42755 55275 42761
rect 55217 42752 55229 42755
rect 54803 42724 55229 42752
rect 54803 42721 54815 42724
rect 54757 42715 54815 42721
rect 55217 42721 55229 42724
rect 55263 42721 55275 42755
rect 55324 42752 55352 42792
rect 56980 42792 57284 42820
rect 56980 42761 57008 42792
rect 56965 42755 57023 42761
rect 56965 42752 56977 42755
rect 55324 42724 56977 42752
rect 55217 42715 55275 42721
rect 56965 42721 56977 42724
rect 57011 42721 57023 42755
rect 57146 42752 57152 42764
rect 57107 42724 57152 42752
rect 56965 42715 57023 42721
rect 57146 42712 57152 42724
rect 57204 42712 57210 42764
rect 57256 42752 57284 42792
rect 58820 42792 60004 42820
rect 57330 42752 57336 42764
rect 57243 42724 57336 42752
rect 57330 42712 57336 42724
rect 57388 42712 57394 42764
rect 58342 42712 58348 42764
rect 58400 42752 58406 42764
rect 58820 42761 58848 42792
rect 59998 42780 60004 42792
rect 60056 42780 60062 42832
rect 68480 42792 68692 42820
rect 58529 42755 58587 42761
rect 58529 42752 58541 42755
rect 58400 42724 58541 42752
rect 58400 42712 58406 42724
rect 58529 42721 58541 42724
rect 58575 42721 58587 42755
rect 58529 42715 58587 42721
rect 58805 42755 58863 42761
rect 58805 42721 58817 42755
rect 58851 42721 58863 42755
rect 60369 42755 60427 42761
rect 60369 42752 60381 42755
rect 58805 42715 58863 42721
rect 58912 42724 60381 42752
rect 54846 42684 54852 42696
rect 54588 42656 54852 42684
rect 53561 42647 53619 42653
rect 54846 42644 54852 42656
rect 54904 42684 54910 42696
rect 56873 42687 56931 42693
rect 56873 42684 56885 42687
rect 54904 42656 56885 42684
rect 54904 42644 54910 42656
rect 56873 42653 56885 42656
rect 56919 42653 56931 42687
rect 56873 42647 56931 42653
rect 57701 42687 57759 42693
rect 57701 42653 57713 42687
rect 57747 42684 57759 42687
rect 58912 42684 58940 42724
rect 60369 42721 60381 42724
rect 60415 42721 60427 42755
rect 60369 42715 60427 42721
rect 60458 42712 60464 42764
rect 60516 42752 60522 42764
rect 60516 42724 60561 42752
rect 60516 42712 60522 42724
rect 61010 42712 61016 42764
rect 61068 42752 61074 42764
rect 61749 42755 61807 42761
rect 61749 42752 61761 42755
rect 61068 42724 61761 42752
rect 61068 42712 61074 42724
rect 61749 42721 61761 42724
rect 61795 42721 61807 42755
rect 61749 42715 61807 42721
rect 63405 42755 63463 42761
rect 63405 42721 63417 42755
rect 63451 42752 63463 42755
rect 63770 42752 63776 42764
rect 63451 42724 63776 42752
rect 63451 42721 63463 42724
rect 63405 42715 63463 42721
rect 63770 42712 63776 42724
rect 63828 42712 63834 42764
rect 66165 42755 66223 42761
rect 66165 42721 66177 42755
rect 66211 42752 66223 42755
rect 66254 42752 66260 42764
rect 66211 42724 66260 42752
rect 66211 42721 66223 42724
rect 66165 42715 66223 42721
rect 66254 42712 66260 42724
rect 66312 42712 66318 42764
rect 67358 42712 67364 42764
rect 67416 42752 67422 42764
rect 68480 42752 68508 42792
rect 67416 42724 68508 42752
rect 68557 42755 68615 42761
rect 67416 42712 67422 42724
rect 68557 42721 68569 42755
rect 68603 42721 68615 42755
rect 68664 42752 68692 42792
rect 71516 42792 71728 42820
rect 68925 42755 68983 42761
rect 68925 42752 68937 42755
rect 68664 42724 68937 42752
rect 68557 42715 68615 42721
rect 68925 42721 68937 42724
rect 68971 42721 68983 42755
rect 69198 42752 69204 42764
rect 69159 42724 69204 42752
rect 68925 42715 68983 42721
rect 57747 42656 58940 42684
rect 58989 42687 59047 42693
rect 57747 42653 57759 42656
rect 57701 42647 57759 42653
rect 58989 42653 59001 42687
rect 59035 42653 59047 42687
rect 58989 42647 59047 42653
rect 58434 42616 58440 42628
rect 50908 42588 51028 42616
rect 52196 42588 58440 42616
rect 39724 42520 43668 42548
rect 39724 42508 39730 42520
rect 43714 42508 43720 42560
rect 43772 42548 43778 42560
rect 50908 42548 50936 42588
rect 43772 42520 50936 42548
rect 43772 42508 43778 42520
rect 50982 42508 50988 42560
rect 51040 42548 51046 42560
rect 52196 42548 52224 42588
rect 58434 42576 58440 42588
rect 58492 42576 58498 42628
rect 58621 42619 58679 42625
rect 58621 42585 58633 42619
rect 58667 42616 58679 42619
rect 58894 42616 58900 42628
rect 58667 42588 58900 42616
rect 58667 42585 58679 42588
rect 58621 42579 58679 42585
rect 58894 42576 58900 42588
rect 58952 42576 58958 42628
rect 52362 42548 52368 42560
rect 51040 42520 52224 42548
rect 52323 42520 52368 42548
rect 51040 42508 51046 42520
rect 52362 42508 52368 42520
rect 52420 42508 52426 42560
rect 53098 42508 53104 42560
rect 53156 42548 53162 42560
rect 54849 42551 54907 42557
rect 54849 42548 54861 42551
rect 53156 42520 54861 42548
rect 53156 42508 53162 42520
rect 54849 42517 54861 42520
rect 54895 42548 54907 42551
rect 55674 42548 55680 42560
rect 54895 42520 55680 42548
rect 54895 42517 54907 42520
rect 54849 42511 54907 42517
rect 55674 42508 55680 42520
rect 55732 42508 55738 42560
rect 56873 42551 56931 42557
rect 56873 42517 56885 42551
rect 56919 42548 56931 42551
rect 59004 42548 59032 42647
rect 59354 42644 59360 42696
rect 59412 42684 59418 42696
rect 60921 42687 60979 42693
rect 60921 42684 60933 42687
rect 59412 42656 60933 42684
rect 59412 42644 59418 42656
rect 60921 42653 60933 42656
rect 60967 42653 60979 42687
rect 60921 42647 60979 42653
rect 61102 42644 61108 42696
rect 61160 42684 61166 42696
rect 63037 42687 63095 42693
rect 63037 42684 63049 42687
rect 61160 42656 63049 42684
rect 61160 42644 61166 42656
rect 63037 42653 63049 42656
rect 63083 42684 63095 42687
rect 63129 42687 63187 42693
rect 63129 42684 63141 42687
rect 63083 42656 63141 42684
rect 63083 42653 63095 42656
rect 63037 42647 63095 42653
rect 63129 42653 63141 42656
rect 63175 42684 63187 42687
rect 65889 42687 65947 42693
rect 65889 42684 65901 42687
rect 63175 42656 65901 42684
rect 63175 42653 63187 42656
rect 63129 42647 63187 42653
rect 59630 42576 59636 42628
rect 59688 42616 59694 42628
rect 61841 42619 61899 42625
rect 61841 42616 61853 42619
rect 59688 42588 61853 42616
rect 59688 42576 59694 42588
rect 61841 42585 61853 42588
rect 61887 42585 61899 42619
rect 61841 42579 61899 42585
rect 65536 42560 65564 42656
rect 65889 42653 65901 42656
rect 65935 42653 65947 42687
rect 68572 42684 68600 42715
rect 69198 42712 69204 42724
rect 69256 42712 69262 42764
rect 71222 42712 71228 42764
rect 71280 42752 71286 42764
rect 71516 42752 71544 42792
rect 71280 42724 71544 42752
rect 71593 42755 71651 42761
rect 71280 42712 71286 42724
rect 71593 42721 71605 42755
rect 71639 42721 71651 42755
rect 71700 42752 71728 42792
rect 75546 42780 75552 42832
rect 75604 42820 75610 42832
rect 81268 42820 81296 42860
rect 81434 42848 81440 42860
rect 81492 42848 81498 42900
rect 85206 42888 85212 42900
rect 81636 42860 85212 42888
rect 81636 42820 81664 42860
rect 85206 42848 85212 42860
rect 85264 42848 85270 42900
rect 75604 42792 77064 42820
rect 81268 42792 81664 42820
rect 75604 42780 75610 42792
rect 71961 42755 72019 42761
rect 71961 42752 71973 42755
rect 71700 42724 71973 42752
rect 71593 42715 71651 42721
rect 71961 42721 71973 42724
rect 72007 42721 72019 42755
rect 73890 42752 73896 42764
rect 73851 42724 73896 42752
rect 71961 42715 72019 42721
rect 71608 42684 71636 42715
rect 73890 42712 73896 42724
rect 73948 42752 73954 42764
rect 74077 42755 74135 42761
rect 74077 42752 74089 42755
rect 73948 42724 74089 42752
rect 73948 42712 73954 42724
rect 74077 42721 74089 42724
rect 74123 42721 74135 42755
rect 74077 42715 74135 42721
rect 74353 42755 74411 42761
rect 74353 42721 74365 42755
rect 74399 42752 74411 42755
rect 74626 42752 74632 42764
rect 74399 42724 74632 42752
rect 74399 42721 74411 42724
rect 74353 42715 74411 42721
rect 74626 42712 74632 42724
rect 74684 42712 74690 42764
rect 77036 42761 77064 42792
rect 77021 42755 77079 42761
rect 77021 42721 77033 42755
rect 77067 42752 77079 42755
rect 77297 42755 77355 42761
rect 77297 42752 77309 42755
rect 77067 42724 77309 42752
rect 77067 42721 77079 42724
rect 77021 42715 77079 42721
rect 77297 42721 77309 42724
rect 77343 42721 77355 42755
rect 77297 42715 77355 42721
rect 81161 42755 81219 42761
rect 81161 42721 81173 42755
rect 81207 42721 81219 42755
rect 81161 42715 81219 42721
rect 81345 42755 81403 42761
rect 81345 42721 81357 42755
rect 81391 42752 81403 42755
rect 81434 42752 81440 42764
rect 81391 42724 81440 42752
rect 81391 42721 81403 42724
rect 81345 42715 81403 42721
rect 65889 42647 65947 42653
rect 68480 42656 68600 42684
rect 69676 42656 71636 42684
rect 56919 42520 59032 42548
rect 56919 42517 56931 42520
rect 56873 42511 56931 42517
rect 60090 42508 60096 42560
rect 60148 42548 60154 42560
rect 60185 42551 60243 42557
rect 60185 42548 60197 42551
rect 60148 42520 60197 42548
rect 60148 42508 60154 42520
rect 60185 42517 60197 42520
rect 60231 42548 60243 42551
rect 61013 42551 61071 42557
rect 61013 42548 61025 42551
rect 60231 42520 61025 42548
rect 60231 42517 60243 42520
rect 60185 42511 60243 42517
rect 61013 42517 61025 42520
rect 61059 42548 61071 42551
rect 63586 42548 63592 42560
rect 61059 42520 63592 42548
rect 61059 42517 61071 42520
rect 61013 42511 61071 42517
rect 63586 42508 63592 42520
rect 63644 42508 63650 42560
rect 64230 42508 64236 42560
rect 64288 42548 64294 42560
rect 64509 42551 64567 42557
rect 64509 42548 64521 42551
rect 64288 42520 64521 42548
rect 64288 42508 64294 42520
rect 64509 42517 64521 42520
rect 64555 42517 64567 42551
rect 65518 42548 65524 42560
rect 65479 42520 65524 42548
rect 64509 42511 64567 42517
rect 65518 42508 65524 42520
rect 65576 42508 65582 42560
rect 67266 42548 67272 42560
rect 67227 42520 67272 42548
rect 67266 42508 67272 42520
rect 67324 42508 67330 42560
rect 68480 42548 68508 42656
rect 69569 42551 69627 42557
rect 69569 42548 69581 42551
rect 68480 42520 69581 42548
rect 69569 42517 69581 42520
rect 69615 42548 69627 42551
rect 69676 42548 69704 42656
rect 71498 42616 71504 42628
rect 71459 42588 71504 42616
rect 71498 42576 71504 42588
rect 71556 42576 71562 42628
rect 71222 42548 71228 42560
rect 69615 42520 69704 42548
rect 71183 42520 71228 42548
rect 69615 42517 69627 42520
rect 69569 42511 69627 42517
rect 71222 42508 71228 42520
rect 71280 42508 71286 42560
rect 71608 42548 71636 42656
rect 72421 42687 72479 42693
rect 72421 42653 72433 42687
rect 72467 42684 72479 42687
rect 73246 42684 73252 42696
rect 72467 42656 73252 42684
rect 72467 42653 72479 42656
rect 72421 42647 72479 42653
rect 73246 42644 73252 42656
rect 73304 42644 73310 42696
rect 78585 42687 78643 42693
rect 78585 42684 78597 42687
rect 78416 42656 78597 42684
rect 77113 42619 77171 42625
rect 77113 42585 77125 42619
rect 77159 42616 77171 42619
rect 77662 42616 77668 42628
rect 77159 42588 77668 42616
rect 77159 42585 77171 42588
rect 77113 42579 77171 42585
rect 77662 42576 77668 42588
rect 77720 42576 77726 42628
rect 72694 42548 72700 42560
rect 71608 42520 72700 42548
rect 72694 42508 72700 42520
rect 72752 42508 72758 42560
rect 73430 42508 73436 42560
rect 73488 42548 73494 42560
rect 74074 42548 74080 42560
rect 73488 42520 74080 42548
rect 73488 42508 73494 42520
rect 74074 42508 74080 42520
rect 74132 42548 74138 42560
rect 75457 42551 75515 42557
rect 75457 42548 75469 42551
rect 74132 42520 75469 42548
rect 74132 42508 74138 42520
rect 75457 42517 75469 42520
rect 75503 42517 75515 42551
rect 75457 42511 75515 42517
rect 78306 42508 78312 42560
rect 78364 42548 78370 42560
rect 78416 42557 78444 42656
rect 78585 42653 78597 42656
rect 78631 42653 78643 42687
rect 78585 42647 78643 42653
rect 78766 42644 78772 42696
rect 78824 42684 78830 42696
rect 78861 42687 78919 42693
rect 78861 42684 78873 42687
rect 78824 42656 78873 42684
rect 78824 42644 78830 42656
rect 78861 42653 78873 42656
rect 78907 42653 78919 42687
rect 81176 42684 81204 42715
rect 81434 42712 81440 42724
rect 81492 42712 81498 42764
rect 82814 42712 82820 42764
rect 82872 42752 82878 42764
rect 83001 42755 83059 42761
rect 83001 42752 83013 42755
rect 82872 42724 83013 42752
rect 82872 42712 82878 42724
rect 83001 42721 83013 42724
rect 83047 42721 83059 42755
rect 83001 42715 83059 42721
rect 81986 42684 81992 42696
rect 81176 42656 81992 42684
rect 78861 42647 78919 42653
rect 81986 42644 81992 42656
rect 82044 42644 82050 42696
rect 82449 42687 82507 42693
rect 82449 42653 82461 42687
rect 82495 42684 82507 42687
rect 82722 42684 82728 42696
rect 82495 42656 82728 42684
rect 82495 42653 82507 42656
rect 82449 42647 82507 42653
rect 82464 42616 82492 42647
rect 82722 42644 82728 42656
rect 82780 42644 82786 42696
rect 79520 42588 82492 42616
rect 78401 42551 78459 42557
rect 78401 42548 78413 42551
rect 78364 42520 78413 42548
rect 78364 42508 78370 42520
rect 78401 42517 78413 42520
rect 78447 42548 78459 42551
rect 79520 42548 79548 42588
rect 78447 42520 79548 42548
rect 78447 42517 78459 42520
rect 78401 42511 78459 42517
rect 79870 42508 79876 42560
rect 79928 42548 79934 42560
rect 79965 42551 80023 42557
rect 79965 42548 79977 42551
rect 79928 42520 79977 42548
rect 79928 42508 79934 42520
rect 79965 42517 79977 42520
rect 80011 42517 80023 42551
rect 79965 42511 80023 42517
rect 82998 42508 83004 42560
rect 83056 42548 83062 42560
rect 83826 42548 83832 42560
rect 83056 42520 83832 42548
rect 83056 42508 83062 42520
rect 83826 42508 83832 42520
rect 83884 42548 83890 42560
rect 84289 42551 84347 42557
rect 84289 42548 84301 42551
rect 83884 42520 84301 42548
rect 83884 42508 83890 42520
rect 84289 42517 84301 42520
rect 84335 42517 84347 42551
rect 84289 42511 84347 42517
rect 1104 42458 105616 42480
rect 1104 42406 4246 42458
rect 4298 42406 4310 42458
rect 4362 42406 4374 42458
rect 4426 42406 4438 42458
rect 4490 42406 34966 42458
rect 35018 42406 35030 42458
rect 35082 42406 35094 42458
rect 35146 42406 35158 42458
rect 35210 42406 65686 42458
rect 65738 42406 65750 42458
rect 65802 42406 65814 42458
rect 65866 42406 65878 42458
rect 65930 42406 96406 42458
rect 96458 42406 96470 42458
rect 96522 42406 96534 42458
rect 96586 42406 96598 42458
rect 96650 42406 105616 42458
rect 1104 42384 105616 42406
rect 4062 42304 4068 42356
rect 4120 42344 4126 42356
rect 4157 42347 4215 42353
rect 4157 42344 4169 42347
rect 4120 42316 4169 42344
rect 4120 42304 4126 42316
rect 4157 42313 4169 42316
rect 4203 42313 4215 42347
rect 11790 42344 11796 42356
rect 4157 42307 4215 42313
rect 4264 42316 11796 42344
rect 3050 42208 3056 42220
rect 3011 42180 3056 42208
rect 3050 42168 3056 42180
rect 3108 42168 3114 42220
rect 3694 42168 3700 42220
rect 3752 42208 3758 42220
rect 4264 42208 4292 42316
rect 11790 42304 11796 42316
rect 11848 42304 11854 42356
rect 21818 42344 21824 42356
rect 15396 42316 21824 42344
rect 8570 42208 8576 42220
rect 3752 42180 4292 42208
rect 8531 42180 8576 42208
rect 3752 42168 3758 42180
rect 8570 42168 8576 42180
rect 8628 42168 8634 42220
rect 8846 42208 8852 42220
rect 8807 42180 8852 42208
rect 8846 42168 8852 42180
rect 8904 42168 8910 42220
rect 10042 42168 10048 42220
rect 10100 42208 10106 42220
rect 10229 42211 10287 42217
rect 10229 42208 10241 42211
rect 10100 42180 10241 42208
rect 10100 42168 10106 42180
rect 10229 42177 10241 42180
rect 10275 42208 10287 42211
rect 15396 42208 15424 42316
rect 21818 42304 21824 42316
rect 21876 42304 21882 42356
rect 21910 42304 21916 42356
rect 21968 42344 21974 42356
rect 38654 42344 38660 42356
rect 21968 42316 38660 42344
rect 21968 42304 21974 42316
rect 38654 42304 38660 42316
rect 38712 42304 38718 42356
rect 38749 42347 38807 42353
rect 38749 42313 38761 42347
rect 38795 42344 38807 42347
rect 38933 42347 38991 42353
rect 38933 42344 38945 42347
rect 38795 42316 38945 42344
rect 38795 42313 38807 42316
rect 38749 42307 38807 42313
rect 38933 42313 38945 42316
rect 38979 42344 38991 42347
rect 39022 42344 39028 42356
rect 38979 42316 39028 42344
rect 38979 42313 38991 42316
rect 38933 42307 38991 42313
rect 16666 42276 16672 42288
rect 16627 42248 16672 42276
rect 16666 42236 16672 42248
rect 16724 42236 16730 42288
rect 21174 42276 21180 42288
rect 18156 42248 21180 42276
rect 10275 42180 15424 42208
rect 15473 42211 15531 42217
rect 10275 42177 10287 42180
rect 10229 42171 10287 42177
rect 15473 42177 15485 42211
rect 15519 42208 15531 42211
rect 15654 42208 15660 42220
rect 15519 42180 15660 42208
rect 15519 42177 15531 42180
rect 15473 42171 15531 42177
rect 15654 42168 15660 42180
rect 15712 42168 15718 42220
rect 16758 42168 16764 42220
rect 16816 42208 16822 42220
rect 17129 42211 17187 42217
rect 17129 42208 17141 42211
rect 16816 42180 17141 42208
rect 16816 42168 16822 42180
rect 17129 42177 17141 42180
rect 17175 42208 17187 42211
rect 18046 42208 18052 42220
rect 17175 42180 18052 42208
rect 17175 42177 17187 42180
rect 17129 42171 17187 42177
rect 18046 42168 18052 42180
rect 18104 42168 18110 42220
rect 2777 42143 2835 42149
rect 2777 42109 2789 42143
rect 2823 42109 2835 42143
rect 8588 42140 8616 42168
rect 10321 42143 10379 42149
rect 10321 42140 10333 42143
rect 8588 42112 10333 42140
rect 2777 42103 2835 42109
rect 10321 42109 10333 42112
rect 10367 42140 10379 42143
rect 10778 42140 10784 42152
rect 10367 42112 10784 42140
rect 10367 42109 10379 42112
rect 10321 42103 10379 42109
rect 2792 42004 2820 42103
rect 10778 42100 10784 42112
rect 10836 42100 10842 42152
rect 11057 42143 11115 42149
rect 11057 42109 11069 42143
rect 11103 42140 11115 42143
rect 15749 42143 15807 42149
rect 11103 42112 11468 42140
rect 11103 42109 11115 42112
rect 11057 42103 11115 42109
rect 11440 42016 11468 42112
rect 15749 42109 15761 42143
rect 15795 42109 15807 42143
rect 16206 42140 16212 42152
rect 16167 42112 16212 42140
rect 15749 42103 15807 42109
rect 15764 42072 15792 42103
rect 16206 42100 16212 42112
rect 16264 42100 16270 42152
rect 16301 42143 16359 42149
rect 16301 42109 16313 42143
rect 16347 42140 16359 42143
rect 18156 42140 18184 42248
rect 21174 42236 21180 42248
rect 21232 42236 21238 42288
rect 21358 42236 21364 42288
rect 21416 42276 21422 42288
rect 36817 42279 36875 42285
rect 36817 42276 36829 42279
rect 21416 42248 36829 42276
rect 21416 42236 21422 42248
rect 36817 42245 36829 42248
rect 36863 42276 36875 42279
rect 37001 42279 37059 42285
rect 37001 42276 37013 42279
rect 36863 42248 37013 42276
rect 36863 42245 36875 42248
rect 36817 42239 36875 42245
rect 37001 42245 37013 42248
rect 37047 42276 37059 42279
rect 37047 42248 37228 42276
rect 37047 42245 37059 42248
rect 37001 42239 37059 42245
rect 18414 42208 18420 42220
rect 18375 42180 18420 42208
rect 18414 42168 18420 42180
rect 18472 42168 18478 42220
rect 27154 42208 27160 42220
rect 18892 42180 20300 42208
rect 27115 42180 27160 42208
rect 18322 42140 18328 42152
rect 16347 42112 18184 42140
rect 18283 42112 18328 42140
rect 16347 42109 16359 42112
rect 16301 42103 16359 42109
rect 16316 42072 16344 42103
rect 18322 42100 18328 42112
rect 18380 42100 18386 42152
rect 15764 42044 16344 42072
rect 16942 42032 16948 42084
rect 17000 42072 17006 42084
rect 18432 42072 18460 42168
rect 17000 42044 18460 42072
rect 17000 42032 17006 42044
rect 4617 42007 4675 42013
rect 4617 42004 4629 42007
rect 2792 41976 4629 42004
rect 4617 41973 4629 41976
rect 4663 42004 4675 42007
rect 4798 42004 4804 42016
rect 4663 41976 4804 42004
rect 4663 41973 4675 41976
rect 4617 41967 4675 41973
rect 4798 41964 4804 41976
rect 4856 41964 4862 42016
rect 10502 41964 10508 42016
rect 10560 42004 10566 42016
rect 11241 42007 11299 42013
rect 11241 42004 11253 42007
rect 10560 41976 11253 42004
rect 10560 41964 10566 41976
rect 11241 41973 11253 41976
rect 11287 41973 11299 42007
rect 11422 42004 11428 42016
rect 11383 41976 11428 42004
rect 11241 41967 11299 41973
rect 11422 41964 11428 41976
rect 11480 41964 11486 42016
rect 16206 41964 16212 42016
rect 16264 42004 16270 42016
rect 16758 42004 16764 42016
rect 16264 41976 16764 42004
rect 16264 41964 16270 41976
rect 16758 41964 16764 41976
rect 16816 41964 16822 42016
rect 17862 41964 17868 42016
rect 17920 42004 17926 42016
rect 18892 42004 18920 42180
rect 20272 42149 20300 42180
rect 27154 42168 27160 42180
rect 27212 42168 27218 42220
rect 32125 42211 32183 42217
rect 32125 42177 32137 42211
rect 32171 42208 32183 42211
rect 32214 42208 32220 42220
rect 32171 42180 32220 42208
rect 32171 42177 32183 42180
rect 32125 42171 32183 42177
rect 32214 42168 32220 42180
rect 32272 42168 32278 42220
rect 32582 42208 32588 42220
rect 32543 42180 32588 42208
rect 32582 42168 32588 42180
rect 32640 42168 32646 42220
rect 32784 42180 32996 42208
rect 20073 42143 20131 42149
rect 20073 42109 20085 42143
rect 20119 42109 20131 42143
rect 20073 42103 20131 42109
rect 20257 42143 20315 42149
rect 20257 42109 20269 42143
rect 20303 42140 20315 42143
rect 20809 42143 20867 42149
rect 20809 42140 20821 42143
rect 20303 42112 20821 42140
rect 20303 42109 20315 42112
rect 20257 42103 20315 42109
rect 20809 42109 20821 42112
rect 20855 42109 20867 42143
rect 20809 42103 20867 42109
rect 20993 42143 21051 42149
rect 20993 42109 21005 42143
rect 21039 42140 21051 42143
rect 22554 42140 22560 42152
rect 21039 42112 21680 42140
rect 22515 42112 22560 42140
rect 21039 42109 21051 42112
rect 20993 42103 21051 42109
rect 17920 41976 18920 42004
rect 19981 42007 20039 42013
rect 17920 41964 17926 41976
rect 19981 41973 19993 42007
rect 20027 42004 20039 42007
rect 20088 42004 20116 42103
rect 20824 42072 20852 42103
rect 21542 42072 21548 42084
rect 20824 42044 21548 42072
rect 21542 42032 21548 42044
rect 21600 42032 21606 42084
rect 20162 42004 20168 42016
rect 20027 41976 20168 42004
rect 20027 41973 20039 41976
rect 19981 41967 20039 41973
rect 20162 41964 20168 41976
rect 20220 41964 20226 42016
rect 21174 41964 21180 42016
rect 21232 42004 21238 42016
rect 21652 42013 21680 42112
rect 22554 42100 22560 42112
rect 22612 42100 22618 42152
rect 24026 42100 24032 42152
rect 24084 42140 24090 42152
rect 25777 42143 25835 42149
rect 25777 42140 25789 42143
rect 24084 42112 25789 42140
rect 24084 42100 24090 42112
rect 25777 42109 25789 42112
rect 25823 42140 25835 42143
rect 25961 42143 26019 42149
rect 25961 42140 25973 42143
rect 25823 42112 25973 42140
rect 25823 42109 25835 42112
rect 25777 42103 25835 42109
rect 25961 42109 25973 42112
rect 26007 42109 26019 42143
rect 25961 42103 26019 42109
rect 26050 42100 26056 42152
rect 26108 42140 26114 42152
rect 26145 42143 26203 42149
rect 26145 42140 26157 42143
rect 26108 42112 26157 42140
rect 26108 42100 26114 42112
rect 26145 42109 26157 42112
rect 26191 42109 26203 42143
rect 26602 42140 26608 42152
rect 26563 42112 26608 42140
rect 26145 42103 26203 42109
rect 26602 42100 26608 42112
rect 26660 42100 26666 42152
rect 26694 42100 26700 42152
rect 26752 42140 26758 42152
rect 32232 42140 32260 42168
rect 32784 42149 32812 42180
rect 32769 42143 32827 42149
rect 32769 42140 32781 42143
rect 26752 42112 32781 42140
rect 26752 42100 26758 42112
rect 32769 42109 32781 42112
rect 32815 42109 32827 42143
rect 32968 42140 32996 42180
rect 34146 42168 34152 42220
rect 34204 42208 34210 42220
rect 37090 42208 37096 42220
rect 34204 42180 37096 42208
rect 34204 42168 34210 42180
rect 37090 42168 37096 42180
rect 37148 42168 37154 42220
rect 37200 42217 37228 42248
rect 37366 42236 37372 42288
rect 37424 42276 37430 42288
rect 38764 42276 38792 42307
rect 39022 42304 39028 42316
rect 39080 42304 39086 42356
rect 39114 42304 39120 42356
rect 39172 42344 39178 42356
rect 39485 42347 39543 42353
rect 39485 42344 39497 42347
rect 39172 42316 39497 42344
rect 39172 42304 39178 42316
rect 39485 42313 39497 42316
rect 39531 42344 39543 42347
rect 39531 42316 40632 42344
rect 39531 42313 39543 42316
rect 39485 42307 39543 42313
rect 37424 42248 38792 42276
rect 37424 42236 37430 42248
rect 37185 42211 37243 42217
rect 37185 42177 37197 42211
rect 37231 42208 37243 42211
rect 37231 42180 37504 42208
rect 37231 42177 37243 42180
rect 37185 42171 37243 42177
rect 33321 42143 33379 42149
rect 33321 42140 33333 42143
rect 32968 42112 33333 42140
rect 32769 42103 32827 42109
rect 33321 42109 33333 42112
rect 33367 42109 33379 42143
rect 33502 42140 33508 42152
rect 33463 42112 33508 42140
rect 33321 42103 33379 42109
rect 33502 42100 33508 42112
rect 33560 42140 33566 42152
rect 34333 42143 34391 42149
rect 34333 42140 34345 42143
rect 33560 42112 34345 42140
rect 33560 42100 33566 42112
rect 34333 42109 34345 42112
rect 34379 42140 34391 42143
rect 34422 42140 34428 42152
rect 34379 42112 34428 42140
rect 34379 42109 34391 42112
rect 34333 42103 34391 42109
rect 34422 42100 34428 42112
rect 34480 42100 34486 42152
rect 37366 42140 37372 42152
rect 37327 42112 37372 42140
rect 37366 42100 37372 42112
rect 37424 42100 37430 42152
rect 37476 42140 37504 42180
rect 37829 42143 37887 42149
rect 37829 42140 37841 42143
rect 37476 42112 37841 42140
rect 37829 42109 37841 42112
rect 37875 42109 37887 42143
rect 37829 42103 37887 42109
rect 37921 42143 37979 42149
rect 37921 42109 37933 42143
rect 37967 42140 37979 42143
rect 38396 42140 38424 42248
rect 39390 42236 39396 42288
rect 39448 42276 39454 42288
rect 40604 42276 40632 42316
rect 40954 42304 40960 42356
rect 41012 42344 41018 42356
rect 41969 42347 42027 42353
rect 41969 42344 41981 42347
rect 41012 42316 41981 42344
rect 41012 42304 41018 42316
rect 41969 42313 41981 42316
rect 42015 42344 42027 42347
rect 42015 42316 43024 42344
rect 42015 42313 42027 42316
rect 41969 42307 42027 42313
rect 41874 42276 41880 42288
rect 39448 42248 40540 42276
rect 40604 42248 41880 42276
rect 39448 42236 39454 42248
rect 38473 42211 38531 42217
rect 38473 42177 38485 42211
rect 38519 42208 38531 42211
rect 40402 42208 40408 42220
rect 38519 42180 40408 42208
rect 38519 42177 38531 42180
rect 38473 42171 38531 42177
rect 40402 42168 40408 42180
rect 40460 42168 40466 42220
rect 40512 42208 40540 42248
rect 41874 42236 41880 42248
rect 41932 42236 41938 42288
rect 41966 42208 41972 42220
rect 40512 42180 41972 42208
rect 41966 42168 41972 42180
rect 42024 42168 42030 42220
rect 42076 42217 42104 42316
rect 42996 42276 43024 42316
rect 43530 42304 43536 42356
rect 43588 42344 43594 42356
rect 48866 42344 48872 42356
rect 43588 42316 48872 42344
rect 43588 42304 43594 42316
rect 48866 42304 48872 42316
rect 48924 42304 48930 42356
rect 53742 42344 53748 42356
rect 53703 42316 53748 42344
rect 53742 42304 53748 42316
rect 53800 42304 53806 42356
rect 81069 42347 81127 42353
rect 53852 42316 81020 42344
rect 46106 42276 46112 42288
rect 42996 42248 46112 42276
rect 46106 42236 46112 42248
rect 46164 42236 46170 42288
rect 53852 42276 53880 42316
rect 46216 42248 53880 42276
rect 42061 42211 42119 42217
rect 42061 42177 42073 42211
rect 42107 42177 42119 42211
rect 42061 42171 42119 42177
rect 42242 42168 42248 42220
rect 42300 42208 42306 42220
rect 46216 42208 46244 42248
rect 58526 42236 58532 42288
rect 58584 42276 58590 42288
rect 59081 42279 59139 42285
rect 59081 42276 59093 42279
rect 58584 42248 59093 42276
rect 58584 42236 58590 42248
rect 59081 42245 59093 42248
rect 59127 42245 59139 42279
rect 59081 42239 59139 42245
rect 59170 42236 59176 42288
rect 59228 42276 59234 42288
rect 61194 42276 61200 42288
rect 59228 42248 61200 42276
rect 59228 42236 59234 42248
rect 61194 42236 61200 42248
rect 61252 42236 61258 42288
rect 66714 42276 66720 42288
rect 63696 42248 65380 42276
rect 66627 42248 66720 42276
rect 42300 42180 46244 42208
rect 42300 42168 42306 42180
rect 49142 42168 49148 42220
rect 49200 42208 49206 42220
rect 63696 42208 63724 42248
rect 63862 42208 63868 42220
rect 49200 42180 63724 42208
rect 63823 42180 63868 42208
rect 49200 42168 49206 42180
rect 63862 42168 63868 42180
rect 63920 42168 63926 42220
rect 64414 42168 64420 42220
rect 64472 42208 64478 42220
rect 64472 42180 65288 42208
rect 64472 42168 64478 42180
rect 37967 42112 38424 42140
rect 37967 42109 37979 42112
rect 37921 42103 37979 42109
rect 39298 42100 39304 42152
rect 39356 42140 39362 42152
rect 39393 42143 39451 42149
rect 39393 42140 39405 42143
rect 39356 42112 39405 42140
rect 39356 42100 39362 42112
rect 39393 42109 39405 42112
rect 39439 42109 39451 42143
rect 39393 42103 39451 42109
rect 39574 42100 39580 42152
rect 39632 42140 39638 42152
rect 39850 42140 39856 42152
rect 39632 42112 39856 42140
rect 39632 42100 39638 42112
rect 39850 42100 39856 42112
rect 39908 42140 39914 42152
rect 40497 42143 40555 42149
rect 40497 42140 40509 42143
rect 39908 42112 40509 42140
rect 39908 42100 39914 42112
rect 40497 42109 40509 42112
rect 40543 42109 40555 42143
rect 42337 42143 42395 42149
rect 42337 42140 42349 42143
rect 40497 42103 40555 42109
rect 40604 42112 42349 42140
rect 30742 42032 30748 42084
rect 30800 42072 30806 42084
rect 33134 42072 33140 42084
rect 30800 42044 33140 42072
rect 30800 42032 30806 42044
rect 33134 42032 33140 42044
rect 33192 42032 33198 42084
rect 33873 42075 33931 42081
rect 33873 42041 33885 42075
rect 33919 42072 33931 42075
rect 40604 42072 40632 42112
rect 42337 42109 42349 42112
rect 42383 42109 42395 42143
rect 42337 42103 42395 42109
rect 43717 42143 43775 42149
rect 43717 42109 43729 42143
rect 43763 42140 43775 42143
rect 43898 42140 43904 42152
rect 43763 42112 43904 42140
rect 43763 42109 43775 42112
rect 43717 42103 43775 42109
rect 43898 42100 43904 42112
rect 43956 42140 43962 42152
rect 44545 42143 44603 42149
rect 44545 42140 44557 42143
rect 43956 42112 44557 42140
rect 43956 42100 43962 42112
rect 44545 42109 44557 42112
rect 44591 42109 44603 42143
rect 44545 42103 44603 42109
rect 44910 42100 44916 42152
rect 44968 42140 44974 42152
rect 47581 42143 47639 42149
rect 47581 42140 47593 42143
rect 44968 42112 47593 42140
rect 44968 42100 44974 42112
rect 47581 42109 47593 42112
rect 47627 42140 47639 42143
rect 47949 42143 48007 42149
rect 47949 42140 47961 42143
rect 47627 42112 47961 42140
rect 47627 42109 47639 42112
rect 47581 42103 47639 42109
rect 47949 42109 47961 42112
rect 47995 42109 48007 42143
rect 47949 42103 48007 42109
rect 48133 42143 48191 42149
rect 48133 42109 48145 42143
rect 48179 42140 48191 42143
rect 48314 42140 48320 42152
rect 48179 42112 48320 42140
rect 48179 42109 48191 42112
rect 48133 42103 48191 42109
rect 48314 42100 48320 42112
rect 48372 42100 48378 42152
rect 48590 42140 48596 42152
rect 48503 42112 48596 42140
rect 47762 42072 47768 42084
rect 33919 42044 40632 42072
rect 44100 42044 47768 42072
rect 33919 42041 33931 42044
rect 33873 42035 33931 42041
rect 21269 42007 21327 42013
rect 21269 42004 21281 42007
rect 21232 41976 21281 42004
rect 21232 41964 21238 41976
rect 21269 41973 21281 41976
rect 21315 41973 21327 42007
rect 21269 41967 21327 41973
rect 21637 42007 21695 42013
rect 21637 41973 21649 42007
rect 21683 42004 21695 42007
rect 21726 42004 21732 42016
rect 21683 41976 21732 42004
rect 21683 41973 21695 41976
rect 21637 41967 21695 41973
rect 21726 41964 21732 41976
rect 21784 41964 21790 42016
rect 22094 41964 22100 42016
rect 22152 42004 22158 42016
rect 22649 42007 22707 42013
rect 22649 42004 22661 42007
rect 22152 41976 22661 42004
rect 22152 41964 22158 41976
rect 22649 41973 22661 41976
rect 22695 41973 22707 42007
rect 22649 41967 22707 41973
rect 22830 41964 22836 42016
rect 22888 42004 22894 42016
rect 25682 42004 25688 42016
rect 22888 41976 25688 42004
rect 22888 41964 22894 41976
rect 25682 41964 25688 41976
rect 25740 41964 25746 42016
rect 25774 41964 25780 42016
rect 25832 42004 25838 42016
rect 26602 42004 26608 42016
rect 25832 41976 26608 42004
rect 25832 41964 25838 41976
rect 26602 41964 26608 41976
rect 26660 42004 26666 42016
rect 27525 42007 27583 42013
rect 27525 42004 27537 42007
rect 26660 41976 27537 42004
rect 26660 41964 26666 41976
rect 27525 41973 27537 41976
rect 27571 42004 27583 42007
rect 29362 42004 29368 42016
rect 27571 41976 29368 42004
rect 27571 41973 27583 41976
rect 27525 41967 27583 41973
rect 29362 41964 29368 41976
rect 29420 41964 29426 42016
rect 32122 41964 32128 42016
rect 32180 42004 32186 42016
rect 32401 42007 32459 42013
rect 32401 42004 32413 42007
rect 32180 41976 32413 42004
rect 32180 41964 32186 41976
rect 32401 41973 32413 41976
rect 32447 42004 32459 42007
rect 32582 42004 32588 42016
rect 32447 41976 32588 42004
rect 32447 41973 32459 41976
rect 32401 41967 32459 41973
rect 32582 41964 32588 41976
rect 32640 42004 32646 42016
rect 34149 42007 34207 42013
rect 34149 42004 34161 42007
rect 32640 41976 34161 42004
rect 32640 41964 32646 41976
rect 34149 41973 34161 41976
rect 34195 42004 34207 42007
rect 34330 42004 34336 42016
rect 34195 41976 34336 42004
rect 34195 41973 34207 41976
rect 34149 41967 34207 41973
rect 34330 41964 34336 41976
rect 34388 41964 34394 42016
rect 35526 41964 35532 42016
rect 35584 42004 35590 42016
rect 40034 42004 40040 42016
rect 35584 41976 40040 42004
rect 35584 41964 35590 41976
rect 40034 41964 40040 41976
rect 40092 41964 40098 42016
rect 40126 41964 40132 42016
rect 40184 42004 40190 42016
rect 40586 42004 40592 42016
rect 40184 41976 40592 42004
rect 40184 41964 40190 41976
rect 40586 41964 40592 41976
rect 40644 41964 40650 42016
rect 41874 41964 41880 42016
rect 41932 42004 41938 42016
rect 44100 42004 44128 42044
rect 47762 42032 47768 42044
rect 47820 42032 47826 42084
rect 48516 42072 48544 42112
rect 48590 42100 48596 42112
rect 48648 42100 48654 42152
rect 48685 42143 48743 42149
rect 48685 42109 48697 42143
rect 48731 42140 48743 42143
rect 49605 42143 49663 42149
rect 49605 42140 49617 42143
rect 48731 42112 49617 42140
rect 48731 42109 48743 42112
rect 48685 42103 48743 42109
rect 49605 42109 49617 42112
rect 49651 42140 49663 42143
rect 50062 42140 50068 42152
rect 49651 42112 50068 42140
rect 49651 42109 49663 42112
rect 49605 42103 49663 42109
rect 48424 42044 48544 42072
rect 41932 41976 44128 42004
rect 41932 41964 41938 41976
rect 44174 41964 44180 42016
rect 44232 42004 44238 42016
rect 44637 42007 44695 42013
rect 44637 42004 44649 42007
rect 44232 41976 44649 42004
rect 44232 41964 44238 41976
rect 44637 41973 44649 41976
rect 44683 42004 44695 42007
rect 45186 42004 45192 42016
rect 44683 41976 45192 42004
rect 44683 41973 44695 41976
rect 44637 41967 44695 41973
rect 45186 41964 45192 41976
rect 45244 41964 45250 42016
rect 47857 42007 47915 42013
rect 47857 41973 47869 42007
rect 47903 42004 47915 42007
rect 48424 42004 48452 42044
rect 47903 41976 48452 42004
rect 47903 41973 47915 41976
rect 47857 41967 47915 41973
rect 48498 41964 48504 42016
rect 48556 42004 48562 42016
rect 48700 42004 48728 42103
rect 50062 42100 50068 42112
rect 50120 42100 50126 42152
rect 51721 42143 51779 42149
rect 51721 42140 51733 42143
rect 50264 42112 51733 42140
rect 49237 42075 49295 42081
rect 49237 42041 49249 42075
rect 49283 42072 49295 42075
rect 49694 42072 49700 42084
rect 49283 42044 49700 42072
rect 49283 42041 49295 42044
rect 49237 42035 49295 42041
rect 49694 42032 49700 42044
rect 49752 42032 49758 42084
rect 49510 42004 49516 42016
rect 48556 41976 48728 42004
rect 49471 41976 49516 42004
rect 48556 41964 48562 41976
rect 49510 41964 49516 41976
rect 49568 41964 49574 42016
rect 49602 41964 49608 42016
rect 49660 42004 49666 42016
rect 50264 42004 50292 42112
rect 51721 42109 51733 42112
rect 51767 42140 51779 42143
rect 52362 42140 52368 42152
rect 51767 42112 52368 42140
rect 51767 42109 51779 42112
rect 51721 42103 51779 42109
rect 52362 42100 52368 42112
rect 52420 42100 52426 42152
rect 54297 42143 54355 42149
rect 54297 42109 54309 42143
rect 54343 42109 54355 42143
rect 54297 42103 54355 42109
rect 54389 42143 54447 42149
rect 54389 42109 54401 42143
rect 54435 42109 54447 42143
rect 54389 42103 54447 42109
rect 49660 41976 50292 42004
rect 49660 41964 49666 41976
rect 51074 41964 51080 42016
rect 51132 42004 51138 42016
rect 51813 42007 51871 42013
rect 51813 42004 51825 42007
rect 51132 41976 51825 42004
rect 51132 41964 51138 41976
rect 51813 41973 51825 41976
rect 51859 42004 51871 42007
rect 53469 42007 53527 42013
rect 53469 42004 53481 42007
rect 51859 41976 53481 42004
rect 51859 41973 51871 41976
rect 51813 41967 51871 41973
rect 53469 41973 53481 41976
rect 53515 42004 53527 42007
rect 54202 42004 54208 42016
rect 53515 41976 54208 42004
rect 53515 41973 53527 41976
rect 53469 41967 53527 41973
rect 54202 41964 54208 41976
rect 54260 41964 54266 42016
rect 54312 42004 54340 42103
rect 54404 42072 54432 42103
rect 54478 42100 54484 42152
rect 54536 42140 54542 42152
rect 54662 42140 54668 42152
rect 54536 42112 54668 42140
rect 54536 42100 54542 42112
rect 54662 42100 54668 42112
rect 54720 42100 54726 42152
rect 54846 42140 54852 42152
rect 54807 42112 54852 42140
rect 54846 42100 54852 42112
rect 54904 42100 54910 42152
rect 55674 42140 55680 42152
rect 55635 42112 55680 42140
rect 55674 42100 55680 42112
rect 55732 42100 55738 42152
rect 57146 42100 57152 42152
rect 57204 42140 57210 42152
rect 59630 42140 59636 42152
rect 57204 42112 59636 42140
rect 57204 42100 57210 42112
rect 59630 42100 59636 42112
rect 59688 42100 59694 42152
rect 59725 42143 59783 42149
rect 59725 42109 59737 42143
rect 59771 42109 59783 42143
rect 59998 42140 60004 42152
rect 59959 42112 60004 42140
rect 59725 42103 59783 42109
rect 54941 42075 54999 42081
rect 54941 42072 54953 42075
rect 54404 42044 54953 42072
rect 54941 42041 54953 42044
rect 54987 42072 54999 42075
rect 59740 42072 59768 42103
rect 59998 42100 60004 42112
rect 60056 42100 60062 42152
rect 60182 42140 60188 42152
rect 60095 42112 60188 42140
rect 60182 42100 60188 42112
rect 60240 42140 60246 42152
rect 60642 42140 60648 42152
rect 60240 42112 60648 42140
rect 60240 42100 60246 42112
rect 60642 42100 60648 42112
rect 60700 42100 60706 42152
rect 61010 42140 61016 42152
rect 60971 42112 61016 42140
rect 61010 42100 61016 42112
rect 61068 42100 61074 42152
rect 61194 42140 61200 42152
rect 61155 42112 61200 42140
rect 61194 42100 61200 42112
rect 61252 42100 61258 42152
rect 64506 42140 64512 42152
rect 64467 42112 64512 42140
rect 64506 42100 64512 42112
rect 64564 42100 64570 42152
rect 64601 42143 64659 42149
rect 64601 42109 64613 42143
rect 64647 42109 64659 42143
rect 64874 42140 64880 42152
rect 64835 42112 64880 42140
rect 64601 42103 64659 42109
rect 60277 42075 60335 42081
rect 60277 42072 60289 42075
rect 54987 42044 60289 42072
rect 54987 42041 54999 42044
rect 54941 42035 54999 42041
rect 60277 42041 60289 42044
rect 60323 42072 60335 42075
rect 64616 42072 64644 42103
rect 64874 42100 64880 42112
rect 64932 42100 64938 42152
rect 65058 42140 65064 42152
rect 65019 42112 65064 42140
rect 65058 42100 65064 42112
rect 65116 42100 65122 42152
rect 60323 42044 64644 42072
rect 65260 42072 65288 42180
rect 65352 42140 65380 42248
rect 66714 42236 66720 42248
rect 66772 42276 66778 42288
rect 67358 42276 67364 42288
rect 66772 42248 67364 42276
rect 66772 42236 66778 42248
rect 67358 42236 67364 42248
rect 67416 42236 67422 42288
rect 72694 42236 72700 42288
rect 72752 42276 72758 42288
rect 77849 42279 77907 42285
rect 77849 42276 77861 42279
rect 72752 42248 77861 42276
rect 72752 42236 72758 42248
rect 77849 42245 77861 42248
rect 77895 42276 77907 42279
rect 78582 42276 78588 42288
rect 77895 42248 78588 42276
rect 77895 42245 77907 42248
rect 77849 42239 77907 42245
rect 78582 42236 78588 42248
rect 78640 42236 78646 42288
rect 70578 42208 70584 42220
rect 70539 42180 70584 42208
rect 70578 42168 70584 42180
rect 70636 42168 70642 42220
rect 71133 42211 71191 42217
rect 71133 42177 71145 42211
rect 71179 42208 71191 42211
rect 71498 42208 71504 42220
rect 71179 42180 71504 42208
rect 71179 42177 71191 42180
rect 71133 42171 71191 42177
rect 71498 42168 71504 42180
rect 71556 42168 71562 42220
rect 73246 42208 73252 42220
rect 72712 42180 73252 42208
rect 66625 42143 66683 42149
rect 66625 42140 66637 42143
rect 65352 42112 66637 42140
rect 66625 42109 66637 42112
rect 66671 42140 66683 42143
rect 66901 42143 66959 42149
rect 66901 42140 66913 42143
rect 66671 42112 66913 42140
rect 66671 42109 66683 42112
rect 66625 42103 66683 42109
rect 66901 42109 66913 42112
rect 66947 42140 66959 42143
rect 67266 42140 67272 42152
rect 66947 42112 67272 42140
rect 66947 42109 66959 42112
rect 66901 42103 66959 42109
rect 67266 42100 67272 42112
rect 67324 42100 67330 42152
rect 69477 42143 69535 42149
rect 69477 42109 69489 42143
rect 69523 42109 69535 42143
rect 71222 42140 71228 42152
rect 69477 42103 69535 42109
rect 70412 42112 71228 42140
rect 69492 42072 69520 42103
rect 69842 42072 69848 42084
rect 65260 42044 69848 42072
rect 60323 42041 60335 42044
rect 60277 42035 60335 42041
rect 54662 42004 54668 42016
rect 54312 41976 54668 42004
rect 54662 41964 54668 41976
rect 54720 42004 54726 42016
rect 55769 42007 55827 42013
rect 55769 42004 55781 42007
rect 54720 41976 55781 42004
rect 54720 41964 54726 41976
rect 55769 41973 55781 41976
rect 55815 41973 55827 42007
rect 55769 41967 55827 41973
rect 55950 41964 55956 42016
rect 56008 42004 56014 42016
rect 60090 42004 60096 42016
rect 56008 41976 60096 42004
rect 56008 41964 56014 41976
rect 60090 41964 60096 41976
rect 60148 41964 60154 42016
rect 60458 41964 60464 42016
rect 60516 42004 60522 42016
rect 61289 42007 61347 42013
rect 61289 42004 61301 42007
rect 60516 41976 61301 42004
rect 60516 41964 60522 41976
rect 61289 41973 61301 41976
rect 61335 41973 61347 42007
rect 64616 42004 64644 42044
rect 69842 42032 69848 42044
rect 69900 42032 69906 42084
rect 65245 42007 65303 42013
rect 65245 42004 65257 42007
rect 64616 41976 65257 42004
rect 61289 41967 61347 41973
rect 65245 41973 65257 41976
rect 65291 42004 65303 42007
rect 66346 42004 66352 42016
rect 65291 41976 66352 42004
rect 65291 41973 65303 41976
rect 65245 41967 65303 41973
rect 66346 41964 66352 41976
rect 66404 41964 66410 42016
rect 69658 42004 69664 42016
rect 69619 41976 69664 42004
rect 69658 41964 69664 41976
rect 69716 42004 69722 42016
rect 70412 42013 70440 42112
rect 71222 42100 71228 42112
rect 71280 42149 71286 42152
rect 71280 42143 71329 42149
rect 71280 42109 71283 42143
rect 71317 42109 71329 42143
rect 71280 42103 71329 42109
rect 71409 42143 71467 42149
rect 71409 42109 71421 42143
rect 71455 42109 71467 42143
rect 72712 42140 72740 42180
rect 73246 42168 73252 42180
rect 73304 42168 73310 42220
rect 74350 42208 74356 42220
rect 74184 42180 74356 42208
rect 74184 42149 74212 42180
rect 74350 42168 74356 42180
rect 74408 42168 74414 42220
rect 74534 42168 74540 42220
rect 74592 42208 74598 42220
rect 74592 42180 74637 42208
rect 74592 42168 74598 42180
rect 75914 42168 75920 42220
rect 75972 42208 75978 42220
rect 80992 42208 81020 42316
rect 81069 42313 81081 42347
rect 81115 42344 81127 42347
rect 82078 42344 82084 42356
rect 81115 42316 82084 42344
rect 81115 42313 81127 42316
rect 81069 42307 81127 42313
rect 82078 42304 82084 42316
rect 82136 42344 82142 42356
rect 82354 42344 82360 42356
rect 82136 42316 82360 42344
rect 82136 42304 82142 42316
rect 82354 42304 82360 42316
rect 82412 42304 82418 42356
rect 85758 42208 85764 42220
rect 75972 42180 80928 42208
rect 80992 42180 85764 42208
rect 75972 42168 75978 42180
rect 71409 42103 71467 42109
rect 71700 42112 72740 42140
rect 72881 42143 72939 42149
rect 71280 42100 71286 42103
rect 71424 42072 71452 42103
rect 71700 42072 71728 42112
rect 72881 42109 72893 42143
rect 72927 42109 72939 42143
rect 72881 42103 72939 42109
rect 74169 42143 74227 42149
rect 74169 42109 74181 42143
rect 74215 42109 74227 42143
rect 74169 42103 74227 42109
rect 71424 42044 71728 42072
rect 72697 42075 72755 42081
rect 72697 42041 72709 42075
rect 72743 42041 72755 42075
rect 72896 42072 72924 42103
rect 74258 42100 74264 42152
rect 74316 42140 74322 42152
rect 74721 42143 74779 42149
rect 74721 42140 74733 42143
rect 74316 42112 74733 42140
rect 74316 42100 74322 42112
rect 74721 42109 74733 42112
rect 74767 42109 74779 42143
rect 74721 42103 74779 42109
rect 76561 42143 76619 42149
rect 76561 42109 76573 42143
rect 76607 42140 76619 42143
rect 77662 42140 77668 42152
rect 76607 42112 77668 42140
rect 76607 42109 76619 42112
rect 76561 42103 76619 42109
rect 77662 42100 77668 42112
rect 77720 42140 77726 42152
rect 78398 42140 78404 42152
rect 77720 42112 78404 42140
rect 77720 42100 77726 42112
rect 78398 42100 78404 42112
rect 78456 42100 78462 42152
rect 79870 42140 79876 42152
rect 79831 42112 79876 42140
rect 79870 42100 79876 42112
rect 79928 42100 79934 42152
rect 80900 42149 80928 42180
rect 85758 42168 85764 42180
rect 85816 42168 85822 42220
rect 80891 42143 80949 42149
rect 80891 42109 80903 42143
rect 80937 42109 80949 42143
rect 80891 42103 80949 42109
rect 82722 42100 82728 42152
rect 82780 42140 82786 42152
rect 82817 42143 82875 42149
rect 82817 42140 82829 42143
rect 82780 42112 82829 42140
rect 82780 42100 82786 42112
rect 82817 42109 82829 42112
rect 82863 42109 82875 42143
rect 83090 42140 83096 42152
rect 83051 42112 83096 42140
rect 82817 42103 82875 42109
rect 73246 42072 73252 42084
rect 72896 42044 73252 42072
rect 72697 42035 72755 42041
rect 70397 42007 70455 42013
rect 70397 42004 70409 42007
rect 69716 41976 70409 42004
rect 69716 41964 69722 41976
rect 70397 41973 70409 41976
rect 70443 41973 70455 42007
rect 72712 42004 72740 42035
rect 73246 42032 73252 42044
rect 73304 42072 73310 42084
rect 74276 42072 74304 42100
rect 73304 42044 74304 42072
rect 73304 42032 73310 42044
rect 74350 42004 74356 42016
rect 72712 41976 74356 42004
rect 70397 41967 70455 41973
rect 74350 41964 74356 41976
rect 74408 41964 74414 42016
rect 76742 42004 76748 42016
rect 76703 41976 76748 42004
rect 76742 41964 76748 41976
rect 76800 41964 76806 42016
rect 79962 42004 79968 42016
rect 79923 41976 79968 42004
rect 79962 41964 79968 41976
rect 80020 41964 80026 42016
rect 82725 42007 82783 42013
rect 82725 41973 82737 42007
rect 82771 42004 82783 42007
rect 82832 42004 82860 42103
rect 83090 42100 83096 42112
rect 83148 42100 83154 42152
rect 87138 42072 87144 42084
rect 83752 42044 87144 42072
rect 83752 42004 83780 42044
rect 87138 42032 87144 42044
rect 87196 42032 87202 42084
rect 82771 41976 83780 42004
rect 82771 41973 82783 41976
rect 82725 41967 82783 41973
rect 84102 41964 84108 42016
rect 84160 42004 84166 42016
rect 84197 42007 84255 42013
rect 84197 42004 84209 42007
rect 84160 41976 84209 42004
rect 84160 41964 84166 41976
rect 84197 41973 84209 41976
rect 84243 41973 84255 42007
rect 84197 41967 84255 41973
rect 1104 41914 105616 41936
rect 1104 41862 19606 41914
rect 19658 41862 19670 41914
rect 19722 41862 19734 41914
rect 19786 41862 19798 41914
rect 19850 41862 50326 41914
rect 50378 41862 50390 41914
rect 50442 41862 50454 41914
rect 50506 41862 50518 41914
rect 50570 41862 81046 41914
rect 81098 41862 81110 41914
rect 81162 41862 81174 41914
rect 81226 41862 81238 41914
rect 81290 41862 105616 41914
rect 1104 41840 105616 41862
rect 7834 41760 7840 41812
rect 7892 41800 7898 41812
rect 8021 41803 8079 41809
rect 8021 41800 8033 41803
rect 7892 41772 8033 41800
rect 7892 41760 7898 41772
rect 8021 41769 8033 41772
rect 8067 41769 8079 41803
rect 11514 41800 11520 41812
rect 11475 41772 11520 41800
rect 8021 41763 8079 41769
rect 11514 41760 11520 41772
rect 11572 41760 11578 41812
rect 11885 41803 11943 41809
rect 11885 41800 11897 41803
rect 11716 41772 11897 41800
rect 7024 41704 7604 41732
rect 7024 41673 7052 41704
rect 7009 41667 7067 41673
rect 7009 41633 7021 41667
rect 7055 41633 7067 41667
rect 7466 41664 7472 41676
rect 7427 41636 7472 41664
rect 7009 41627 7067 41633
rect 7466 41624 7472 41636
rect 7524 41624 7530 41676
rect 7576 41673 7604 41704
rect 9122 41692 9128 41744
rect 9180 41732 9186 41744
rect 11716 41732 11744 41772
rect 11885 41769 11897 41772
rect 11931 41800 11943 41803
rect 12526 41800 12532 41812
rect 11931 41772 12532 41800
rect 11931 41769 11943 41772
rect 11885 41763 11943 41769
rect 12526 41760 12532 41772
rect 12584 41800 12590 41812
rect 13722 41800 13728 41812
rect 12584 41772 13728 41800
rect 12584 41760 12590 41772
rect 13722 41760 13728 41772
rect 13780 41760 13786 41812
rect 16758 41800 16764 41812
rect 16719 41772 16764 41800
rect 16758 41760 16764 41772
rect 16816 41760 16822 41812
rect 16942 41800 16948 41812
rect 16903 41772 16948 41800
rect 16942 41760 16948 41772
rect 17000 41760 17006 41812
rect 26605 41803 26663 41809
rect 26605 41800 26617 41803
rect 17236 41772 26617 41800
rect 9180 41704 11744 41732
rect 9180 41692 9186 41704
rect 7561 41667 7619 41673
rect 7561 41633 7573 41667
rect 7607 41664 7619 41667
rect 7926 41664 7932 41676
rect 7607 41636 7932 41664
rect 7607 41633 7619 41636
rect 7561 41627 7619 41633
rect 7926 41624 7932 41636
rect 7984 41624 7990 41676
rect 8110 41624 8116 41676
rect 8168 41664 8174 41676
rect 10502 41664 10508 41676
rect 8168 41636 10508 41664
rect 8168 41624 8174 41636
rect 10502 41624 10508 41636
rect 10560 41624 10566 41676
rect 10980 41673 11008 41704
rect 11790 41692 11796 41744
rect 11848 41732 11854 41744
rect 17236 41732 17264 41772
rect 26605 41769 26617 41772
rect 26651 41769 26663 41803
rect 27890 41800 27896 41812
rect 27851 41772 27896 41800
rect 26605 41763 26663 41769
rect 27890 41760 27896 41772
rect 27948 41760 27954 41812
rect 28077 41803 28135 41809
rect 28077 41800 28089 41803
rect 28000 41772 28089 41800
rect 25774 41732 25780 41744
rect 11848 41704 17264 41732
rect 25332 41704 25544 41732
rect 11848 41692 11854 41704
rect 10965 41667 11023 41673
rect 10965 41633 10977 41667
rect 11011 41633 11023 41667
rect 10965 41627 11023 41633
rect 11054 41624 11060 41676
rect 11112 41664 11118 41676
rect 14182 41664 14188 41676
rect 11112 41636 11157 41664
rect 14143 41636 14188 41664
rect 11112 41624 11118 41636
rect 14182 41624 14188 41636
rect 14240 41624 14246 41676
rect 16022 41664 16028 41676
rect 15983 41636 16028 41664
rect 16022 41624 16028 41636
rect 16080 41624 16086 41676
rect 16393 41667 16451 41673
rect 16393 41633 16405 41667
rect 16439 41664 16451 41667
rect 16482 41664 16488 41676
rect 16439 41636 16488 41664
rect 16439 41633 16451 41636
rect 16393 41627 16451 41633
rect 16482 41624 16488 41636
rect 16540 41624 16546 41676
rect 16577 41667 16635 41673
rect 16577 41633 16589 41667
rect 16623 41664 16635 41667
rect 16758 41664 16764 41676
rect 16623 41636 16764 41664
rect 16623 41633 16635 41636
rect 16577 41627 16635 41633
rect 16758 41624 16764 41636
rect 16816 41624 16822 41676
rect 21174 41664 21180 41676
rect 17236 41636 21036 41664
rect 21135 41636 21180 41664
rect 6914 41556 6920 41608
rect 6972 41596 6978 41608
rect 10229 41599 10287 41605
rect 6972 41568 7017 41596
rect 6972 41556 6978 41568
rect 10229 41565 10241 41599
rect 10275 41596 10287 41599
rect 10318 41596 10324 41608
rect 10275 41568 10324 41596
rect 10275 41565 10287 41568
rect 10229 41559 10287 41565
rect 10318 41556 10324 41568
rect 10376 41556 10382 41608
rect 12526 41556 12532 41608
rect 12584 41596 12590 41608
rect 15381 41599 15439 41605
rect 15381 41596 15393 41599
rect 12584 41568 15393 41596
rect 12584 41556 12590 41568
rect 15381 41565 15393 41568
rect 15427 41565 15439 41599
rect 15381 41559 15439 41565
rect 16117 41599 16175 41605
rect 16117 41565 16129 41599
rect 16163 41596 16175 41599
rect 16942 41596 16948 41608
rect 16163 41568 16948 41596
rect 16163 41565 16175 41568
rect 16117 41559 16175 41565
rect 16942 41556 16948 41568
rect 17000 41556 17006 41608
rect 5074 41488 5080 41540
rect 5132 41528 5138 41540
rect 17236 41528 17264 41636
rect 20898 41596 20904 41608
rect 20859 41568 20904 41596
rect 20898 41556 20904 41568
rect 20956 41556 20962 41608
rect 21008 41596 21036 41636
rect 21174 41624 21180 41636
rect 21232 41624 21238 41676
rect 25038 41664 25044 41676
rect 24999 41636 25044 41664
rect 25038 41624 25044 41636
rect 25096 41624 25102 41676
rect 24397 41599 24455 41605
rect 24397 41596 24409 41599
rect 21008 41568 24409 41596
rect 24397 41565 24409 41568
rect 24443 41565 24455 41599
rect 24397 41559 24455 41565
rect 25133 41599 25191 41605
rect 25133 41565 25145 41599
rect 25179 41596 25191 41599
rect 25332 41596 25360 41704
rect 25409 41667 25467 41673
rect 25409 41633 25421 41667
rect 25455 41633 25467 41667
rect 25409 41627 25467 41633
rect 25179 41568 25360 41596
rect 25179 41565 25191 41568
rect 25133 41559 25191 41565
rect 5132 41500 17264 41528
rect 5132 41488 5138 41500
rect 18138 41488 18144 41540
rect 18196 41528 18202 41540
rect 18196 41500 20944 41528
rect 18196 41488 18202 41500
rect 2958 41420 2964 41472
rect 3016 41460 3022 41472
rect 6641 41463 6699 41469
rect 6641 41460 6653 41463
rect 3016 41432 6653 41460
rect 3016 41420 3022 41432
rect 6641 41429 6653 41432
rect 6687 41460 6699 41463
rect 6914 41460 6920 41472
rect 6687 41432 6920 41460
rect 6687 41429 6699 41432
rect 6641 41423 6699 41429
rect 6914 41420 6920 41432
rect 6972 41420 6978 41472
rect 11054 41420 11060 41472
rect 11112 41460 11118 41472
rect 13078 41460 13084 41472
rect 11112 41432 13084 41460
rect 11112 41420 11118 41432
rect 13078 41420 13084 41432
rect 13136 41420 13142 41472
rect 14274 41460 14280 41472
rect 14235 41432 14280 41460
rect 14274 41420 14280 41432
rect 14332 41420 14338 41472
rect 16482 41420 16488 41472
rect 16540 41460 16546 41472
rect 17129 41463 17187 41469
rect 17129 41460 17141 41463
rect 16540 41432 17141 41460
rect 16540 41420 16546 41432
rect 17129 41429 17141 41432
rect 17175 41460 17187 41463
rect 20714 41460 20720 41472
rect 17175 41432 20720 41460
rect 17175 41429 17187 41432
rect 17129 41423 17187 41429
rect 20714 41420 20720 41432
rect 20772 41420 20778 41472
rect 20916 41460 20944 41500
rect 21910 41488 21916 41540
rect 21968 41528 21974 41540
rect 24213 41531 24271 41537
rect 24213 41528 24225 41531
rect 21968 41500 24225 41528
rect 21968 41488 21974 41500
rect 24213 41497 24225 41500
rect 24259 41528 24271 41531
rect 25424 41528 25452 41627
rect 25516 41596 25544 41704
rect 25608 41704 25780 41732
rect 25608 41673 25636 41704
rect 25774 41692 25780 41704
rect 25832 41692 25838 41744
rect 26694 41732 26700 41744
rect 25884 41704 26700 41732
rect 25593 41667 25651 41673
rect 25593 41633 25605 41667
rect 25639 41633 25651 41667
rect 25593 41627 25651 41633
rect 25682 41624 25688 41676
rect 25740 41664 25746 41676
rect 25884 41664 25912 41704
rect 26694 41692 26700 41704
rect 26752 41692 26758 41744
rect 25740 41636 25912 41664
rect 25740 41624 25746 41636
rect 26142 41624 26148 41676
rect 26200 41664 26206 41676
rect 27157 41667 27215 41673
rect 27157 41664 27169 41667
rect 26200 41636 27169 41664
rect 26200 41624 26206 41636
rect 27157 41633 27169 41636
rect 27203 41633 27215 41667
rect 27157 41627 27215 41633
rect 27338 41624 27344 41676
rect 27396 41664 27402 41676
rect 27525 41667 27583 41673
rect 27525 41664 27537 41667
rect 27396 41636 27537 41664
rect 27396 41624 27402 41636
rect 27525 41633 27537 41636
rect 27571 41633 27583 41667
rect 27525 41627 27583 41633
rect 27709 41667 27767 41673
rect 27709 41633 27721 41667
rect 27755 41664 27767 41667
rect 27890 41664 27896 41676
rect 27755 41636 27896 41664
rect 27755 41633 27767 41636
rect 27709 41627 27767 41633
rect 27890 41624 27896 41636
rect 27948 41624 27954 41676
rect 25961 41599 26019 41605
rect 25961 41596 25973 41599
rect 25516 41568 25973 41596
rect 25961 41565 25973 41568
rect 26007 41596 26019 41599
rect 26326 41596 26332 41608
rect 26007 41568 26332 41596
rect 26007 41565 26019 41568
rect 25961 41559 26019 41565
rect 26326 41556 26332 41568
rect 26384 41556 26390 41608
rect 27249 41599 27307 41605
rect 27249 41565 27261 41599
rect 27295 41596 27307 41599
rect 28000 41596 28028 41772
rect 28077 41769 28089 41772
rect 28123 41800 28135 41803
rect 29270 41800 29276 41812
rect 28123 41772 29276 41800
rect 28123 41769 28135 41772
rect 28077 41763 28135 41769
rect 29270 41760 29276 41772
rect 29328 41760 29334 41812
rect 31570 41760 31576 41812
rect 31628 41800 31634 41812
rect 35526 41800 35532 41812
rect 31628 41772 35388 41800
rect 35487 41772 35532 41800
rect 31628 41760 31634 41772
rect 28166 41692 28172 41744
rect 28224 41732 28230 41744
rect 34054 41732 34060 41744
rect 28224 41704 34060 41732
rect 28224 41692 28230 41704
rect 34054 41692 34060 41704
rect 34112 41692 34118 41744
rect 34698 41692 34704 41744
rect 34756 41732 34762 41744
rect 35360 41732 35388 41772
rect 35526 41760 35532 41772
rect 35584 41760 35590 41812
rect 38010 41760 38016 41812
rect 38068 41800 38074 41812
rect 39390 41800 39396 41812
rect 38068 41772 39396 41800
rect 38068 41760 38074 41772
rect 39390 41760 39396 41772
rect 39448 41760 39454 41812
rect 39577 41803 39635 41809
rect 39577 41769 39589 41803
rect 39623 41800 39635 41803
rect 39666 41800 39672 41812
rect 39623 41772 39672 41800
rect 39623 41769 39635 41772
rect 39577 41763 39635 41769
rect 39666 41760 39672 41772
rect 39724 41760 39730 41812
rect 43162 41800 43168 41812
rect 39776 41772 43168 41800
rect 37461 41735 37519 41741
rect 37461 41732 37473 41735
rect 34756 41704 35296 41732
rect 35360 41704 37473 41732
rect 34756 41692 34762 41704
rect 30926 41664 30932 41676
rect 30887 41636 30932 41664
rect 30926 41624 30932 41636
rect 30984 41624 30990 41676
rect 32309 41667 32367 41673
rect 32309 41633 32321 41667
rect 32355 41664 32367 41667
rect 32398 41664 32404 41676
rect 32355 41636 32404 41664
rect 32355 41633 32367 41636
rect 32309 41627 32367 41633
rect 32398 41624 32404 41636
rect 32456 41624 32462 41676
rect 32674 41624 32680 41676
rect 32732 41664 32738 41676
rect 32769 41667 32827 41673
rect 32769 41664 32781 41667
rect 32732 41636 32781 41664
rect 32732 41624 32738 41636
rect 32769 41633 32781 41636
rect 32815 41633 32827 41667
rect 32769 41627 32827 41633
rect 32861 41667 32919 41673
rect 32861 41633 32873 41667
rect 32907 41664 32919 41667
rect 33870 41664 33876 41676
rect 32907 41636 33876 41664
rect 32907 41633 32919 41636
rect 32861 41627 32919 41633
rect 33870 41624 33876 41636
rect 33928 41624 33934 41676
rect 33962 41624 33968 41676
rect 34020 41664 34026 41676
rect 34149 41667 34207 41673
rect 34149 41664 34161 41667
rect 34020 41636 34161 41664
rect 34020 41624 34026 41636
rect 34149 41633 34161 41636
rect 34195 41633 34207 41667
rect 34330 41664 34336 41676
rect 34291 41636 34336 41664
rect 34149 41627 34207 41633
rect 27295 41568 28028 41596
rect 27295 41565 27307 41568
rect 27249 41559 27307 41565
rect 31754 41556 31760 41608
rect 31812 41596 31818 41608
rect 31849 41599 31907 41605
rect 31849 41596 31861 41599
rect 31812 41568 31861 41596
rect 31812 41556 31818 41568
rect 31849 41565 31861 41568
rect 31895 41596 31907 41599
rect 32125 41599 32183 41605
rect 32125 41596 32137 41599
rect 31895 41568 32137 41596
rect 31895 41565 31907 41568
rect 31849 41559 31907 41565
rect 32125 41565 32137 41568
rect 32171 41565 32183 41599
rect 34164 41596 34192 41627
rect 34330 41624 34336 41636
rect 34388 41624 34394 41676
rect 35268 41673 35296 41704
rect 37461 41701 37473 41704
rect 37507 41732 37519 41735
rect 37507 41704 38516 41732
rect 37507 41701 37519 41704
rect 37461 41695 37519 41701
rect 34517 41667 34575 41673
rect 34517 41633 34529 41667
rect 34563 41664 34575 41667
rect 35069 41667 35127 41673
rect 35069 41664 35081 41667
rect 34563 41636 35081 41664
rect 34563 41633 34575 41636
rect 34517 41627 34575 41633
rect 35069 41633 35081 41636
rect 35115 41633 35127 41667
rect 35069 41627 35127 41633
rect 35253 41667 35311 41673
rect 35253 41633 35265 41667
rect 35299 41664 35311 41667
rect 38010 41664 38016 41676
rect 35299 41636 35940 41664
rect 37971 41636 38016 41664
rect 35299 41633 35311 41636
rect 35253 41627 35311 41633
rect 34532 41596 34560 41627
rect 34164 41568 34560 41596
rect 32125 41559 32183 41565
rect 26234 41528 26240 41540
rect 24259 41500 26240 41528
rect 24259 41497 24271 41500
rect 24213 41491 24271 41497
rect 26234 41488 26240 41500
rect 26292 41528 26298 41540
rect 27154 41528 27160 41540
rect 26292 41500 27160 41528
rect 26292 41488 26298 41500
rect 27154 41488 27160 41500
rect 27212 41488 27218 41540
rect 30742 41528 30748 41540
rect 30703 41500 30748 41528
rect 30742 41488 30748 41500
rect 30800 41488 30806 41540
rect 32214 41488 32220 41540
rect 32272 41528 32278 41540
rect 32272 41500 32812 41528
rect 32272 41488 32278 41500
rect 21358 41460 21364 41472
rect 20916 41432 21364 41460
rect 21358 41420 21364 41432
rect 21416 41420 21422 41472
rect 22278 41460 22284 41472
rect 22239 41432 22284 41460
rect 22278 41420 22284 41432
rect 22336 41420 22342 41472
rect 22741 41463 22799 41469
rect 22741 41429 22753 41463
rect 22787 41460 22799 41463
rect 23106 41460 23112 41472
rect 22787 41432 23112 41460
rect 22787 41429 22799 41432
rect 22741 41423 22799 41429
rect 23106 41420 23112 41432
rect 23164 41460 23170 41472
rect 30760 41460 30788 41488
rect 23164 41432 30788 41460
rect 23164 41420 23170 41432
rect 31478 41420 31484 41472
rect 31536 41460 31542 41472
rect 31573 41463 31631 41469
rect 31573 41460 31585 41463
rect 31536 41432 31585 41460
rect 31536 41420 31542 41432
rect 31573 41429 31585 41432
rect 31619 41460 31631 41463
rect 32674 41460 32680 41472
rect 31619 41432 32680 41460
rect 31619 41429 31631 41432
rect 31573 41423 31631 41429
rect 32674 41420 32680 41432
rect 32732 41420 32738 41472
rect 32784 41460 32812 41500
rect 32858 41488 32864 41540
rect 32916 41528 32922 41540
rect 33229 41531 33287 41537
rect 33229 41528 33241 41531
rect 32916 41500 33241 41528
rect 32916 41488 32922 41500
rect 33229 41497 33241 41500
rect 33275 41497 33287 41531
rect 33686 41528 33692 41540
rect 33647 41500 33692 41528
rect 33229 41491 33287 41497
rect 33686 41488 33692 41500
rect 33744 41488 33750 41540
rect 35912 41537 35940 41636
rect 38010 41624 38016 41636
rect 38068 41624 38074 41676
rect 38488 41673 38516 41704
rect 38654 41692 38660 41744
rect 38712 41732 38718 41744
rect 39776 41732 39804 41772
rect 43162 41760 43168 41772
rect 43220 41800 43226 41812
rect 43717 41803 43775 41809
rect 43717 41800 43729 41803
rect 43220 41772 43729 41800
rect 43220 41760 43226 41772
rect 43717 41769 43729 41772
rect 43763 41769 43775 41803
rect 43717 41763 43775 41769
rect 38712 41704 39804 41732
rect 38712 41692 38718 41704
rect 40586 41692 40592 41744
rect 40644 41732 40650 41744
rect 43622 41732 43628 41744
rect 40644 41704 43628 41732
rect 40644 41692 40650 41704
rect 43622 41692 43628 41704
rect 43680 41692 43686 41744
rect 38473 41667 38531 41673
rect 38473 41633 38485 41667
rect 38519 41633 38531 41667
rect 38473 41627 38531 41633
rect 38562 41624 38568 41676
rect 38620 41664 38626 41676
rect 39666 41664 39672 41676
rect 38620 41636 39672 41664
rect 38620 41624 38626 41636
rect 39666 41624 39672 41636
rect 39724 41624 39730 41676
rect 42245 41667 42303 41673
rect 42245 41633 42257 41667
rect 42291 41664 42303 41667
rect 42610 41664 42616 41676
rect 42291 41636 42616 41664
rect 42291 41633 42303 41636
rect 42245 41627 42303 41633
rect 42610 41624 42616 41636
rect 42668 41664 42674 41676
rect 43530 41664 43536 41676
rect 42668 41636 43536 41664
rect 42668 41624 42674 41636
rect 43530 41624 43536 41636
rect 43588 41624 43594 41676
rect 43732 41664 43760 41763
rect 44818 41760 44824 41812
rect 44876 41800 44882 41812
rect 45465 41803 45523 41809
rect 45465 41800 45477 41803
rect 44876 41772 45477 41800
rect 44876 41760 44882 41772
rect 45465 41769 45477 41772
rect 45511 41800 45523 41803
rect 45922 41800 45928 41812
rect 45511 41772 45928 41800
rect 45511 41769 45523 41772
rect 45465 41763 45523 41769
rect 45922 41760 45928 41772
rect 45980 41800 45986 41812
rect 48222 41800 48228 41812
rect 45980 41772 48228 41800
rect 45980 41760 45986 41772
rect 48222 41760 48228 41772
rect 48280 41760 48286 41812
rect 48501 41803 48559 41809
rect 48501 41769 48513 41803
rect 48547 41800 48559 41803
rect 48590 41800 48596 41812
rect 48547 41772 48596 41800
rect 48547 41769 48559 41772
rect 48501 41763 48559 41769
rect 44100 41704 45600 41732
rect 44100 41673 44128 41704
rect 45572 41676 45600 41704
rect 45646 41692 45652 41744
rect 45704 41732 45710 41744
rect 46109 41735 46167 41741
rect 46109 41732 46121 41735
rect 45704 41704 46121 41732
rect 45704 41692 45710 41704
rect 46109 41701 46121 41704
rect 46155 41701 46167 41735
rect 46109 41695 46167 41701
rect 47762 41692 47768 41744
rect 47820 41732 47826 41744
rect 48516 41732 48544 41763
rect 48590 41760 48596 41772
rect 48648 41760 48654 41812
rect 49528 41772 50568 41800
rect 47820 41704 48544 41732
rect 47820 41692 47826 41704
rect 43901 41667 43959 41673
rect 43901 41664 43913 41667
rect 43732 41636 43913 41664
rect 43901 41633 43913 41636
rect 43947 41633 43959 41667
rect 43901 41627 43959 41633
rect 44085 41667 44143 41673
rect 44085 41633 44097 41667
rect 44131 41633 44143 41667
rect 44542 41664 44548 41676
rect 44503 41636 44548 41664
rect 44085 41627 44143 41633
rect 44542 41624 44548 41636
rect 44600 41624 44606 41676
rect 44637 41667 44695 41673
rect 44637 41633 44649 41667
rect 44683 41664 44695 41667
rect 44818 41664 44824 41676
rect 44683 41636 44824 41664
rect 44683 41633 44695 41636
rect 44637 41627 44695 41633
rect 44818 41624 44824 41636
rect 44876 41624 44882 41676
rect 45554 41664 45560 41676
rect 45467 41636 45560 41664
rect 45554 41624 45560 41636
rect 45612 41664 45618 41676
rect 48498 41664 48504 41676
rect 45612 41636 48504 41664
rect 45612 41624 45618 41636
rect 48498 41624 48504 41636
rect 48556 41624 48562 41676
rect 49145 41667 49203 41673
rect 49145 41633 49157 41667
rect 49191 41664 49203 41667
rect 49528 41664 49556 41772
rect 50540 41741 50568 41772
rect 51258 41760 51264 41812
rect 51316 41800 51322 41812
rect 69658 41800 69664 41812
rect 51316 41772 69664 41800
rect 51316 41760 51322 41772
rect 69658 41760 69664 41772
rect 69716 41760 69722 41812
rect 71682 41800 71688 41812
rect 69768 41772 71688 41800
rect 50525 41735 50583 41741
rect 50525 41701 50537 41735
rect 50571 41732 50583 41735
rect 64414 41732 64420 41744
rect 50571 41704 64420 41732
rect 50571 41701 50583 41704
rect 50525 41695 50583 41701
rect 64414 41692 64420 41704
rect 64472 41692 64478 41744
rect 64874 41732 64880 41744
rect 64524 41704 64880 41732
rect 49191 41636 49556 41664
rect 49191 41633 49203 41636
rect 49145 41627 49203 41633
rect 49602 41624 49608 41676
rect 49660 41664 49666 41676
rect 49697 41667 49755 41673
rect 49697 41664 49709 41667
rect 49660 41636 49709 41664
rect 49660 41624 49666 41636
rect 49697 41633 49709 41636
rect 49743 41633 49755 41667
rect 49878 41664 49884 41676
rect 49839 41636 49884 41664
rect 49697 41627 49755 41633
rect 49878 41624 49884 41636
rect 49936 41624 49942 41676
rect 53098 41664 53104 41676
rect 53059 41636 53104 41664
rect 53098 41624 53104 41636
rect 53156 41624 53162 41676
rect 53282 41664 53288 41676
rect 53243 41636 53288 41664
rect 53282 41624 53288 41636
rect 53340 41624 53346 41676
rect 55030 41664 55036 41676
rect 54991 41636 55036 41664
rect 55030 41624 55036 41636
rect 55088 41624 55094 41676
rect 55122 41624 55128 41676
rect 55180 41673 55186 41676
rect 55180 41667 55195 41673
rect 55183 41633 55195 41667
rect 55237 41667 55295 41673
rect 55237 41664 55249 41667
rect 55180 41627 55195 41633
rect 55232 41633 55249 41664
rect 55283 41633 55295 41667
rect 55232 41627 55295 41633
rect 55769 41667 55827 41673
rect 55769 41633 55781 41667
rect 55815 41664 55827 41667
rect 55950 41664 55956 41676
rect 55815 41636 55956 41664
rect 55815 41633 55827 41636
rect 55769 41627 55827 41633
rect 55180 41624 55186 41627
rect 37918 41596 37924 41608
rect 37879 41568 37924 41596
rect 37918 41556 37924 41568
rect 37976 41556 37982 41608
rect 39022 41556 39028 41608
rect 39080 41596 39086 41608
rect 42334 41596 42340 41608
rect 39080 41568 39125 41596
rect 42247 41568 42340 41596
rect 39080 41556 39086 41568
rect 42334 41556 42340 41568
rect 42392 41596 42398 41608
rect 43714 41596 43720 41608
rect 42392 41568 43720 41596
rect 42392 41556 42398 41568
rect 43714 41556 43720 41568
rect 43772 41556 43778 41608
rect 45189 41599 45247 41605
rect 45189 41565 45201 41599
rect 45235 41596 45247 41599
rect 45830 41596 45836 41608
rect 45235 41568 45836 41596
rect 45235 41565 45247 41568
rect 45189 41559 45247 41565
rect 45830 41556 45836 41568
rect 45888 41556 45894 41608
rect 46014 41556 46020 41608
rect 46072 41596 46078 41608
rect 46477 41599 46535 41605
rect 46477 41596 46489 41599
rect 46072 41568 46489 41596
rect 46072 41556 46078 41568
rect 46477 41565 46489 41568
rect 46523 41565 46535 41599
rect 46477 41559 46535 41565
rect 48685 41599 48743 41605
rect 48685 41565 48697 41599
rect 48731 41596 48743 41599
rect 48958 41596 48964 41608
rect 48731 41568 48964 41596
rect 48731 41565 48743 41568
rect 48685 41559 48743 41565
rect 48958 41556 48964 41568
rect 49016 41556 49022 41608
rect 53653 41599 53711 41605
rect 53653 41565 53665 41599
rect 53699 41596 53711 41599
rect 55232 41596 55260 41627
rect 55950 41624 55956 41636
rect 56008 41624 56014 41676
rect 57330 41624 57336 41676
rect 57388 41664 57394 41676
rect 58713 41667 58771 41673
rect 58713 41664 58725 41667
rect 57388 41636 58725 41664
rect 57388 41624 57394 41636
rect 58713 41633 58725 41636
rect 58759 41664 58771 41667
rect 58897 41667 58955 41673
rect 58897 41664 58909 41667
rect 58759 41636 58909 41664
rect 58759 41633 58771 41636
rect 58713 41627 58771 41633
rect 58897 41633 58909 41636
rect 58943 41633 58955 41667
rect 58897 41627 58955 41633
rect 58989 41667 59047 41673
rect 58989 41633 59001 41667
rect 59035 41664 59047 41667
rect 59170 41664 59176 41676
rect 59035 41636 59176 41664
rect 59035 41633 59047 41636
rect 58989 41627 59047 41633
rect 59170 41624 59176 41636
rect 59228 41624 59234 41676
rect 59906 41624 59912 41676
rect 59964 41664 59970 41676
rect 60185 41667 60243 41673
rect 60185 41664 60197 41667
rect 59964 41636 60197 41664
rect 59964 41624 59970 41636
rect 60185 41633 60197 41636
rect 60231 41664 60243 41667
rect 60461 41667 60519 41673
rect 60461 41664 60473 41667
rect 60231 41636 60473 41664
rect 60231 41633 60243 41636
rect 60185 41627 60243 41633
rect 60461 41633 60473 41636
rect 60507 41633 60519 41667
rect 60461 41627 60519 41633
rect 63221 41667 63279 41673
rect 63221 41633 63233 41667
rect 63267 41664 63279 41667
rect 63313 41667 63371 41673
rect 63313 41664 63325 41667
rect 63267 41636 63325 41664
rect 63267 41633 63279 41636
rect 63221 41627 63279 41633
rect 63313 41633 63325 41636
rect 63359 41633 63371 41667
rect 64322 41664 64328 41676
rect 64283 41636 64328 41664
rect 63313 41627 63371 41633
rect 64322 41624 64328 41636
rect 64380 41624 64386 41676
rect 64524 41673 64552 41704
rect 64874 41692 64880 41704
rect 64932 41692 64938 41744
rect 66346 41692 66352 41744
rect 66404 41732 66410 41744
rect 69768 41732 69796 41772
rect 71682 41760 71688 41772
rect 71740 41760 71746 41812
rect 74350 41760 74356 41812
rect 74408 41800 74414 41812
rect 74721 41803 74779 41809
rect 74721 41800 74733 41803
rect 74408 41772 74733 41800
rect 74408 41760 74414 41772
rect 74721 41769 74733 41772
rect 74767 41769 74779 41803
rect 74721 41763 74779 41769
rect 66404 41704 69796 41732
rect 66404 41692 66410 41704
rect 69842 41692 69848 41744
rect 69900 41732 69906 41744
rect 71869 41735 71927 41741
rect 71869 41732 71881 41735
rect 69900 41704 71881 41732
rect 69900 41692 69906 41704
rect 71869 41701 71881 41704
rect 71915 41732 71927 41735
rect 72697 41735 72755 41741
rect 72697 41732 72709 41735
rect 71915 41704 72709 41732
rect 71915 41701 71927 41704
rect 71869 41695 71927 41701
rect 72697 41701 72709 41704
rect 72743 41732 72755 41735
rect 72881 41735 72939 41741
rect 72881 41732 72893 41735
rect 72743 41704 72893 41732
rect 72743 41701 72755 41704
rect 72697 41695 72755 41701
rect 72881 41701 72893 41704
rect 72927 41701 72939 41735
rect 73246 41732 73252 41744
rect 72881 41695 72939 41701
rect 73080 41704 73252 41732
rect 64509 41667 64567 41673
rect 64509 41633 64521 41667
rect 64555 41633 64567 41667
rect 64509 41627 64567 41633
rect 53699 41568 55260 41596
rect 53699 41565 53711 41568
rect 53653 41559 53711 41565
rect 55858 41556 55864 41608
rect 55916 41596 55922 41608
rect 60001 41599 60059 41605
rect 60001 41596 60013 41599
rect 55916 41568 60013 41596
rect 55916 41556 55922 41568
rect 60001 41565 60013 41568
rect 60047 41565 60059 41599
rect 60001 41559 60059 41565
rect 60090 41556 60096 41608
rect 60148 41596 60154 41608
rect 60277 41599 60335 41605
rect 60277 41596 60289 41599
rect 60148 41568 60289 41596
rect 60148 41556 60154 41568
rect 60277 41565 60289 41568
rect 60323 41565 60335 41599
rect 60277 41559 60335 41565
rect 63405 41599 63463 41605
rect 63405 41565 63417 41599
rect 63451 41596 63463 41599
rect 64524 41596 64552 41627
rect 65058 41624 65064 41676
rect 65116 41664 65122 41676
rect 65797 41667 65855 41673
rect 65797 41664 65809 41667
rect 65116 41636 65809 41664
rect 65116 41624 65122 41636
rect 65797 41633 65809 41636
rect 65843 41664 65855 41667
rect 67542 41664 67548 41676
rect 65843 41636 67548 41664
rect 65843 41633 65855 41636
rect 65797 41627 65855 41633
rect 67542 41624 67548 41636
rect 67600 41624 67606 41676
rect 71774 41664 71780 41676
rect 71735 41636 71780 41664
rect 71774 41624 71780 41636
rect 71832 41624 71838 41676
rect 73080 41673 73108 41704
rect 73246 41692 73252 41704
rect 73304 41692 73310 41744
rect 74166 41692 74172 41744
rect 74224 41732 74230 41744
rect 81713 41735 81771 41741
rect 74224 41704 81664 41732
rect 74224 41692 74230 41704
rect 73028 41667 73108 41673
rect 73028 41633 73040 41667
rect 73074 41636 73108 41667
rect 73074 41633 73086 41636
rect 73028 41627 73086 41633
rect 73154 41624 73160 41676
rect 73212 41664 73218 41676
rect 74445 41667 74503 41673
rect 74445 41664 74457 41667
rect 73212 41636 74457 41664
rect 73212 41624 73218 41636
rect 74445 41633 74457 41636
rect 74491 41633 74503 41667
rect 74445 41627 74503 41633
rect 74629 41667 74687 41673
rect 74629 41633 74641 41667
rect 74675 41633 74687 41667
rect 74629 41627 74687 41633
rect 77941 41667 77999 41673
rect 77941 41633 77953 41667
rect 77987 41664 77999 41667
rect 78401 41667 78459 41673
rect 78401 41664 78413 41667
rect 77987 41636 78413 41664
rect 77987 41633 77999 41636
rect 77941 41627 77999 41633
rect 78401 41633 78413 41636
rect 78447 41664 78459 41667
rect 78674 41664 78680 41676
rect 78447 41636 78680 41664
rect 78447 41633 78459 41636
rect 78401 41627 78459 41633
rect 63451 41568 64552 41596
rect 63451 41565 63463 41568
rect 63405 41559 63463 41565
rect 65426 41556 65432 41608
rect 65484 41596 65490 41608
rect 65521 41599 65579 41605
rect 65521 41596 65533 41599
rect 65484 41568 65533 41596
rect 65484 41556 65490 41568
rect 65521 41565 65533 41568
rect 65567 41596 65579 41599
rect 66165 41599 66223 41605
rect 66165 41596 66177 41599
rect 65567 41568 66177 41596
rect 65567 41565 65579 41568
rect 65521 41559 65579 41565
rect 66165 41565 66177 41568
rect 66211 41565 66223 41599
rect 66346 41596 66352 41608
rect 66307 41568 66352 41596
rect 66165 41559 66223 41565
rect 66346 41556 66352 41568
rect 66404 41556 66410 41608
rect 73246 41596 73252 41608
rect 73207 41568 73252 41596
rect 73246 41556 73252 41568
rect 73304 41556 73310 41608
rect 73338 41556 73344 41608
rect 73396 41596 73402 41608
rect 74644 41596 74672 41627
rect 78674 41624 78680 41636
rect 78732 41624 78738 41676
rect 81158 41664 81164 41676
rect 81119 41636 81164 41664
rect 81158 41624 81164 41636
rect 81216 41624 81222 41676
rect 81345 41667 81403 41673
rect 81345 41633 81357 41667
rect 81391 41633 81403 41667
rect 81636 41664 81664 41704
rect 81713 41701 81725 41735
rect 81759 41732 81771 41735
rect 81986 41732 81992 41744
rect 81759 41704 81992 41732
rect 81759 41701 81771 41704
rect 81713 41695 81771 41701
rect 81986 41692 81992 41704
rect 82044 41732 82050 41744
rect 82817 41735 82875 41741
rect 82817 41732 82829 41735
rect 82044 41704 82829 41732
rect 82044 41692 82050 41704
rect 82817 41701 82829 41704
rect 82863 41701 82875 41735
rect 82817 41695 82875 41701
rect 82354 41664 82360 41676
rect 81636 41636 82360 41664
rect 81345 41627 81403 41633
rect 73396 41568 74672 41596
rect 73396 41556 73402 41568
rect 80882 41556 80888 41608
rect 80940 41596 80946 41608
rect 81360 41596 81388 41627
rect 82354 41624 82360 41636
rect 82412 41664 82418 41676
rect 82633 41667 82691 41673
rect 82633 41664 82645 41667
rect 82412 41636 82645 41664
rect 82412 41624 82418 41636
rect 82633 41633 82645 41636
rect 82679 41633 82691 41667
rect 82633 41627 82691 41633
rect 82906 41624 82912 41676
rect 82964 41664 82970 41676
rect 82964 41636 83009 41664
rect 82964 41624 82970 41636
rect 83642 41624 83648 41676
rect 83700 41664 83706 41676
rect 84102 41664 84108 41676
rect 83700 41636 84108 41664
rect 83700 41624 83706 41636
rect 84102 41624 84108 41636
rect 84160 41664 84166 41676
rect 84197 41667 84255 41673
rect 84197 41664 84209 41667
rect 84160 41636 84209 41664
rect 84160 41624 84166 41636
rect 84197 41633 84209 41636
rect 84243 41633 84255 41667
rect 84197 41627 84255 41633
rect 84289 41599 84347 41605
rect 84289 41596 84301 41599
rect 80940 41568 84301 41596
rect 80940 41556 80946 41568
rect 84289 41565 84301 41568
rect 84335 41565 84347 41599
rect 84289 41559 84347 41565
rect 35897 41531 35955 41537
rect 35897 41497 35909 41531
rect 35943 41528 35955 41531
rect 35943 41500 39068 41528
rect 35943 41497 35955 41500
rect 35897 41491 35955 41497
rect 33502 41460 33508 41472
rect 32784 41432 33508 41460
rect 33502 41420 33508 41432
rect 33560 41420 33566 41472
rect 33870 41460 33876 41472
rect 33831 41432 33876 41460
rect 33870 41420 33876 41432
rect 33928 41420 33934 41472
rect 34054 41420 34060 41472
rect 34112 41460 34118 41472
rect 38930 41460 38936 41472
rect 34112 41432 38936 41460
rect 34112 41420 34118 41432
rect 38930 41420 38936 41432
rect 38988 41420 38994 41472
rect 39040 41460 39068 41500
rect 39114 41488 39120 41540
rect 39172 41528 39178 41540
rect 78125 41531 78183 41537
rect 78125 41528 78137 41531
rect 39172 41500 78137 41528
rect 39172 41488 39178 41500
rect 78125 41497 78137 41500
rect 78171 41528 78183 41531
rect 78858 41528 78864 41540
rect 78171 41500 78864 41528
rect 78171 41497 78183 41500
rect 78125 41491 78183 41497
rect 78858 41488 78864 41500
rect 78916 41488 78922 41540
rect 42334 41460 42340 41472
rect 39040 41432 42340 41460
rect 42334 41420 42340 41432
rect 42392 41420 42398 41472
rect 43438 41420 43444 41472
rect 43496 41460 43502 41472
rect 43533 41463 43591 41469
rect 43533 41460 43545 41463
rect 43496 41432 43545 41460
rect 43496 41420 43502 41432
rect 43533 41429 43545 41432
rect 43579 41460 43591 41463
rect 44542 41460 44548 41472
rect 43579 41432 44548 41460
rect 43579 41429 43591 41432
rect 43533 41423 43591 41429
rect 44542 41420 44548 41432
rect 44600 41420 44606 41472
rect 45922 41420 45928 41472
rect 45980 41460 45986 41472
rect 46247 41463 46305 41469
rect 46247 41460 46259 41463
rect 45980 41432 46259 41460
rect 45980 41420 45986 41432
rect 46247 41429 46259 41432
rect 46293 41429 46305 41463
rect 46382 41460 46388 41472
rect 46343 41432 46388 41460
rect 46247 41423 46305 41429
rect 46382 41420 46388 41432
rect 46440 41420 46446 41472
rect 46566 41460 46572 41472
rect 46527 41432 46572 41460
rect 46566 41420 46572 41432
rect 46624 41420 46630 41472
rect 50154 41460 50160 41472
rect 50115 41432 50160 41460
rect 50154 41420 50160 41432
rect 50212 41420 50218 41472
rect 55030 41420 55036 41472
rect 55088 41460 55094 41472
rect 55401 41463 55459 41469
rect 55401 41460 55413 41463
rect 55088 41432 55413 41460
rect 55088 41420 55094 41432
rect 55401 41429 55413 41432
rect 55447 41429 55459 41463
rect 55401 41423 55459 41429
rect 60001 41463 60059 41469
rect 60001 41429 60013 41463
rect 60047 41460 60059 41463
rect 63221 41463 63279 41469
rect 63221 41460 63233 41463
rect 60047 41432 63233 41460
rect 60047 41429 60059 41432
rect 60001 41423 60059 41429
rect 63221 41429 63233 41432
rect 63267 41460 63279 41463
rect 63589 41463 63647 41469
rect 63589 41460 63601 41463
rect 63267 41432 63601 41460
rect 63267 41429 63279 41432
rect 63221 41423 63279 41429
rect 63589 41429 63601 41432
rect 63635 41460 63647 41463
rect 64230 41460 64236 41472
rect 63635 41432 64236 41460
rect 63635 41429 63647 41432
rect 63589 41423 63647 41429
rect 64230 41420 64236 41432
rect 64288 41420 64294 41472
rect 64601 41463 64659 41469
rect 64601 41429 64613 41463
rect 64647 41460 64659 41463
rect 65935 41463 65993 41469
rect 65935 41460 65947 41463
rect 64647 41432 65947 41460
rect 64647 41429 64659 41432
rect 64601 41423 64659 41429
rect 65935 41429 65947 41432
rect 65981 41429 65993 41463
rect 65935 41423 65993 41429
rect 66073 41463 66131 41469
rect 66073 41429 66085 41463
rect 66119 41460 66131 41463
rect 66714 41460 66720 41472
rect 66119 41432 66720 41460
rect 66119 41429 66131 41432
rect 66073 41423 66131 41429
rect 66714 41420 66720 41432
rect 66772 41420 66778 41472
rect 72602 41420 72608 41472
rect 72660 41460 72666 41472
rect 73157 41463 73215 41469
rect 73157 41460 73169 41463
rect 72660 41432 73169 41460
rect 72660 41420 72666 41432
rect 73157 41429 73169 41432
rect 73203 41460 73215 41463
rect 73338 41460 73344 41472
rect 73203 41432 73344 41460
rect 73203 41429 73215 41432
rect 73157 41423 73215 41429
rect 73338 41420 73344 41432
rect 73396 41420 73402 41472
rect 73522 41460 73528 41472
rect 73483 41432 73528 41460
rect 73522 41420 73528 41432
rect 73580 41420 73586 41472
rect 83090 41460 83096 41472
rect 83051 41432 83096 41460
rect 83090 41420 83096 41432
rect 83148 41420 83154 41472
rect 1104 41370 105616 41392
rect 1104 41318 4246 41370
rect 4298 41318 4310 41370
rect 4362 41318 4374 41370
rect 4426 41318 4438 41370
rect 4490 41318 34966 41370
rect 35018 41318 35030 41370
rect 35082 41318 35094 41370
rect 35146 41318 35158 41370
rect 35210 41318 65686 41370
rect 65738 41318 65750 41370
rect 65802 41318 65814 41370
rect 65866 41318 65878 41370
rect 65930 41318 96406 41370
rect 96458 41318 96470 41370
rect 96522 41318 96534 41370
rect 96586 41318 96598 41370
rect 96650 41318 105616 41370
rect 1104 41296 105616 41318
rect 4617 41259 4675 41265
rect 4617 41256 4629 41259
rect 2792 41228 4629 41256
rect 2792 41129 2820 41228
rect 4617 41225 4629 41228
rect 4663 41256 4675 41259
rect 4798 41256 4804 41268
rect 4663 41228 4804 41256
rect 4663 41225 4675 41228
rect 4617 41219 4675 41225
rect 4798 41216 4804 41228
rect 4856 41216 4862 41268
rect 8386 41216 8392 41268
rect 8444 41256 8450 41268
rect 8757 41259 8815 41265
rect 8757 41256 8769 41259
rect 8444 41228 8769 41256
rect 8444 41216 8450 41228
rect 8757 41225 8769 41228
rect 8803 41256 8815 41259
rect 8938 41256 8944 41268
rect 8803 41228 8944 41256
rect 8803 41225 8815 41228
rect 8757 41219 8815 41225
rect 8938 41216 8944 41228
rect 8996 41256 9002 41268
rect 45005 41259 45063 41265
rect 8996 41228 44956 41256
rect 8996 41216 9002 41228
rect 14093 41191 14151 41197
rect 14093 41157 14105 41191
rect 14139 41188 14151 41191
rect 14182 41188 14188 41200
rect 14139 41160 14188 41188
rect 14139 41157 14151 41160
rect 14093 41151 14151 41157
rect 14182 41148 14188 41160
rect 14240 41148 14246 41200
rect 25317 41191 25375 41197
rect 25317 41157 25329 41191
rect 25363 41188 25375 41191
rect 26050 41188 26056 41200
rect 25363 41160 26056 41188
rect 25363 41157 25375 41160
rect 25317 41151 25375 41157
rect 26050 41148 26056 41160
rect 26108 41148 26114 41200
rect 26145 41191 26203 41197
rect 26145 41157 26157 41191
rect 26191 41188 26203 41191
rect 26234 41188 26240 41200
rect 26191 41160 26240 41188
rect 26191 41157 26203 41160
rect 26145 41151 26203 41157
rect 26234 41148 26240 41160
rect 26292 41148 26298 41200
rect 27798 41188 27804 41200
rect 26896 41160 27804 41188
rect 2777 41123 2835 41129
rect 2777 41089 2789 41123
rect 2823 41089 2835 41123
rect 2777 41083 2835 41089
rect 9674 41080 9680 41132
rect 9732 41120 9738 41132
rect 26694 41120 26700 41132
rect 9732 41092 26700 41120
rect 9732 41080 9738 41092
rect 26694 41080 26700 41092
rect 26752 41080 26758 41132
rect 26789 41123 26847 41129
rect 26789 41089 26801 41123
rect 26835 41120 26847 41123
rect 26896 41120 26924 41160
rect 27798 41148 27804 41160
rect 27856 41148 27862 41200
rect 30926 41148 30932 41200
rect 30984 41188 30990 41200
rect 33965 41191 34023 41197
rect 33965 41188 33977 41191
rect 30984 41160 33977 41188
rect 30984 41148 30990 41160
rect 33965 41157 33977 41160
rect 34011 41157 34023 41191
rect 33965 41151 34023 41157
rect 34422 41148 34428 41200
rect 34480 41188 34486 41200
rect 44174 41188 44180 41200
rect 34480 41160 38884 41188
rect 34480 41148 34486 41160
rect 26835 41092 26924 41120
rect 26835 41089 26847 41092
rect 26789 41083 26847 41089
rect 26970 41080 26976 41132
rect 27028 41120 27034 41132
rect 32122 41120 32128 41132
rect 27028 41092 32128 41120
rect 27028 41080 27034 41092
rect 32122 41080 32128 41092
rect 32180 41080 32186 41132
rect 33410 41080 33416 41132
rect 33468 41120 33474 41132
rect 38289 41123 38347 41129
rect 33468 41092 37136 41120
rect 33468 41080 33474 41092
rect 3053 41055 3111 41061
rect 3053 41021 3065 41055
rect 3099 41052 3111 41055
rect 3786 41052 3792 41064
rect 3099 41024 3792 41052
rect 3099 41021 3111 41024
rect 3053 41015 3111 41021
rect 3786 41012 3792 41024
rect 3844 41012 3850 41064
rect 8386 41052 8392 41064
rect 8347 41024 8392 41052
rect 8386 41012 8392 41024
rect 8444 41012 8450 41064
rect 12713 41055 12771 41061
rect 12713 41021 12725 41055
rect 12759 41021 12771 41055
rect 12986 41052 12992 41064
rect 12947 41024 12992 41052
rect 12713 41015 12771 41021
rect 4433 40987 4491 40993
rect 4433 40953 4445 40987
rect 4479 40984 4491 40987
rect 5626 40984 5632 40996
rect 4479 40956 5632 40984
rect 4479 40953 4491 40956
rect 4433 40947 4491 40953
rect 5626 40944 5632 40956
rect 5684 40944 5690 40996
rect 7466 40876 7472 40928
rect 7524 40916 7530 40928
rect 8481 40919 8539 40925
rect 8481 40916 8493 40919
rect 7524 40888 8493 40916
rect 7524 40876 7530 40888
rect 8481 40885 8493 40888
rect 8527 40885 8539 40919
rect 12728 40916 12756 41015
rect 12986 41012 12992 41024
rect 13044 41012 13050 41064
rect 13722 41012 13728 41064
rect 13780 41052 13786 41064
rect 15197 41055 15255 41061
rect 15197 41052 15209 41055
rect 13780 41024 15209 41052
rect 13780 41012 13786 41024
rect 15197 41021 15209 41024
rect 15243 41021 15255 41055
rect 15197 41015 15255 41021
rect 19334 41012 19340 41064
rect 19392 41052 19398 41064
rect 19705 41055 19763 41061
rect 19705 41052 19717 41055
rect 19392 41024 19717 41052
rect 19392 41012 19398 41024
rect 19705 41021 19717 41024
rect 19751 41021 19763 41055
rect 19978 41052 19984 41064
rect 19939 41024 19984 41052
rect 19705 41015 19763 41021
rect 19978 41012 19984 41024
rect 20036 41012 20042 41064
rect 22278 41052 22284 41064
rect 21284 41024 21772 41052
rect 22239 41024 22284 41052
rect 14274 40944 14280 40996
rect 14332 40984 14338 40996
rect 14332 40956 15516 40984
rect 14332 40944 14338 40956
rect 13630 40916 13636 40928
rect 12728 40888 13636 40916
rect 8481 40879 8539 40885
rect 13630 40876 13636 40888
rect 13688 40916 13694 40928
rect 14461 40919 14519 40925
rect 14461 40916 14473 40919
rect 13688 40888 14473 40916
rect 13688 40876 13694 40888
rect 14461 40885 14473 40888
rect 14507 40885 14519 40919
rect 15378 40916 15384 40928
rect 15339 40888 15384 40916
rect 14461 40879 14519 40885
rect 15378 40876 15384 40888
rect 15436 40876 15442 40928
rect 15488 40916 15516 40956
rect 21284 40916 21312 41024
rect 21361 40987 21419 40993
rect 21361 40953 21373 40987
rect 21407 40984 21419 40987
rect 21634 40984 21640 40996
rect 21407 40956 21640 40984
rect 21407 40953 21419 40956
rect 21361 40947 21419 40953
rect 21634 40944 21640 40956
rect 21692 40944 21698 40996
rect 21744 40984 21772 41024
rect 22278 41012 22284 41024
rect 22336 41012 22342 41064
rect 24854 41012 24860 41064
rect 24912 41052 24918 41064
rect 25133 41055 25191 41061
rect 25133 41052 25145 41055
rect 24912 41024 25145 41052
rect 24912 41012 24918 41024
rect 25133 41021 25145 41024
rect 25179 41021 25191 41055
rect 25133 41015 25191 41021
rect 26142 41012 26148 41064
rect 26200 41052 26206 41064
rect 26881 41055 26939 41061
rect 26881 41052 26893 41055
rect 26200 41024 26893 41052
rect 26200 41012 26206 41024
rect 26881 41021 26893 41024
rect 26927 41021 26939 41055
rect 27246 41052 27252 41064
rect 27207 41024 27252 41052
rect 26881 41015 26939 41021
rect 27246 41012 27252 41024
rect 27304 41012 27310 41064
rect 27433 41055 27491 41061
rect 27433 41021 27445 41055
rect 27479 41052 27491 41055
rect 27614 41052 27620 41064
rect 27479 41024 27620 41052
rect 27479 41021 27491 41024
rect 27433 41015 27491 41021
rect 27614 41012 27620 41024
rect 27672 41012 27678 41064
rect 27706 41012 27712 41064
rect 27764 41052 27770 41064
rect 31478 41052 31484 41064
rect 27764 41024 31484 41052
rect 27764 41012 27770 41024
rect 31478 41012 31484 41024
rect 31536 41012 31542 41064
rect 31570 41012 31576 41064
rect 31628 41052 31634 41064
rect 31757 41055 31815 41061
rect 31757 41052 31769 41055
rect 31628 41024 31769 41052
rect 31628 41012 31634 41024
rect 31757 41021 31769 41024
rect 31803 41021 31815 41055
rect 31938 41052 31944 41064
rect 31899 41024 31944 41052
rect 31757 41015 31815 41021
rect 31938 41012 31944 41024
rect 31996 41012 32002 41064
rect 32398 41052 32404 41064
rect 32359 41024 32404 41052
rect 32398 41012 32404 41024
rect 32456 41012 32462 41064
rect 32490 41012 32496 41064
rect 32548 41052 32554 41064
rect 32548 41024 32593 41052
rect 32548 41012 32554 41024
rect 32674 41012 32680 41064
rect 32732 41052 32738 41064
rect 34149 41055 34207 41061
rect 32732 41024 33548 41052
rect 32732 41012 32738 41024
rect 33410 40984 33416 40996
rect 21744 40956 33416 40984
rect 33410 40944 33416 40956
rect 33468 40944 33474 40996
rect 33520 40984 33548 41024
rect 34149 41021 34161 41055
rect 34195 41052 34207 41055
rect 34790 41052 34796 41064
rect 34195 41024 34796 41052
rect 34195 41021 34207 41024
rect 34149 41015 34207 41021
rect 34790 41012 34796 41024
rect 34848 41012 34854 41064
rect 37001 41055 37059 41061
rect 37001 41021 37013 41055
rect 37047 41021 37059 41055
rect 37001 41015 37059 41021
rect 36817 40987 36875 40993
rect 36817 40984 36829 40987
rect 33520 40956 33640 40984
rect 21450 40916 21456 40928
rect 15488 40888 21312 40916
rect 21411 40888 21456 40916
rect 21450 40876 21456 40888
rect 21508 40876 21514 40928
rect 22370 40916 22376 40928
rect 22331 40888 22376 40916
rect 22370 40876 22376 40888
rect 22428 40876 22434 40928
rect 24854 40876 24860 40928
rect 24912 40916 24918 40928
rect 24949 40919 25007 40925
rect 24949 40916 24961 40919
rect 24912 40888 24961 40916
rect 24912 40876 24918 40888
rect 24949 40885 24961 40888
rect 24995 40885 25007 40919
rect 24949 40879 25007 40885
rect 25038 40876 25044 40928
rect 25096 40916 25102 40928
rect 26142 40916 26148 40928
rect 25096 40888 26148 40916
rect 25096 40876 25102 40888
rect 26142 40876 26148 40888
rect 26200 40876 26206 40928
rect 26326 40916 26332 40928
rect 26287 40888 26332 40916
rect 26326 40876 26332 40888
rect 26384 40876 26390 40928
rect 26418 40876 26424 40928
rect 26476 40916 26482 40928
rect 27430 40916 27436 40928
rect 26476 40888 27436 40916
rect 26476 40876 26482 40888
rect 27430 40876 27436 40888
rect 27488 40876 27494 40928
rect 27614 40916 27620 40928
rect 27575 40888 27620 40916
rect 27614 40876 27620 40888
rect 27672 40876 27678 40928
rect 27798 40916 27804 40928
rect 27759 40888 27804 40916
rect 27798 40876 27804 40888
rect 27856 40876 27862 40928
rect 30282 40876 30288 40928
rect 30340 40916 30346 40928
rect 31389 40919 31447 40925
rect 31389 40916 31401 40919
rect 30340 40888 31401 40916
rect 30340 40876 30346 40888
rect 31389 40885 31401 40888
rect 31435 40916 31447 40919
rect 31754 40916 31760 40928
rect 31435 40888 31760 40916
rect 31435 40885 31447 40888
rect 31389 40879 31447 40885
rect 31754 40876 31760 40888
rect 31812 40916 31818 40928
rect 32398 40916 32404 40928
rect 31812 40888 32404 40916
rect 31812 40876 31818 40888
rect 32398 40876 32404 40888
rect 32456 40876 32462 40928
rect 32953 40919 33011 40925
rect 32953 40885 32965 40919
rect 32999 40916 33011 40919
rect 33134 40916 33140 40928
rect 32999 40888 33140 40916
rect 32999 40885 33011 40888
rect 32953 40879 33011 40885
rect 33134 40876 33140 40888
rect 33192 40876 33198 40928
rect 33318 40916 33324 40928
rect 33279 40888 33324 40916
rect 33318 40876 33324 40888
rect 33376 40876 33382 40928
rect 33502 40916 33508 40928
rect 33463 40888 33508 40916
rect 33502 40876 33508 40888
rect 33560 40876 33566 40928
rect 33612 40916 33640 40956
rect 34256 40956 36829 40984
rect 34256 40916 34284 40956
rect 36817 40953 36829 40956
rect 36863 40984 36875 40987
rect 37016 40984 37044 41015
rect 36863 40956 37044 40984
rect 37108 40984 37136 41092
rect 38289 41089 38301 41123
rect 38335 41120 38347 41123
rect 38746 41120 38752 41132
rect 38335 41092 38752 41120
rect 38335 41089 38347 41092
rect 38289 41083 38347 41089
rect 38746 41080 38752 41092
rect 38804 41080 38810 41132
rect 38856 41120 38884 41160
rect 42812 41160 44180 41188
rect 42812 41120 42840 41160
rect 44174 41148 44180 41160
rect 44232 41148 44238 41200
rect 44928 41188 44956 41228
rect 45005 41225 45017 41259
rect 45051 41256 45063 41259
rect 45922 41256 45928 41268
rect 45051 41228 45928 41256
rect 45051 41225 45063 41228
rect 45005 41219 45063 41225
rect 45922 41216 45928 41228
rect 45980 41216 45986 41268
rect 48958 41256 48964 41268
rect 47964 41228 48964 41256
rect 47964 41197 47992 41228
rect 48958 41216 48964 41228
rect 49016 41216 49022 41268
rect 49050 41216 49056 41268
rect 49108 41256 49114 41268
rect 49881 41259 49939 41265
rect 49881 41256 49893 41259
rect 49108 41228 49893 41256
rect 49108 41216 49114 41228
rect 49881 41225 49893 41228
rect 49927 41256 49939 41259
rect 51258 41256 51264 41268
rect 49927 41228 51264 41256
rect 49927 41225 49939 41228
rect 49881 41219 49939 41225
rect 51258 41216 51264 41228
rect 51316 41216 51322 41268
rect 52457 41259 52515 41265
rect 52457 41225 52469 41259
rect 52503 41256 52515 41259
rect 52733 41259 52791 41265
rect 52733 41256 52745 41259
rect 52503 41228 52745 41256
rect 52503 41225 52515 41228
rect 52457 41219 52515 41225
rect 52733 41225 52745 41228
rect 52779 41256 52791 41259
rect 53282 41256 53288 41268
rect 52779 41228 53288 41256
rect 52779 41225 52791 41228
rect 52733 41219 52791 41225
rect 53282 41216 53288 41228
rect 53340 41216 53346 41268
rect 55858 41256 55864 41268
rect 53392 41228 55864 41256
rect 47949 41191 48007 41197
rect 47949 41188 47961 41191
rect 44928 41160 47961 41188
rect 47949 41157 47961 41160
rect 47995 41157 48007 41191
rect 50062 41188 50068 41200
rect 49975 41160 50068 41188
rect 47949 41151 48007 41157
rect 50062 41148 50068 41160
rect 50120 41188 50126 41200
rect 53392 41188 53420 41228
rect 55858 41216 55864 41228
rect 55916 41216 55922 41268
rect 63770 41256 63776 41268
rect 63683 41228 63776 41256
rect 63770 41216 63776 41228
rect 63828 41256 63834 41268
rect 64506 41256 64512 41268
rect 63828 41228 64512 41256
rect 63828 41216 63834 41228
rect 64506 41216 64512 41228
rect 64564 41216 64570 41268
rect 67542 41216 67548 41268
rect 67600 41256 67606 41268
rect 71222 41256 71228 41268
rect 67600 41228 71228 41256
rect 67600 41216 67606 41228
rect 71222 41216 71228 41228
rect 71280 41216 71286 41268
rect 76742 41256 76748 41268
rect 73080 41228 76748 41256
rect 73080 41200 73108 41228
rect 76742 41216 76748 41228
rect 76800 41216 76806 41268
rect 78674 41216 78680 41268
rect 78732 41256 78738 41268
rect 79962 41256 79968 41268
rect 78732 41228 79968 41256
rect 78732 41216 78738 41228
rect 79962 41216 79968 41228
rect 80020 41256 80026 41268
rect 80241 41259 80299 41265
rect 80241 41256 80253 41259
rect 80020 41228 80253 41256
rect 80020 41216 80026 41228
rect 80241 41225 80253 41228
rect 80287 41225 80299 41259
rect 80882 41256 80888 41268
rect 80843 41228 80888 41256
rect 80241 41219 80299 41225
rect 50120 41160 53420 41188
rect 62776 41160 66392 41188
rect 50120 41148 50126 41160
rect 43898 41120 43904 41132
rect 38856 41092 42840 41120
rect 43859 41092 43904 41120
rect 43898 41080 43904 41092
rect 43956 41080 43962 41132
rect 45094 41080 45100 41132
rect 45152 41120 45158 41132
rect 45281 41123 45339 41129
rect 45281 41120 45293 41123
rect 45152 41092 45293 41120
rect 45152 41080 45158 41092
rect 45281 41089 45293 41092
rect 45327 41089 45339 41123
rect 48409 41123 48467 41129
rect 48409 41120 48421 41123
rect 45281 41083 45339 41089
rect 48148 41092 48421 41120
rect 37185 41055 37243 41061
rect 37185 41021 37197 41055
rect 37231 41052 37243 41055
rect 37366 41052 37372 41064
rect 37231 41024 37372 41052
rect 37231 41021 37243 41024
rect 37185 41015 37243 41021
rect 37366 41012 37372 41024
rect 37424 41012 37430 41064
rect 37642 41052 37648 41064
rect 37603 41024 37648 41052
rect 37642 41012 37648 41024
rect 37700 41012 37706 41064
rect 37737 41055 37795 41061
rect 37737 41021 37749 41055
rect 37783 41052 37795 41055
rect 38102 41052 38108 41064
rect 37783 41024 38108 41052
rect 37783 41021 37795 41024
rect 37737 41015 37795 41021
rect 38102 41012 38108 41024
rect 38160 41052 38166 41064
rect 38473 41055 38531 41061
rect 38473 41052 38485 41055
rect 38160 41024 38485 41052
rect 38160 41012 38166 41024
rect 38473 41021 38485 41024
rect 38519 41021 38531 41055
rect 43990 41052 43996 41064
rect 43951 41024 43996 41052
rect 38473 41015 38531 41021
rect 43990 41012 43996 41024
rect 44048 41012 44054 41064
rect 44082 41012 44088 41064
rect 44140 41052 44146 41064
rect 44453 41055 44511 41061
rect 44453 41052 44465 41055
rect 44140 41024 44465 41052
rect 44140 41012 44146 41024
rect 44453 41021 44465 41024
rect 44499 41021 44511 41055
rect 44453 41015 44511 41021
rect 44545 41055 44603 41061
rect 44545 41021 44557 41055
rect 44591 41052 44603 41055
rect 45112 41052 45140 41080
rect 44591 41024 45140 41052
rect 44591 41021 44603 41024
rect 44545 41015 44603 41021
rect 45186 41012 45192 41064
rect 45244 41052 45250 41064
rect 45462 41052 45468 41064
rect 45244 41024 45468 41052
rect 45244 41012 45250 41024
rect 45462 41012 45468 41024
rect 45520 41012 45526 41064
rect 48148 40993 48176 41092
rect 48409 41089 48421 41092
rect 48455 41120 48467 41123
rect 48682 41120 48688 41132
rect 48455 41092 48688 41120
rect 48455 41089 48467 41092
rect 48409 41083 48467 41089
rect 48682 41080 48688 41092
rect 48740 41080 48746 41132
rect 49510 41080 49516 41132
rect 49568 41120 49574 41132
rect 62776 41120 62804 41160
rect 65153 41123 65211 41129
rect 65153 41120 65165 41123
rect 49568 41092 62804 41120
rect 63696 41092 65165 41120
rect 49568 41080 49574 41092
rect 48498 41052 48504 41064
rect 48459 41024 48504 41052
rect 48498 41012 48504 41024
rect 48556 41012 48562 41064
rect 48958 41052 48964 41064
rect 48919 41024 48964 41052
rect 48958 41012 48964 41024
rect 49016 41012 49022 41064
rect 49050 41012 49056 41064
rect 49108 41052 49114 41064
rect 52638 41052 52644 41064
rect 49108 41024 49153 41052
rect 52599 41024 52644 41052
rect 49108 41012 49114 41024
rect 52638 41012 52644 41024
rect 52696 41012 52702 41064
rect 54757 41055 54815 41061
rect 54757 41052 54769 41055
rect 54588 41024 54769 41052
rect 48133 40987 48191 40993
rect 48133 40984 48145 40987
rect 37108 40956 48145 40984
rect 36863 40953 36875 40956
rect 36817 40947 36875 40953
rect 48133 40953 48145 40956
rect 48179 40953 48191 40987
rect 48133 40947 48191 40953
rect 48314 40944 48320 40996
rect 48372 40984 48378 40996
rect 49068 40984 49096 41012
rect 52457 40987 52515 40993
rect 52457 40984 52469 40987
rect 48372 40956 49096 40984
rect 49160 40956 52469 40984
rect 48372 40944 48378 40956
rect 33612 40888 34284 40916
rect 38749 40919 38807 40925
rect 38749 40885 38761 40919
rect 38795 40916 38807 40919
rect 38930 40916 38936 40928
rect 38795 40888 38936 40916
rect 38795 40885 38807 40888
rect 38749 40879 38807 40885
rect 38930 40876 38936 40888
rect 38988 40916 38994 40928
rect 45186 40916 45192 40928
rect 38988 40888 45192 40916
rect 38988 40876 38994 40888
rect 45186 40876 45192 40888
rect 45244 40876 45250 40928
rect 45370 40876 45376 40928
rect 45428 40916 45434 40928
rect 49160 40916 49188 40956
rect 52457 40953 52469 40956
rect 52503 40953 52515 40987
rect 52457 40947 52515 40953
rect 54588 40928 54616 41024
rect 54757 41021 54769 41024
rect 54803 41021 54815 41055
rect 55030 41052 55036 41064
rect 54991 41024 55036 41052
rect 54757 41015 54815 41021
rect 55030 41012 55036 41024
rect 55088 41012 55094 41064
rect 63696 41061 63724 41092
rect 65153 41089 65165 41092
rect 65199 41120 65211 41123
rect 65199 41092 65288 41120
rect 65199 41089 65211 41092
rect 65153 41083 65211 41089
rect 63681 41055 63739 41061
rect 63681 41021 63693 41055
rect 63727 41021 63739 41055
rect 64874 41052 64880 41064
rect 64835 41024 64880 41052
rect 63681 41015 63739 41021
rect 64874 41012 64880 41024
rect 64932 41012 64938 41064
rect 64693 40987 64751 40993
rect 64693 40953 64705 40987
rect 64739 40984 64751 40987
rect 65058 40984 65064 40996
rect 64739 40956 65064 40984
rect 64739 40953 64751 40956
rect 64693 40947 64751 40953
rect 65058 40944 65064 40956
rect 65116 40944 65122 40996
rect 65260 40984 65288 41092
rect 66257 41055 66315 41061
rect 66257 41052 66269 41055
rect 66180 41024 66269 41052
rect 66073 40987 66131 40993
rect 66073 40984 66085 40987
rect 65260 40956 66085 40984
rect 66073 40953 66085 40956
rect 66119 40953 66131 40987
rect 66073 40947 66131 40953
rect 45428 40888 49188 40916
rect 45428 40876 45434 40888
rect 49326 40876 49332 40928
rect 49384 40916 49390 40928
rect 49513 40919 49571 40925
rect 49513 40916 49525 40919
rect 49384 40888 49525 40916
rect 49384 40876 49390 40888
rect 49513 40885 49525 40888
rect 49559 40885 49571 40919
rect 54570 40916 54576 40928
rect 54531 40888 54576 40916
rect 49513 40879 49571 40885
rect 54570 40876 54576 40888
rect 54628 40876 54634 40928
rect 54846 40876 54852 40928
rect 54904 40916 54910 40928
rect 56137 40919 56195 40925
rect 56137 40916 56149 40919
rect 54904 40888 56149 40916
rect 54904 40876 54910 40888
rect 56137 40885 56149 40888
rect 56183 40885 56195 40919
rect 56137 40879 56195 40885
rect 63494 40876 63500 40928
rect 63552 40916 63558 40928
rect 64322 40916 64328 40928
rect 63552 40888 64328 40916
rect 63552 40876 63558 40888
rect 64322 40876 64328 40888
rect 64380 40916 64386 40928
rect 66180 40916 66208 41024
rect 66257 41021 66269 41024
rect 66303 41021 66315 41055
rect 66257 41015 66315 41021
rect 66364 40984 66392 41160
rect 71682 41148 71688 41200
rect 71740 41188 71746 41200
rect 73062 41188 73068 41200
rect 71740 41160 73068 41188
rect 71740 41148 71746 41160
rect 73062 41148 73068 41160
rect 73120 41148 73126 41200
rect 73522 41148 73528 41200
rect 73580 41188 73586 41200
rect 74445 41191 74503 41197
rect 74445 41188 74457 41191
rect 73580 41160 74457 41188
rect 73580 41148 73586 41160
rect 74445 41157 74457 41160
rect 74491 41157 74503 41191
rect 74445 41151 74503 41157
rect 74644 41092 79272 41120
rect 71685 41055 71743 41061
rect 71685 41021 71697 41055
rect 71731 41021 71743 41055
rect 71685 41015 71743 41021
rect 71777 41055 71835 41061
rect 71777 41021 71789 41055
rect 71823 41052 71835 41055
rect 72881 41055 72939 41061
rect 72881 41052 72893 41055
rect 71823 41024 72893 41052
rect 71823 41021 71835 41024
rect 71777 41015 71835 41021
rect 72881 41021 72893 41024
rect 72927 41052 72939 41055
rect 73246 41052 73252 41064
rect 72927 41024 73252 41052
rect 72927 41021 72939 41024
rect 72881 41015 72939 41021
rect 71700 40984 71728 41015
rect 73246 41012 73252 41024
rect 73304 41052 73310 41064
rect 73430 41052 73436 41064
rect 73304 41024 73436 41052
rect 73304 41012 73310 41024
rect 73430 41012 73436 41024
rect 73488 41012 73494 41064
rect 74644 41061 74672 41092
rect 74353 41055 74411 41061
rect 74353 41021 74365 41055
rect 74399 41021 74411 41055
rect 74353 41015 74411 41021
rect 74629 41055 74687 41061
rect 74629 41021 74641 41055
rect 74675 41052 74687 41055
rect 74718 41052 74724 41064
rect 74675 41024 74724 41052
rect 74675 41021 74687 41024
rect 74629 41015 74687 41021
rect 72697 40987 72755 40993
rect 66364 40956 72096 40984
rect 64380 40888 66208 40916
rect 64380 40876 64386 40888
rect 66254 40876 66260 40928
rect 66312 40916 66318 40928
rect 66349 40919 66407 40925
rect 66349 40916 66361 40919
rect 66312 40888 66361 40916
rect 66312 40876 66318 40888
rect 66349 40885 66361 40888
rect 66395 40916 66407 40919
rect 67358 40916 67364 40928
rect 66395 40888 67364 40916
rect 66395 40885 66407 40888
rect 66349 40879 66407 40885
rect 67358 40876 67364 40888
rect 67416 40876 67422 40928
rect 72068 40925 72096 40956
rect 72697 40953 72709 40987
rect 72743 40984 72755 40987
rect 73522 40984 73528 40996
rect 72743 40956 73528 40984
rect 72743 40953 72755 40956
rect 72697 40947 72755 40953
rect 73522 40944 73528 40956
rect 73580 40944 73586 40996
rect 74368 40984 74396 41015
rect 74718 41012 74724 41024
rect 74776 41012 74782 41064
rect 78398 41052 78404 41064
rect 78359 41024 78404 41052
rect 78398 41012 78404 41024
rect 78456 41012 78462 41064
rect 79244 41052 79272 41092
rect 80256 41052 80284 41219
rect 80882 41216 80888 41228
rect 80940 41216 80946 41268
rect 87138 41256 87144 41268
rect 87099 41228 87144 41256
rect 87138 41216 87144 41228
rect 87196 41216 87202 41268
rect 80774 41191 80832 41197
rect 80774 41157 80786 41191
rect 80820 41188 80832 41191
rect 81434 41188 81440 41200
rect 80820 41160 81440 41188
rect 80820 41157 80832 41160
rect 80774 41151 80832 41157
rect 81434 41148 81440 41160
rect 81492 41148 81498 41200
rect 80977 41123 81035 41129
rect 80977 41089 80989 41123
rect 81023 41089 81035 41123
rect 87156 41120 87184 41216
rect 87325 41123 87383 41129
rect 87325 41120 87337 41123
rect 87156 41092 87337 41120
rect 80977 41083 81035 41089
rect 87325 41089 87337 41092
rect 87371 41120 87383 41123
rect 88978 41120 88984 41132
rect 87371 41092 88984 41120
rect 87371 41089 87383 41092
rect 87325 41083 87383 41089
rect 80609 41055 80667 41061
rect 80609 41052 80621 41055
rect 79244 41024 80100 41052
rect 80256 41024 80621 41052
rect 74902 40984 74908 40996
rect 74368 40956 74908 40984
rect 74902 40944 74908 40956
rect 74960 40984 74966 40996
rect 75181 40987 75239 40993
rect 75181 40984 75193 40987
rect 74960 40956 75193 40984
rect 74960 40944 74966 40956
rect 75181 40953 75193 40956
rect 75227 40953 75239 40987
rect 80072 40984 80100 41024
rect 80609 41021 80621 41024
rect 80655 41021 80667 41055
rect 80609 41015 80667 41021
rect 80790 41012 80796 41064
rect 80848 41052 80854 41064
rect 80992 41052 81020 41083
rect 88978 41080 88984 41092
rect 89036 41080 89042 41132
rect 80848 41024 81020 41052
rect 82633 41055 82691 41061
rect 80848 41012 80854 41024
rect 82633 41021 82645 41055
rect 82679 41052 82691 41055
rect 83642 41052 83648 41064
rect 82679 41024 83648 41052
rect 82679 41021 82691 41024
rect 82633 41015 82691 41021
rect 83642 41012 83648 41024
rect 83700 41012 83706 41064
rect 87598 41052 87604 41064
rect 87559 41024 87604 41052
rect 87598 41012 87604 41024
rect 87656 41012 87662 41064
rect 81345 40987 81403 40993
rect 81345 40984 81357 40987
rect 80072 40956 81357 40984
rect 75181 40947 75239 40953
rect 81345 40953 81357 40956
rect 81391 40953 81403 40987
rect 81345 40947 81403 40953
rect 72053 40919 72111 40925
rect 72053 40885 72065 40919
rect 72099 40916 72111 40919
rect 72142 40916 72148 40928
rect 72099 40888 72148 40916
rect 72099 40885 72111 40888
rect 72053 40879 72111 40885
rect 72142 40876 72148 40888
rect 72200 40876 72206 40928
rect 72970 40916 72976 40928
rect 72931 40888 72976 40916
rect 72970 40876 72976 40888
rect 73028 40916 73034 40928
rect 73154 40916 73160 40928
rect 73028 40888 73160 40916
rect 73028 40876 73034 40888
rect 73154 40876 73160 40888
rect 73212 40876 73218 40928
rect 74810 40916 74816 40928
rect 74771 40888 74816 40916
rect 74810 40876 74816 40888
rect 74868 40876 74874 40928
rect 78585 40919 78643 40925
rect 78585 40885 78597 40919
rect 78631 40916 78643 40919
rect 79410 40916 79416 40928
rect 78631 40888 79416 40916
rect 78631 40885 78643 40888
rect 78585 40879 78643 40885
rect 79410 40876 79416 40888
rect 79468 40876 79474 40928
rect 80517 40919 80575 40925
rect 80517 40885 80529 40919
rect 80563 40916 80575 40919
rect 80790 40916 80796 40928
rect 80563 40888 80796 40916
rect 80563 40885 80575 40888
rect 80517 40879 80575 40885
rect 80790 40876 80796 40888
rect 80848 40876 80854 40928
rect 82722 40876 82728 40928
rect 82780 40916 82786 40928
rect 82817 40919 82875 40925
rect 82817 40916 82829 40919
rect 82780 40888 82829 40916
rect 82780 40876 82786 40888
rect 82817 40885 82829 40888
rect 82863 40885 82875 40919
rect 82817 40879 82875 40885
rect 88518 40876 88524 40928
rect 88576 40916 88582 40928
rect 88705 40919 88763 40925
rect 88705 40916 88717 40919
rect 88576 40888 88717 40916
rect 88576 40876 88582 40888
rect 88705 40885 88717 40888
rect 88751 40885 88763 40919
rect 88705 40879 88763 40885
rect 1104 40826 105616 40848
rect 1104 40774 19606 40826
rect 19658 40774 19670 40826
rect 19722 40774 19734 40826
rect 19786 40774 19798 40826
rect 19850 40774 50326 40826
rect 50378 40774 50390 40826
rect 50442 40774 50454 40826
rect 50506 40774 50518 40826
rect 50570 40774 81046 40826
rect 81098 40774 81110 40826
rect 81162 40774 81174 40826
rect 81226 40774 81238 40826
rect 81290 40774 105616 40826
rect 1104 40752 105616 40774
rect 2866 40672 2872 40724
rect 2924 40712 2930 40724
rect 4157 40715 4215 40721
rect 4157 40712 4169 40715
rect 2924 40684 4169 40712
rect 2924 40672 2930 40684
rect 4157 40681 4169 40684
rect 4203 40681 4215 40715
rect 4157 40675 4215 40681
rect 4982 40672 4988 40724
rect 5040 40712 5046 40724
rect 12529 40715 12587 40721
rect 5040 40684 8340 40712
rect 5040 40672 5046 40684
rect 8202 40644 8208 40656
rect 7760 40616 8208 40644
rect 4341 40579 4399 40585
rect 4341 40545 4353 40579
rect 4387 40545 4399 40579
rect 4341 40539 4399 40545
rect 4617 40579 4675 40585
rect 4617 40545 4629 40579
rect 4663 40576 4675 40579
rect 5626 40576 5632 40588
rect 4663 40548 5028 40576
rect 5587 40548 5632 40576
rect 4663 40545 4675 40548
rect 4617 40539 4675 40545
rect 4356 40508 4384 40539
rect 4798 40508 4804 40520
rect 4356 40480 4804 40508
rect 4798 40468 4804 40480
rect 4856 40468 4862 40520
rect 5000 40449 5028 40548
rect 5626 40536 5632 40548
rect 5684 40536 5690 40588
rect 7466 40536 7472 40588
rect 7524 40576 7530 40588
rect 7760 40585 7788 40616
rect 8202 40604 8208 40616
rect 8260 40604 8266 40656
rect 8312 40644 8340 40684
rect 12529 40681 12541 40715
rect 12575 40712 12587 40715
rect 12986 40712 12992 40724
rect 12575 40684 12992 40712
rect 12575 40681 12587 40684
rect 12529 40675 12587 40681
rect 12986 40672 12992 40684
rect 13044 40672 13050 40724
rect 16669 40715 16727 40721
rect 16669 40681 16681 40715
rect 16715 40712 16727 40715
rect 17862 40712 17868 40724
rect 16715 40684 17868 40712
rect 16715 40681 16727 40684
rect 16669 40675 16727 40681
rect 17862 40672 17868 40684
rect 17920 40672 17926 40724
rect 20714 40712 20720 40724
rect 20627 40684 20720 40712
rect 20714 40672 20720 40684
rect 20772 40712 20778 40724
rect 21910 40712 21916 40724
rect 20772 40684 21916 40712
rect 20772 40672 20778 40684
rect 21910 40672 21916 40684
rect 21968 40672 21974 40724
rect 24946 40672 24952 40724
rect 25004 40712 25010 40724
rect 26418 40712 26424 40724
rect 25004 40684 26424 40712
rect 25004 40672 25010 40684
rect 26418 40672 26424 40684
rect 26476 40672 26482 40724
rect 27798 40672 27804 40724
rect 27856 40712 27862 40724
rect 31754 40712 31760 40724
rect 27856 40684 31760 40712
rect 27856 40672 27862 40684
rect 31754 40672 31760 40684
rect 31812 40672 31818 40724
rect 31941 40715 31999 40721
rect 31941 40681 31953 40715
rect 31987 40712 31999 40715
rect 31987 40684 37596 40712
rect 31987 40681 31999 40684
rect 31941 40675 31999 40681
rect 26326 40644 26332 40656
rect 8312 40616 26332 40644
rect 26326 40604 26332 40616
rect 26384 40604 26390 40656
rect 27522 40604 27528 40656
rect 27580 40644 27586 40656
rect 27580 40616 31064 40644
rect 27580 40604 27586 40616
rect 7561 40579 7619 40585
rect 7561 40576 7573 40579
rect 7524 40548 7573 40576
rect 7524 40536 7530 40548
rect 7561 40545 7573 40548
rect 7607 40545 7619 40579
rect 7561 40539 7619 40545
rect 7745 40579 7803 40585
rect 7745 40545 7757 40579
rect 7791 40545 7803 40579
rect 7745 40539 7803 40545
rect 8113 40579 8171 40585
rect 8113 40545 8125 40579
rect 8159 40576 8171 40579
rect 8478 40576 8484 40588
rect 8159 40548 8484 40576
rect 8159 40545 8171 40548
rect 8113 40539 8171 40545
rect 8478 40536 8484 40548
rect 8536 40536 8542 40588
rect 11517 40579 11575 40585
rect 11517 40545 11529 40579
rect 11563 40576 11575 40579
rect 11974 40576 11980 40588
rect 11563 40548 11980 40576
rect 11563 40545 11575 40548
rect 11517 40539 11575 40545
rect 11974 40536 11980 40548
rect 12032 40536 12038 40588
rect 12066 40536 12072 40588
rect 12124 40576 12130 40588
rect 12253 40579 12311 40585
rect 12124 40548 12169 40576
rect 12124 40536 12130 40548
rect 12253 40545 12265 40579
rect 12299 40576 12311 40579
rect 12710 40576 12716 40588
rect 12299 40548 12716 40576
rect 12299 40545 12311 40548
rect 12253 40539 12311 40545
rect 12710 40536 12716 40548
rect 12768 40576 12774 40588
rect 13538 40576 13544 40588
rect 12768 40548 12940 40576
rect 13451 40548 13544 40576
rect 12768 40536 12774 40548
rect 8018 40508 8024 40520
rect 7979 40480 8024 40508
rect 8018 40468 8024 40480
rect 8076 40468 8082 40520
rect 10962 40468 10968 40520
rect 11020 40508 11026 40520
rect 12912 40517 12940 40548
rect 13538 40536 13544 40548
rect 13596 40576 13602 40588
rect 13722 40576 13728 40588
rect 13596 40548 13728 40576
rect 13596 40536 13602 40548
rect 13722 40536 13728 40548
rect 13780 40536 13786 40588
rect 16393 40579 16451 40585
rect 16393 40545 16405 40579
rect 16439 40576 16451 40579
rect 16485 40579 16543 40585
rect 16485 40576 16497 40579
rect 16439 40548 16497 40576
rect 16439 40545 16451 40548
rect 16393 40539 16451 40545
rect 16485 40545 16497 40548
rect 16531 40576 16543 40579
rect 16574 40576 16580 40588
rect 16531 40548 16580 40576
rect 16531 40545 16543 40548
rect 16485 40539 16543 40545
rect 16574 40536 16580 40548
rect 16632 40536 16638 40588
rect 21545 40579 21603 40585
rect 21545 40576 21557 40579
rect 20824 40548 21557 40576
rect 11333 40511 11391 40517
rect 11333 40508 11345 40511
rect 11020 40480 11345 40508
rect 11020 40468 11026 40480
rect 11333 40477 11345 40480
rect 11379 40477 11391 40511
rect 11333 40471 11391 40477
rect 12897 40511 12955 40517
rect 12897 40477 12909 40511
rect 12943 40508 12955 40511
rect 14274 40508 14280 40520
rect 12943 40480 14280 40508
rect 12943 40477 12955 40480
rect 12897 40471 12955 40477
rect 14274 40468 14280 40480
rect 14332 40468 14338 40520
rect 16022 40468 16028 40520
rect 16080 40508 16086 40520
rect 20824 40508 20852 40548
rect 21545 40545 21557 40548
rect 21591 40545 21603 40579
rect 21910 40576 21916 40588
rect 21871 40548 21916 40576
rect 21545 40539 21603 40545
rect 16080 40480 20852 40508
rect 20901 40511 20959 40517
rect 16080 40468 16086 40480
rect 20901 40477 20913 40511
rect 20947 40477 20959 40511
rect 20901 40471 20959 40477
rect 4985 40443 5043 40449
rect 4985 40409 4997 40443
rect 5031 40440 5043 40443
rect 20916 40440 20944 40471
rect 5031 40412 20944 40440
rect 21560 40440 21588 40539
rect 21910 40536 21916 40548
rect 21968 40536 21974 40588
rect 22094 40576 22100 40588
rect 22055 40548 22100 40576
rect 22094 40536 22100 40548
rect 22152 40536 22158 40588
rect 22370 40536 22376 40588
rect 22428 40576 22434 40588
rect 22465 40579 22523 40585
rect 22465 40576 22477 40579
rect 22428 40548 22477 40576
rect 22428 40536 22434 40548
rect 22465 40545 22477 40548
rect 22511 40576 22523 40579
rect 30469 40579 30527 40585
rect 22511 40548 26924 40576
rect 22511 40545 22523 40548
rect 22465 40539 22523 40545
rect 21637 40511 21695 40517
rect 21637 40477 21649 40511
rect 21683 40508 21695 40511
rect 21726 40508 21732 40520
rect 21683 40480 21732 40508
rect 21683 40477 21695 40480
rect 21637 40471 21695 40477
rect 21726 40468 21732 40480
rect 21784 40508 21790 40520
rect 22388 40508 22416 40536
rect 26510 40508 26516 40520
rect 21784 40480 22416 40508
rect 26471 40480 26516 40508
rect 21784 40468 21790 40480
rect 26510 40468 26516 40480
rect 26568 40468 26574 40520
rect 26786 40508 26792 40520
rect 26747 40480 26792 40508
rect 26786 40468 26792 40480
rect 26844 40468 26850 40520
rect 26896 40508 26924 40548
rect 30469 40545 30481 40579
rect 30515 40576 30527 40579
rect 30926 40576 30932 40588
rect 30515 40548 30932 40576
rect 30515 40545 30527 40548
rect 30469 40539 30527 40545
rect 30926 40536 30932 40548
rect 30984 40536 30990 40588
rect 31036 40576 31064 40616
rect 31956 40576 31984 40675
rect 32030 40604 32036 40656
rect 32088 40644 32094 40656
rect 33686 40644 33692 40656
rect 32088 40616 33692 40644
rect 32088 40604 32094 40616
rect 32125 40579 32183 40585
rect 32125 40576 32137 40579
rect 31036 40548 32137 40576
rect 32125 40545 32137 40548
rect 32171 40545 32183 40579
rect 32125 40539 32183 40545
rect 32309 40579 32367 40585
rect 32309 40545 32321 40579
rect 32355 40576 32367 40579
rect 32766 40576 32772 40588
rect 32355 40548 32536 40576
rect 32727 40548 32772 40576
rect 32355 40545 32367 40548
rect 32309 40539 32367 40545
rect 31570 40508 31576 40520
rect 26896 40480 31576 40508
rect 31570 40468 31576 40480
rect 31628 40468 31634 40520
rect 31938 40468 31944 40520
rect 31996 40508 32002 40520
rect 32508 40508 32536 40548
rect 32766 40536 32772 40548
rect 32824 40536 32830 40588
rect 32876 40585 32904 40616
rect 33686 40604 33692 40616
rect 33744 40604 33750 40656
rect 37568 40653 37596 40684
rect 37642 40672 37648 40724
rect 37700 40712 37706 40724
rect 38470 40712 38476 40724
rect 37700 40684 38476 40712
rect 37700 40672 37706 40684
rect 38470 40672 38476 40684
rect 38528 40672 38534 40724
rect 43162 40712 43168 40724
rect 43123 40684 43168 40712
rect 43162 40672 43168 40684
rect 43220 40712 43226 40724
rect 43438 40712 43444 40724
rect 43220 40684 43444 40712
rect 43220 40672 43226 40684
rect 43438 40672 43444 40684
rect 43496 40672 43502 40724
rect 44174 40672 44180 40724
rect 44232 40712 44238 40724
rect 45097 40715 45155 40721
rect 45097 40712 45109 40715
rect 44232 40684 45109 40712
rect 44232 40672 44238 40684
rect 45097 40681 45109 40684
rect 45143 40712 45155 40715
rect 45554 40712 45560 40724
rect 45143 40684 45560 40712
rect 45143 40681 45155 40684
rect 45097 40675 45155 40681
rect 45554 40672 45560 40684
rect 45612 40672 45618 40724
rect 45922 40672 45928 40724
rect 45980 40712 45986 40724
rect 82722 40712 82728 40724
rect 45980 40684 82728 40712
rect 45980 40672 45986 40684
rect 82722 40672 82728 40684
rect 82780 40672 82786 40724
rect 82906 40712 82912 40724
rect 82867 40684 82912 40712
rect 82906 40672 82912 40684
rect 82964 40672 82970 40724
rect 88978 40712 88984 40724
rect 88939 40684 88984 40712
rect 88978 40672 88984 40684
rect 89036 40672 89042 40724
rect 37553 40647 37611 40653
rect 37553 40613 37565 40647
rect 37599 40644 37611 40647
rect 37599 40616 38424 40644
rect 37599 40613 37611 40616
rect 37553 40607 37611 40613
rect 32861 40579 32919 40585
rect 32861 40545 32873 40579
rect 32907 40545 32919 40579
rect 32861 40539 32919 40545
rect 37921 40579 37979 40585
rect 37921 40545 37933 40579
rect 37967 40576 37979 40579
rect 38102 40576 38108 40588
rect 37967 40548 38108 40576
rect 37967 40545 37979 40548
rect 37921 40539 37979 40545
rect 38102 40536 38108 40548
rect 38160 40536 38166 40588
rect 38396 40585 38424 40616
rect 38488 40585 38516 40672
rect 44637 40647 44695 40653
rect 43548 40616 44312 40644
rect 38381 40579 38439 40585
rect 38381 40545 38393 40579
rect 38427 40545 38439 40579
rect 38381 40539 38439 40545
rect 38473 40579 38531 40585
rect 38473 40545 38485 40579
rect 38519 40576 38531 40579
rect 39393 40579 39451 40585
rect 39393 40576 39405 40579
rect 38519 40548 39405 40576
rect 38519 40545 38531 40548
rect 38473 40539 38531 40545
rect 39393 40545 39405 40548
rect 39439 40545 39451 40579
rect 39393 40539 39451 40545
rect 42702 40536 42708 40588
rect 42760 40576 42766 40588
rect 43548 40585 43576 40616
rect 43533 40579 43591 40585
rect 43533 40576 43545 40579
rect 42760 40548 43545 40576
rect 42760 40536 42766 40548
rect 43533 40545 43545 40548
rect 43579 40545 43591 40579
rect 43993 40579 44051 40585
rect 43993 40576 44005 40579
rect 43533 40539 43591 40545
rect 43640 40548 44005 40576
rect 31996 40480 32536 40508
rect 31996 40468 32002 40480
rect 25038 40440 25044 40452
rect 21560 40412 25044 40440
rect 5031 40409 5043 40412
rect 4985 40403 5043 40409
rect 25038 40400 25044 40412
rect 25096 40400 25102 40452
rect 27614 40400 27620 40452
rect 27672 40440 27678 40452
rect 32214 40440 32220 40452
rect 27672 40412 32220 40440
rect 27672 40400 27678 40412
rect 32214 40400 32220 40412
rect 32272 40400 32278 40452
rect 32508 40440 32536 40480
rect 33413 40511 33471 40517
rect 33413 40477 33425 40511
rect 33459 40508 33471 40511
rect 34606 40508 34612 40520
rect 33459 40480 34612 40508
rect 33459 40477 33471 40480
rect 33413 40471 33471 40477
rect 34606 40468 34612 40480
rect 34664 40468 34670 40520
rect 37829 40511 37887 40517
rect 37829 40477 37841 40511
rect 37875 40508 37887 40511
rect 38010 40508 38016 40520
rect 37875 40480 38016 40508
rect 37875 40477 37887 40480
rect 37829 40471 37887 40477
rect 38010 40468 38016 40480
rect 38068 40468 38074 40520
rect 39025 40511 39083 40517
rect 39025 40477 39037 40511
rect 39071 40508 39083 40511
rect 40586 40508 40592 40520
rect 39071 40480 40592 40508
rect 39071 40477 39083 40480
rect 39025 40471 39083 40477
rect 40586 40468 40592 40480
rect 40644 40468 40650 40520
rect 42886 40468 42892 40520
rect 42944 40508 42950 40520
rect 43349 40511 43407 40517
rect 43349 40508 43361 40511
rect 42944 40480 43361 40508
rect 42944 40468 42950 40480
rect 43349 40477 43361 40480
rect 43395 40477 43407 40511
rect 43349 40471 43407 40477
rect 43438 40468 43444 40520
rect 43496 40508 43502 40520
rect 43640 40508 43668 40548
rect 43993 40545 44005 40548
rect 44039 40545 44051 40579
rect 43993 40539 44051 40545
rect 44085 40579 44143 40585
rect 44085 40545 44097 40579
rect 44131 40576 44143 40579
rect 44174 40576 44180 40588
rect 44131 40548 44180 40576
rect 44131 40545 44143 40548
rect 44085 40539 44143 40545
rect 44174 40536 44180 40548
rect 44232 40536 44238 40588
rect 44284 40576 44312 40616
rect 44637 40613 44649 40647
rect 44683 40644 44695 40647
rect 46382 40644 46388 40656
rect 44683 40616 46388 40644
rect 44683 40613 44695 40616
rect 44637 40607 44695 40613
rect 46382 40604 46388 40616
rect 46440 40604 46446 40656
rect 49421 40647 49479 40653
rect 49421 40613 49433 40647
rect 49467 40644 49479 40647
rect 50154 40644 50160 40656
rect 49467 40616 50160 40644
rect 49467 40613 49479 40616
rect 49421 40607 49479 40613
rect 50154 40604 50160 40616
rect 50212 40604 50218 40656
rect 54662 40644 54668 40656
rect 54623 40616 54668 40644
rect 54662 40604 54668 40616
rect 54720 40604 54726 40656
rect 81342 40644 81348 40656
rect 54772 40616 81204 40644
rect 81303 40616 81348 40644
rect 44284 40548 44956 40576
rect 44928 40517 44956 40548
rect 45186 40536 45192 40588
rect 45244 40576 45250 40588
rect 54772 40576 54800 40616
rect 45244 40548 54800 40576
rect 45244 40536 45250 40548
rect 54846 40536 54852 40588
rect 54904 40576 54910 40588
rect 57790 40576 57796 40588
rect 54904 40548 54949 40576
rect 57751 40548 57796 40576
rect 54904 40536 54910 40548
rect 57790 40536 57796 40548
rect 57848 40536 57854 40588
rect 58802 40576 58808 40588
rect 58763 40548 58808 40576
rect 58802 40536 58808 40548
rect 58860 40536 58866 40588
rect 62761 40579 62819 40585
rect 62761 40545 62773 40579
rect 62807 40545 62819 40579
rect 62942 40576 62948 40588
rect 62903 40548 62948 40576
rect 62761 40539 62819 40545
rect 43496 40480 43668 40508
rect 44913 40511 44971 40517
rect 43496 40468 43502 40480
rect 44913 40477 44925 40511
rect 44959 40508 44971 40511
rect 49510 40508 49516 40520
rect 44959 40480 49516 40508
rect 44959 40477 44971 40480
rect 44913 40471 44971 40477
rect 49510 40468 49516 40480
rect 49568 40468 49574 40520
rect 49786 40508 49792 40520
rect 49747 40480 49792 40508
rect 49786 40468 49792 40480
rect 49844 40468 49850 40520
rect 52638 40468 52644 40520
rect 52696 40508 52702 40520
rect 52914 40508 52920 40520
rect 52696 40480 52920 40508
rect 52696 40468 52702 40480
rect 52914 40468 52920 40480
rect 52972 40508 52978 40520
rect 54864 40508 54892 40536
rect 55122 40508 55128 40520
rect 52972 40480 54892 40508
rect 55083 40480 55128 40508
rect 52972 40468 52978 40480
rect 55122 40468 55128 40480
rect 55180 40468 55186 40520
rect 62776 40508 62804 40539
rect 62942 40536 62948 40548
rect 63000 40536 63006 40588
rect 63770 40576 63776 40588
rect 63052 40548 63776 40576
rect 63052 40508 63080 40548
rect 63770 40536 63776 40548
rect 63828 40536 63834 40588
rect 64322 40576 64328 40588
rect 64283 40548 64328 40576
rect 64322 40536 64328 40548
rect 64380 40536 64386 40588
rect 64417 40579 64475 40585
rect 64417 40545 64429 40579
rect 64463 40545 64475 40579
rect 64417 40539 64475 40545
rect 62776 40480 63080 40508
rect 63313 40511 63371 40517
rect 63313 40477 63325 40511
rect 63359 40508 63371 40511
rect 64432 40508 64460 40539
rect 64690 40536 64696 40588
rect 64748 40576 64754 40588
rect 65797 40579 65855 40585
rect 65797 40576 65809 40579
rect 64748 40548 65809 40576
rect 64748 40536 64754 40548
rect 65797 40545 65809 40548
rect 65843 40576 65855 40579
rect 66070 40576 66076 40588
rect 65843 40548 66076 40576
rect 65843 40545 65855 40548
rect 65797 40539 65855 40545
rect 66070 40536 66076 40548
rect 66128 40536 66134 40588
rect 66165 40579 66223 40585
rect 66165 40545 66177 40579
rect 66211 40576 66223 40579
rect 66254 40576 66260 40588
rect 66211 40548 66260 40576
rect 66211 40545 66223 40548
rect 66165 40539 66223 40545
rect 66254 40536 66260 40548
rect 66312 40536 66318 40588
rect 66346 40536 66352 40588
rect 66404 40576 66410 40588
rect 67358 40576 67364 40588
rect 66404 40548 66449 40576
rect 67319 40548 67364 40576
rect 66404 40536 66410 40548
rect 67358 40536 67364 40548
rect 67416 40536 67422 40588
rect 67450 40536 67456 40588
rect 67508 40576 67514 40588
rect 67545 40579 67603 40585
rect 67545 40576 67557 40579
rect 67508 40548 67557 40576
rect 67508 40536 67514 40548
rect 67545 40545 67557 40548
rect 67591 40545 67603 40579
rect 67910 40576 67916 40588
rect 67871 40548 67916 40576
rect 67545 40539 67603 40545
rect 67910 40536 67916 40548
rect 67968 40536 67974 40588
rect 71409 40579 71467 40585
rect 71409 40545 71421 40579
rect 71455 40576 71467 40579
rect 72970 40576 72976 40588
rect 71455 40548 72976 40576
rect 71455 40545 71467 40548
rect 71409 40539 71467 40545
rect 72970 40536 72976 40548
rect 73028 40536 73034 40588
rect 73062 40536 73068 40588
rect 73120 40576 73126 40588
rect 73430 40576 73436 40588
rect 73120 40548 73165 40576
rect 73391 40548 73436 40576
rect 73120 40536 73126 40548
rect 73430 40536 73436 40548
rect 73488 40536 73494 40588
rect 74718 40576 74724 40588
rect 74679 40548 74724 40576
rect 74718 40536 74724 40548
rect 74776 40536 74782 40588
rect 74902 40576 74908 40588
rect 74863 40548 74908 40576
rect 74902 40536 74908 40548
rect 74960 40576 74966 40588
rect 75365 40579 75423 40585
rect 75365 40576 75377 40579
rect 74960 40548 75377 40576
rect 74960 40536 74966 40548
rect 75365 40545 75377 40548
rect 75411 40545 75423 40579
rect 80793 40579 80851 40585
rect 80793 40576 80805 40579
rect 75365 40539 75423 40545
rect 80716 40548 80805 40576
rect 63359 40480 64460 40508
rect 63359 40477 63371 40480
rect 63313 40471 63371 40477
rect 64598 40468 64604 40520
rect 64656 40508 64662 40520
rect 64877 40511 64935 40517
rect 64877 40508 64889 40511
rect 64656 40480 64889 40508
rect 64656 40468 64662 40480
rect 64877 40477 64889 40480
rect 64923 40477 64935 40511
rect 64877 40471 64935 40477
rect 64966 40468 64972 40520
rect 65024 40508 65030 40520
rect 71038 40508 71044 40520
rect 65024 40480 71044 40508
rect 65024 40468 65030 40480
rect 71038 40468 71044 40480
rect 71096 40468 71102 40520
rect 71501 40511 71559 40517
rect 71501 40477 71513 40511
rect 71547 40508 71559 40511
rect 73080 40508 73108 40536
rect 71547 40480 73108 40508
rect 71547 40477 71559 40480
rect 71501 40471 71559 40477
rect 73154 40468 73160 40520
rect 73212 40508 73218 40520
rect 73522 40508 73528 40520
rect 73212 40480 73257 40508
rect 73435 40480 73528 40508
rect 73212 40468 73218 40480
rect 73522 40468 73528 40480
rect 73580 40508 73586 40520
rect 75181 40511 75239 40517
rect 75181 40508 75193 40511
rect 73580 40480 75193 40508
rect 73580 40468 73586 40480
rect 75181 40477 75193 40480
rect 75227 40477 75239 40511
rect 75380 40508 75408 40539
rect 80716 40508 80744 40548
rect 80793 40545 80805 40548
rect 80839 40576 80851 40579
rect 80882 40576 80888 40588
rect 80839 40548 80888 40576
rect 80839 40545 80851 40548
rect 80793 40539 80851 40545
rect 80882 40536 80888 40548
rect 80940 40536 80946 40588
rect 80977 40579 81035 40585
rect 80977 40545 80989 40579
rect 81023 40545 81035 40579
rect 80977 40539 81035 40545
rect 80992 40508 81020 40539
rect 75380 40480 80744 40508
rect 80808 40480 81020 40508
rect 81176 40508 81204 40616
rect 81342 40604 81348 40616
rect 81400 40604 81406 40656
rect 81434 40536 81440 40588
rect 81492 40576 81498 40588
rect 82633 40579 82691 40585
rect 82633 40576 82645 40579
rect 81492 40548 82645 40576
rect 81492 40536 81498 40548
rect 82633 40545 82645 40548
rect 82679 40545 82691 40579
rect 82740 40576 82768 40672
rect 85669 40647 85727 40653
rect 85669 40613 85681 40647
rect 85715 40644 85727 40647
rect 87598 40644 87604 40656
rect 85715 40616 87604 40644
rect 85715 40613 85727 40616
rect 85669 40607 85727 40613
rect 87598 40604 87604 40616
rect 87656 40604 87662 40656
rect 82817 40579 82875 40585
rect 82817 40576 82829 40579
rect 82740 40548 82829 40576
rect 82633 40539 82691 40545
rect 82817 40545 82829 40548
rect 82863 40576 82875 40579
rect 83277 40579 83335 40585
rect 83277 40576 83289 40579
rect 82863 40548 83289 40576
rect 82863 40545 82875 40548
rect 82817 40539 82875 40545
rect 83277 40545 83289 40548
rect 83323 40545 83335 40579
rect 86494 40576 86500 40588
rect 86455 40548 86500 40576
rect 83277 40539 83335 40545
rect 86494 40536 86500 40548
rect 86552 40536 86558 40588
rect 88996 40576 89024 40672
rect 89165 40579 89223 40585
rect 89165 40576 89177 40579
rect 88996 40548 89177 40576
rect 89165 40545 89177 40548
rect 89211 40545 89223 40579
rect 89165 40539 89223 40545
rect 82998 40508 83004 40520
rect 81176 40480 83004 40508
rect 75181 40471 75239 40477
rect 33226 40440 33232 40452
rect 32508 40412 33232 40440
rect 33226 40400 33232 40412
rect 33284 40400 33290 40452
rect 33318 40400 33324 40452
rect 33376 40440 33382 40452
rect 67266 40440 67272 40452
rect 33376 40412 67272 40440
rect 33376 40400 33382 40412
rect 67266 40400 67272 40412
rect 67324 40400 67330 40452
rect 75822 40400 75828 40452
rect 75880 40440 75886 40452
rect 78674 40440 78680 40452
rect 75880 40412 78680 40440
rect 75880 40400 75886 40412
rect 78674 40400 78680 40412
rect 78732 40400 78738 40452
rect 80808 40384 80836 40480
rect 82998 40468 83004 40480
rect 83056 40468 83062 40520
rect 86218 40508 86224 40520
rect 86179 40480 86224 40508
rect 86218 40468 86224 40480
rect 86276 40468 86282 40520
rect 86678 40508 86684 40520
rect 86639 40480 86684 40508
rect 86678 40468 86684 40480
rect 86736 40508 86742 40520
rect 86773 40511 86831 40517
rect 86773 40508 86785 40511
rect 86736 40480 86785 40508
rect 86736 40468 86742 40480
rect 86773 40477 86785 40480
rect 86819 40477 86831 40511
rect 89438 40508 89444 40520
rect 89399 40480 89444 40508
rect 86773 40471 86831 40477
rect 89438 40468 89444 40480
rect 89496 40468 89502 40520
rect 5718 40372 5724 40384
rect 5631 40344 5724 40372
rect 5718 40332 5724 40344
rect 5776 40372 5782 40384
rect 6362 40372 6368 40384
rect 5776 40344 6368 40372
rect 5776 40332 5782 40344
rect 6362 40332 6368 40344
rect 6420 40332 6426 40384
rect 7282 40332 7288 40384
rect 7340 40372 7346 40384
rect 7377 40375 7435 40381
rect 7377 40372 7389 40375
rect 7340 40344 7389 40372
rect 7340 40332 7346 40344
rect 7377 40341 7389 40344
rect 7423 40341 7435 40375
rect 7377 40335 7435 40341
rect 10318 40332 10324 40384
rect 10376 40372 10382 40384
rect 10962 40372 10968 40384
rect 10376 40344 10968 40372
rect 10376 40332 10382 40344
rect 10962 40332 10968 40344
rect 11020 40372 11026 40384
rect 11149 40375 11207 40381
rect 11149 40372 11161 40375
rect 11020 40344 11161 40372
rect 11020 40332 11026 40344
rect 11149 40341 11161 40344
rect 11195 40341 11207 40375
rect 13722 40372 13728 40384
rect 13683 40344 13728 40372
rect 11149 40335 11207 40341
rect 13722 40332 13728 40344
rect 13780 40332 13786 40384
rect 22094 40332 22100 40384
rect 22152 40372 22158 40384
rect 22281 40375 22339 40381
rect 22281 40372 22293 40375
rect 22152 40344 22293 40372
rect 22152 40332 22158 40344
rect 22281 40341 22293 40344
rect 22327 40372 22339 40375
rect 27522 40372 27528 40384
rect 22327 40344 27528 40372
rect 22327 40341 22339 40344
rect 22281 40335 22339 40341
rect 27522 40332 27528 40344
rect 27580 40332 27586 40384
rect 27890 40372 27896 40384
rect 27851 40344 27896 40372
rect 27890 40332 27896 40344
rect 27948 40332 27954 40384
rect 28258 40372 28264 40384
rect 28219 40344 28264 40372
rect 28258 40332 28264 40344
rect 28316 40372 28322 40384
rect 30285 40375 30343 40381
rect 30285 40372 30297 40375
rect 28316 40344 30297 40372
rect 28316 40332 28322 40344
rect 30285 40341 30297 40344
rect 30331 40341 30343 40375
rect 30285 40335 30343 40341
rect 33502 40332 33508 40384
rect 33560 40372 33566 40384
rect 33873 40375 33931 40381
rect 33873 40372 33885 40375
rect 33560 40344 33885 40372
rect 33560 40332 33566 40344
rect 33873 40341 33885 40344
rect 33919 40372 33931 40375
rect 37642 40372 37648 40384
rect 33919 40344 37648 40372
rect 33919 40341 33931 40344
rect 33873 40335 33931 40341
rect 37642 40332 37648 40344
rect 37700 40332 37706 40384
rect 39298 40372 39304 40384
rect 39259 40344 39304 40372
rect 39298 40332 39304 40344
rect 39356 40332 39362 40384
rect 42886 40372 42892 40384
rect 42847 40344 42892 40372
rect 42886 40332 42892 40344
rect 42944 40332 42950 40384
rect 43990 40332 43996 40384
rect 44048 40372 44054 40384
rect 45370 40372 45376 40384
rect 44048 40344 45376 40372
rect 44048 40332 44054 40344
rect 45370 40332 45376 40344
rect 45428 40332 45434 40384
rect 48314 40332 48320 40384
rect 48372 40372 48378 40384
rect 49559 40375 49617 40381
rect 49559 40372 49571 40375
rect 48372 40344 49571 40372
rect 48372 40332 48378 40344
rect 49559 40341 49571 40344
rect 49605 40341 49617 40375
rect 49559 40335 49617 40341
rect 49694 40332 49700 40384
rect 49752 40372 49758 40384
rect 50065 40375 50123 40381
rect 49752 40344 49797 40372
rect 49752 40332 49758 40344
rect 50065 40341 50077 40375
rect 50111 40372 50123 40375
rect 51442 40372 51448 40384
rect 50111 40344 51448 40372
rect 50111 40341 50123 40344
rect 50065 40335 50123 40341
rect 51442 40332 51448 40344
rect 51500 40332 51506 40384
rect 57698 40332 57704 40384
rect 57756 40372 57762 40384
rect 57885 40375 57943 40381
rect 57885 40372 57897 40375
rect 57756 40344 57897 40372
rect 57756 40332 57762 40344
rect 57885 40341 57897 40344
rect 57931 40341 57943 40375
rect 57885 40335 57943 40341
rect 58897 40375 58955 40381
rect 58897 40341 58909 40375
rect 58943 40372 58955 40375
rect 59170 40372 59176 40384
rect 58943 40344 59176 40372
rect 58943 40341 58955 40344
rect 58897 40335 58955 40341
rect 59170 40332 59176 40344
rect 59228 40332 59234 40384
rect 63586 40332 63592 40384
rect 63644 40372 63650 40384
rect 64141 40375 64199 40381
rect 64141 40372 64153 40375
rect 63644 40344 64153 40372
rect 63644 40332 63650 40344
rect 64141 40341 64153 40344
rect 64187 40372 64199 40375
rect 64966 40372 64972 40384
rect 64187 40344 64972 40372
rect 64187 40341 64199 40344
rect 64141 40335 64199 40341
rect 64966 40332 64972 40344
rect 65024 40332 65030 40384
rect 65426 40332 65432 40384
rect 65484 40372 65490 40384
rect 65521 40375 65579 40381
rect 65521 40372 65533 40375
rect 65484 40344 65533 40372
rect 65484 40332 65490 40344
rect 65521 40341 65533 40344
rect 65567 40372 65579 40375
rect 66346 40372 66352 40384
rect 65567 40344 66352 40372
rect 65567 40341 65579 40344
rect 65521 40335 65579 40341
rect 66346 40332 66352 40344
rect 66404 40372 66410 40384
rect 67177 40375 67235 40381
rect 67177 40372 67189 40375
rect 66404 40344 67189 40372
rect 66404 40332 66410 40344
rect 67177 40341 67189 40344
rect 67223 40372 67235 40375
rect 67358 40372 67364 40384
rect 67223 40344 67364 40372
rect 67223 40341 67235 40344
rect 67177 40335 67235 40341
rect 67358 40332 67364 40344
rect 67416 40332 67422 40384
rect 71958 40332 71964 40384
rect 72016 40372 72022 40384
rect 72513 40375 72571 40381
rect 72513 40372 72525 40375
rect 72016 40344 72525 40372
rect 72016 40332 72022 40344
rect 72513 40341 72525 40344
rect 72559 40341 72571 40375
rect 72513 40335 72571 40341
rect 73154 40332 73160 40384
rect 73212 40372 73218 40384
rect 73709 40375 73767 40381
rect 73709 40372 73721 40375
rect 73212 40344 73721 40372
rect 73212 40332 73218 40344
rect 73709 40341 73721 40344
rect 73755 40341 73767 40375
rect 73709 40335 73767 40341
rect 80701 40375 80759 40381
rect 80701 40341 80713 40375
rect 80747 40372 80759 40375
rect 80790 40372 80796 40384
rect 80747 40344 80796 40372
rect 80747 40341 80759 40344
rect 80701 40335 80759 40341
rect 80790 40332 80796 40344
rect 80848 40332 80854 40384
rect 80882 40332 80888 40384
rect 80940 40372 80946 40384
rect 81437 40375 81495 40381
rect 81437 40372 81449 40375
rect 80940 40344 81449 40372
rect 80940 40332 80946 40344
rect 81437 40341 81449 40344
rect 81483 40341 81495 40375
rect 81437 40335 81495 40341
rect 89898 40332 89904 40384
rect 89956 40372 89962 40384
rect 90545 40375 90603 40381
rect 90545 40372 90557 40375
rect 89956 40344 90557 40372
rect 89956 40332 89962 40344
rect 90545 40341 90557 40344
rect 90591 40341 90603 40375
rect 90545 40335 90603 40341
rect 1104 40282 105616 40304
rect 1104 40230 4246 40282
rect 4298 40230 4310 40282
rect 4362 40230 4374 40282
rect 4426 40230 4438 40282
rect 4490 40230 34966 40282
rect 35018 40230 35030 40282
rect 35082 40230 35094 40282
rect 35146 40230 35158 40282
rect 35210 40230 65686 40282
rect 65738 40230 65750 40282
rect 65802 40230 65814 40282
rect 65866 40230 65878 40282
rect 65930 40230 96406 40282
rect 96458 40230 96470 40282
rect 96522 40230 96534 40282
rect 96586 40230 96598 40282
rect 96650 40230 105616 40282
rect 1104 40208 105616 40230
rect 1486 40128 1492 40180
rect 1544 40168 1550 40180
rect 9674 40168 9680 40180
rect 1544 40140 9680 40168
rect 1544 40128 1550 40140
rect 9674 40128 9680 40140
rect 9732 40128 9738 40180
rect 12434 40128 12440 40180
rect 12492 40168 12498 40180
rect 13538 40168 13544 40180
rect 12492 40140 13544 40168
rect 12492 40128 12498 40140
rect 13538 40128 13544 40140
rect 13596 40128 13602 40180
rect 15378 40128 15384 40180
rect 15436 40168 15442 40180
rect 23842 40168 23848 40180
rect 15436 40140 23848 40168
rect 15436 40128 15442 40140
rect 23842 40128 23848 40140
rect 23900 40128 23906 40180
rect 26421 40171 26479 40177
rect 26421 40137 26433 40171
rect 26467 40168 26479 40171
rect 26786 40168 26792 40180
rect 26467 40140 26792 40168
rect 26467 40137 26479 40140
rect 26421 40131 26479 40137
rect 26786 40128 26792 40140
rect 26844 40128 26850 40180
rect 27338 40128 27344 40180
rect 27396 40168 27402 40180
rect 27525 40171 27583 40177
rect 27525 40168 27537 40171
rect 27396 40140 27537 40168
rect 27396 40128 27402 40140
rect 27525 40137 27537 40140
rect 27571 40168 27583 40171
rect 27982 40168 27988 40180
rect 27571 40140 27988 40168
rect 27571 40137 27583 40140
rect 27525 40131 27583 40137
rect 27982 40128 27988 40140
rect 28040 40128 28046 40180
rect 31754 40128 31760 40180
rect 31812 40168 31818 40180
rect 34698 40168 34704 40180
rect 31812 40140 34704 40168
rect 31812 40128 31818 40140
rect 34698 40128 34704 40140
rect 34756 40128 34762 40180
rect 38102 40128 38108 40180
rect 38160 40168 38166 40180
rect 38841 40171 38899 40177
rect 38841 40168 38853 40171
rect 38160 40140 38853 40168
rect 38160 40128 38166 40140
rect 38841 40137 38853 40140
rect 38887 40168 38899 40171
rect 39298 40168 39304 40180
rect 38887 40140 39304 40168
rect 38887 40137 38899 40140
rect 38841 40131 38899 40137
rect 39298 40128 39304 40140
rect 39356 40128 39362 40180
rect 40773 40171 40831 40177
rect 40773 40137 40785 40171
rect 40819 40168 40831 40171
rect 40819 40140 44588 40168
rect 40819 40137 40831 40140
rect 40773 40131 40831 40137
rect 3786 40100 3792 40112
rect 3747 40072 3792 40100
rect 3786 40060 3792 40072
rect 3844 40060 3850 40112
rect 4249 40103 4307 40109
rect 4249 40069 4261 40103
rect 4295 40100 4307 40103
rect 5718 40100 5724 40112
rect 4295 40072 5724 40100
rect 4295 40069 4307 40072
rect 4249 40063 4307 40069
rect 2593 40035 2651 40041
rect 2593 40001 2605 40035
rect 2639 40032 2651 40035
rect 2774 40032 2780 40044
rect 2639 40004 2780 40032
rect 2639 40001 2651 40004
rect 2593 39995 2651 40001
rect 2774 39992 2780 40004
rect 2832 40032 2838 40044
rect 2832 40004 3004 40032
rect 2832 39992 2838 40004
rect 2976 39976 3004 40004
rect 2869 39967 2927 39973
rect 2869 39933 2881 39967
rect 2915 39933 2927 39967
rect 2869 39927 2927 39933
rect 2884 39896 2912 39927
rect 2958 39924 2964 39976
rect 3016 39964 3022 39976
rect 3418 39964 3424 39976
rect 3016 39936 3061 39964
rect 3160 39936 3424 39964
rect 3016 39924 3022 39936
rect 3160 39896 3188 39936
rect 3418 39924 3424 39936
rect 3476 39924 3482 39976
rect 3605 39967 3663 39973
rect 3605 39933 3617 39967
rect 3651 39964 3663 39967
rect 4264 39964 4292 40063
rect 5718 40060 5724 40072
rect 5776 40060 5782 40112
rect 9122 40100 9128 40112
rect 8864 40072 9128 40100
rect 8297 40035 8355 40041
rect 8297 40001 8309 40035
rect 8343 40032 8355 40035
rect 8570 40032 8576 40044
rect 8343 40004 8576 40032
rect 8343 40001 8355 40004
rect 8297 39995 8355 40001
rect 8570 39992 8576 40004
rect 8628 39992 8634 40044
rect 3651 39936 4292 39964
rect 3651 39933 3663 39936
rect 3605 39927 3663 39933
rect 4798 39924 4804 39976
rect 4856 39964 4862 39976
rect 4893 39967 4951 39973
rect 4893 39964 4905 39967
rect 4856 39936 4905 39964
rect 4856 39924 4862 39936
rect 4893 39933 4905 39936
rect 4939 39933 4951 39967
rect 4893 39927 4951 39933
rect 5445 39967 5503 39973
rect 5445 39933 5457 39967
rect 5491 39933 5503 39967
rect 5445 39927 5503 39933
rect 2884 39868 3188 39896
rect 3234 39856 3240 39908
rect 3292 39896 3298 39908
rect 5460 39896 5488 39927
rect 8202 39924 8208 39976
rect 8260 39964 8266 39976
rect 8379 39967 8437 39973
rect 8379 39964 8391 39967
rect 8260 39936 8391 39964
rect 8260 39924 8266 39936
rect 8379 39933 8391 39936
rect 8425 39933 8437 39967
rect 8379 39927 8437 39933
rect 8478 39924 8484 39976
rect 8536 39964 8542 39976
rect 8864 39973 8892 40072
rect 9122 40060 9128 40072
rect 9180 40060 9186 40112
rect 12710 40100 12716 40112
rect 9784 40072 12716 40100
rect 8938 39992 8944 40044
rect 8996 40032 9002 40044
rect 9217 40035 9275 40041
rect 9217 40032 9229 40035
rect 8996 40004 9229 40032
rect 8996 39992 9002 40004
rect 9217 40001 9229 40004
rect 9263 40032 9275 40035
rect 9784 40032 9812 40072
rect 12710 40060 12716 40072
rect 12768 40060 12774 40112
rect 13722 40100 13728 40112
rect 13188 40072 13728 40100
rect 9263 40004 9812 40032
rect 9263 40001 9275 40004
rect 9217 39995 9275 40001
rect 12802 39992 12808 40044
rect 12860 40032 12866 40044
rect 12989 40035 13047 40041
rect 12989 40032 13001 40035
rect 12860 40004 13001 40032
rect 12860 39992 12866 40004
rect 12989 40001 13001 40004
rect 13035 40001 13047 40035
rect 12989 39995 13047 40001
rect 8757 39967 8815 39973
rect 8757 39964 8769 39967
rect 8536 39936 8769 39964
rect 8536 39924 8542 39936
rect 8757 39933 8769 39936
rect 8803 39933 8815 39967
rect 8757 39927 8815 39933
rect 8849 39967 8907 39973
rect 8849 39933 8861 39967
rect 8895 39933 8907 39967
rect 8849 39927 8907 39933
rect 12066 39924 12072 39976
rect 12124 39964 12130 39976
rect 13188 39973 13216 40072
rect 13722 40060 13728 40072
rect 13780 40060 13786 40112
rect 26510 40060 26516 40112
rect 26568 40100 26574 40112
rect 28258 40100 28264 40112
rect 26568 40072 28264 40100
rect 26568 40060 26574 40072
rect 28258 40060 28264 40072
rect 28316 40060 28322 40112
rect 31662 40060 31668 40112
rect 31720 40100 31726 40112
rect 32030 40100 32036 40112
rect 31720 40072 31800 40100
rect 31720 40060 31726 40072
rect 17773 40035 17831 40041
rect 17773 40032 17785 40035
rect 14476 40004 17785 40032
rect 13173 39967 13231 39973
rect 13173 39964 13185 39967
rect 12124 39936 13185 39964
rect 12124 39924 12130 39936
rect 13173 39933 13185 39936
rect 13219 39933 13231 39967
rect 13173 39927 13231 39933
rect 13722 39924 13728 39976
rect 13780 39964 13786 39976
rect 13906 39973 13912 39976
rect 13780 39936 13825 39964
rect 13780 39924 13786 39936
rect 13900 39927 13912 39973
rect 13964 39964 13970 39976
rect 14476 39973 14504 40004
rect 17773 40001 17785 40004
rect 17819 40001 17831 40035
rect 21450 40032 21456 40044
rect 17773 39995 17831 40001
rect 19996 40004 21456 40032
rect 14461 39967 14519 39973
rect 14461 39964 14473 39967
rect 13964 39936 14000 39964
rect 14384 39936 14473 39964
rect 13906 39924 13912 39927
rect 13964 39924 13970 39936
rect 12526 39896 12532 39908
rect 3292 39868 5028 39896
rect 5460 39868 12532 39896
rect 3292 39856 3298 39868
rect 5000 39837 5028 39868
rect 12526 39856 12532 39868
rect 12584 39856 12590 39908
rect 12618 39856 12624 39908
rect 12676 39896 12682 39908
rect 14274 39896 14280 39908
rect 12676 39868 13584 39896
rect 14235 39868 14280 39896
rect 12676 39856 12682 39868
rect 4985 39831 5043 39837
rect 4985 39797 4997 39831
rect 5031 39797 5043 39831
rect 4985 39791 5043 39797
rect 5902 39788 5908 39840
rect 5960 39828 5966 39840
rect 7837 39831 7895 39837
rect 7837 39828 7849 39831
rect 5960 39800 7849 39828
rect 5960 39788 5966 39800
rect 7837 39797 7849 39800
rect 7883 39797 7895 39831
rect 7837 39791 7895 39797
rect 7926 39788 7932 39840
rect 7984 39828 7990 39840
rect 11974 39828 11980 39840
rect 7984 39800 11980 39828
rect 7984 39788 7990 39800
rect 11974 39788 11980 39800
rect 12032 39788 12038 39840
rect 12710 39788 12716 39840
rect 12768 39828 12774 39840
rect 12805 39831 12863 39837
rect 12805 39828 12817 39831
rect 12768 39800 12817 39828
rect 12768 39788 12774 39800
rect 12805 39797 12817 39800
rect 12851 39797 12863 39831
rect 13556 39828 13584 39868
rect 14274 39856 14280 39868
rect 14332 39856 14338 39908
rect 13906 39828 13912 39840
rect 13556 39800 13912 39828
rect 12805 39791 12863 39797
rect 13906 39788 13912 39800
rect 13964 39828 13970 39840
rect 14384 39828 14412 39936
rect 14461 39933 14473 39936
rect 14507 39933 14519 39967
rect 15194 39964 15200 39976
rect 15155 39936 15200 39964
rect 14461 39927 14519 39933
rect 15194 39924 15200 39936
rect 15252 39924 15258 39976
rect 19334 39924 19340 39976
rect 19392 39964 19398 39976
rect 19996 39973 20024 40004
rect 21450 39992 21456 40004
rect 21508 40032 21514 40044
rect 31772 40041 31800 40072
rect 31956 40072 32036 40100
rect 21729 40035 21787 40041
rect 21729 40032 21741 40035
rect 21508 40004 21741 40032
rect 21508 39992 21514 40004
rect 21729 40001 21741 40004
rect 21775 40001 21787 40035
rect 21729 39995 21787 40001
rect 25133 40035 25191 40041
rect 25133 40001 25145 40035
rect 25179 40032 25191 40035
rect 31757 40035 31815 40041
rect 25179 40004 25544 40032
rect 25179 40001 25191 40004
rect 25133 39995 25191 40001
rect 19981 39967 20039 39973
rect 19981 39964 19993 39967
rect 19392 39936 19993 39964
rect 19392 39924 19398 39936
rect 19981 39933 19993 39936
rect 20027 39933 20039 39967
rect 19981 39927 20039 39933
rect 20257 39967 20315 39973
rect 20257 39933 20269 39967
rect 20303 39964 20315 39967
rect 21174 39964 21180 39976
rect 20303 39936 21180 39964
rect 20303 39933 20315 39936
rect 20257 39927 20315 39933
rect 21174 39924 21180 39936
rect 21232 39924 21238 39976
rect 25406 39964 25412 39976
rect 25367 39936 25412 39964
rect 25406 39924 25412 39936
rect 25464 39924 25470 39976
rect 25516 39973 25544 40004
rect 31757 40001 31769 40035
rect 31803 40001 31815 40035
rect 31757 39995 31815 40001
rect 25501 39967 25559 39973
rect 25501 39933 25513 39967
rect 25547 39964 25559 39967
rect 25774 39964 25780 39976
rect 25547 39936 25780 39964
rect 25547 39933 25559 39936
rect 25501 39927 25559 39933
rect 25774 39924 25780 39936
rect 25832 39924 25838 39976
rect 25958 39924 25964 39976
rect 26016 39964 26022 39976
rect 26016 39936 26061 39964
rect 26016 39924 26022 39936
rect 26142 39924 26148 39976
rect 26200 39964 26206 39976
rect 26789 39967 26847 39973
rect 26789 39964 26801 39967
rect 26200 39936 26801 39964
rect 26200 39924 26206 39936
rect 26789 39933 26801 39936
rect 26835 39964 26847 39967
rect 27338 39964 27344 39976
rect 26835 39936 27344 39964
rect 26835 39933 26847 39936
rect 26789 39927 26847 39933
rect 27338 39924 27344 39936
rect 27396 39924 27402 39976
rect 27433 39967 27491 39973
rect 27433 39933 27445 39967
rect 27479 39964 27491 39967
rect 27890 39964 27896 39976
rect 27479 39936 27896 39964
rect 27479 39933 27491 39936
rect 27433 39927 27491 39933
rect 27890 39924 27896 39936
rect 27948 39924 27954 39976
rect 28074 39924 28080 39976
rect 28132 39964 28138 39976
rect 28994 39964 29000 39976
rect 28132 39936 29000 39964
rect 28132 39924 28138 39936
rect 28994 39924 29000 39936
rect 29052 39924 29058 39976
rect 31956 39973 31984 40072
rect 32030 40060 32036 40072
rect 32088 40060 32094 40112
rect 33505 40103 33563 40109
rect 33505 40069 33517 40103
rect 33551 40100 33563 40103
rect 33870 40100 33876 40112
rect 33551 40072 33876 40100
rect 33551 40069 33563 40072
rect 33505 40063 33563 40069
rect 33520 40032 33548 40063
rect 33870 40060 33876 40072
rect 33928 40100 33934 40112
rect 37366 40100 37372 40112
rect 33928 40072 37372 40100
rect 33928 40060 33934 40072
rect 37366 40060 37372 40072
rect 37424 40060 37430 40112
rect 38930 40100 38936 40112
rect 38891 40072 38936 40100
rect 38930 40060 38936 40072
rect 38988 40060 38994 40112
rect 40494 40060 40500 40112
rect 40552 40060 40558 40112
rect 42245 40103 42303 40109
rect 42245 40069 42257 40103
rect 42291 40069 42303 40103
rect 44560 40100 44588 40140
rect 48222 40128 48228 40180
rect 48280 40168 48286 40180
rect 64874 40168 64880 40180
rect 48280 40140 64880 40168
rect 48280 40128 48286 40140
rect 64874 40128 64880 40140
rect 64932 40128 64938 40180
rect 64966 40128 64972 40180
rect 65024 40168 65030 40180
rect 66717 40171 66775 40177
rect 66717 40168 66729 40171
rect 65024 40140 66729 40168
rect 65024 40128 65030 40140
rect 66717 40137 66729 40140
rect 66763 40137 66775 40171
rect 66717 40131 66775 40137
rect 49142 40100 49148 40112
rect 44560 40072 49148 40100
rect 42245 40063 42303 40069
rect 32876 40004 33548 40032
rect 31941 39967 31999 39973
rect 31941 39933 31953 39967
rect 31987 39933 31999 39967
rect 32398 39964 32404 39976
rect 32359 39936 32404 39964
rect 31941 39927 31999 39933
rect 32398 39924 32404 39936
rect 32456 39924 32462 39976
rect 32493 39967 32551 39973
rect 32493 39933 32505 39967
rect 32539 39964 32551 39967
rect 32876 39964 32904 40004
rect 34422 39992 34428 40044
rect 34480 40032 34486 40044
rect 34480 40004 37688 40032
rect 34480 39992 34486 40004
rect 32539 39936 32904 39964
rect 33321 39967 33379 39973
rect 32539 39933 32551 39936
rect 32493 39927 32551 39933
rect 33321 39933 33333 39967
rect 33367 39964 33379 39967
rect 33686 39964 33692 39976
rect 33367 39936 33692 39964
rect 33367 39933 33379 39936
rect 33321 39927 33379 39933
rect 33686 39924 33692 39936
rect 33744 39924 33750 39976
rect 37277 39967 37335 39973
rect 37277 39964 37289 39967
rect 37108 39936 37289 39964
rect 20990 39856 20996 39908
rect 21048 39896 21054 39908
rect 31570 39896 31576 39908
rect 21048 39868 30420 39896
rect 31531 39868 31576 39896
rect 21048 39856 21054 39868
rect 13964 39800 14412 39828
rect 15381 39831 15439 39837
rect 13964 39788 13970 39800
rect 15381 39797 15393 39831
rect 15427 39828 15439 39831
rect 16022 39828 16028 39840
rect 15427 39800 16028 39828
rect 15427 39797 15439 39800
rect 15381 39791 15439 39797
rect 16022 39788 16028 39800
rect 16080 39788 16086 39840
rect 17773 39831 17831 39837
rect 17773 39797 17785 39831
rect 17819 39828 17831 39831
rect 21358 39828 21364 39840
rect 17819 39800 21364 39828
rect 17819 39797 17831 39800
rect 17773 39791 17831 39797
rect 21358 39788 21364 39800
rect 21416 39788 21422 39840
rect 21542 39828 21548 39840
rect 21455 39800 21548 39828
rect 21542 39788 21548 39800
rect 21600 39828 21606 39840
rect 30282 39828 30288 39840
rect 21600 39800 30288 39828
rect 21600 39788 21606 39800
rect 30282 39788 30288 39800
rect 30340 39788 30346 39840
rect 30392 39828 30420 39868
rect 31570 39856 31576 39868
rect 31628 39856 31634 39908
rect 32306 39828 32312 39840
rect 30392 39800 32312 39828
rect 32306 39788 32312 39800
rect 32364 39788 32370 39840
rect 32416 39828 32444 39924
rect 33045 39899 33103 39905
rect 33045 39865 33057 39899
rect 33091 39896 33103 39899
rect 34330 39896 34336 39908
rect 33091 39868 34336 39896
rect 33091 39865 33103 39868
rect 33045 39859 33103 39865
rect 34330 39856 34336 39868
rect 34388 39856 34394 39908
rect 37108 39837 37136 39936
rect 37277 39933 37289 39936
rect 37323 39933 37335 39967
rect 37277 39927 37335 39933
rect 37366 39924 37372 39976
rect 37424 39964 37430 39976
rect 37461 39967 37519 39973
rect 37461 39964 37473 39967
rect 37424 39936 37473 39964
rect 37424 39924 37430 39936
rect 37461 39933 37473 39936
rect 37507 39964 37519 39967
rect 37550 39964 37556 39976
rect 37507 39936 37556 39964
rect 37507 39933 37519 39936
rect 37461 39927 37519 39933
rect 37550 39924 37556 39936
rect 37608 39924 37614 39976
rect 37660 39964 37688 40004
rect 38654 39992 38660 40044
rect 38712 40032 38718 40044
rect 40512 40032 40540 40060
rect 38712 40004 40540 40032
rect 38712 39992 38718 40004
rect 40586 39992 40592 40044
rect 40644 40041 40650 40044
rect 40644 40035 40702 40041
rect 40644 40001 40656 40035
rect 40690 40001 40702 40035
rect 40644 39995 40702 40001
rect 40865 40035 40923 40041
rect 40865 40001 40877 40035
rect 40911 40001 40923 40035
rect 40865 39995 40923 40001
rect 40644 39992 40650 39995
rect 37918 39964 37924 39976
rect 37660 39936 37924 39964
rect 37918 39924 37924 39936
rect 37976 39924 37982 39976
rect 38013 39967 38071 39973
rect 38013 39933 38025 39967
rect 38059 39964 38071 39967
rect 38102 39964 38108 39976
rect 38059 39936 38108 39964
rect 38059 39933 38071 39936
rect 38013 39927 38071 39933
rect 38102 39924 38108 39936
rect 38160 39924 38166 39976
rect 40402 39924 40408 39976
rect 40460 39964 40466 39976
rect 40497 39967 40555 39973
rect 40497 39964 40509 39967
rect 40460 39936 40509 39964
rect 40460 39924 40466 39936
rect 40497 39933 40509 39936
rect 40543 39933 40555 39967
rect 40497 39927 40555 39933
rect 38565 39899 38623 39905
rect 38565 39865 38577 39899
rect 38611 39896 38623 39899
rect 40880 39896 40908 39995
rect 40954 39924 40960 39976
rect 41012 39964 41018 39976
rect 42260 39964 42288 40063
rect 49142 40060 49148 40072
rect 49200 40060 49206 40112
rect 49467 40103 49525 40109
rect 49467 40100 49479 40103
rect 49344 40072 49479 40100
rect 49344 40044 49372 40072
rect 49467 40069 49479 40072
rect 49513 40069 49525 40103
rect 49467 40063 49525 40069
rect 49605 40103 49663 40109
rect 49605 40069 49617 40103
rect 49651 40069 49663 40103
rect 49605 40063 49663 40069
rect 43530 40032 43536 40044
rect 43491 40004 43536 40032
rect 43530 39992 43536 40004
rect 43588 39992 43594 40044
rect 44821 40035 44879 40041
rect 44821 40001 44833 40035
rect 44867 40032 44879 40035
rect 48314 40032 48320 40044
rect 44867 40004 48320 40032
rect 44867 40001 44879 40004
rect 44821 39995 44879 40001
rect 48314 39992 48320 40004
rect 48372 39992 48378 40044
rect 49326 39992 49332 40044
rect 49384 39992 49390 40044
rect 49620 40032 49648 40063
rect 49786 40060 49792 40112
rect 49844 40100 49850 40112
rect 52917 40103 52975 40109
rect 52917 40100 52929 40103
rect 49844 40072 52929 40100
rect 49844 40060 49850 40072
rect 52917 40069 52929 40072
rect 52963 40069 52975 40103
rect 66732 40100 66760 40131
rect 77202 40128 77208 40180
rect 77260 40168 77266 40180
rect 79870 40168 79876 40180
rect 77260 40140 79876 40168
rect 77260 40128 77266 40140
rect 79870 40128 79876 40140
rect 79928 40128 79934 40180
rect 67542 40100 67548 40112
rect 66732 40072 67548 40100
rect 52917 40063 52975 40069
rect 67542 40060 67548 40072
rect 67600 40060 67606 40112
rect 70762 40100 70768 40112
rect 70504 40072 70768 40100
rect 49436 40004 49648 40032
rect 49697 40035 49755 40041
rect 41012 39936 42288 39964
rect 42429 39967 42487 39973
rect 41012 39924 41018 39936
rect 42429 39933 42441 39967
rect 42475 39964 42487 39967
rect 43717 39967 43775 39973
rect 42475 39936 42656 39964
rect 42475 39933 42487 39936
rect 42429 39927 42487 39933
rect 38611 39868 40908 39896
rect 38611 39865 38623 39868
rect 38565 39859 38623 39865
rect 37093 39831 37151 39837
rect 37093 39828 37105 39831
rect 32416 39800 37105 39828
rect 37093 39797 37105 39800
rect 37139 39797 37151 39831
rect 37093 39791 37151 39797
rect 37734 39788 37740 39840
rect 37792 39828 37798 39840
rect 38930 39828 38936 39840
rect 37792 39800 38936 39828
rect 37792 39788 37798 39800
rect 38930 39788 38936 39800
rect 38988 39788 38994 39840
rect 40310 39788 40316 39840
rect 40368 39828 40374 39840
rect 40954 39828 40960 39840
rect 40368 39800 40960 39828
rect 40368 39788 40374 39800
rect 40954 39788 40960 39800
rect 41012 39788 41018 39840
rect 41138 39828 41144 39840
rect 41099 39800 41144 39828
rect 41138 39788 41144 39800
rect 41196 39788 41202 39840
rect 42628 39837 42656 39936
rect 43717 39933 43729 39967
rect 43763 39964 43775 39967
rect 43898 39964 43904 39976
rect 43763 39936 43904 39964
rect 43763 39933 43775 39936
rect 43717 39927 43775 39933
rect 43898 39924 43904 39936
rect 43956 39924 43962 39976
rect 44174 39964 44180 39976
rect 44135 39936 44180 39964
rect 44174 39924 44180 39936
rect 44232 39924 44238 39976
rect 44269 39967 44327 39973
rect 44269 39933 44281 39967
rect 44315 39964 44327 39967
rect 45094 39964 45100 39976
rect 44315 39936 45100 39964
rect 44315 39933 44327 39936
rect 44269 39927 44327 39933
rect 45094 39924 45100 39936
rect 45152 39924 45158 39976
rect 49234 39964 49240 39976
rect 45204 39936 49240 39964
rect 42794 39856 42800 39908
rect 42852 39896 42858 39908
rect 45204 39896 45232 39936
rect 49234 39924 49240 39936
rect 49292 39924 49298 39976
rect 49326 39896 49332 39908
rect 42852 39868 45232 39896
rect 49287 39868 49332 39896
rect 42852 39856 42858 39868
rect 49326 39856 49332 39868
rect 49384 39856 49390 39908
rect 42613 39831 42671 39837
rect 42613 39797 42625 39831
rect 42659 39828 42671 39831
rect 44266 39828 44272 39840
rect 42659 39800 44272 39828
rect 42659 39797 42671 39800
rect 42613 39791 42671 39797
rect 44266 39788 44272 39800
rect 44324 39788 44330 39840
rect 45094 39788 45100 39840
rect 45152 39828 45158 39840
rect 49436 39828 49464 40004
rect 49697 40001 49709 40035
rect 49743 40001 49755 40035
rect 49697 39995 49755 40001
rect 45152 39800 49464 39828
rect 45152 39788 45158 39800
rect 49602 39788 49608 39840
rect 49660 39828 49666 39840
rect 49712 39828 49740 39995
rect 53098 39992 53104 40044
rect 53156 40032 53162 40044
rect 70504 40032 70532 40072
rect 70762 40060 70768 40072
rect 70820 40060 70826 40112
rect 72142 40100 72148 40112
rect 72103 40072 72148 40100
rect 72142 40060 72148 40072
rect 72200 40060 72206 40112
rect 80146 40060 80152 40112
rect 80204 40100 80210 40112
rect 85669 40103 85727 40109
rect 80204 40072 85528 40100
rect 80204 40060 80210 40072
rect 73338 40032 73344 40044
rect 53156 40004 64736 40032
rect 53156 39992 53162 40004
rect 50065 39967 50123 39973
rect 50065 39933 50077 39967
rect 50111 39964 50123 39967
rect 51810 39964 51816 39976
rect 50111 39936 51816 39964
rect 50111 39933 50123 39936
rect 50065 39927 50123 39933
rect 51810 39924 51816 39936
rect 51868 39924 51874 39976
rect 51994 39964 52000 39976
rect 51955 39936 52000 39964
rect 51994 39924 52000 39936
rect 52052 39924 52058 39976
rect 52089 39967 52147 39973
rect 52089 39933 52101 39967
rect 52135 39964 52147 39967
rect 52362 39964 52368 39976
rect 52135 39936 52368 39964
rect 52135 39933 52147 39936
rect 52089 39927 52147 39933
rect 52362 39924 52368 39936
rect 52420 39924 52426 39976
rect 52457 39967 52515 39973
rect 52457 39933 52469 39967
rect 52503 39933 52515 39967
rect 52457 39927 52515 39933
rect 52549 39967 52607 39973
rect 52549 39933 52561 39967
rect 52595 39933 52607 39967
rect 52549 39927 52607 39933
rect 51537 39899 51595 39905
rect 51537 39865 51549 39899
rect 51583 39896 51595 39899
rect 52472 39896 52500 39927
rect 52564 39896 52592 39927
rect 53282 39924 53288 39976
rect 53340 39964 53346 39976
rect 54297 39967 54355 39973
rect 54297 39964 54309 39967
rect 53340 39936 54309 39964
rect 53340 39924 53346 39936
rect 54297 39933 54309 39936
rect 54343 39964 54355 39967
rect 54570 39964 54576 39976
rect 54343 39936 54576 39964
rect 54343 39933 54355 39936
rect 54297 39927 54355 39933
rect 54570 39924 54576 39936
rect 54628 39924 54634 39976
rect 57057 39967 57115 39973
rect 57057 39964 57069 39967
rect 55968 39936 57069 39964
rect 52638 39896 52644 39908
rect 51583 39868 52500 39896
rect 52551 39868 52644 39896
rect 51583 39865 51595 39868
rect 51537 39859 51595 39865
rect 49660 39800 49740 39828
rect 49660 39788 49666 39800
rect 50062 39788 50068 39840
rect 50120 39828 50126 39840
rect 51552 39828 51580 39859
rect 52638 39856 52644 39868
rect 52696 39896 52702 39908
rect 52696 39868 53604 39896
rect 52696 39856 52702 39868
rect 53576 39840 53604 39868
rect 50120 39800 51580 39828
rect 50120 39788 50126 39800
rect 52086 39788 52092 39840
rect 52144 39828 52150 39840
rect 53374 39828 53380 39840
rect 52144 39800 53380 39828
rect 52144 39788 52150 39800
rect 53374 39788 53380 39800
rect 53432 39788 53438 39840
rect 53558 39828 53564 39840
rect 53519 39800 53564 39828
rect 53558 39788 53564 39800
rect 53616 39788 53622 39840
rect 54113 39831 54171 39837
rect 54113 39797 54125 39831
rect 54159 39828 54171 39831
rect 54662 39828 54668 39840
rect 54159 39800 54668 39828
rect 54159 39797 54171 39800
rect 54113 39791 54171 39797
rect 54662 39788 54668 39800
rect 54720 39828 54726 39840
rect 55968 39828 55996 39936
rect 57057 39933 57069 39936
rect 57103 39964 57115 39967
rect 57333 39967 57391 39973
rect 57333 39964 57345 39967
rect 57103 39936 57345 39964
rect 57103 39933 57115 39936
rect 57057 39927 57115 39933
rect 57333 39933 57345 39936
rect 57379 39933 57391 39967
rect 57609 39967 57667 39973
rect 57609 39964 57621 39967
rect 57333 39927 57391 39933
rect 57440 39936 57621 39964
rect 57440 39896 57468 39936
rect 57609 39933 57621 39936
rect 57655 39933 57667 39967
rect 57609 39927 57667 39933
rect 58066 39924 58072 39976
rect 58124 39964 58130 39976
rect 58618 39964 58624 39976
rect 58124 39936 58624 39964
rect 58124 39924 58130 39936
rect 58618 39924 58624 39936
rect 58676 39964 58682 39976
rect 62942 39964 62948 39976
rect 58676 39936 62948 39964
rect 58676 39924 58682 39936
rect 62942 39924 62948 39936
rect 63000 39964 63006 39976
rect 63221 39967 63279 39973
rect 63221 39964 63233 39967
rect 63000 39936 63233 39964
rect 63000 39924 63006 39936
rect 63221 39933 63233 39936
rect 63267 39964 63279 39967
rect 64138 39964 64144 39976
rect 63267 39936 64144 39964
rect 63267 39933 63279 39936
rect 63221 39927 63279 39933
rect 64138 39924 64144 39936
rect 64196 39924 64202 39976
rect 64233 39967 64291 39973
rect 64233 39933 64245 39967
rect 64279 39933 64291 39967
rect 64233 39927 64291 39933
rect 64509 39967 64567 39973
rect 64509 39933 64521 39967
rect 64555 39964 64567 39967
rect 64598 39964 64604 39976
rect 64555 39936 64604 39964
rect 64555 39933 64567 39936
rect 64509 39927 64567 39933
rect 56796 39868 57468 39896
rect 56796 39840 56824 39868
rect 58802 39856 58808 39908
rect 58860 39896 58866 39908
rect 58989 39899 59047 39905
rect 58989 39896 59001 39899
rect 58860 39868 59001 39896
rect 58860 39856 58866 39868
rect 58989 39865 59001 39868
rect 59035 39896 59047 39899
rect 61194 39896 61200 39908
rect 59035 39868 61200 39896
rect 59035 39865 59047 39868
rect 58989 39859 59047 39865
rect 61194 39856 61200 39868
rect 61252 39856 61258 39908
rect 63313 39899 63371 39905
rect 63313 39865 63325 39899
rect 63359 39896 63371 39899
rect 63494 39896 63500 39908
rect 63359 39868 63500 39896
rect 63359 39865 63371 39868
rect 63313 39859 63371 39865
rect 63494 39856 63500 39868
rect 63552 39856 63558 39908
rect 64248 39896 64276 39927
rect 64598 39924 64604 39936
rect 64656 39924 64662 39976
rect 64708 39964 64736 40004
rect 66824 40004 70532 40032
rect 70596 40004 73344 40032
rect 66824 39964 66852 40004
rect 66990 39964 66996 39976
rect 64708 39936 66852 39964
rect 66951 39936 66996 39964
rect 66990 39924 66996 39936
rect 67048 39924 67054 39976
rect 67910 39964 67916 39976
rect 67284 39936 67916 39964
rect 64156 39868 64276 39896
rect 66901 39899 66959 39905
rect 64156 39840 64184 39868
rect 66901 39865 66913 39899
rect 66947 39896 66959 39899
rect 67284 39896 67312 39936
rect 67910 39924 67916 39936
rect 67968 39924 67974 39976
rect 67450 39896 67456 39908
rect 66947 39868 67312 39896
rect 67411 39868 67456 39896
rect 66947 39865 66959 39868
rect 66901 39859 66959 39865
rect 67450 39856 67456 39868
rect 67508 39856 67514 39908
rect 70596 39896 70624 40004
rect 73338 39992 73344 40004
rect 73396 39992 73402 40044
rect 74166 40032 74172 40044
rect 74127 40004 74172 40032
rect 74166 39992 74172 40004
rect 74224 39992 74230 40044
rect 79410 40032 79416 40044
rect 79371 40004 79416 40032
rect 79410 39992 79416 40004
rect 79468 39992 79474 40044
rect 79502 39992 79508 40044
rect 79560 40032 79566 40044
rect 82354 40032 82360 40044
rect 79560 40004 81572 40032
rect 82315 40004 82360 40032
rect 79560 39992 79566 40004
rect 70673 39967 70731 39973
rect 70673 39933 70685 39967
rect 70719 39964 70731 39967
rect 70765 39967 70823 39973
rect 70765 39964 70777 39967
rect 70719 39936 70777 39964
rect 70719 39933 70731 39936
rect 70673 39927 70731 39933
rect 70765 39933 70777 39936
rect 70811 39933 70823 39967
rect 71038 39964 71044 39976
rect 70999 39936 71044 39964
rect 70765 39927 70823 39933
rect 67560 39868 70624 39896
rect 56778 39828 56784 39840
rect 54720 39800 55996 39828
rect 56739 39800 56784 39828
rect 54720 39788 54726 39800
rect 56778 39788 56784 39800
rect 56836 39788 56842 39840
rect 57882 39788 57888 39840
rect 57940 39828 57946 39840
rect 61654 39828 61660 39840
rect 57940 39800 61660 39828
rect 57940 39788 57946 39800
rect 61654 39788 61660 39800
rect 61712 39788 61718 39840
rect 64138 39828 64144 39840
rect 64099 39800 64144 39828
rect 64138 39788 64144 39800
rect 64196 39788 64202 39840
rect 64230 39788 64236 39840
rect 64288 39828 64294 39840
rect 65613 39831 65671 39837
rect 65613 39828 65625 39831
rect 64288 39800 65625 39828
rect 64288 39788 64294 39800
rect 65613 39797 65625 39800
rect 65659 39797 65671 39831
rect 65613 39791 65671 39797
rect 65702 39788 65708 39840
rect 65760 39828 65766 39840
rect 67560 39828 67588 39868
rect 65760 39800 67588 39828
rect 65760 39788 65766 39800
rect 67634 39788 67640 39840
rect 67692 39828 67698 39840
rect 70688 39828 70716 39927
rect 71038 39924 71044 39936
rect 71096 39924 71102 39976
rect 73982 39964 73988 39976
rect 73943 39936 73988 39964
rect 73982 39924 73988 39936
rect 74040 39924 74046 39976
rect 74442 39964 74448 39976
rect 74403 39936 74448 39964
rect 74442 39924 74448 39936
rect 74500 39924 74506 39976
rect 77478 39964 77484 39976
rect 77439 39936 77484 39964
rect 77478 39924 77484 39936
rect 77536 39964 77542 39976
rect 77757 39967 77815 39973
rect 77757 39964 77769 39967
rect 77536 39936 77769 39964
rect 77536 39924 77542 39936
rect 77757 39933 77769 39936
rect 77803 39933 77815 39967
rect 79428 39964 79456 39992
rect 80330 39964 80336 39976
rect 79428 39936 80336 39964
rect 77757 39927 77815 39933
rect 80330 39924 80336 39936
rect 80388 39924 80394 39976
rect 80425 39967 80483 39973
rect 80425 39933 80437 39967
rect 80471 39933 80483 39967
rect 80425 39927 80483 39933
rect 74350 39896 74356 39908
rect 73724 39868 74212 39896
rect 74311 39868 74356 39896
rect 67692 39800 70716 39828
rect 67692 39788 67698 39800
rect 70762 39788 70768 39840
rect 70820 39828 70826 39840
rect 73724 39828 73752 39868
rect 70820 39800 73752 39828
rect 73801 39831 73859 39837
rect 70820 39788 70826 39800
rect 73801 39797 73813 39831
rect 73847 39828 73859 39831
rect 73890 39828 73896 39840
rect 73847 39800 73896 39828
rect 73847 39797 73859 39800
rect 73801 39791 73859 39797
rect 73890 39788 73896 39800
rect 73948 39788 73954 39840
rect 74184 39828 74212 39868
rect 74350 39856 74356 39868
rect 74408 39856 74414 39908
rect 74902 39896 74908 39908
rect 74863 39868 74908 39896
rect 74902 39856 74908 39868
rect 74960 39856 74966 39908
rect 79781 39899 79839 39905
rect 79781 39865 79793 39899
rect 79827 39896 79839 39899
rect 79870 39896 79876 39908
rect 79827 39868 79876 39896
rect 79827 39865 79839 39868
rect 79781 39859 79839 39865
rect 79870 39856 79876 39868
rect 79928 39856 79934 39908
rect 80440 39896 80468 39927
rect 80514 39924 80520 39976
rect 80572 39964 80578 39976
rect 80790 39964 80796 39976
rect 80572 39936 80617 39964
rect 80751 39936 80796 39964
rect 80572 39924 80578 39936
rect 80790 39924 80796 39936
rect 80848 39924 80854 39976
rect 80882 39924 80888 39976
rect 80940 39964 80946 39976
rect 81544 39964 81572 40004
rect 82354 39992 82360 40004
rect 82412 39992 82418 40044
rect 83093 40035 83151 40041
rect 83093 40032 83105 40035
rect 82464 40004 83105 40032
rect 82464 39964 82492 40004
rect 83093 40001 83105 40004
rect 83139 40001 83151 40035
rect 84565 40035 84623 40041
rect 84565 40032 84577 40035
rect 83093 39995 83151 40001
rect 84212 40004 84577 40032
rect 80940 39936 80985 39964
rect 81544 39936 82492 39964
rect 82633 39967 82691 39973
rect 80940 39924 80946 39936
rect 82633 39933 82645 39967
rect 82679 39964 82691 39967
rect 82722 39964 82728 39976
rect 82679 39936 82728 39964
rect 82679 39933 82691 39936
rect 82633 39927 82691 39933
rect 82722 39924 82728 39936
rect 82780 39924 82786 39976
rect 84102 39924 84108 39976
rect 84160 39964 84166 39976
rect 84212 39973 84240 40004
rect 84565 40001 84577 40004
rect 84611 40032 84623 40035
rect 84930 40032 84936 40044
rect 84611 40004 84936 40032
rect 84611 40001 84623 40004
rect 84565 39995 84623 40001
rect 84930 39992 84936 40004
rect 84988 39992 84994 40044
rect 85206 40032 85212 40044
rect 85167 40004 85212 40032
rect 85206 39992 85212 40004
rect 85264 40032 85270 40044
rect 85264 40004 85436 40032
rect 85264 39992 85270 40004
rect 85408 39973 85436 40004
rect 84197 39967 84255 39973
rect 84197 39964 84209 39967
rect 84160 39936 84209 39964
rect 84160 39924 84166 39936
rect 84197 39933 84209 39936
rect 84243 39933 84255 39967
rect 85393 39967 85451 39973
rect 84197 39927 84255 39933
rect 84304 39936 85344 39964
rect 81434 39896 81440 39908
rect 80440 39868 81440 39896
rect 81434 39856 81440 39868
rect 81492 39856 81498 39908
rect 82553 39899 82611 39905
rect 82553 39865 82565 39899
rect 82599 39896 82611 39899
rect 84304 39896 84332 39936
rect 82599 39868 84332 39896
rect 85316 39896 85344 39936
rect 85393 39933 85405 39967
rect 85439 39933 85451 39967
rect 85500 39964 85528 40072
rect 85669 40069 85681 40103
rect 85715 40100 85727 40103
rect 86218 40100 86224 40112
rect 85715 40072 86224 40100
rect 85715 40069 85727 40072
rect 85669 40063 85727 40069
rect 86218 40060 86224 40072
rect 86276 40060 86282 40112
rect 85758 39992 85764 40044
rect 85816 40032 85822 40044
rect 88426 40032 88432 40044
rect 85816 40004 88432 40032
rect 85816 39992 85822 40004
rect 88426 39992 88432 40004
rect 88484 40032 88490 40044
rect 88613 40035 88671 40041
rect 88613 40032 88625 40035
rect 88484 40004 88625 40032
rect 88484 39992 88490 40004
rect 88613 40001 88625 40004
rect 88659 40001 88671 40035
rect 88613 39995 88671 40001
rect 88978 39992 88984 40044
rect 89036 40032 89042 40044
rect 90729 40035 90787 40041
rect 90729 40032 90741 40035
rect 89036 40004 90741 40032
rect 89036 39992 89042 40004
rect 90729 40001 90741 40004
rect 90775 40032 90787 40035
rect 91005 40035 91063 40041
rect 91005 40032 91017 40035
rect 90775 40004 91017 40032
rect 90775 40001 90787 40004
rect 90729 39995 90787 40001
rect 91005 40001 91017 40004
rect 91051 40001 91063 40035
rect 91005 39995 91063 40001
rect 85942 39964 85948 39976
rect 85500 39936 85948 39964
rect 85393 39927 85451 39933
rect 85942 39924 85948 39936
rect 86000 39924 86006 39976
rect 86221 39967 86279 39973
rect 86221 39933 86233 39967
rect 86267 39964 86279 39967
rect 86494 39964 86500 39976
rect 86267 39936 86500 39964
rect 86267 39933 86279 39936
rect 86221 39927 86279 39933
rect 86236 39896 86264 39927
rect 86494 39924 86500 39936
rect 86552 39924 86558 39976
rect 88518 39964 88524 39976
rect 88479 39936 88524 39964
rect 88518 39924 88524 39936
rect 88576 39924 88582 39976
rect 91094 39924 91100 39976
rect 91152 39964 91158 39976
rect 91281 39967 91339 39973
rect 91281 39964 91293 39967
rect 91152 39936 91293 39964
rect 91152 39924 91158 39936
rect 91281 39933 91293 39936
rect 91327 39933 91339 39967
rect 91281 39927 91339 39933
rect 85316 39868 86264 39896
rect 82599 39865 82611 39868
rect 82553 39859 82611 39865
rect 77386 39828 77392 39840
rect 74184 39800 77392 39828
rect 77386 39788 77392 39800
rect 77444 39788 77450 39840
rect 77570 39828 77576 39840
rect 77531 39800 77576 39828
rect 77570 39788 77576 39800
rect 77628 39828 77634 39840
rect 79229 39831 79287 39837
rect 79229 39828 79241 39831
rect 77628 39800 79241 39828
rect 77628 39788 77634 39800
rect 79229 39797 79241 39800
rect 79275 39828 79287 39831
rect 80790 39828 80796 39840
rect 79275 39800 80796 39828
rect 79275 39797 79287 39800
rect 79229 39791 79287 39797
rect 80790 39788 80796 39800
rect 80848 39788 80854 39840
rect 80882 39788 80888 39840
rect 80940 39828 80946 39840
rect 81069 39831 81127 39837
rect 81069 39828 81081 39831
rect 80940 39800 81081 39828
rect 80940 39788 80946 39800
rect 81069 39797 81081 39800
rect 81115 39797 81127 39831
rect 84120 39828 84148 39868
rect 84194 39828 84200 39840
rect 84120 39800 84200 39828
rect 81069 39791 81127 39797
rect 84194 39788 84200 39800
rect 84252 39788 84258 39840
rect 84381 39831 84439 39837
rect 84381 39797 84393 39831
rect 84427 39828 84439 39831
rect 84562 39828 84568 39840
rect 84427 39800 84568 39828
rect 84427 39797 84439 39800
rect 84381 39791 84439 39797
rect 84562 39788 84568 39800
rect 84620 39788 84626 39840
rect 85942 39788 85948 39840
rect 86000 39828 86006 39840
rect 86589 39831 86647 39837
rect 86589 39828 86601 39831
rect 86000 39800 86601 39828
rect 86000 39788 86006 39800
rect 86589 39797 86601 39800
rect 86635 39828 86647 39831
rect 86678 39828 86684 39840
rect 86635 39800 86684 39828
rect 86635 39797 86647 39800
rect 86589 39791 86647 39797
rect 86678 39788 86684 39800
rect 86736 39788 86742 39840
rect 86862 39788 86868 39840
rect 86920 39828 86926 39840
rect 92385 39831 92443 39837
rect 92385 39828 92397 39831
rect 86920 39800 92397 39828
rect 86920 39788 86926 39800
rect 92385 39797 92397 39800
rect 92431 39797 92443 39831
rect 92385 39791 92443 39797
rect 1104 39738 105616 39760
rect 1104 39686 19606 39738
rect 19658 39686 19670 39738
rect 19722 39686 19734 39738
rect 19786 39686 19798 39738
rect 19850 39686 50326 39738
rect 50378 39686 50390 39738
rect 50442 39686 50454 39738
rect 50506 39686 50518 39738
rect 50570 39686 81046 39738
rect 81098 39686 81110 39738
rect 81162 39686 81174 39738
rect 81226 39686 81238 39738
rect 81290 39686 105616 39738
rect 1104 39664 105616 39686
rect 2774 39584 2780 39636
rect 2832 39624 2838 39636
rect 4157 39627 4215 39633
rect 4157 39624 4169 39627
rect 2832 39596 4169 39624
rect 2832 39584 2838 39596
rect 4157 39593 4169 39596
rect 4203 39593 4215 39627
rect 15473 39627 15531 39633
rect 4157 39587 4215 39593
rect 4264 39596 15424 39624
rect 3329 39559 3387 39565
rect 3329 39525 3341 39559
rect 3375 39556 3387 39559
rect 3694 39556 3700 39568
rect 3375 39528 3700 39556
rect 3375 39525 3387 39528
rect 3329 39519 3387 39525
rect 2593 39491 2651 39497
rect 2593 39457 2605 39491
rect 2639 39457 2651 39491
rect 2593 39451 2651 39457
rect 2961 39491 3019 39497
rect 2961 39457 2973 39491
rect 3007 39488 3019 39491
rect 3344 39488 3372 39519
rect 3694 39516 3700 39528
rect 3752 39516 3758 39568
rect 3970 39516 3976 39568
rect 4028 39556 4034 39568
rect 4264 39556 4292 39596
rect 4798 39556 4804 39568
rect 4028 39528 4292 39556
rect 4356 39528 4804 39556
rect 4028 39516 4034 39528
rect 4356 39497 4384 39528
rect 4798 39516 4804 39528
rect 4856 39516 4862 39568
rect 4982 39556 4988 39568
rect 4943 39528 4988 39556
rect 4982 39516 4988 39528
rect 5040 39516 5046 39568
rect 8202 39556 8208 39568
rect 7300 39528 8208 39556
rect 3007 39460 3372 39488
rect 4341 39491 4399 39497
rect 3007 39457 3019 39460
rect 2961 39451 3019 39457
rect 4341 39457 4353 39491
rect 4387 39457 4399 39491
rect 4341 39451 4399 39457
rect 4525 39491 4583 39497
rect 4525 39457 4537 39491
rect 4571 39488 4583 39491
rect 5000 39488 5028 39516
rect 7300 39497 7328 39528
rect 8202 39516 8208 39528
rect 8260 39516 8266 39568
rect 8294 39516 8300 39568
rect 8352 39556 8358 39568
rect 15396 39556 15424 39596
rect 15473 39593 15485 39627
rect 15519 39624 15531 39627
rect 16482 39624 16488 39636
rect 15519 39596 16488 39624
rect 15519 39593 15531 39596
rect 15473 39587 15531 39593
rect 16482 39584 16488 39596
rect 16540 39584 16546 39636
rect 19705 39627 19763 39633
rect 19705 39593 19717 39627
rect 19751 39624 19763 39627
rect 20165 39627 20223 39633
rect 20165 39624 20177 39627
rect 19751 39596 20177 39624
rect 19751 39593 19763 39596
rect 19705 39587 19763 39593
rect 20165 39593 20177 39596
rect 20211 39624 20223 39627
rect 21542 39624 21548 39636
rect 20211 39596 21548 39624
rect 20211 39593 20223 39596
rect 20165 39587 20223 39593
rect 21542 39584 21548 39596
rect 21600 39584 21606 39636
rect 24118 39584 24124 39636
rect 24176 39624 24182 39636
rect 31941 39627 31999 39633
rect 31941 39624 31953 39627
rect 24176 39596 31953 39624
rect 24176 39584 24182 39596
rect 31941 39593 31953 39596
rect 31987 39593 31999 39627
rect 31941 39587 31999 39593
rect 32214 39584 32220 39636
rect 32272 39624 32278 39636
rect 33962 39624 33968 39636
rect 32272 39596 33968 39624
rect 32272 39584 32278 39596
rect 33962 39584 33968 39596
rect 34020 39584 34026 39636
rect 43622 39624 43628 39636
rect 34072 39596 43628 39624
rect 20990 39556 20996 39568
rect 8352 39528 15240 39556
rect 15396 39528 20996 39556
rect 8352 39516 8358 39528
rect 4571 39460 5028 39488
rect 7285 39491 7343 39497
rect 4571 39457 4583 39460
rect 4525 39451 4583 39457
rect 7285 39457 7297 39491
rect 7331 39457 7343 39491
rect 7285 39451 7343 39457
rect 2608 39420 2636 39451
rect 7466 39448 7472 39500
rect 7524 39488 7530 39500
rect 7607 39491 7665 39497
rect 7607 39488 7619 39491
rect 7524 39460 7619 39488
rect 7524 39448 7530 39460
rect 7607 39457 7619 39460
rect 7653 39457 7665 39491
rect 7607 39451 7665 39457
rect 7834 39448 7840 39500
rect 7892 39488 7898 39500
rect 9674 39488 9680 39500
rect 7892 39460 7937 39488
rect 9635 39460 9680 39488
rect 7892 39448 7898 39460
rect 9674 39448 9680 39460
rect 9732 39488 9738 39500
rect 9953 39491 10011 39497
rect 9953 39488 9965 39491
rect 9732 39460 9965 39488
rect 9732 39448 9738 39460
rect 9953 39457 9965 39460
rect 9999 39457 10011 39491
rect 11790 39488 11796 39500
rect 9953 39451 10011 39457
rect 11716 39460 11796 39488
rect 3145 39423 3203 39429
rect 2608 39392 2728 39420
rect 2700 39284 2728 39392
rect 3145 39389 3157 39423
rect 3191 39420 3203 39423
rect 4614 39420 4620 39432
rect 3191 39392 4620 39420
rect 3191 39389 3203 39392
rect 3145 39383 3203 39389
rect 4614 39380 4620 39392
rect 4672 39380 4678 39432
rect 5718 39380 5724 39432
rect 5776 39420 5782 39432
rect 6641 39423 6699 39429
rect 6641 39420 6653 39423
rect 5776 39392 6653 39420
rect 5776 39380 5782 39392
rect 6641 39389 6653 39392
rect 6687 39389 6699 39423
rect 7374 39420 7380 39432
rect 7335 39392 7380 39420
rect 6641 39383 6699 39389
rect 7374 39380 7380 39392
rect 7432 39380 7438 39432
rect 11716 39420 11744 39460
rect 11790 39448 11796 39460
rect 11848 39448 11854 39500
rect 13078 39448 13084 39500
rect 13136 39488 13142 39500
rect 13538 39488 13544 39500
rect 13136 39460 13544 39488
rect 13136 39448 13142 39460
rect 13538 39448 13544 39460
rect 13596 39488 13602 39500
rect 13633 39491 13691 39497
rect 13633 39488 13645 39491
rect 13596 39460 13645 39488
rect 13596 39448 13602 39460
rect 13633 39457 13645 39460
rect 13679 39457 13691 39491
rect 13814 39488 13820 39500
rect 13727 39460 13820 39488
rect 13633 39451 13691 39457
rect 13814 39448 13820 39460
rect 13872 39488 13878 39500
rect 14458 39488 14464 39500
rect 13872 39460 14464 39488
rect 13872 39448 13878 39460
rect 14458 39448 14464 39460
rect 14516 39448 14522 39500
rect 12161 39423 12219 39429
rect 12161 39420 12173 39423
rect 11716 39392 12173 39420
rect 12161 39389 12173 39392
rect 12207 39389 12219 39423
rect 12161 39383 12219 39389
rect 12710 39380 12716 39432
rect 12768 39420 12774 39432
rect 12897 39423 12955 39429
rect 12897 39420 12909 39423
rect 12768 39392 12909 39420
rect 12768 39380 12774 39392
rect 12897 39389 12909 39392
rect 12943 39389 12955 39423
rect 15212 39420 15240 39528
rect 20990 39516 20996 39528
rect 21048 39516 21054 39568
rect 25406 39516 25412 39568
rect 25464 39556 25470 39568
rect 25958 39556 25964 39568
rect 25464 39528 25964 39556
rect 25464 39516 25470 39528
rect 25958 39516 25964 39528
rect 26016 39516 26022 39568
rect 31570 39556 31576 39568
rect 26068 39528 31576 39556
rect 15289 39491 15347 39497
rect 15289 39457 15301 39491
rect 15335 39488 15347 39491
rect 15562 39488 15568 39500
rect 15335 39460 15568 39488
rect 15335 39457 15347 39460
rect 15289 39451 15347 39457
rect 15562 39448 15568 39460
rect 15620 39448 15626 39500
rect 19705 39491 19763 39497
rect 19705 39457 19717 39491
rect 19751 39488 19763 39491
rect 19797 39491 19855 39497
rect 19797 39488 19809 39491
rect 19751 39460 19809 39488
rect 19751 39457 19763 39460
rect 19705 39451 19763 39457
rect 19797 39457 19809 39460
rect 19843 39457 19855 39491
rect 19797 39451 19855 39457
rect 20714 39448 20720 39500
rect 20772 39488 20778 39500
rect 20901 39491 20959 39497
rect 20901 39488 20913 39491
rect 20772 39460 20913 39488
rect 20772 39448 20778 39460
rect 20901 39457 20913 39460
rect 20947 39457 20959 39491
rect 20901 39451 20959 39457
rect 25590 39448 25596 39500
rect 25648 39488 25654 39500
rect 26068 39488 26096 39528
rect 31570 39516 31576 39528
rect 31628 39516 31634 39568
rect 31754 39516 31760 39568
rect 31812 39556 31818 39568
rect 34072 39556 34100 39596
rect 43622 39584 43628 39596
rect 43680 39584 43686 39636
rect 43717 39627 43775 39633
rect 43717 39593 43729 39627
rect 43763 39624 43775 39627
rect 49050 39624 49056 39636
rect 43763 39596 49056 39624
rect 43763 39593 43775 39596
rect 43717 39587 43775 39593
rect 49050 39584 49056 39596
rect 49108 39584 49114 39636
rect 49786 39624 49792 39636
rect 49160 39596 49792 39624
rect 46106 39556 46112 39568
rect 31812 39528 34100 39556
rect 38120 39528 46112 39556
rect 31812 39516 31818 39528
rect 25648 39460 26096 39488
rect 27525 39491 27583 39497
rect 25648 39448 25654 39460
rect 27525 39457 27537 39491
rect 27571 39488 27583 39491
rect 27614 39488 27620 39500
rect 27571 39460 27620 39488
rect 27571 39457 27583 39460
rect 27525 39451 27583 39457
rect 27614 39448 27620 39460
rect 27672 39448 27678 39500
rect 32306 39488 32312 39500
rect 32267 39460 32312 39488
rect 32306 39448 32312 39460
rect 32364 39448 32370 39500
rect 32766 39448 32772 39500
rect 32824 39488 32830 39500
rect 32861 39491 32919 39497
rect 32861 39488 32873 39491
rect 32824 39460 32873 39488
rect 32824 39448 32830 39460
rect 32861 39457 32873 39460
rect 32907 39457 32919 39491
rect 33042 39488 33048 39500
rect 33003 39460 33048 39488
rect 32861 39451 32919 39457
rect 33042 39448 33048 39460
rect 33100 39448 33106 39500
rect 34330 39488 34336 39500
rect 34291 39460 34336 39488
rect 34330 39448 34336 39460
rect 34388 39448 34394 39500
rect 35069 39491 35127 39497
rect 34440 39460 34836 39488
rect 27706 39420 27712 39432
rect 15212 39392 27712 39420
rect 12897 39383 12955 39389
rect 27706 39380 27712 39392
rect 27764 39380 27770 39432
rect 27798 39380 27804 39432
rect 27856 39420 27862 39432
rect 31754 39420 31760 39432
rect 27856 39392 31760 39420
rect 27856 39380 27862 39392
rect 31754 39380 31760 39392
rect 31812 39380 31818 39432
rect 31849 39423 31907 39429
rect 31849 39389 31861 39423
rect 31895 39420 31907 39423
rect 31941 39423 31999 39429
rect 31941 39420 31953 39423
rect 31895 39392 31953 39420
rect 31895 39389 31907 39392
rect 31849 39383 31907 39389
rect 31941 39389 31953 39392
rect 31987 39420 31999 39423
rect 32125 39423 32183 39429
rect 32125 39420 32137 39423
rect 31987 39392 32137 39420
rect 31987 39389 31999 39392
rect 31941 39383 31999 39389
rect 32125 39389 32137 39392
rect 32171 39389 32183 39423
rect 32125 39383 32183 39389
rect 33502 39380 33508 39432
rect 33560 39420 33566 39432
rect 33689 39423 33747 39429
rect 33689 39420 33701 39423
rect 33560 39392 33701 39420
rect 33560 39380 33566 39392
rect 33689 39389 33701 39392
rect 33735 39420 33747 39423
rect 34440 39420 34468 39460
rect 33735 39392 34468 39420
rect 33735 39389 33747 39392
rect 33689 39383 33747 39389
rect 34514 39380 34520 39432
rect 34572 39420 34578 39432
rect 34701 39423 34759 39429
rect 34701 39420 34713 39423
rect 34572 39392 34713 39420
rect 34572 39380 34578 39392
rect 34701 39389 34713 39392
rect 34747 39389 34759 39423
rect 34808 39420 34836 39460
rect 35069 39457 35081 39491
rect 35115 39488 35127 39491
rect 38120 39488 38148 39528
rect 46106 39516 46112 39528
rect 46164 39516 46170 39568
rect 48317 39559 48375 39565
rect 48317 39556 48329 39559
rect 46308 39528 48329 39556
rect 35115 39460 38148 39488
rect 35115 39457 35127 39460
rect 35069 39451 35127 39457
rect 39114 39448 39120 39500
rect 39172 39488 39178 39500
rect 39393 39491 39451 39497
rect 39393 39488 39405 39491
rect 39172 39460 39405 39488
rect 39172 39448 39178 39460
rect 39393 39457 39405 39460
rect 39439 39457 39451 39491
rect 39393 39451 39451 39457
rect 39482 39448 39488 39500
rect 39540 39488 39546 39500
rect 39850 39488 39856 39500
rect 39540 39460 39585 39488
rect 39811 39460 39856 39488
rect 39540 39448 39546 39460
rect 39850 39448 39856 39460
rect 39908 39448 39914 39500
rect 39942 39448 39948 39500
rect 40000 39488 40006 39500
rect 40773 39491 40831 39497
rect 40773 39488 40785 39491
rect 40000 39460 40785 39488
rect 40000 39448 40006 39460
rect 40773 39457 40785 39460
rect 40819 39488 40831 39491
rect 43717 39491 43775 39497
rect 43717 39488 43729 39491
rect 40819 39460 43729 39488
rect 40819 39457 40831 39460
rect 40773 39451 40831 39457
rect 43717 39457 43729 39460
rect 43763 39457 43775 39491
rect 43717 39451 43775 39457
rect 43898 39448 43904 39500
rect 43956 39488 43962 39500
rect 44177 39491 44235 39497
rect 44177 39488 44189 39491
rect 43956 39460 44189 39488
rect 43956 39448 43962 39460
rect 44177 39457 44189 39460
rect 44223 39457 44235 39491
rect 44358 39488 44364 39500
rect 44319 39460 44364 39488
rect 44177 39451 44235 39457
rect 39574 39420 39580 39432
rect 34808 39392 39580 39420
rect 34701 39383 34759 39389
rect 39574 39380 39580 39392
rect 39632 39380 39638 39432
rect 40862 39380 40868 39432
rect 40920 39420 40926 39432
rect 40957 39423 41015 39429
rect 40957 39420 40969 39423
rect 40920 39392 40969 39420
rect 40920 39380 40926 39392
rect 40957 39389 40969 39392
rect 41003 39420 41015 39423
rect 42794 39420 42800 39432
rect 41003 39392 42800 39420
rect 41003 39389 41015 39392
rect 40957 39383 41015 39389
rect 42794 39380 42800 39392
rect 42852 39380 42858 39432
rect 44192 39420 44220 39451
rect 44358 39448 44364 39460
rect 44416 39448 44422 39500
rect 44821 39491 44879 39497
rect 44821 39488 44833 39491
rect 44468 39460 44833 39488
rect 44468 39420 44496 39460
rect 44821 39457 44833 39460
rect 44867 39457 44879 39491
rect 44821 39451 44879 39457
rect 44910 39448 44916 39500
rect 44968 39488 44974 39500
rect 46308 39488 46336 39528
rect 48317 39525 48329 39528
rect 48363 39525 48375 39559
rect 48317 39519 48375 39525
rect 48590 39516 48596 39568
rect 48648 39556 48654 39568
rect 48685 39559 48743 39565
rect 48685 39556 48697 39559
rect 48648 39528 48697 39556
rect 48648 39516 48654 39528
rect 48685 39525 48697 39528
rect 48731 39556 48743 39559
rect 48774 39556 48780 39568
rect 48731 39528 48780 39556
rect 48731 39525 48743 39528
rect 48685 39519 48743 39525
rect 48774 39516 48780 39528
rect 48832 39516 48838 39568
rect 48866 39516 48872 39568
rect 48924 39556 48930 39568
rect 49160 39556 49188 39596
rect 49786 39584 49792 39596
rect 49844 39584 49850 39636
rect 50154 39624 50160 39636
rect 50115 39596 50160 39624
rect 50154 39584 50160 39596
rect 50212 39584 50218 39636
rect 50706 39624 50712 39636
rect 50667 39596 50712 39624
rect 50706 39584 50712 39596
rect 50764 39584 50770 39636
rect 50798 39584 50804 39636
rect 50856 39624 50862 39636
rect 51353 39627 51411 39633
rect 51353 39624 51365 39627
rect 50856 39596 51365 39624
rect 50856 39584 50862 39596
rect 51353 39593 51365 39596
rect 51399 39624 51411 39627
rect 51534 39624 51540 39636
rect 51399 39596 51540 39624
rect 51399 39593 51411 39596
rect 51353 39587 51411 39593
rect 51534 39584 51540 39596
rect 51592 39584 51598 39636
rect 53650 39584 53656 39636
rect 53708 39624 53714 39636
rect 53708 39596 70992 39624
rect 53708 39584 53714 39596
rect 48924 39528 49188 39556
rect 48924 39516 48930 39528
rect 49160 39497 49188 39528
rect 49418 39516 49424 39568
rect 49476 39556 49482 39568
rect 50430 39556 50436 39568
rect 49476 39528 50436 39556
rect 49476 39516 49482 39528
rect 44968 39460 45013 39488
rect 45296 39460 46336 39488
rect 46385 39491 46443 39497
rect 44968 39448 44974 39460
rect 44192 39392 44496 39420
rect 6362 39352 6368 39364
rect 6275 39324 6368 39352
rect 6362 39312 6368 39324
rect 6420 39352 6426 39364
rect 7392 39352 7420 39380
rect 6420 39324 7420 39352
rect 6420 39312 6426 39324
rect 7742 39312 7748 39364
rect 7800 39352 7806 39364
rect 45296 39352 45324 39460
rect 46385 39457 46397 39491
rect 46431 39488 46443 39491
rect 49145 39491 49203 39497
rect 46431 39460 49096 39488
rect 46431 39457 46443 39460
rect 46385 39451 46443 39457
rect 45830 39380 45836 39432
rect 45888 39420 45894 39432
rect 46532 39423 46590 39429
rect 46532 39420 46544 39423
rect 45888 39392 46544 39420
rect 45888 39380 45894 39392
rect 46532 39389 46544 39392
rect 46578 39389 46590 39423
rect 46750 39420 46756 39432
rect 46711 39392 46756 39420
rect 46532 39383 46590 39389
rect 46750 39380 46756 39392
rect 46808 39380 46814 39432
rect 48317 39423 48375 39429
rect 48317 39389 48329 39423
rect 48363 39420 48375 39423
rect 48501 39423 48559 39429
rect 48501 39420 48513 39423
rect 48363 39392 48513 39420
rect 48363 39389 48375 39392
rect 48317 39383 48375 39389
rect 48501 39389 48513 39392
rect 48547 39420 48559 39423
rect 48958 39420 48964 39432
rect 48547 39392 48964 39420
rect 48547 39389 48559 39392
rect 48501 39383 48559 39389
rect 48958 39380 48964 39392
rect 49016 39380 49022 39432
rect 7800 39324 45324 39352
rect 45373 39355 45431 39361
rect 7800 39312 7806 39324
rect 45373 39321 45385 39355
rect 45419 39352 45431 39355
rect 46661 39355 46719 39361
rect 46661 39352 46673 39355
rect 45419 39324 46673 39352
rect 45419 39321 45431 39324
rect 45373 39315 45431 39321
rect 46661 39321 46673 39324
rect 46707 39321 46719 39355
rect 49068 39352 49096 39460
rect 49145 39457 49157 39491
rect 49191 39457 49203 39491
rect 49145 39451 49203 39457
rect 49326 39448 49332 39500
rect 49384 39488 49390 39500
rect 49712 39497 49740 39528
rect 50430 39516 50436 39528
rect 50488 39516 50494 39568
rect 54662 39556 54668 39568
rect 54623 39528 54668 39556
rect 54662 39516 54668 39528
rect 54720 39516 54726 39568
rect 56413 39559 56471 39565
rect 56413 39525 56425 39559
rect 56459 39556 56471 39559
rect 57790 39556 57796 39568
rect 56459 39528 57796 39556
rect 56459 39525 56471 39528
rect 56413 39519 56471 39525
rect 57790 39516 57796 39528
rect 57848 39516 57854 39568
rect 59078 39556 59084 39568
rect 58636 39528 59084 39556
rect 49605 39491 49663 39497
rect 49605 39488 49617 39491
rect 49384 39460 49617 39488
rect 49384 39448 49390 39460
rect 49605 39457 49617 39460
rect 49651 39457 49663 39491
rect 49605 39451 49663 39457
rect 49697 39491 49755 39497
rect 49697 39457 49709 39491
rect 49743 39457 49755 39491
rect 49697 39451 49755 39457
rect 49786 39448 49792 39500
rect 49844 39488 49850 39500
rect 50706 39488 50712 39500
rect 49844 39460 50712 39488
rect 49844 39448 49850 39460
rect 50706 39448 50712 39460
rect 50764 39448 50770 39500
rect 51537 39491 51595 39497
rect 51537 39457 51549 39491
rect 51583 39488 51595 39491
rect 51813 39491 51871 39497
rect 51813 39488 51825 39491
rect 51583 39460 51825 39488
rect 51583 39457 51595 39460
rect 51537 39451 51595 39457
rect 51813 39457 51825 39460
rect 51859 39488 51871 39491
rect 51859 39460 52040 39488
rect 51859 39457 51871 39460
rect 51813 39451 51871 39457
rect 50430 39380 50436 39432
rect 50488 39420 50494 39432
rect 50525 39423 50583 39429
rect 50525 39420 50537 39423
rect 50488 39392 50537 39420
rect 50488 39380 50494 39392
rect 50525 39389 50537 39392
rect 50571 39420 50583 39423
rect 51626 39420 51632 39432
rect 50571 39392 51632 39420
rect 50571 39389 50583 39392
rect 50525 39383 50583 39389
rect 51626 39380 51632 39392
rect 51684 39380 51690 39432
rect 51902 39420 51908 39432
rect 51863 39392 51908 39420
rect 51902 39380 51908 39392
rect 51960 39380 51966 39432
rect 52012 39420 52040 39460
rect 52086 39448 52092 39500
rect 52144 39488 52150 39500
rect 52144 39460 52189 39488
rect 52144 39448 52150 39460
rect 52638 39448 52644 39500
rect 52696 39488 52702 39500
rect 52696 39460 52741 39488
rect 52696 39448 52702 39460
rect 52822 39448 52828 39500
rect 52880 39488 52886 39500
rect 52880 39460 52925 39488
rect 52880 39448 52886 39460
rect 54294 39448 54300 39500
rect 54352 39488 54358 39500
rect 55033 39491 55091 39497
rect 55033 39488 55045 39491
rect 54352 39460 55045 39488
rect 54352 39448 54358 39460
rect 55033 39457 55045 39460
rect 55079 39457 55091 39491
rect 58066 39488 58072 39500
rect 58027 39460 58072 39488
rect 55033 39451 55091 39457
rect 58066 39448 58072 39460
rect 58124 39448 58130 39500
rect 58158 39448 58164 39500
rect 58216 39488 58222 39500
rect 58636 39497 58664 39528
rect 59078 39516 59084 39528
rect 59136 39516 59142 39568
rect 59170 39516 59176 39568
rect 59228 39556 59234 39568
rect 59541 39559 59599 39565
rect 59541 39556 59553 39559
rect 59228 39528 59553 39556
rect 59228 39516 59234 39528
rect 59541 39525 59553 39528
rect 59587 39525 59599 39559
rect 65702 39556 65708 39568
rect 59541 39519 59599 39525
rect 61028 39528 65708 39556
rect 58529 39491 58587 39497
rect 58529 39488 58541 39491
rect 58216 39460 58541 39488
rect 58216 39448 58222 39460
rect 58529 39457 58541 39460
rect 58575 39457 58587 39491
rect 58529 39451 58587 39457
rect 58621 39491 58679 39497
rect 58621 39457 58633 39491
rect 58667 39457 58679 39491
rect 60185 39491 60243 39497
rect 60185 39488 60197 39491
rect 58621 39451 58679 39457
rect 59004 39460 60197 39488
rect 52178 39420 52184 39432
rect 52012 39392 52184 39420
rect 52178 39380 52184 39392
rect 52236 39380 52242 39432
rect 54662 39380 54668 39432
rect 54720 39420 54726 39432
rect 54757 39423 54815 39429
rect 54757 39420 54769 39423
rect 54720 39392 54769 39420
rect 54720 39380 54726 39392
rect 54757 39389 54769 39392
rect 54803 39389 54815 39423
rect 57974 39420 57980 39432
rect 57935 39392 57980 39420
rect 54757 39383 54815 39389
rect 57974 39380 57980 39392
rect 58032 39380 58038 39432
rect 49878 39352 49884 39364
rect 46661 39315 46719 39321
rect 46768 39324 49004 39352
rect 49068 39324 49884 39352
rect 4798 39284 4804 39296
rect 2700 39256 4804 39284
rect 4798 39244 4804 39256
rect 4856 39244 4862 39296
rect 6546 39284 6552 39296
rect 6459 39256 6552 39284
rect 6546 39244 6552 39256
rect 6604 39284 6610 39296
rect 7834 39284 7840 39296
rect 6604 39256 7840 39284
rect 6604 39244 6610 39256
rect 7834 39244 7840 39256
rect 7892 39244 7898 39296
rect 8294 39244 8300 39296
rect 8352 39284 8358 39296
rect 9769 39287 9827 39293
rect 9769 39284 9781 39287
rect 8352 39256 9781 39284
rect 8352 39244 8358 39256
rect 9769 39253 9781 39256
rect 9815 39253 9827 39287
rect 11974 39284 11980 39296
rect 11935 39256 11980 39284
rect 9769 39247 9827 39253
rect 11974 39244 11980 39256
rect 12032 39244 12038 39296
rect 12710 39284 12716 39296
rect 12671 39256 12716 39284
rect 12710 39244 12716 39256
rect 12768 39244 12774 39296
rect 14090 39284 14096 39296
rect 14051 39256 14096 39284
rect 14090 39244 14096 39256
rect 14148 39244 14154 39296
rect 14458 39284 14464 39296
rect 14419 39256 14464 39284
rect 14458 39244 14464 39256
rect 14516 39244 14522 39296
rect 19886 39284 19892 39296
rect 19847 39256 19892 39284
rect 19886 39244 19892 39256
rect 19944 39244 19950 39296
rect 20806 39244 20812 39296
rect 20864 39284 20870 39296
rect 20993 39287 21051 39293
rect 20993 39284 21005 39287
rect 20864 39256 21005 39284
rect 20864 39244 20870 39256
rect 20993 39253 21005 39256
rect 21039 39253 21051 39287
rect 27798 39284 27804 39296
rect 27759 39256 27804 39284
rect 20993 39247 21051 39253
rect 27798 39244 27804 39256
rect 27856 39244 27862 39296
rect 27982 39244 27988 39296
rect 28040 39284 28046 39296
rect 31665 39287 31723 39293
rect 31665 39284 31677 39287
rect 28040 39256 31677 39284
rect 28040 39244 28046 39256
rect 31665 39253 31677 39256
rect 31711 39284 31723 39287
rect 33042 39284 33048 39296
rect 31711 39256 33048 39284
rect 31711 39253 31723 39256
rect 31665 39247 31723 39253
rect 33042 39244 33048 39256
rect 33100 39244 33106 39296
rect 33226 39244 33232 39296
rect 33284 39284 33290 39296
rect 33321 39287 33379 39293
rect 33321 39284 33333 39287
rect 33284 39256 33333 39284
rect 33284 39244 33290 39256
rect 33321 39253 33333 39256
rect 33367 39253 33379 39287
rect 33870 39284 33876 39296
rect 33831 39256 33876 39284
rect 33321 39247 33379 39253
rect 33870 39244 33876 39256
rect 33928 39244 33934 39296
rect 33962 39244 33968 39296
rect 34020 39284 34026 39296
rect 34471 39287 34529 39293
rect 34471 39284 34483 39287
rect 34020 39256 34483 39284
rect 34020 39244 34026 39256
rect 34471 39253 34483 39256
rect 34517 39253 34529 39287
rect 34606 39284 34612 39296
rect 34567 39256 34612 39284
rect 34471 39247 34529 39253
rect 34606 39244 34612 39256
rect 34664 39244 34670 39296
rect 34790 39244 34796 39296
rect 34848 39284 34854 39296
rect 40310 39284 40316 39296
rect 34848 39256 40316 39284
rect 34848 39244 34854 39256
rect 40310 39244 40316 39256
rect 40368 39244 40374 39296
rect 40405 39287 40463 39293
rect 40405 39253 40417 39287
rect 40451 39284 40463 39287
rect 40678 39284 40684 39296
rect 40451 39256 40684 39284
rect 40451 39253 40463 39256
rect 40405 39247 40463 39253
rect 40678 39244 40684 39256
rect 40736 39244 40742 39296
rect 40954 39244 40960 39296
rect 41012 39284 41018 39296
rect 42702 39284 42708 39296
rect 41012 39256 42708 39284
rect 41012 39244 41018 39256
rect 42702 39244 42708 39256
rect 42760 39244 42766 39296
rect 43438 39244 43444 39296
rect 43496 39284 43502 39296
rect 43809 39287 43867 39293
rect 43809 39284 43821 39287
rect 43496 39256 43821 39284
rect 43496 39244 43502 39256
rect 43809 39253 43821 39256
rect 43855 39284 43867 39287
rect 43898 39284 43904 39296
rect 43855 39256 43904 39284
rect 43855 39253 43867 39256
rect 43809 39247 43867 39253
rect 43898 39244 43904 39256
rect 43956 39284 43962 39296
rect 43993 39287 44051 39293
rect 43993 39284 44005 39287
rect 43956 39256 44005 39284
rect 43956 39244 43962 39256
rect 43993 39253 44005 39256
rect 44039 39253 44051 39287
rect 43993 39247 44051 39253
rect 44082 39244 44088 39296
rect 44140 39284 44146 39296
rect 44358 39284 44364 39296
rect 44140 39256 44364 39284
rect 44140 39244 44146 39256
rect 44358 39244 44364 39256
rect 44416 39284 44422 39296
rect 44910 39284 44916 39296
rect 44416 39256 44916 39284
rect 44416 39244 44422 39256
rect 44910 39244 44916 39256
rect 44968 39244 44974 39296
rect 45741 39287 45799 39293
rect 45741 39253 45753 39287
rect 45787 39284 45799 39287
rect 45922 39284 45928 39296
rect 45787 39256 45928 39284
rect 45787 39253 45799 39256
rect 45741 39247 45799 39253
rect 45922 39244 45928 39256
rect 45980 39244 45986 39296
rect 46198 39244 46204 39296
rect 46256 39284 46262 39296
rect 46768 39284 46796 39324
rect 47026 39284 47032 39296
rect 46256 39256 46796 39284
rect 46987 39256 47032 39284
rect 46256 39244 46262 39256
rect 47026 39244 47032 39256
rect 47084 39244 47090 39296
rect 48976 39284 49004 39324
rect 49878 39312 49884 39324
rect 49936 39312 49942 39364
rect 53009 39355 53067 39361
rect 53009 39352 53021 39355
rect 49988 39324 53021 39352
rect 49988 39284 50016 39324
rect 53009 39321 53021 39324
rect 53055 39321 53067 39355
rect 53009 39315 53067 39321
rect 53558 39312 53564 39364
rect 53616 39352 53622 39364
rect 53653 39355 53711 39361
rect 53653 39352 53665 39355
rect 53616 39324 53665 39352
rect 53616 39312 53622 39324
rect 53653 39321 53665 39324
rect 53699 39352 53711 39355
rect 53699 39324 54708 39352
rect 53699 39321 53711 39324
rect 53653 39315 53711 39321
rect 54680 39296 54708 39324
rect 56686 39312 56692 39364
rect 56744 39352 56750 39364
rect 59004 39352 59032 39460
rect 60185 39457 60197 39460
rect 60231 39457 60243 39491
rect 60185 39451 60243 39457
rect 60829 39491 60887 39497
rect 60829 39457 60841 39491
rect 60875 39488 60887 39491
rect 60918 39488 60924 39500
rect 60875 39460 60924 39488
rect 60875 39457 60887 39460
rect 60829 39451 60887 39457
rect 60918 39448 60924 39460
rect 60976 39448 60982 39500
rect 59173 39423 59231 39429
rect 59173 39389 59185 39423
rect 59219 39420 59231 39423
rect 60737 39423 60795 39429
rect 60737 39420 60749 39423
rect 59219 39392 60749 39420
rect 59219 39389 59231 39392
rect 59173 39383 59231 39389
rect 60737 39389 60749 39392
rect 60783 39389 60795 39423
rect 60737 39383 60795 39389
rect 56744 39324 59032 39352
rect 56744 39312 56750 39324
rect 59078 39312 59084 39364
rect 59136 39352 59142 39364
rect 59136 39324 59400 39352
rect 59136 39312 59142 39324
rect 59372 39296 59400 39324
rect 59446 39312 59452 39364
rect 59504 39352 59510 39364
rect 61028 39352 61056 39528
rect 65702 39516 65708 39528
rect 65760 39516 65766 39568
rect 70964 39556 70992 39596
rect 71038 39584 71044 39636
rect 71096 39624 71102 39636
rect 71593 39627 71651 39633
rect 71593 39624 71605 39627
rect 71096 39596 71605 39624
rect 71096 39584 71102 39596
rect 71593 39593 71605 39596
rect 71639 39593 71651 39627
rect 72602 39624 72608 39636
rect 72563 39596 72608 39624
rect 71593 39587 71651 39593
rect 72602 39584 72608 39596
rect 72660 39584 72666 39636
rect 77478 39624 77484 39636
rect 72712 39596 77484 39624
rect 72712 39556 72740 39596
rect 77478 39584 77484 39596
rect 77536 39624 77542 39636
rect 78769 39627 78827 39633
rect 78769 39624 78781 39627
rect 77536 39596 78781 39624
rect 77536 39584 77542 39596
rect 78769 39593 78781 39596
rect 78815 39593 78827 39627
rect 78769 39587 78827 39593
rect 81345 39627 81403 39633
rect 81345 39593 81357 39627
rect 81391 39624 81403 39627
rect 81434 39624 81440 39636
rect 81391 39596 81440 39624
rect 81391 39593 81403 39596
rect 81345 39587 81403 39593
rect 81434 39584 81440 39596
rect 81492 39584 81498 39636
rect 82998 39624 83004 39636
rect 82740 39596 83004 39624
rect 70964 39528 72740 39556
rect 61194 39488 61200 39500
rect 61155 39460 61200 39488
rect 61194 39448 61200 39460
rect 61252 39448 61258 39500
rect 62025 39491 62083 39497
rect 62025 39457 62037 39491
rect 62071 39488 62083 39491
rect 62485 39491 62543 39497
rect 62485 39488 62497 39491
rect 62071 39460 62497 39488
rect 62071 39457 62083 39460
rect 62025 39451 62083 39457
rect 62485 39457 62497 39460
rect 62531 39457 62543 39491
rect 66257 39491 66315 39497
rect 62485 39451 62543 39457
rect 64432 39460 66116 39488
rect 61289 39423 61347 39429
rect 61289 39389 61301 39423
rect 61335 39420 61347 39423
rect 61838 39420 61844 39432
rect 61335 39392 61844 39420
rect 61335 39389 61347 39392
rect 61289 39383 61347 39389
rect 61838 39380 61844 39392
rect 61896 39420 61902 39432
rect 63494 39420 63500 39432
rect 61896 39392 63500 39420
rect 61896 39380 61902 39392
rect 63494 39380 63500 39392
rect 63552 39380 63558 39432
rect 59504 39324 61056 39352
rect 59504 39312 59510 39324
rect 61102 39312 61108 39364
rect 61160 39352 61166 39364
rect 62301 39355 62359 39361
rect 62301 39352 62313 39355
rect 61160 39324 62313 39352
rect 61160 39312 61166 39324
rect 62301 39321 62313 39324
rect 62347 39352 62359 39355
rect 64432 39352 64460 39460
rect 65981 39423 66039 39429
rect 65981 39420 65993 39423
rect 62347 39324 64460 39352
rect 65812 39392 65993 39420
rect 62347 39321 62359 39324
rect 62301 39315 62359 39321
rect 48976 39256 50016 39284
rect 51629 39287 51687 39293
rect 51629 39253 51641 39287
rect 51675 39284 51687 39287
rect 53282 39284 53288 39296
rect 51675 39256 53288 39284
rect 51675 39253 51687 39256
rect 51629 39247 51687 39253
rect 53282 39244 53288 39256
rect 53340 39244 53346 39296
rect 53374 39244 53380 39296
rect 53432 39284 53438 39296
rect 53469 39287 53527 39293
rect 53469 39284 53481 39287
rect 53432 39256 53481 39284
rect 53432 39244 53438 39256
rect 53469 39253 53481 39256
rect 53515 39284 53527 39287
rect 54110 39284 54116 39296
rect 53515 39256 54116 39284
rect 53515 39253 53527 39256
rect 53469 39247 53527 39253
rect 54110 39244 54116 39256
rect 54168 39244 54174 39296
rect 54294 39284 54300 39296
rect 54255 39256 54300 39284
rect 54294 39244 54300 39256
rect 54352 39244 54358 39296
rect 54662 39244 54668 39296
rect 54720 39244 54726 39296
rect 57974 39244 57980 39296
rect 58032 39284 58038 39296
rect 59170 39284 59176 39296
rect 58032 39256 59176 39284
rect 58032 39244 58038 39256
rect 59170 39244 59176 39256
rect 59228 39244 59234 39296
rect 59354 39284 59360 39296
rect 59315 39256 59360 39284
rect 59354 39244 59360 39256
rect 59412 39244 59418 39296
rect 59538 39244 59544 39296
rect 59596 39284 59602 39296
rect 62025 39287 62083 39293
rect 62025 39284 62037 39287
rect 59596 39256 62037 39284
rect 59596 39244 59602 39256
rect 62025 39253 62037 39256
rect 62071 39284 62083 39287
rect 62117 39287 62175 39293
rect 62117 39284 62129 39287
rect 62071 39256 62129 39284
rect 62071 39253 62083 39256
rect 62025 39247 62083 39253
rect 62117 39253 62129 39256
rect 62163 39253 62175 39287
rect 62117 39247 62175 39253
rect 65334 39244 65340 39296
rect 65392 39284 65398 39296
rect 65812 39293 65840 39392
rect 65981 39389 65993 39392
rect 66027 39389 66039 39423
rect 66088 39420 66116 39460
rect 66257 39457 66269 39491
rect 66303 39488 66315 39491
rect 67450 39488 67456 39500
rect 66303 39460 67456 39488
rect 66303 39457 66315 39460
rect 66257 39451 66315 39457
rect 67450 39448 67456 39460
rect 67508 39448 67514 39500
rect 71501 39491 71559 39497
rect 71501 39457 71513 39491
rect 71547 39488 71559 39491
rect 71958 39488 71964 39500
rect 71547 39460 71964 39488
rect 71547 39457 71559 39460
rect 71501 39451 71559 39457
rect 71958 39448 71964 39460
rect 72016 39448 72022 39500
rect 72326 39448 72332 39500
rect 72384 39488 72390 39500
rect 72513 39491 72571 39497
rect 72513 39488 72525 39491
rect 72384 39460 72525 39488
rect 72384 39448 72390 39460
rect 72513 39457 72525 39460
rect 72559 39488 72571 39491
rect 73801 39491 73859 39497
rect 72559 39460 73292 39488
rect 72559 39457 72571 39460
rect 72513 39451 72571 39457
rect 72418 39420 72424 39432
rect 66088 39392 72424 39420
rect 65981 39383 66039 39389
rect 72418 39380 72424 39392
rect 72476 39380 72482 39432
rect 67542 39312 67548 39364
rect 67600 39352 67606 39364
rect 73154 39352 73160 39364
rect 67600 39324 73160 39352
rect 67600 39312 67606 39324
rect 73154 39312 73160 39324
rect 73212 39312 73218 39364
rect 65797 39287 65855 39293
rect 65797 39284 65809 39287
rect 65392 39256 65809 39284
rect 65392 39244 65398 39256
rect 65797 39253 65809 39256
rect 65843 39253 65855 39287
rect 65797 39247 65855 39253
rect 66162 39244 66168 39296
rect 66220 39284 66226 39296
rect 67361 39287 67419 39293
rect 67361 39284 67373 39287
rect 66220 39256 67373 39284
rect 66220 39244 66226 39256
rect 67361 39253 67373 39256
rect 67407 39253 67419 39287
rect 73264 39284 73292 39460
rect 73801 39457 73813 39491
rect 73847 39488 73859 39491
rect 74902 39488 74908 39500
rect 73847 39460 74908 39488
rect 73847 39457 73859 39460
rect 73801 39451 73859 39457
rect 74902 39448 74908 39460
rect 74960 39448 74966 39500
rect 75365 39491 75423 39497
rect 75365 39457 75377 39491
rect 75411 39488 75423 39491
rect 77294 39488 77300 39500
rect 75411 39460 77300 39488
rect 75411 39457 75423 39460
rect 75365 39451 75423 39457
rect 73525 39423 73583 39429
rect 73525 39389 73537 39423
rect 73571 39420 73583 39423
rect 73890 39420 73896 39432
rect 73571 39392 73896 39420
rect 73571 39389 73583 39392
rect 73525 39383 73583 39389
rect 73890 39380 73896 39392
rect 73948 39420 73954 39432
rect 75380 39420 75408 39451
rect 77294 39448 77300 39460
rect 77352 39488 77358 39500
rect 77389 39491 77447 39497
rect 77389 39488 77401 39491
rect 77352 39460 77401 39488
rect 77352 39448 77358 39460
rect 77389 39457 77401 39460
rect 77435 39488 77447 39491
rect 78306 39488 78312 39500
rect 77435 39460 78312 39488
rect 77435 39457 77447 39460
rect 77389 39451 77447 39457
rect 78306 39448 78312 39460
rect 78364 39448 78370 39500
rect 79870 39488 79876 39500
rect 79831 39460 79876 39488
rect 79870 39448 79876 39460
rect 79928 39448 79934 39500
rect 81253 39491 81311 39497
rect 81253 39457 81265 39491
rect 81299 39488 81311 39491
rect 81342 39488 81348 39500
rect 81299 39460 81348 39488
rect 81299 39457 81311 39460
rect 81253 39451 81311 39457
rect 81342 39448 81348 39460
rect 81400 39448 81406 39500
rect 82740 39497 82768 39596
rect 82998 39584 83004 39596
rect 83056 39624 83062 39636
rect 85666 39624 85672 39636
rect 83056 39596 85672 39624
rect 83056 39584 83062 39596
rect 85666 39584 85672 39596
rect 85724 39584 85730 39636
rect 85942 39624 85948 39636
rect 85903 39596 85948 39624
rect 85942 39584 85948 39596
rect 86000 39584 86006 39636
rect 88797 39627 88855 39633
rect 88797 39593 88809 39627
rect 88843 39624 88855 39627
rect 89438 39624 89444 39636
rect 88843 39596 89444 39624
rect 88843 39593 88855 39596
rect 88797 39587 88855 39593
rect 89438 39584 89444 39596
rect 89496 39584 89502 39636
rect 91094 39624 91100 39636
rect 91055 39596 91100 39624
rect 91094 39584 91100 39596
rect 91152 39584 91158 39636
rect 83737 39559 83795 39565
rect 83737 39525 83749 39559
rect 83783 39556 83795 39559
rect 83783 39528 88748 39556
rect 83783 39525 83795 39528
rect 83737 39519 83795 39525
rect 82725 39491 82783 39497
rect 82725 39457 82737 39491
rect 82771 39457 82783 39491
rect 82725 39451 82783 39457
rect 82817 39491 82875 39497
rect 82817 39457 82829 39491
rect 82863 39488 82875 39491
rect 83826 39488 83832 39500
rect 82863 39460 83832 39488
rect 82863 39457 82875 39460
rect 82817 39451 82875 39457
rect 83826 39448 83832 39460
rect 83884 39488 83890 39500
rect 84381 39491 84439 39497
rect 84381 39488 84393 39491
rect 83884 39460 84393 39488
rect 83884 39448 83890 39460
rect 84381 39457 84393 39460
rect 84427 39457 84439 39491
rect 84381 39451 84439 39457
rect 84562 39448 84568 39500
rect 84620 39488 84626 39500
rect 84749 39491 84807 39497
rect 84749 39488 84761 39491
rect 84620 39460 84761 39488
rect 84620 39448 84626 39460
rect 84749 39457 84761 39460
rect 84795 39488 84807 39491
rect 85025 39491 85083 39497
rect 85025 39488 85037 39491
rect 84795 39460 85037 39488
rect 84795 39457 84807 39460
rect 84749 39451 84807 39457
rect 85025 39457 85037 39460
rect 85071 39457 85083 39491
rect 85758 39488 85764 39500
rect 85719 39460 85764 39488
rect 85025 39451 85083 39457
rect 85758 39448 85764 39460
rect 85816 39488 85822 39500
rect 86129 39491 86187 39497
rect 86129 39488 86141 39491
rect 85816 39460 86141 39488
rect 85816 39448 85822 39460
rect 86129 39457 86141 39460
rect 86175 39457 86187 39491
rect 86862 39488 86868 39500
rect 86823 39460 86868 39488
rect 86129 39451 86187 39457
rect 86862 39448 86868 39460
rect 86920 39488 86926 39500
rect 88720 39497 88748 39528
rect 87141 39491 87199 39497
rect 87141 39488 87153 39491
rect 86920 39460 87153 39488
rect 86920 39448 86926 39460
rect 87141 39457 87153 39460
rect 87187 39457 87199 39491
rect 87141 39451 87199 39457
rect 88705 39491 88763 39497
rect 88705 39457 88717 39491
rect 88751 39457 88763 39491
rect 89898 39488 89904 39500
rect 89859 39460 89904 39488
rect 88705 39451 88763 39457
rect 89898 39448 89904 39460
rect 89956 39448 89962 39500
rect 91002 39488 91008 39500
rect 90963 39460 91008 39488
rect 91002 39448 91008 39460
rect 91060 39448 91066 39500
rect 73948 39392 75408 39420
rect 77665 39423 77723 39429
rect 73948 39380 73954 39392
rect 77665 39389 77677 39423
rect 77711 39420 77723 39423
rect 79965 39423 80023 39429
rect 79965 39420 79977 39423
rect 77711 39392 79977 39420
rect 77711 39389 77723 39392
rect 77665 39383 77723 39389
rect 79965 39389 79977 39392
rect 80011 39389 80023 39423
rect 79965 39383 80023 39389
rect 82354 39380 82360 39432
rect 82412 39420 82418 39432
rect 84102 39420 84108 39432
rect 82412 39392 84108 39420
rect 82412 39380 82418 39392
rect 84102 39380 84108 39392
rect 84160 39380 84166 39432
rect 84473 39423 84531 39429
rect 84473 39389 84485 39423
rect 84519 39389 84531 39423
rect 84838 39420 84844 39432
rect 84799 39392 84844 39420
rect 84473 39383 84531 39389
rect 80514 39312 80520 39364
rect 80572 39352 80578 39364
rect 83274 39352 83280 39364
rect 80572 39324 83280 39352
rect 80572 39312 80578 39324
rect 83274 39312 83280 39324
rect 83332 39352 83338 39364
rect 83645 39355 83703 39361
rect 83645 39352 83657 39355
rect 83332 39324 83657 39352
rect 83332 39312 83338 39324
rect 83645 39321 83657 39324
rect 83691 39352 83703 39355
rect 84488 39352 84516 39383
rect 84838 39380 84844 39392
rect 84896 39380 84902 39432
rect 84930 39380 84936 39432
rect 84988 39420 84994 39432
rect 88518 39420 88524 39432
rect 84988 39392 88524 39420
rect 84988 39380 84994 39392
rect 88518 39380 88524 39392
rect 88576 39380 88582 39432
rect 90082 39352 90088 39364
rect 83691 39324 90088 39352
rect 83691 39321 83703 39324
rect 83645 39315 83703 39321
rect 90082 39312 90088 39324
rect 90140 39312 90146 39364
rect 74902 39284 74908 39296
rect 73264 39256 74908 39284
rect 67361 39247 67419 39253
rect 74902 39244 74908 39256
rect 74960 39244 74966 39296
rect 83734 39244 83740 39296
rect 83792 39284 83798 39296
rect 84562 39284 84568 39296
rect 83792 39256 84568 39284
rect 83792 39244 83798 39256
rect 84562 39244 84568 39256
rect 84620 39244 84626 39296
rect 86218 39244 86224 39296
rect 86276 39284 86282 39296
rect 86957 39287 87015 39293
rect 86957 39284 86969 39287
rect 86276 39256 86969 39284
rect 86276 39244 86282 39256
rect 86957 39253 86969 39256
rect 87003 39253 87015 39287
rect 86957 39247 87015 39253
rect 88518 39244 88524 39296
rect 88576 39284 88582 39296
rect 89993 39287 90051 39293
rect 89993 39284 90005 39287
rect 88576 39256 90005 39284
rect 88576 39244 88582 39256
rect 89993 39253 90005 39256
rect 90039 39253 90051 39287
rect 89993 39247 90051 39253
rect 1104 39194 105616 39216
rect 1104 39142 4246 39194
rect 4298 39142 4310 39194
rect 4362 39142 4374 39194
rect 4426 39142 4438 39194
rect 4490 39142 34966 39194
rect 35018 39142 35030 39194
rect 35082 39142 35094 39194
rect 35146 39142 35158 39194
rect 35210 39142 65686 39194
rect 65738 39142 65750 39194
rect 65802 39142 65814 39194
rect 65866 39142 65878 39194
rect 65930 39142 96406 39194
rect 96458 39142 96470 39194
rect 96522 39142 96534 39194
rect 96586 39142 96598 39194
rect 96650 39142 105616 39194
rect 1104 39120 105616 39142
rect 3418 39040 3424 39092
rect 3476 39080 3482 39092
rect 7926 39080 7932 39092
rect 3476 39052 7932 39080
rect 3476 39040 3482 39052
rect 7926 39040 7932 39052
rect 7984 39040 7990 39092
rect 8941 39083 8999 39089
rect 8941 39049 8953 39083
rect 8987 39080 8999 39083
rect 13814 39080 13820 39092
rect 8987 39052 13820 39080
rect 8987 39049 8999 39052
rect 8941 39043 8999 39049
rect 2774 38904 2780 38956
rect 2832 38944 2838 38956
rect 2832 38916 2877 38944
rect 2832 38904 2838 38916
rect 7466 38904 7472 38956
rect 7524 38944 7530 38956
rect 7524 38916 8524 38944
rect 7524 38904 7530 38916
rect 8496 38888 8524 38916
rect 2501 38879 2559 38885
rect 2501 38845 2513 38879
rect 2547 38876 2559 38879
rect 8021 38879 8079 38885
rect 2547 38848 4384 38876
rect 2547 38845 2559 38848
rect 2501 38839 2559 38845
rect 3878 38740 3884 38752
rect 3839 38712 3884 38740
rect 3878 38700 3884 38712
rect 3936 38700 3942 38752
rect 4356 38749 4384 38848
rect 8021 38845 8033 38879
rect 8067 38845 8079 38879
rect 8202 38876 8208 38888
rect 8163 38848 8208 38876
rect 8021 38839 8079 38845
rect 6270 38768 6276 38820
rect 6328 38808 6334 38820
rect 7561 38811 7619 38817
rect 7561 38808 7573 38811
rect 6328 38780 7573 38808
rect 6328 38768 6334 38780
rect 7561 38777 7573 38780
rect 7607 38777 7619 38811
rect 8036 38808 8064 38839
rect 8202 38836 8208 38848
rect 8260 38836 8266 38888
rect 8478 38836 8484 38888
rect 8536 38876 8542 38888
rect 8573 38879 8631 38885
rect 8573 38876 8585 38879
rect 8536 38848 8585 38876
rect 8536 38836 8542 38848
rect 8573 38845 8585 38848
rect 8619 38845 8631 38879
rect 8573 38839 8631 38845
rect 8757 38879 8815 38885
rect 8757 38845 8769 38879
rect 8803 38876 8815 38879
rect 8956 38876 8984 39043
rect 13814 39040 13820 39052
rect 13872 39040 13878 39092
rect 20714 39080 20720 39092
rect 20675 39052 20720 39080
rect 20714 39040 20720 39052
rect 20772 39040 20778 39092
rect 21358 39040 21364 39092
rect 21416 39080 21422 39092
rect 38654 39080 38660 39092
rect 21416 39052 38660 39080
rect 21416 39040 21422 39052
rect 38654 39040 38660 39052
rect 38712 39040 38718 39092
rect 48314 39040 48320 39092
rect 48372 39080 48378 39092
rect 48372 39052 50844 39080
rect 48372 39040 48378 39052
rect 9125 39015 9183 39021
rect 9125 38981 9137 39015
rect 9171 39012 9183 39015
rect 12618 39012 12624 39024
rect 9171 38984 12624 39012
rect 9171 38981 9183 38984
rect 9125 38975 9183 38981
rect 8803 38848 8984 38876
rect 8803 38845 8815 38848
rect 8757 38839 8815 38845
rect 9140 38808 9168 38975
rect 12618 38972 12624 38984
rect 12676 38972 12682 39024
rect 15289 39015 15347 39021
rect 15289 39012 15301 39015
rect 13832 38984 15301 39012
rect 13832 38956 13860 38984
rect 15289 38981 15301 38984
rect 15335 38981 15347 39015
rect 15289 38975 15347 38981
rect 20806 38972 20812 39024
rect 20864 39012 20870 39024
rect 22002 39012 22008 39024
rect 20864 38984 22008 39012
rect 20864 38972 20870 38984
rect 22002 38972 22008 38984
rect 22060 38972 22066 39024
rect 31849 39015 31907 39021
rect 31849 38981 31861 39015
rect 31895 39012 31907 39015
rect 32766 39012 32772 39024
rect 31895 38984 32260 39012
rect 31895 38981 31907 38984
rect 31849 38975 31907 38981
rect 11425 38947 11483 38953
rect 11425 38913 11437 38947
rect 11471 38944 11483 38947
rect 12989 38947 13047 38953
rect 12989 38944 13001 38947
rect 11471 38916 13001 38944
rect 11471 38913 11483 38916
rect 11425 38907 11483 38913
rect 12989 38913 13001 38916
rect 13035 38913 13047 38947
rect 12989 38907 13047 38913
rect 13814 38904 13820 38956
rect 13872 38904 13878 38956
rect 14369 38947 14427 38953
rect 14369 38913 14381 38947
rect 14415 38944 14427 38947
rect 15105 38947 15163 38953
rect 15105 38944 15117 38947
rect 14415 38916 15117 38944
rect 14415 38913 14427 38916
rect 14369 38907 14427 38913
rect 15105 38913 15117 38916
rect 15151 38944 15163 38947
rect 24118 38944 24124 38956
rect 15151 38916 24124 38944
rect 15151 38913 15163 38916
rect 15105 38907 15163 38913
rect 10137 38879 10195 38885
rect 10137 38876 10149 38879
rect 8036 38780 9168 38808
rect 9968 38848 10149 38876
rect 7561 38771 7619 38777
rect 9968 38752 9996 38848
rect 10137 38845 10149 38848
rect 10183 38845 10195 38879
rect 10137 38839 10195 38845
rect 10321 38879 10379 38885
rect 10321 38845 10333 38879
rect 10367 38845 10379 38879
rect 10778 38876 10784 38888
rect 10739 38848 10784 38876
rect 10321 38839 10379 38845
rect 10336 38808 10364 38839
rect 10778 38836 10784 38848
rect 10836 38836 10842 38888
rect 10873 38879 10931 38885
rect 10873 38845 10885 38879
rect 10919 38876 10931 38879
rect 12066 38876 12072 38888
rect 10919 38848 12072 38876
rect 10919 38845 10931 38848
rect 10873 38839 10931 38845
rect 10888 38808 10916 38839
rect 12066 38836 12072 38848
rect 12124 38836 12130 38888
rect 12713 38879 12771 38885
rect 12713 38845 12725 38879
rect 12759 38876 12771 38879
rect 13630 38876 13636 38888
rect 12759 38848 13636 38876
rect 12759 38845 12771 38848
rect 12713 38839 12771 38845
rect 13630 38836 13636 38848
rect 13688 38876 13694 38888
rect 15212 38885 15240 38916
rect 24118 38904 24124 38916
rect 24176 38904 24182 38956
rect 26326 38904 26332 38956
rect 26384 38944 26390 38956
rect 31573 38947 31631 38953
rect 31573 38944 31585 38947
rect 26384 38916 31585 38944
rect 26384 38904 26390 38916
rect 31573 38913 31585 38916
rect 31619 38944 31631 38947
rect 31941 38947 31999 38953
rect 31941 38944 31953 38947
rect 31619 38916 31953 38944
rect 31619 38913 31631 38916
rect 31573 38907 31631 38913
rect 31941 38913 31953 38916
rect 31987 38913 31999 38947
rect 32232 38944 32260 38984
rect 31941 38907 31999 38913
rect 32048 38916 32260 38944
rect 14461 38879 14519 38885
rect 14461 38876 14473 38879
rect 13688 38848 14473 38876
rect 13688 38836 13694 38848
rect 14461 38845 14473 38848
rect 14507 38845 14519 38879
rect 14461 38839 14519 38845
rect 15197 38879 15255 38885
rect 15197 38845 15209 38879
rect 15243 38876 15255 38879
rect 19153 38879 19211 38885
rect 15243 38848 15277 38876
rect 15243 38845 15255 38848
rect 15197 38839 15255 38845
rect 19153 38845 19165 38879
rect 19199 38876 19211 38879
rect 19242 38876 19248 38888
rect 19199 38848 19248 38876
rect 19199 38845 19211 38848
rect 19153 38839 19211 38845
rect 10336 38780 10916 38808
rect 14476 38808 14504 38839
rect 19168 38808 19196 38839
rect 19242 38836 19248 38848
rect 19300 38836 19306 38888
rect 19426 38876 19432 38888
rect 19387 38848 19432 38876
rect 19426 38836 19432 38848
rect 19484 38836 19490 38888
rect 19886 38836 19892 38888
rect 19944 38876 19950 38888
rect 20346 38876 20352 38888
rect 19944 38848 20352 38876
rect 19944 38836 19950 38848
rect 20346 38836 20352 38848
rect 20404 38836 20410 38888
rect 21634 38876 21640 38888
rect 21595 38848 21640 38876
rect 21634 38836 21640 38848
rect 21692 38836 21698 38888
rect 26145 38879 26203 38885
rect 26145 38845 26157 38879
rect 26191 38845 26203 38879
rect 26418 38876 26424 38888
rect 26379 38848 26424 38876
rect 26145 38839 26203 38845
rect 26160 38808 26188 38839
rect 26418 38836 26424 38848
rect 26476 38836 26482 38888
rect 27801 38879 27859 38885
rect 27801 38845 27813 38879
rect 27847 38876 27859 38879
rect 29273 38879 29331 38885
rect 29273 38876 29285 38879
rect 27847 38848 29285 38876
rect 27847 38845 27859 38848
rect 27801 38839 27859 38845
rect 29273 38845 29285 38848
rect 29319 38845 29331 38879
rect 29273 38839 29331 38845
rect 14476 38780 19196 38808
rect 4341 38743 4399 38749
rect 4341 38709 4353 38743
rect 4387 38740 4399 38743
rect 4706 38740 4712 38752
rect 4387 38712 4712 38740
rect 4387 38709 4399 38712
rect 4341 38703 4399 38709
rect 4706 38700 4712 38712
rect 4764 38700 4770 38752
rect 9950 38740 9956 38752
rect 9911 38712 9956 38740
rect 9950 38700 9956 38712
rect 10008 38700 10014 38752
rect 10778 38700 10784 38752
rect 10836 38740 10842 38752
rect 13814 38740 13820 38752
rect 10836 38712 13820 38740
rect 10836 38700 10842 38712
rect 13814 38700 13820 38712
rect 13872 38700 13878 38752
rect 19168 38740 19196 38780
rect 20916 38780 26188 38808
rect 20916 38749 20944 38780
rect 20901 38743 20959 38749
rect 20901 38740 20913 38743
rect 19168 38712 20913 38740
rect 20901 38709 20913 38712
rect 20947 38709 20959 38743
rect 20901 38703 20959 38709
rect 20990 38700 20996 38752
rect 21048 38740 21054 38752
rect 21729 38743 21787 38749
rect 21729 38740 21741 38743
rect 21048 38712 21741 38740
rect 21048 38700 21054 38712
rect 21729 38709 21741 38712
rect 21775 38709 21787 38743
rect 26160 38740 26188 38780
rect 27154 38768 27160 38820
rect 27212 38808 27218 38820
rect 27212 38780 29408 38808
rect 27212 38768 27218 38780
rect 27893 38743 27951 38749
rect 27893 38740 27905 38743
rect 26160 38712 27905 38740
rect 21729 38703 21787 38709
rect 27893 38709 27905 38712
rect 27939 38740 27951 38743
rect 28258 38740 28264 38752
rect 27939 38712 28264 38740
rect 27939 38709 27951 38712
rect 27893 38703 27951 38709
rect 28258 38700 28264 38712
rect 28316 38700 28322 38752
rect 29380 38749 29408 38780
rect 29365 38743 29423 38749
rect 29365 38709 29377 38743
rect 29411 38740 29423 38743
rect 32048 38740 32076 38916
rect 32125 38879 32183 38885
rect 32125 38845 32137 38879
rect 32171 38845 32183 38879
rect 32125 38839 32183 38845
rect 29411 38712 32076 38740
rect 32140 38740 32168 38839
rect 32232 38808 32260 38916
rect 32324 38984 32772 39012
rect 32324 38876 32352 38984
rect 32766 38972 32772 38984
rect 32824 39012 32830 39024
rect 33137 39015 33195 39021
rect 32824 38984 33088 39012
rect 32824 38972 32830 38984
rect 33060 38944 33088 38984
rect 33137 38981 33149 39015
rect 33183 39012 33195 39015
rect 34514 39012 34520 39024
rect 33183 38984 34520 39012
rect 33183 38981 33195 38984
rect 33137 38975 33195 38981
rect 34514 38972 34520 38984
rect 34572 38972 34578 39024
rect 39022 39021 39028 39024
rect 39006 39015 39028 39021
rect 39006 38981 39018 39015
rect 39006 38975 39028 38981
rect 39022 38972 39028 38975
rect 39080 38972 39086 39024
rect 39117 39015 39175 39021
rect 39117 38981 39129 39015
rect 39163 39012 39175 39015
rect 39761 39015 39819 39021
rect 39761 39012 39773 39015
rect 39163 38984 39773 39012
rect 39163 38981 39175 38984
rect 39117 38975 39175 38981
rect 39761 38981 39773 38984
rect 39807 39012 39819 39015
rect 46198 39012 46204 39024
rect 39807 38984 46204 39012
rect 39807 38981 39819 38984
rect 39761 38975 39819 38981
rect 46198 38972 46204 38984
rect 46256 38972 46262 39024
rect 46385 39015 46443 39021
rect 46385 38981 46397 39015
rect 46431 39012 46443 39015
rect 46431 38984 49832 39012
rect 46431 38981 46443 38984
rect 46385 38975 46443 38981
rect 33689 38947 33747 38953
rect 33689 38944 33701 38947
rect 33060 38916 33701 38944
rect 33689 38913 33701 38916
rect 33735 38944 33747 38947
rect 33870 38944 33876 38956
rect 33735 38916 33876 38944
rect 33735 38913 33747 38916
rect 33689 38907 33747 38913
rect 33870 38904 33876 38916
rect 33928 38944 33934 38956
rect 33928 38916 34468 38944
rect 33928 38904 33934 38916
rect 32677 38879 32735 38885
rect 32677 38876 32689 38879
rect 32324 38848 32689 38876
rect 32677 38845 32689 38848
rect 32723 38845 32735 38879
rect 32677 38839 32735 38845
rect 32861 38879 32919 38885
rect 32861 38845 32873 38879
rect 32907 38876 32919 38879
rect 32907 38848 34376 38876
rect 32907 38845 32919 38848
rect 32861 38839 32919 38845
rect 32876 38808 32904 38839
rect 33502 38808 33508 38820
rect 32232 38780 32904 38808
rect 33463 38780 33508 38808
rect 33502 38768 33508 38780
rect 33560 38768 33566 38820
rect 32306 38740 32312 38752
rect 32140 38712 32312 38740
rect 29411 38709 29423 38712
rect 29365 38703 29423 38709
rect 32306 38700 32312 38712
rect 32364 38740 32370 38752
rect 33520 38740 33548 38768
rect 32364 38712 33548 38740
rect 34348 38740 34376 38848
rect 34440 38808 34468 38916
rect 38746 38904 38752 38956
rect 38804 38944 38810 38956
rect 39209 38947 39267 38953
rect 39209 38944 39221 38947
rect 38804 38916 39221 38944
rect 38804 38904 38810 38916
rect 39209 38913 39221 38916
rect 39255 38913 39267 38947
rect 39209 38907 39267 38913
rect 39574 38904 39580 38956
rect 39632 38944 39638 38956
rect 45094 38944 45100 38956
rect 39632 38916 41092 38944
rect 39632 38904 39638 38916
rect 38838 38876 38844 38888
rect 38799 38848 38844 38876
rect 38838 38836 38844 38848
rect 38896 38836 38902 38888
rect 40954 38876 40960 38888
rect 38948 38848 40960 38876
rect 38948 38808 38976 38848
rect 40954 38836 40960 38848
rect 41012 38836 41018 38888
rect 34440 38780 38976 38808
rect 39577 38811 39635 38817
rect 39577 38777 39589 38811
rect 39623 38808 39635 38811
rect 40218 38808 40224 38820
rect 39623 38780 40224 38808
rect 39623 38777 39635 38780
rect 39577 38771 39635 38777
rect 40218 38768 40224 38780
rect 40276 38768 40282 38820
rect 41064 38808 41092 38916
rect 43824 38916 44220 38944
rect 45055 38916 45100 38944
rect 43824 38888 43852 38916
rect 43806 38876 43812 38888
rect 43767 38848 43812 38876
rect 43806 38836 43812 38848
rect 43864 38836 43870 38888
rect 43993 38879 44051 38885
rect 43993 38845 44005 38879
rect 44039 38876 44051 38879
rect 44082 38876 44088 38888
rect 44039 38848 44088 38876
rect 44039 38845 44051 38848
rect 43993 38839 44051 38845
rect 44082 38836 44088 38848
rect 44140 38836 44146 38888
rect 44192 38876 44220 38916
rect 45094 38904 45100 38916
rect 45152 38904 45158 38956
rect 45373 38947 45431 38953
rect 45373 38913 45385 38947
rect 45419 38944 45431 38947
rect 45557 38947 45615 38953
rect 45557 38944 45569 38947
rect 45419 38916 45569 38944
rect 45419 38913 45431 38916
rect 45373 38907 45431 38913
rect 45557 38913 45569 38916
rect 45603 38944 45615 38947
rect 45922 38944 45928 38956
rect 45603 38916 45928 38944
rect 45603 38913 45615 38916
rect 45557 38907 45615 38913
rect 44453 38879 44511 38885
rect 44453 38876 44465 38879
rect 44192 38848 44465 38876
rect 44453 38845 44465 38848
rect 44499 38845 44511 38879
rect 44453 38839 44511 38845
rect 44545 38879 44603 38885
rect 44545 38845 44557 38879
rect 44591 38876 44603 38879
rect 44910 38876 44916 38888
rect 44591 38848 44916 38876
rect 44591 38845 44603 38848
rect 44545 38839 44603 38845
rect 44910 38836 44916 38848
rect 44968 38876 44974 38888
rect 45388 38876 45416 38907
rect 45922 38904 45928 38916
rect 45980 38904 45986 38956
rect 46477 38947 46535 38953
rect 46477 38913 46489 38947
rect 46523 38944 46535 38947
rect 47026 38944 47032 38956
rect 46523 38916 47032 38944
rect 46523 38913 46535 38916
rect 46477 38907 46535 38913
rect 47026 38904 47032 38916
rect 47084 38904 47090 38956
rect 48958 38944 48964 38956
rect 48700 38916 48964 38944
rect 46106 38876 46112 38888
rect 44968 38848 45416 38876
rect 46067 38848 46112 38876
rect 44968 38836 44974 38848
rect 46106 38836 46112 38848
rect 46164 38836 46170 38888
rect 46256 38879 46314 38885
rect 46256 38845 46268 38879
rect 46302 38876 46314 38879
rect 46566 38876 46572 38888
rect 46302 38848 46572 38876
rect 46302 38845 46314 38848
rect 46256 38839 46314 38845
rect 46566 38836 46572 38848
rect 46624 38836 46630 38888
rect 46658 38836 46664 38888
rect 46716 38876 46722 38888
rect 48700 38885 48728 38916
rect 48958 38904 48964 38916
rect 49016 38904 49022 38956
rect 49804 38944 49832 38984
rect 49878 38972 49884 39024
rect 49936 39012 49942 39024
rect 50430 39012 50436 39024
rect 49936 38984 49981 39012
rect 50391 38984 50436 39012
rect 49936 38972 49942 38984
rect 50430 38972 50436 38984
rect 50488 38972 50494 39024
rect 50617 39015 50675 39021
rect 50617 38981 50629 39015
rect 50663 39012 50675 39015
rect 50706 39012 50712 39024
rect 50663 38984 50712 39012
rect 50663 38981 50675 38984
rect 50617 38975 50675 38981
rect 50706 38972 50712 38984
rect 50764 38972 50770 39024
rect 50816 39012 50844 39052
rect 51442 39040 51448 39092
rect 51500 39080 51506 39092
rect 51859 39083 51917 39089
rect 51859 39080 51871 39083
rect 51500 39052 51871 39080
rect 51500 39040 51506 39052
rect 51859 39049 51871 39052
rect 51905 39049 51917 39083
rect 51859 39043 51917 39049
rect 52178 39040 52184 39092
rect 52236 39080 52242 39092
rect 61102 39080 61108 39092
rect 52236 39052 61108 39080
rect 52236 39040 52242 39052
rect 61102 39040 61108 39052
rect 61160 39040 61166 39092
rect 83734 39080 83740 39092
rect 61212 39052 83740 39080
rect 51997 39015 52055 39021
rect 50816 38984 51948 39012
rect 51074 38944 51080 38956
rect 49804 38916 51080 38944
rect 51074 38904 51080 38916
rect 51132 38904 51138 38956
rect 48501 38879 48559 38885
rect 48501 38876 48513 38879
rect 46716 38848 48513 38876
rect 46716 38836 46722 38848
rect 48501 38845 48513 38848
rect 48547 38876 48559 38879
rect 48685 38879 48743 38885
rect 48685 38876 48697 38879
rect 48547 38848 48697 38876
rect 48547 38845 48559 38848
rect 48501 38839 48559 38845
rect 48685 38845 48697 38848
rect 48731 38845 48743 38879
rect 48866 38876 48872 38888
rect 48827 38848 48872 38876
rect 48685 38839 48743 38845
rect 48866 38836 48872 38848
rect 48924 38836 48930 38888
rect 49418 38876 49424 38888
rect 49379 38848 49424 38876
rect 49418 38836 49424 38848
rect 49476 38836 49482 38888
rect 49510 38836 49516 38888
rect 49568 38876 49574 38888
rect 49605 38879 49663 38885
rect 49605 38876 49617 38879
rect 49568 38848 49617 38876
rect 49568 38836 49574 38848
rect 49605 38845 49617 38848
rect 49651 38845 49663 38879
rect 51920 38876 51948 38984
rect 51997 38981 52009 39015
rect 52043 39012 52055 39015
rect 52546 39012 52552 39024
rect 52043 38984 52552 39012
rect 52043 38981 52055 38984
rect 51997 38975 52055 38981
rect 52546 38972 52552 38984
rect 52604 38972 52610 39024
rect 54202 38972 54208 39024
rect 54260 39012 54266 39024
rect 60642 39012 60648 39024
rect 54260 38984 60648 39012
rect 54260 38972 54266 38984
rect 60642 38972 60648 38984
rect 60700 38972 60706 39024
rect 60734 38972 60740 39024
rect 60792 39012 60798 39024
rect 60792 38984 60837 39012
rect 60792 38972 60798 38984
rect 61010 38972 61016 39024
rect 61068 39012 61074 39024
rect 61212 39012 61240 39052
rect 83734 39040 83740 39052
rect 83792 39040 83798 39092
rect 84013 39083 84071 39089
rect 84013 39080 84025 39083
rect 83936 39052 84025 39080
rect 61068 38984 61240 39012
rect 61068 38972 61074 38984
rect 64138 38972 64144 39024
rect 64196 39012 64202 39024
rect 65518 39012 65524 39024
rect 64196 38984 65524 39012
rect 64196 38972 64202 38984
rect 65518 38972 65524 38984
rect 65576 39012 65582 39024
rect 67634 39012 67640 39024
rect 65576 38984 67640 39012
rect 65576 38972 65582 38984
rect 67634 38972 67640 38984
rect 67692 38972 67698 39024
rect 80882 38972 80888 39024
rect 80940 39012 80946 39024
rect 80940 38984 83044 39012
rect 80940 38972 80946 38984
rect 52086 38944 52092 38956
rect 52047 38916 52092 38944
rect 52086 38904 52092 38916
rect 52144 38904 52150 38956
rect 52454 38944 52460 38956
rect 52415 38916 52460 38944
rect 52454 38904 52460 38916
rect 52512 38904 52518 38956
rect 52564 38916 54616 38944
rect 52564 38876 52592 38916
rect 49605 38839 49663 38845
rect 49712 38848 51856 38876
rect 51920 38848 52592 38876
rect 49712 38808 49740 38848
rect 51721 38811 51779 38817
rect 51721 38808 51733 38811
rect 41064 38780 49740 38808
rect 51460 38780 51733 38808
rect 51460 38752 51488 38780
rect 51721 38777 51733 38780
rect 51767 38777 51779 38811
rect 51828 38808 51856 38848
rect 54202 38836 54208 38888
rect 54260 38836 54266 38888
rect 54305 38879 54363 38885
rect 54305 38845 54317 38879
rect 54351 38876 54363 38879
rect 54588 38876 54616 38916
rect 54662 38904 54668 38956
rect 54720 38944 54726 38956
rect 54720 38916 58848 38944
rect 54720 38904 54726 38916
rect 57974 38876 57980 38888
rect 54351 38848 54432 38876
rect 54588 38848 57980 38876
rect 54351 38845 54363 38848
rect 54305 38839 54363 38845
rect 54220 38808 54248 38836
rect 51828 38780 54248 38808
rect 51721 38771 51779 38777
rect 42886 38740 42892 38752
rect 34348 38712 42892 38740
rect 32364 38700 32370 38712
rect 42886 38700 42892 38712
rect 42944 38700 42950 38752
rect 43254 38700 43260 38752
rect 43312 38740 43318 38752
rect 43441 38743 43499 38749
rect 43441 38740 43453 38743
rect 43312 38712 43453 38740
rect 43312 38700 43318 38712
rect 43441 38709 43453 38712
rect 43487 38740 43499 38743
rect 43625 38743 43683 38749
rect 43625 38740 43637 38743
rect 43487 38712 43637 38740
rect 43487 38709 43499 38712
rect 43441 38703 43499 38709
rect 43625 38709 43637 38712
rect 43671 38740 43683 38743
rect 43806 38740 43812 38752
rect 43671 38712 43812 38740
rect 43671 38709 43683 38712
rect 43625 38703 43683 38709
rect 43806 38700 43812 38712
rect 43864 38700 43870 38752
rect 43898 38700 43904 38752
rect 43956 38740 43962 38752
rect 46658 38740 46664 38752
rect 43956 38712 46664 38740
rect 43956 38700 43962 38712
rect 46658 38700 46664 38712
rect 46716 38700 46722 38752
rect 46753 38743 46811 38749
rect 46753 38709 46765 38743
rect 46799 38740 46811 38743
rect 48406 38740 48412 38752
rect 46799 38712 48412 38740
rect 46799 38709 46811 38712
rect 46753 38703 46811 38709
rect 48406 38700 48412 38712
rect 48464 38700 48470 38752
rect 49510 38700 49516 38752
rect 49568 38740 49574 38752
rect 50157 38743 50215 38749
rect 50157 38740 50169 38743
rect 49568 38712 50169 38740
rect 49568 38700 49574 38712
rect 50157 38709 50169 38712
rect 50203 38709 50215 38743
rect 51442 38740 51448 38752
rect 51403 38712 51448 38740
rect 50157 38703 50215 38709
rect 51442 38700 51448 38712
rect 51500 38700 51506 38752
rect 54113 38743 54171 38749
rect 54113 38709 54125 38743
rect 54159 38740 54171 38743
rect 54202 38740 54208 38752
rect 54159 38712 54208 38740
rect 54159 38709 54171 38712
rect 54113 38703 54171 38709
rect 54202 38700 54208 38712
rect 54260 38700 54266 38752
rect 54404 38740 54432 38848
rect 57974 38836 57980 38848
rect 58032 38836 58038 38888
rect 58250 38876 58256 38888
rect 58211 38848 58256 38876
rect 58250 38836 58256 38848
rect 58308 38876 58314 38888
rect 58437 38879 58495 38885
rect 58437 38876 58449 38879
rect 58308 38848 58449 38876
rect 58308 38836 58314 38848
rect 58437 38845 58449 38848
rect 58483 38845 58495 38879
rect 58618 38876 58624 38888
rect 58579 38848 58624 38876
rect 58437 38839 58495 38845
rect 58618 38836 58624 38848
rect 58676 38836 58682 38888
rect 58820 38876 58848 38916
rect 67542 38904 67548 38956
rect 67600 38944 67606 38956
rect 70210 38944 70216 38956
rect 67600 38916 70216 38944
rect 67600 38904 67606 38916
rect 70210 38904 70216 38916
rect 70268 38904 70274 38956
rect 71593 38947 71651 38953
rect 71593 38913 71605 38947
rect 71639 38913 71651 38947
rect 71593 38907 71651 38913
rect 59078 38876 59084 38888
rect 58820 38848 58940 38876
rect 59039 38848 59084 38876
rect 54478 38768 54484 38820
rect 54536 38808 54542 38820
rect 58912 38808 58940 38848
rect 59078 38836 59084 38848
rect 59136 38836 59142 38888
rect 59173 38879 59231 38885
rect 59173 38845 59185 38879
rect 59219 38876 59231 38879
rect 59354 38876 59360 38888
rect 59219 38848 59360 38876
rect 59219 38845 59231 38848
rect 59173 38839 59231 38845
rect 59354 38836 59360 38848
rect 59412 38876 59418 38888
rect 60001 38879 60059 38885
rect 60001 38876 60013 38879
rect 59412 38848 60013 38876
rect 59412 38836 59418 38848
rect 60001 38845 60013 38848
rect 60047 38876 60059 38879
rect 61010 38876 61016 38888
rect 60047 38848 61016 38876
rect 60047 38845 60059 38848
rect 60001 38839 60059 38845
rect 61010 38836 61016 38848
rect 61068 38836 61074 38888
rect 61194 38836 61200 38888
rect 61252 38885 61258 38888
rect 61252 38879 61269 38885
rect 61257 38845 61269 38879
rect 61252 38839 61269 38845
rect 61381 38879 61439 38885
rect 61381 38845 61393 38879
rect 61427 38845 61439 38879
rect 61654 38876 61660 38888
rect 61615 38848 61660 38876
rect 61381 38839 61439 38845
rect 61252 38836 61258 38839
rect 59446 38808 59452 38820
rect 54536 38780 58848 38808
rect 58912 38780 59452 38808
rect 54536 38768 54542 38780
rect 54570 38740 54576 38752
rect 54404 38712 54576 38740
rect 54570 38700 54576 38712
rect 54628 38700 54634 38752
rect 56594 38700 56600 38752
rect 56652 38740 56658 38752
rect 58158 38740 58164 38752
rect 56652 38712 58164 38740
rect 56652 38700 56658 38712
rect 58158 38700 58164 38712
rect 58216 38700 58222 38752
rect 58820 38740 58848 38780
rect 59446 38768 59452 38780
rect 59504 38768 59510 38820
rect 59725 38811 59783 38817
rect 59725 38777 59737 38811
rect 59771 38808 59783 38811
rect 61396 38808 61424 38839
rect 61654 38836 61660 38848
rect 61712 38836 61718 38888
rect 61838 38876 61844 38888
rect 61799 38848 61844 38876
rect 61838 38836 61844 38848
rect 61896 38836 61902 38888
rect 65518 38876 65524 38888
rect 65479 38848 65524 38876
rect 65518 38836 65524 38848
rect 65576 38876 65582 38888
rect 65797 38879 65855 38885
rect 65797 38876 65809 38879
rect 65576 38848 65809 38876
rect 65576 38836 65582 38848
rect 65797 38845 65809 38848
rect 65843 38876 65855 38879
rect 66162 38876 66168 38888
rect 65843 38848 66168 38876
rect 65843 38845 65855 38848
rect 65797 38839 65855 38845
rect 66162 38836 66168 38848
rect 66220 38836 66226 38888
rect 69658 38876 69664 38888
rect 69619 38848 69664 38876
rect 69658 38836 69664 38848
rect 69716 38836 69722 38888
rect 70302 38836 70308 38888
rect 70360 38876 70366 38888
rect 71133 38879 71191 38885
rect 71133 38876 71145 38879
rect 70360 38848 71145 38876
rect 70360 38836 70366 38848
rect 71133 38845 71145 38848
rect 71179 38845 71191 38879
rect 71133 38839 71191 38845
rect 71317 38879 71375 38885
rect 71317 38845 71329 38879
rect 71363 38876 71375 38879
rect 71498 38876 71504 38888
rect 71363 38848 71504 38876
rect 71363 38845 71375 38848
rect 71317 38839 71375 38845
rect 71498 38836 71504 38848
rect 71556 38836 71562 38888
rect 59771 38780 61424 38808
rect 69676 38808 69704 38836
rect 71608 38808 71636 38907
rect 72418 38904 72424 38956
rect 72476 38944 72482 38956
rect 72513 38947 72571 38953
rect 72513 38944 72525 38947
rect 72476 38916 72525 38944
rect 72476 38904 72482 38916
rect 72513 38913 72525 38916
rect 72559 38944 72571 38947
rect 72559 38916 72924 38944
rect 72559 38913 72571 38916
rect 72513 38907 72571 38913
rect 71685 38879 71743 38885
rect 71685 38845 71697 38879
rect 71731 38876 71743 38879
rect 72326 38876 72332 38888
rect 71731 38848 72332 38876
rect 71731 38845 71743 38848
rect 71685 38839 71743 38845
rect 72326 38836 72332 38848
rect 72384 38836 72390 38888
rect 72896 38885 72924 38916
rect 74442 38904 74448 38956
rect 74500 38944 74506 38956
rect 74629 38947 74687 38953
rect 74629 38944 74641 38947
rect 74500 38916 74641 38944
rect 74500 38904 74506 38916
rect 74629 38913 74641 38916
rect 74675 38913 74687 38947
rect 74629 38907 74687 38913
rect 74718 38904 74724 38956
rect 74776 38944 74782 38956
rect 82354 38944 82360 38956
rect 74776 38916 82360 38944
rect 74776 38904 74782 38916
rect 82354 38904 82360 38916
rect 82412 38904 82418 38956
rect 82541 38947 82599 38953
rect 82541 38913 82553 38947
rect 82587 38944 82599 38947
rect 82722 38944 82728 38956
rect 82587 38916 82728 38944
rect 82587 38913 82599 38916
rect 82541 38907 82599 38913
rect 82722 38904 82728 38916
rect 82780 38904 82786 38956
rect 72881 38879 72939 38885
rect 72881 38845 72893 38879
rect 72927 38845 72939 38879
rect 72881 38839 72939 38845
rect 73062 38836 73068 38888
rect 73120 38876 73126 38888
rect 74169 38879 74227 38885
rect 74169 38876 74181 38879
rect 73120 38848 74181 38876
rect 73120 38836 73126 38848
rect 74169 38845 74181 38848
rect 74215 38845 74227 38879
rect 74169 38839 74227 38845
rect 74353 38879 74411 38885
rect 74353 38845 74365 38879
rect 74399 38876 74411 38879
rect 74902 38876 74908 38888
rect 74399 38848 74908 38876
rect 74399 38845 74411 38848
rect 74353 38839 74411 38845
rect 74902 38836 74908 38848
rect 74960 38836 74966 38888
rect 77021 38879 77079 38885
rect 77021 38845 77033 38879
rect 77067 38845 77079 38879
rect 77021 38839 77079 38845
rect 77297 38879 77355 38885
rect 77297 38845 77309 38879
rect 77343 38876 77355 38879
rect 79502 38876 79508 38888
rect 77343 38848 79508 38876
rect 77343 38845 77355 38848
rect 77297 38839 77355 38845
rect 69676 38780 71636 38808
rect 59771 38777 59783 38780
rect 59725 38771 59783 38777
rect 65426 38740 65432 38752
rect 58820 38712 65432 38740
rect 65426 38700 65432 38712
rect 65484 38740 65490 38752
rect 65613 38743 65671 38749
rect 65613 38740 65625 38743
rect 65484 38712 65625 38740
rect 65484 38700 65490 38712
rect 65613 38709 65625 38712
rect 65659 38709 65671 38743
rect 65613 38703 65671 38709
rect 67726 38700 67732 38752
rect 67784 38740 67790 38752
rect 69753 38743 69811 38749
rect 69753 38740 69765 38743
rect 67784 38712 69765 38740
rect 67784 38700 67790 38712
rect 69753 38709 69765 38712
rect 69799 38740 69811 38743
rect 70302 38740 70308 38752
rect 69799 38712 70308 38740
rect 69799 38709 69811 38712
rect 69753 38703 69811 38709
rect 70302 38700 70308 38712
rect 70360 38740 70366 38752
rect 70489 38743 70547 38749
rect 70489 38740 70501 38743
rect 70360 38712 70501 38740
rect 70360 38700 70366 38712
rect 70489 38709 70501 38712
rect 70535 38709 70547 38743
rect 70489 38703 70547 38709
rect 70949 38743 71007 38749
rect 70949 38709 70961 38743
rect 70995 38740 71007 38743
rect 72418 38740 72424 38752
rect 70995 38712 72424 38740
rect 70995 38709 71007 38712
rect 70949 38703 71007 38709
rect 72418 38700 72424 38712
rect 72476 38700 72482 38752
rect 72697 38743 72755 38749
rect 72697 38709 72709 38743
rect 72743 38740 72755 38743
rect 73982 38740 73988 38752
rect 72743 38712 73988 38740
rect 72743 38709 72755 38712
rect 72697 38703 72755 38709
rect 73982 38700 73988 38712
rect 74040 38700 74046 38752
rect 76929 38743 76987 38749
rect 76929 38709 76941 38743
rect 76975 38740 76987 38743
rect 77036 38740 77064 38839
rect 79502 38836 79508 38848
rect 79560 38836 79566 38888
rect 82449 38879 82507 38885
rect 82449 38845 82461 38879
rect 82495 38845 82507 38879
rect 82449 38839 82507 38845
rect 82909 38879 82967 38885
rect 82909 38845 82921 38879
rect 82955 38845 82967 38879
rect 83016 38876 83044 38984
rect 83182 38972 83188 39024
rect 83240 39012 83246 39024
rect 83553 39015 83611 39021
rect 83553 39012 83565 39015
rect 83240 38984 83565 39012
rect 83240 38972 83246 38984
rect 83553 38981 83565 38984
rect 83599 38981 83611 39015
rect 83936 39012 83964 39052
rect 84013 39049 84025 39052
rect 84059 39049 84071 39083
rect 84562 39080 84568 39092
rect 84523 39052 84568 39080
rect 84013 39043 84071 39049
rect 84562 39040 84568 39052
rect 84620 39040 84626 39092
rect 85666 39080 85672 39092
rect 85627 39052 85672 39080
rect 85666 39040 85672 39052
rect 85724 39040 85730 39092
rect 84194 39012 84200 39024
rect 83553 38975 83611 38981
rect 83660 38984 83964 39012
rect 84155 38984 84200 39012
rect 83366 38904 83372 38956
rect 83424 38944 83430 38956
rect 83660 38944 83688 38984
rect 84194 38972 84200 38984
rect 84252 38972 84258 39024
rect 83424 38916 83688 38944
rect 83424 38904 83430 38916
rect 83734 38904 83740 38956
rect 83792 38944 83798 38956
rect 83884 38947 83942 38953
rect 83884 38944 83896 38947
rect 83792 38916 83896 38944
rect 83792 38904 83798 38916
rect 83884 38913 83896 38916
rect 83930 38913 83942 38947
rect 84102 38944 84108 38956
rect 84063 38916 84108 38944
rect 83884 38907 83942 38913
rect 84102 38904 84108 38916
rect 84160 38904 84166 38956
rect 83016 38848 83504 38876
rect 82909 38839 82967 38845
rect 82464 38808 82492 38839
rect 82814 38808 82820 38820
rect 82464 38780 82820 38808
rect 82814 38768 82820 38780
rect 82872 38768 82878 38820
rect 82924 38808 82952 38839
rect 83366 38808 83372 38820
rect 82924 38780 83372 38808
rect 77294 38740 77300 38752
rect 76975 38712 77300 38740
rect 76975 38709 76987 38712
rect 76929 38703 76987 38709
rect 77294 38700 77300 38712
rect 77352 38700 77358 38752
rect 77386 38700 77392 38752
rect 77444 38740 77450 38752
rect 78401 38743 78459 38749
rect 78401 38740 78413 38743
rect 77444 38712 78413 38740
rect 77444 38700 77450 38712
rect 78401 38709 78413 38712
rect 78447 38709 78459 38743
rect 78401 38703 78459 38709
rect 81526 38700 81532 38752
rect 81584 38740 81590 38752
rect 81989 38743 82047 38749
rect 81989 38740 82001 38743
rect 81584 38712 82001 38740
rect 81584 38700 81590 38712
rect 81989 38709 82001 38712
rect 82035 38740 82047 38743
rect 82924 38740 82952 38780
rect 83366 38768 83372 38780
rect 83424 38768 83430 38820
rect 82035 38712 82952 38740
rect 83476 38740 83504 38848
rect 84562 38836 84568 38888
rect 84620 38876 84626 38888
rect 85577 38879 85635 38885
rect 85577 38876 85589 38879
rect 84620 38848 85589 38876
rect 84620 38836 84626 38848
rect 85577 38845 85589 38848
rect 85623 38876 85635 38879
rect 86037 38879 86095 38885
rect 86037 38876 86049 38879
rect 85623 38848 86049 38876
rect 85623 38845 85635 38848
rect 85577 38839 85635 38845
rect 86037 38845 86049 38848
rect 86083 38845 86095 38879
rect 86862 38876 86868 38888
rect 86823 38848 86868 38876
rect 86037 38839 86095 38845
rect 86862 38836 86868 38848
rect 86920 38836 86926 38888
rect 86954 38836 86960 38888
rect 87012 38876 87018 38888
rect 87141 38879 87199 38885
rect 87012 38848 87057 38876
rect 87012 38836 87018 38848
rect 87141 38845 87153 38879
rect 87187 38876 87199 38879
rect 89070 38876 89076 38888
rect 87187 38848 89076 38876
rect 87187 38845 87199 38848
rect 87141 38839 87199 38845
rect 89070 38836 89076 38848
rect 89128 38836 89134 38888
rect 91554 38876 91560 38888
rect 91515 38848 91560 38876
rect 91554 38836 91560 38848
rect 91612 38836 91618 38888
rect 92845 38879 92903 38885
rect 92845 38845 92857 38879
rect 92891 38845 92903 38879
rect 92845 38839 92903 38845
rect 83737 38811 83795 38817
rect 83737 38777 83749 38811
rect 83783 38808 83795 38811
rect 84838 38808 84844 38820
rect 83783 38780 84844 38808
rect 83783 38777 83795 38780
rect 83737 38771 83795 38777
rect 84838 38768 84844 38780
rect 84896 38808 84902 38820
rect 85393 38811 85451 38817
rect 85393 38808 85405 38811
rect 84896 38780 85405 38808
rect 84896 38768 84902 38780
rect 85393 38777 85405 38780
rect 85439 38808 85451 38811
rect 89898 38808 89904 38820
rect 85439 38780 89904 38808
rect 85439 38777 85451 38780
rect 85393 38771 85451 38777
rect 89898 38768 89904 38780
rect 89956 38768 89962 38820
rect 91094 38768 91100 38820
rect 91152 38808 91158 38820
rect 91649 38811 91707 38817
rect 91649 38808 91661 38811
rect 91152 38780 91661 38808
rect 91152 38768 91158 38780
rect 91649 38777 91661 38780
rect 91695 38808 91707 38811
rect 92661 38811 92719 38817
rect 92661 38808 92673 38811
rect 91695 38780 92673 38808
rect 91695 38777 91707 38780
rect 91649 38771 91707 38777
rect 92661 38777 92673 38780
rect 92707 38777 92719 38811
rect 92661 38771 92719 38777
rect 87325 38743 87383 38749
rect 87325 38740 87337 38743
rect 83476 38712 87337 38740
rect 82035 38709 82047 38712
rect 81989 38703 82047 38709
rect 87325 38709 87337 38712
rect 87371 38709 87383 38743
rect 92860 38740 92888 38839
rect 93213 38811 93271 38817
rect 93213 38777 93225 38811
rect 93259 38808 93271 38811
rect 93486 38808 93492 38820
rect 93259 38780 93492 38808
rect 93259 38777 93271 38780
rect 93213 38771 93271 38777
rect 93486 38768 93492 38780
rect 93544 38768 93550 38820
rect 93394 38740 93400 38752
rect 92860 38712 93400 38740
rect 87325 38703 87383 38709
rect 93394 38700 93400 38712
rect 93452 38700 93458 38752
rect 1104 38650 105616 38672
rect 1104 38598 19606 38650
rect 19658 38598 19670 38650
rect 19722 38598 19734 38650
rect 19786 38598 19798 38650
rect 19850 38598 50326 38650
rect 50378 38598 50390 38650
rect 50442 38598 50454 38650
rect 50506 38598 50518 38650
rect 50570 38598 81046 38650
rect 81098 38598 81110 38650
rect 81162 38598 81174 38650
rect 81226 38598 81238 38650
rect 81290 38598 105616 38650
rect 1104 38576 105616 38598
rect 2774 38496 2780 38548
rect 2832 38536 2838 38548
rect 4157 38539 4215 38545
rect 4157 38536 4169 38539
rect 2832 38508 4169 38536
rect 2832 38496 2838 38508
rect 4157 38505 4169 38508
rect 4203 38505 4215 38539
rect 4157 38499 4215 38505
rect 4985 38539 5043 38545
rect 4985 38505 4997 38539
rect 5031 38536 5043 38539
rect 5074 38536 5080 38548
rect 5031 38508 5080 38536
rect 5031 38505 5043 38508
rect 4985 38499 5043 38505
rect 4798 38468 4804 38480
rect 4356 38440 4804 38468
rect 4356 38409 4384 38440
rect 4798 38428 4804 38440
rect 4856 38428 4862 38480
rect 4341 38403 4399 38409
rect 4341 38369 4353 38403
rect 4387 38369 4399 38403
rect 4341 38363 4399 38369
rect 4617 38403 4675 38409
rect 4617 38369 4629 38403
rect 4663 38400 4675 38403
rect 5000 38400 5028 38499
rect 5074 38496 5080 38508
rect 5132 38496 5138 38548
rect 8478 38496 8484 38548
rect 8536 38536 8542 38548
rect 8665 38539 8723 38545
rect 8665 38536 8677 38539
rect 8536 38508 8677 38536
rect 8536 38496 8542 38508
rect 8665 38505 8677 38508
rect 8711 38505 8723 38539
rect 8665 38499 8723 38505
rect 11974 38496 11980 38548
rect 12032 38536 12038 38548
rect 13538 38536 13544 38548
rect 12032 38508 13544 38536
rect 12032 38496 12038 38508
rect 13538 38496 13544 38508
rect 13596 38496 13602 38548
rect 20530 38536 20536 38548
rect 17236 38508 20536 38536
rect 17236 38468 17264 38508
rect 20530 38496 20536 38508
rect 20588 38496 20594 38548
rect 21174 38496 21180 38548
rect 21232 38536 21238 38548
rect 22097 38539 22155 38545
rect 22097 38536 22109 38539
rect 21232 38508 22109 38536
rect 21232 38496 21238 38508
rect 22097 38505 22109 38508
rect 22143 38505 22155 38539
rect 22097 38499 22155 38505
rect 22186 38496 22192 38548
rect 22244 38536 22250 38548
rect 31478 38536 31484 38548
rect 22244 38508 31484 38536
rect 22244 38496 22250 38508
rect 31478 38496 31484 38508
rect 31536 38496 31542 38548
rect 31941 38539 31999 38545
rect 31941 38505 31953 38539
rect 31987 38536 31999 38539
rect 42886 38536 42892 38548
rect 31987 38508 42892 38536
rect 31987 38505 31999 38508
rect 31941 38499 31999 38505
rect 42886 38496 42892 38508
rect 42944 38496 42950 38548
rect 48314 38496 48320 38548
rect 48372 38536 48378 38548
rect 61102 38536 61108 38548
rect 48372 38508 61108 38536
rect 48372 38496 48378 38508
rect 61102 38496 61108 38508
rect 61160 38496 61166 38548
rect 61286 38496 61292 38548
rect 61344 38536 61350 38548
rect 70762 38536 70768 38548
rect 61344 38508 70768 38536
rect 61344 38496 61350 38508
rect 70762 38496 70768 38508
rect 70820 38496 70826 38548
rect 70872 38508 71176 38536
rect 4663 38372 5028 38400
rect 5092 38440 17264 38468
rect 18509 38471 18567 38477
rect 4663 38369 4675 38372
rect 4617 38363 4675 38369
rect 4062 38292 4068 38344
rect 4120 38332 4126 38344
rect 5092 38332 5120 38440
rect 18509 38437 18521 38471
rect 18555 38468 18567 38471
rect 18690 38468 18696 38480
rect 18555 38440 18696 38468
rect 18555 38437 18567 38440
rect 18509 38431 18567 38437
rect 18690 38428 18696 38440
rect 18748 38468 18754 38480
rect 19889 38471 19947 38477
rect 18748 38440 19748 38468
rect 18748 38428 18754 38440
rect 7377 38403 7435 38409
rect 7377 38369 7389 38403
rect 7423 38369 7435 38403
rect 7377 38363 7435 38369
rect 8481 38403 8539 38409
rect 8481 38369 8493 38403
rect 8527 38400 8539 38403
rect 8570 38400 8576 38412
rect 8527 38372 8576 38400
rect 8527 38369 8539 38372
rect 8481 38363 8539 38369
rect 4120 38304 5120 38332
rect 7392 38332 7420 38363
rect 8570 38360 8576 38372
rect 8628 38360 8634 38412
rect 11425 38403 11483 38409
rect 9692 38372 11376 38400
rect 9582 38332 9588 38344
rect 7392 38304 9588 38332
rect 4120 38292 4126 38304
rect 9582 38292 9588 38304
rect 9640 38292 9646 38344
rect 3786 38224 3792 38276
rect 3844 38264 3850 38276
rect 9692 38264 9720 38372
rect 11241 38335 11299 38341
rect 11241 38332 11253 38335
rect 3844 38236 9720 38264
rect 11072 38304 11253 38332
rect 3844 38224 3850 38236
rect 7561 38199 7619 38205
rect 7561 38165 7573 38199
rect 7607 38196 7619 38199
rect 8202 38196 8208 38208
rect 7607 38168 8208 38196
rect 7607 38165 7619 38168
rect 7561 38159 7619 38165
rect 8202 38156 8208 38168
rect 8260 38156 8266 38208
rect 9950 38156 9956 38208
rect 10008 38196 10014 38208
rect 11072 38205 11100 38304
rect 11241 38301 11253 38304
rect 11287 38301 11299 38335
rect 11241 38295 11299 38301
rect 11348 38264 11376 38372
rect 11425 38369 11437 38403
rect 11471 38400 11483 38403
rect 11974 38400 11980 38412
rect 11471 38372 11980 38400
rect 11471 38369 11483 38372
rect 11425 38363 11483 38369
rect 11974 38360 11980 38372
rect 12032 38360 12038 38412
rect 12158 38400 12164 38412
rect 12119 38372 12164 38400
rect 12158 38360 12164 38372
rect 12216 38400 12222 38412
rect 13449 38403 13507 38409
rect 12216 38372 12388 38400
rect 12216 38360 12222 38372
rect 12360 38332 12388 38372
rect 13449 38369 13461 38403
rect 13495 38400 13507 38403
rect 14090 38400 14096 38412
rect 13495 38372 14096 38400
rect 13495 38369 13507 38372
rect 13449 38363 13507 38369
rect 14090 38360 14096 38372
rect 14148 38360 14154 38412
rect 18782 38400 18788 38412
rect 18743 38372 18788 38400
rect 18782 38360 18788 38372
rect 18840 38360 18846 38412
rect 18892 38409 18920 38440
rect 18877 38403 18935 38409
rect 18877 38369 18889 38403
rect 18923 38369 18935 38403
rect 18877 38363 18935 38369
rect 19334 38360 19340 38412
rect 19392 38409 19398 38412
rect 19392 38403 19441 38409
rect 19392 38369 19395 38403
rect 19429 38369 19441 38403
rect 19392 38363 19441 38369
rect 19392 38360 19398 38363
rect 19518 38360 19524 38412
rect 19576 38400 19582 38412
rect 19720 38400 19748 38440
rect 19889 38437 19901 38471
rect 19935 38468 19947 38471
rect 19978 38468 19984 38480
rect 19935 38440 19984 38468
rect 19935 38437 19947 38440
rect 19889 38431 19947 38437
rect 19978 38428 19984 38440
rect 20036 38428 20042 38480
rect 20165 38471 20223 38477
rect 20165 38437 20177 38471
rect 20211 38468 20223 38471
rect 20257 38471 20315 38477
rect 20257 38468 20269 38471
rect 20211 38440 20269 38468
rect 20211 38437 20223 38440
rect 20165 38431 20223 38437
rect 20257 38437 20269 38440
rect 20303 38468 20315 38471
rect 20990 38468 20996 38480
rect 20303 38440 20996 38468
rect 20303 38437 20315 38440
rect 20257 38431 20315 38437
rect 20990 38428 20996 38440
rect 21048 38428 21054 38480
rect 25406 38468 25412 38480
rect 21652 38440 25412 38468
rect 21082 38400 21088 38412
rect 19576 38372 19621 38400
rect 19720 38372 20760 38400
rect 21043 38372 21088 38400
rect 19576 38360 19582 38372
rect 20732 38341 20760 38372
rect 21082 38360 21088 38372
rect 21140 38360 21146 38412
rect 21652 38409 21680 38440
rect 25406 38428 25412 38440
rect 25464 38468 25470 38480
rect 27798 38468 27804 38480
rect 25464 38440 27804 38468
rect 25464 38428 25470 38440
rect 27798 38428 27804 38440
rect 27856 38428 27862 38480
rect 28810 38428 28816 38480
rect 28868 38468 28874 38480
rect 42978 38468 42984 38480
rect 28868 38440 42984 38468
rect 28868 38428 28874 38440
rect 42978 38428 42984 38440
rect 43036 38428 43042 38480
rect 51442 38468 51448 38480
rect 44376 38440 51448 38468
rect 21637 38403 21695 38409
rect 21637 38369 21649 38403
rect 21683 38369 21695 38403
rect 21637 38363 21695 38369
rect 21726 38360 21732 38412
rect 21784 38400 21790 38412
rect 21821 38403 21879 38409
rect 21821 38400 21833 38403
rect 21784 38372 21833 38400
rect 21784 38360 21790 38372
rect 21821 38369 21833 38372
rect 21867 38369 21879 38403
rect 21821 38363 21879 38369
rect 22002 38360 22008 38412
rect 22060 38400 22066 38412
rect 24302 38400 24308 38412
rect 22060 38372 24308 38400
rect 22060 38360 22066 38372
rect 24302 38360 24308 38372
rect 24360 38400 24366 38412
rect 25590 38400 25596 38412
rect 24360 38372 25596 38400
rect 24360 38360 24366 38372
rect 25590 38360 25596 38372
rect 25648 38360 25654 38412
rect 27890 38400 27896 38412
rect 27851 38372 27896 38400
rect 27890 38360 27896 38372
rect 27948 38400 27954 38412
rect 28445 38403 28503 38409
rect 28445 38400 28457 38403
rect 27948 38372 28457 38400
rect 27948 38360 27954 38372
rect 28445 38369 28457 38372
rect 28491 38369 28503 38403
rect 28626 38400 28632 38412
rect 28539 38372 28632 38400
rect 28445 38363 28503 38369
rect 28626 38360 28632 38372
rect 28684 38400 28690 38412
rect 29273 38403 29331 38409
rect 29273 38400 29285 38403
rect 28684 38372 29285 38400
rect 28684 38360 28690 38372
rect 29273 38369 29285 38372
rect 29319 38400 29331 38403
rect 31941 38403 31999 38409
rect 31941 38400 31953 38403
rect 29319 38372 31953 38400
rect 29319 38369 29331 38372
rect 29273 38363 29331 38369
rect 31941 38369 31953 38372
rect 31987 38369 31999 38403
rect 32858 38400 32864 38412
rect 32819 38372 32864 38400
rect 31941 38363 31999 38369
rect 32858 38360 32864 38372
rect 32916 38360 32922 38412
rect 39025 38403 39083 38409
rect 39025 38369 39037 38403
rect 39071 38400 39083 38403
rect 39114 38400 39120 38412
rect 39071 38372 39120 38400
rect 39071 38369 39083 38372
rect 39025 38363 39083 38369
rect 39114 38360 39120 38372
rect 39172 38360 39178 38412
rect 39206 38360 39212 38412
rect 39264 38400 39270 38412
rect 39485 38403 39543 38409
rect 39485 38400 39497 38403
rect 39264 38372 39497 38400
rect 39264 38360 39270 38372
rect 39485 38369 39497 38372
rect 39531 38369 39543 38403
rect 39485 38363 39543 38369
rect 39577 38403 39635 38409
rect 39577 38369 39589 38403
rect 39623 38400 39635 38403
rect 39942 38400 39948 38412
rect 39623 38372 39948 38400
rect 39623 38369 39635 38372
rect 39577 38363 39635 38369
rect 39942 38360 39948 38372
rect 40000 38400 40006 38412
rect 40313 38403 40371 38409
rect 40313 38400 40325 38403
rect 40000 38372 40325 38400
rect 40000 38360 40006 38372
rect 40313 38369 40325 38372
rect 40359 38369 40371 38403
rect 40586 38400 40592 38412
rect 40313 38363 40371 38369
rect 40420 38372 40592 38400
rect 13541 38335 13599 38341
rect 13541 38332 13553 38335
rect 12360 38304 13553 38332
rect 13541 38301 13553 38304
rect 13587 38301 13599 38335
rect 13541 38295 13599 38301
rect 20717 38335 20775 38341
rect 20717 38301 20729 38335
rect 20763 38332 20775 38335
rect 20901 38335 20959 38341
rect 20901 38332 20913 38335
rect 20763 38304 20913 38332
rect 20763 38301 20775 38304
rect 20717 38295 20775 38301
rect 20901 38301 20913 38304
rect 20947 38301 20959 38335
rect 20901 38295 20959 38301
rect 27338 38292 27344 38344
rect 27396 38332 27402 38344
rect 27709 38335 27767 38341
rect 27709 38332 27721 38335
rect 27396 38304 27721 38332
rect 27396 38292 27402 38304
rect 27709 38301 27721 38304
rect 27755 38301 27767 38335
rect 33226 38332 33232 38344
rect 33187 38304 33232 38332
rect 27709 38295 27767 38301
rect 33226 38292 33232 38304
rect 33284 38292 33290 38344
rect 38930 38332 38936 38344
rect 38891 38304 38936 38332
rect 38930 38292 38936 38304
rect 38988 38292 38994 38344
rect 40129 38335 40187 38341
rect 40129 38301 40141 38335
rect 40175 38332 40187 38335
rect 40420 38332 40448 38372
rect 40586 38360 40592 38372
rect 40644 38360 40650 38412
rect 40175 38304 40448 38332
rect 40175 38301 40187 38304
rect 40129 38295 40187 38301
rect 40494 38292 40500 38344
rect 40552 38332 40558 38344
rect 44269 38335 44327 38341
rect 44269 38332 44281 38335
rect 40552 38304 44281 38332
rect 40552 38292 40558 38304
rect 44269 38301 44281 38304
rect 44315 38301 44327 38335
rect 44269 38295 44327 38301
rect 24486 38264 24492 38276
rect 11348 38236 24492 38264
rect 24486 38224 24492 38236
rect 24544 38224 24550 38276
rect 24854 38224 24860 38276
rect 24912 38264 24918 38276
rect 32766 38264 32772 38276
rect 24912 38236 32772 38264
rect 24912 38224 24918 38236
rect 32766 38224 32772 38236
rect 32824 38224 32830 38276
rect 33026 38267 33084 38273
rect 33026 38233 33038 38267
rect 33072 38264 33084 38267
rect 33318 38264 33324 38276
rect 33072 38236 33324 38264
rect 33072 38233 33084 38236
rect 33026 38227 33084 38233
rect 33318 38224 33324 38236
rect 33376 38224 33382 38276
rect 33505 38267 33563 38273
rect 33505 38233 33517 38267
rect 33551 38264 33563 38267
rect 44376 38264 44404 38440
rect 51442 38428 51448 38440
rect 51500 38428 51506 38480
rect 52454 38428 52460 38480
rect 52512 38468 52518 38480
rect 52917 38471 52975 38477
rect 52917 38468 52929 38471
rect 52512 38440 52929 38468
rect 52512 38428 52518 38440
rect 52917 38437 52929 38440
rect 52963 38437 52975 38471
rect 56686 38468 56692 38480
rect 52917 38431 52975 38437
rect 56520 38440 56692 38468
rect 44453 38403 44511 38409
rect 44453 38369 44465 38403
rect 44499 38400 44511 38403
rect 44910 38400 44916 38412
rect 44499 38372 44680 38400
rect 44871 38372 44916 38400
rect 44499 38369 44511 38372
rect 44453 38363 44511 38369
rect 33551 38236 44404 38264
rect 44652 38264 44680 38372
rect 44910 38360 44916 38372
rect 44968 38360 44974 38412
rect 45005 38403 45063 38409
rect 45005 38369 45017 38403
rect 45051 38400 45063 38403
rect 45370 38400 45376 38412
rect 45051 38372 45376 38400
rect 45051 38369 45063 38372
rect 45005 38363 45063 38369
rect 45370 38360 45376 38372
rect 45428 38400 45434 38412
rect 45833 38403 45891 38409
rect 45833 38400 45845 38403
rect 45428 38372 45845 38400
rect 45428 38360 45434 38372
rect 45833 38369 45845 38372
rect 45879 38400 45891 38403
rect 50062 38400 50068 38412
rect 45879 38372 50068 38400
rect 45879 38369 45891 38372
rect 45833 38363 45891 38369
rect 50062 38360 50068 38372
rect 50120 38360 50126 38412
rect 50338 38400 50344 38412
rect 50299 38372 50344 38400
rect 50338 38360 50344 38372
rect 50396 38360 50402 38412
rect 50801 38403 50859 38409
rect 50801 38400 50813 38403
rect 50448 38372 50813 38400
rect 45465 38335 45523 38341
rect 45465 38301 45477 38335
rect 45511 38332 45523 38335
rect 46750 38332 46756 38344
rect 45511 38304 46756 38332
rect 45511 38301 45523 38304
rect 45465 38295 45523 38301
rect 46750 38292 46756 38304
rect 46808 38292 46814 38344
rect 49878 38332 49884 38344
rect 46860 38304 49884 38332
rect 44652 38236 45600 38264
rect 33551 38233 33563 38236
rect 33505 38227 33563 38233
rect 11057 38199 11115 38205
rect 11057 38196 11069 38199
rect 10008 38168 11069 38196
rect 10008 38156 10014 38168
rect 11057 38165 11069 38168
rect 11103 38165 11115 38199
rect 11057 38159 11115 38165
rect 12437 38199 12495 38205
rect 12437 38165 12449 38199
rect 12483 38196 12495 38199
rect 12710 38196 12716 38208
rect 12483 38168 12716 38196
rect 12483 38165 12495 38168
rect 12437 38159 12495 38165
rect 12710 38156 12716 38168
rect 12768 38156 12774 38208
rect 13817 38199 13875 38205
rect 13817 38165 13829 38199
rect 13863 38196 13875 38199
rect 14090 38196 14096 38208
rect 13863 38168 14096 38196
rect 13863 38165 13875 38168
rect 13817 38159 13875 38165
rect 14090 38156 14096 38168
rect 14148 38156 14154 38208
rect 16022 38156 16028 38208
rect 16080 38196 16086 38208
rect 19518 38196 19524 38208
rect 16080 38168 19524 38196
rect 16080 38156 16086 38168
rect 19518 38156 19524 38168
rect 19576 38196 19582 38208
rect 20257 38199 20315 38205
rect 20257 38196 20269 38199
rect 19576 38168 20269 38196
rect 19576 38156 19582 38168
rect 20257 38165 20269 38168
rect 20303 38165 20315 38199
rect 20257 38159 20315 38165
rect 20346 38156 20352 38208
rect 20404 38196 20410 38208
rect 20441 38199 20499 38205
rect 20441 38196 20453 38199
rect 20404 38168 20453 38196
rect 20404 38156 20410 38168
rect 20441 38165 20453 38168
rect 20487 38165 20499 38199
rect 20441 38159 20499 38165
rect 20530 38156 20536 38208
rect 20588 38196 20594 38208
rect 24026 38196 24032 38208
rect 20588 38168 24032 38196
rect 20588 38156 20594 38168
rect 24026 38156 24032 38168
rect 24084 38156 24090 38208
rect 26234 38156 26240 38208
rect 26292 38196 26298 38208
rect 27154 38196 27160 38208
rect 26292 38168 27160 38196
rect 26292 38156 26298 38168
rect 27154 38156 27160 38168
rect 27212 38156 27218 38208
rect 27338 38156 27344 38208
rect 27396 38196 27402 38208
rect 27525 38199 27583 38205
rect 27525 38196 27537 38199
rect 27396 38168 27537 38196
rect 27396 38156 27402 38168
rect 27525 38165 27537 38168
rect 27571 38165 27583 38199
rect 28902 38196 28908 38208
rect 28863 38168 28908 38196
rect 27525 38159 27583 38165
rect 28902 38156 28908 38168
rect 28960 38156 28966 38208
rect 33134 38196 33140 38208
rect 33095 38168 33140 38196
rect 33134 38156 33140 38168
rect 33192 38156 33198 38208
rect 39114 38156 39120 38208
rect 39172 38196 39178 38208
rect 40497 38199 40555 38205
rect 40497 38196 40509 38199
rect 39172 38168 40509 38196
rect 39172 38156 39178 38168
rect 40497 38165 40509 38168
rect 40543 38196 40555 38199
rect 40862 38196 40868 38208
rect 40543 38168 40868 38196
rect 40543 38165 40555 38168
rect 40497 38159 40555 38165
rect 40862 38156 40868 38168
rect 40920 38156 40926 38208
rect 44082 38156 44088 38208
rect 44140 38196 44146 38208
rect 44652 38196 44680 38236
rect 45572 38208 45600 38236
rect 44140 38168 44680 38196
rect 44140 38156 44146 38168
rect 45554 38156 45560 38208
rect 45612 38196 45618 38208
rect 46017 38199 46075 38205
rect 46017 38196 46029 38199
rect 45612 38168 46029 38196
rect 45612 38156 45618 38168
rect 46017 38165 46029 38168
rect 46063 38196 46075 38199
rect 46860 38196 46888 38304
rect 49878 38292 49884 38304
rect 49936 38292 49942 38344
rect 50246 38332 50252 38344
rect 50207 38304 50252 38332
rect 50246 38292 50252 38304
rect 50304 38292 50310 38344
rect 49786 38264 49792 38276
rect 49747 38236 49792 38264
rect 49786 38224 49792 38236
rect 49844 38264 49850 38276
rect 50448 38264 50476 38372
rect 50801 38369 50813 38372
rect 50847 38369 50859 38403
rect 50801 38363 50859 38369
rect 50893 38403 50951 38409
rect 50893 38369 50905 38403
rect 50939 38400 50951 38403
rect 53064 38403 53122 38409
rect 50939 38372 51764 38400
rect 50939 38369 50951 38372
rect 50893 38363 50951 38369
rect 51736 38341 51764 38372
rect 53064 38369 53076 38403
rect 53110 38400 53122 38403
rect 56520 38400 56548 38440
rect 56686 38428 56692 38440
rect 56744 38428 56750 38480
rect 60844 38440 63724 38468
rect 53110 38372 56548 38400
rect 53110 38369 53122 38372
rect 53064 38363 53122 38369
rect 56594 38360 56600 38412
rect 56652 38400 56658 38412
rect 56652 38372 56697 38400
rect 56796 38372 58112 38400
rect 56652 38360 56658 38372
rect 51721 38335 51779 38341
rect 51721 38301 51733 38335
rect 51767 38332 51779 38335
rect 52454 38332 52460 38344
rect 51767 38304 52460 38332
rect 51767 38301 51779 38304
rect 51721 38295 51779 38301
rect 52454 38292 52460 38304
rect 52512 38292 52518 38344
rect 53285 38335 53343 38341
rect 53285 38301 53297 38335
rect 53331 38301 53343 38335
rect 53285 38295 53343 38301
rect 49844 38236 50476 38264
rect 53300 38264 53328 38295
rect 56226 38292 56232 38344
rect 56284 38332 56290 38344
rect 56796 38332 56824 38372
rect 56284 38304 56824 38332
rect 56284 38292 56290 38304
rect 57422 38292 57428 38344
rect 57480 38332 57486 38344
rect 57609 38335 57667 38341
rect 57609 38332 57621 38335
rect 57480 38304 57621 38332
rect 57480 38292 57486 38304
rect 57609 38301 57621 38304
rect 57655 38301 57667 38335
rect 57609 38295 57667 38301
rect 57885 38335 57943 38341
rect 57885 38301 57897 38335
rect 57931 38332 57943 38335
rect 57974 38332 57980 38344
rect 57931 38304 57980 38332
rect 57931 38301 57943 38304
rect 57885 38295 57943 38301
rect 57974 38292 57980 38304
rect 58032 38292 58038 38344
rect 58084 38332 58112 38372
rect 58158 38360 58164 38412
rect 58216 38400 58222 38412
rect 58986 38400 58992 38412
rect 58216 38372 58992 38400
rect 58216 38360 58222 38372
rect 58986 38360 58992 38372
rect 59044 38360 59050 38412
rect 59722 38360 59728 38412
rect 59780 38400 59786 38412
rect 60844 38400 60872 38440
rect 59780 38372 60872 38400
rect 59780 38360 59786 38372
rect 62850 38360 62856 38412
rect 62908 38400 62914 38412
rect 63405 38403 63463 38409
rect 63405 38400 63417 38403
rect 62908 38372 63417 38400
rect 62908 38360 62914 38372
rect 63405 38369 63417 38372
rect 63451 38369 63463 38403
rect 63405 38363 63463 38369
rect 63494 38360 63500 38412
rect 63552 38400 63558 38412
rect 63589 38403 63647 38409
rect 63589 38400 63601 38403
rect 63552 38372 63601 38400
rect 63552 38360 63558 38372
rect 63589 38369 63601 38372
rect 63635 38369 63647 38403
rect 63696 38400 63724 38440
rect 63770 38428 63776 38480
rect 63828 38468 63834 38480
rect 67726 38468 67732 38480
rect 63828 38440 67732 38468
rect 63828 38428 63834 38440
rect 67726 38428 67732 38440
rect 67784 38428 67790 38480
rect 69293 38471 69351 38477
rect 69293 38437 69305 38471
rect 69339 38468 69351 38471
rect 69658 38468 69664 38480
rect 69339 38440 69664 38468
rect 69339 38437 69351 38440
rect 69293 38431 69351 38437
rect 69658 38428 69664 38440
rect 69716 38428 69722 38480
rect 70118 38468 70124 38480
rect 70079 38440 70124 38468
rect 70118 38428 70124 38440
rect 70176 38468 70182 38480
rect 70176 38440 70348 38468
rect 70176 38428 70182 38440
rect 70320 38409 70348 38440
rect 70305 38403 70363 38409
rect 63696 38372 68600 38400
rect 63589 38363 63647 38369
rect 59078 38332 59084 38344
rect 58084 38304 59084 38332
rect 59078 38292 59084 38304
rect 59136 38292 59142 38344
rect 62669 38335 62727 38341
rect 62669 38332 62681 38335
rect 62592 38304 62681 38332
rect 53837 38267 53895 38273
rect 53837 38264 53849 38267
rect 53300 38236 53849 38264
rect 49844 38224 49850 38236
rect 53837 38233 53849 38236
rect 53883 38264 53895 38267
rect 53883 38236 57560 38264
rect 53883 38233 53895 38236
rect 53837 38227 53895 38233
rect 46063 38168 46888 38196
rect 46063 38165 46075 38168
rect 46017 38159 46075 38165
rect 48314 38156 48320 38208
rect 48372 38196 48378 38208
rect 49973 38199 50031 38205
rect 49973 38196 49985 38199
rect 48372 38168 49985 38196
rect 48372 38156 48378 38168
rect 49973 38165 49985 38168
rect 50019 38196 50031 38199
rect 50246 38196 50252 38208
rect 50019 38168 50252 38196
rect 50019 38165 50031 38168
rect 49973 38159 50031 38165
rect 50246 38156 50252 38168
rect 50304 38156 50310 38208
rect 51353 38199 51411 38205
rect 51353 38165 51365 38199
rect 51399 38196 51411 38199
rect 51442 38196 51448 38208
rect 51399 38168 51448 38196
rect 51399 38165 51411 38168
rect 51353 38159 51411 38165
rect 51442 38156 51448 38168
rect 51500 38156 51506 38208
rect 53190 38196 53196 38208
rect 53151 38168 53196 38196
rect 53190 38156 53196 38168
rect 53248 38156 53254 38208
rect 53282 38156 53288 38208
rect 53340 38196 53346 38208
rect 53377 38199 53435 38205
rect 53377 38196 53389 38199
rect 53340 38168 53389 38196
rect 53340 38156 53346 38168
rect 53377 38165 53389 38168
rect 53423 38165 53435 38199
rect 56686 38196 56692 38208
rect 56647 38168 56692 38196
rect 53377 38159 53435 38165
rect 56686 38156 56692 38168
rect 56744 38156 56750 38208
rect 57422 38196 57428 38208
rect 57383 38168 57428 38196
rect 57422 38156 57428 38168
rect 57480 38156 57486 38208
rect 57532 38196 57560 38236
rect 62592 38208 62620 38304
rect 62669 38301 62681 38304
rect 62715 38301 62727 38335
rect 67637 38335 67695 38341
rect 67637 38332 67649 38335
rect 62669 38295 62727 38301
rect 67284 38304 67649 38332
rect 61930 38196 61936 38208
rect 57532 38168 61936 38196
rect 61930 38156 61936 38168
rect 61988 38156 61994 38208
rect 62114 38196 62120 38208
rect 62075 38168 62120 38196
rect 62114 38156 62120 38168
rect 62172 38196 62178 38208
rect 62301 38199 62359 38205
rect 62301 38196 62313 38199
rect 62172 38168 62313 38196
rect 62172 38156 62178 38168
rect 62301 38165 62313 38168
rect 62347 38165 62359 38199
rect 62574 38196 62580 38208
rect 62535 38168 62580 38196
rect 62301 38159 62359 38165
rect 62574 38156 62580 38168
rect 62632 38156 62638 38208
rect 63865 38199 63923 38205
rect 63865 38165 63877 38199
rect 63911 38196 63923 38199
rect 64690 38196 64696 38208
rect 63911 38168 64696 38196
rect 63911 38165 63923 38168
rect 63865 38159 63923 38165
rect 64690 38156 64696 38168
rect 64748 38156 64754 38208
rect 65334 38156 65340 38208
rect 65392 38196 65398 38208
rect 67284 38205 67312 38304
rect 67637 38301 67649 38304
rect 67683 38301 67695 38335
rect 67637 38295 67695 38301
rect 67818 38292 67824 38344
rect 67876 38332 67882 38344
rect 67913 38335 67971 38341
rect 67913 38332 67925 38335
rect 67876 38304 67925 38332
rect 67876 38292 67882 38304
rect 67913 38301 67925 38304
rect 67959 38301 67971 38335
rect 67913 38295 67971 38301
rect 67358 38224 67364 38276
rect 67416 38264 67422 38276
rect 68572 38264 68600 38372
rect 70305 38369 70317 38403
rect 70351 38400 70363 38403
rect 70872 38400 70900 38508
rect 71148 38477 71176 38508
rect 71222 38496 71228 38548
rect 71280 38536 71286 38548
rect 77570 38536 77576 38548
rect 71280 38508 77576 38536
rect 71280 38496 71286 38508
rect 77570 38496 77576 38508
rect 77628 38496 77634 38548
rect 84010 38496 84016 38548
rect 84068 38536 84074 38548
rect 84657 38539 84715 38545
rect 84657 38536 84669 38539
rect 84068 38508 84669 38536
rect 84068 38496 84074 38508
rect 84657 38505 84669 38508
rect 84703 38536 84715 38539
rect 84749 38539 84807 38545
rect 84749 38536 84761 38539
rect 84703 38508 84761 38536
rect 84703 38505 84715 38508
rect 84657 38499 84715 38505
rect 84749 38505 84761 38508
rect 84795 38505 84807 38539
rect 85945 38539 86003 38545
rect 85945 38536 85957 38539
rect 84749 38499 84807 38505
rect 85132 38508 85957 38536
rect 71133 38471 71191 38477
rect 71133 38437 71145 38471
rect 71179 38468 71191 38471
rect 71179 38440 72556 38468
rect 71179 38437 71191 38440
rect 71133 38431 71191 38437
rect 70351 38372 70900 38400
rect 70949 38403 71007 38409
rect 70351 38369 70363 38372
rect 70305 38363 70363 38369
rect 70949 38369 70961 38403
rect 70995 38400 71007 38403
rect 71225 38403 71283 38409
rect 71225 38400 71237 38403
rect 70995 38372 71237 38400
rect 70995 38369 71007 38372
rect 70949 38363 71007 38369
rect 71225 38369 71237 38372
rect 71271 38400 71283 38403
rect 71869 38403 71927 38409
rect 71869 38400 71881 38403
rect 71271 38372 71881 38400
rect 71271 38369 71283 38372
rect 71225 38363 71283 38369
rect 71869 38369 71881 38372
rect 71915 38369 71927 38403
rect 71869 38363 71927 38369
rect 72053 38403 72111 38409
rect 72053 38369 72065 38403
rect 72099 38369 72111 38403
rect 72053 38363 72111 38369
rect 68922 38292 68928 38344
rect 68980 38332 68986 38344
rect 71409 38335 71467 38341
rect 71409 38332 71421 38335
rect 68980 38304 71421 38332
rect 68980 38292 68986 38304
rect 71409 38301 71421 38304
rect 71455 38301 71467 38335
rect 71409 38295 71467 38301
rect 71774 38292 71780 38344
rect 71832 38332 71838 38344
rect 72068 38332 72096 38363
rect 72326 38360 72332 38412
rect 72384 38400 72390 38412
rect 72528 38409 72556 38440
rect 72421 38403 72479 38409
rect 72421 38400 72433 38403
rect 72384 38372 72433 38400
rect 72384 38360 72390 38372
rect 72421 38369 72433 38372
rect 72467 38369 72479 38403
rect 72421 38363 72479 38369
rect 72513 38403 72571 38409
rect 72513 38369 72525 38403
rect 72559 38369 72571 38403
rect 72513 38363 72571 38369
rect 73982 38360 73988 38412
rect 74040 38400 74046 38412
rect 74353 38403 74411 38409
rect 74353 38400 74365 38403
rect 74040 38372 74365 38400
rect 74040 38360 74046 38372
rect 74353 38369 74365 38372
rect 74399 38369 74411 38403
rect 77386 38400 77392 38412
rect 77347 38372 77392 38400
rect 74353 38363 74411 38369
rect 77386 38360 77392 38372
rect 77444 38400 77450 38412
rect 77665 38403 77723 38409
rect 77665 38400 77677 38403
rect 77444 38372 77677 38400
rect 77444 38360 77450 38372
rect 77665 38369 77677 38372
rect 77711 38369 77723 38403
rect 77665 38363 77723 38369
rect 81434 38360 81440 38412
rect 81492 38400 81498 38412
rect 81529 38403 81587 38409
rect 81529 38400 81541 38403
rect 81492 38372 81541 38400
rect 81492 38360 81498 38372
rect 81529 38369 81541 38372
rect 81575 38400 81587 38403
rect 81805 38403 81863 38409
rect 81805 38400 81817 38403
rect 81575 38372 81817 38400
rect 81575 38369 81587 38372
rect 81529 38363 81587 38369
rect 81805 38369 81817 38372
rect 81851 38369 81863 38403
rect 82814 38400 82820 38412
rect 82775 38372 82820 38400
rect 81805 38363 81863 38369
rect 82814 38360 82820 38372
rect 82872 38360 82878 38412
rect 82906 38360 82912 38412
rect 82964 38400 82970 38412
rect 85132 38409 85160 38508
rect 85945 38505 85957 38508
rect 85991 38536 86003 38539
rect 89070 38536 89076 38548
rect 85991 38508 88932 38536
rect 89031 38508 89076 38536
rect 85991 38505 86003 38508
rect 85945 38499 86003 38505
rect 85853 38471 85911 38477
rect 85853 38437 85865 38471
rect 85899 38468 85911 38471
rect 86954 38468 86960 38480
rect 85899 38440 86960 38468
rect 85899 38437 85911 38440
rect 85853 38431 85911 38437
rect 86954 38428 86960 38440
rect 87012 38428 87018 38480
rect 88426 38468 88432 38480
rect 88387 38440 88432 38468
rect 88426 38428 88432 38440
rect 88484 38428 88490 38480
rect 88904 38468 88932 38508
rect 89070 38496 89076 38508
rect 89128 38496 89134 38548
rect 90082 38536 90088 38548
rect 90043 38508 90088 38536
rect 90082 38496 90088 38508
rect 90140 38496 90146 38548
rect 93394 38496 93400 38548
rect 93452 38536 93458 38548
rect 95697 38539 95755 38545
rect 95697 38536 95709 38539
rect 93452 38508 95709 38536
rect 93452 38496 93458 38508
rect 95697 38505 95709 38508
rect 95743 38505 95755 38539
rect 95697 38499 95755 38505
rect 89438 38468 89444 38480
rect 88904 38440 89444 38468
rect 89438 38428 89444 38440
rect 89496 38428 89502 38480
rect 90453 38471 90511 38477
rect 90453 38437 90465 38471
rect 90499 38468 90511 38471
rect 91002 38468 91008 38480
rect 90499 38440 91008 38468
rect 90499 38437 90511 38440
rect 90453 38431 90511 38437
rect 91002 38428 91008 38440
rect 91060 38428 91066 38480
rect 85117 38403 85175 38409
rect 82964 38372 83009 38400
rect 82964 38360 82970 38372
rect 85117 38369 85129 38403
rect 85163 38369 85175 38403
rect 85117 38363 85175 38369
rect 85264 38403 85322 38409
rect 85264 38369 85276 38403
rect 85310 38400 85322 38403
rect 85666 38400 85672 38412
rect 85310 38372 85672 38400
rect 85310 38369 85322 38372
rect 85264 38363 85322 38369
rect 72602 38332 72608 38344
rect 71832 38304 72608 38332
rect 71832 38292 71838 38304
rect 72602 38292 72608 38304
rect 72660 38292 72666 38344
rect 72786 38292 72792 38344
rect 72844 38332 72850 38344
rect 85132 38332 85160 38363
rect 85666 38360 85672 38372
rect 85724 38400 85730 38412
rect 86218 38400 86224 38412
rect 85724 38372 86224 38400
rect 85724 38360 85730 38372
rect 86218 38360 86224 38372
rect 86276 38360 86282 38412
rect 88444 38400 88472 38428
rect 89257 38403 89315 38409
rect 89257 38400 89269 38403
rect 88444 38372 89269 38400
rect 89257 38369 89269 38372
rect 89303 38369 89315 38403
rect 91094 38400 91100 38412
rect 91055 38372 91100 38400
rect 89257 38363 89315 38369
rect 91094 38360 91100 38372
rect 91152 38360 91158 38412
rect 91465 38403 91523 38409
rect 91465 38369 91477 38403
rect 91511 38369 91523 38403
rect 91465 38363 91523 38369
rect 72844 38304 85160 38332
rect 85485 38335 85543 38341
rect 72844 38292 72850 38304
rect 85485 38301 85497 38335
rect 85531 38301 85543 38335
rect 85485 38295 85543 38301
rect 70397 38267 70455 38273
rect 70397 38264 70409 38267
rect 67416 38236 67588 38264
rect 68572 38236 70409 38264
rect 67416 38224 67422 38236
rect 67269 38199 67327 38205
rect 67269 38196 67281 38199
rect 65392 38168 67281 38196
rect 65392 38156 65398 38168
rect 67269 38165 67281 38168
rect 67315 38165 67327 38199
rect 67450 38196 67456 38208
rect 67411 38168 67456 38196
rect 67269 38159 67327 38165
rect 67450 38156 67456 38168
rect 67508 38156 67514 38208
rect 67560 38196 67588 38236
rect 70397 38233 70409 38236
rect 70443 38264 70455 38267
rect 71225 38267 71283 38273
rect 71225 38264 71237 38267
rect 70443 38236 71237 38264
rect 70443 38233 70455 38236
rect 70397 38227 70455 38233
rect 71225 38233 71237 38236
rect 71271 38233 71283 38267
rect 71225 38227 71283 38233
rect 71590 38224 71596 38276
rect 71648 38264 71654 38276
rect 81621 38267 81679 38273
rect 81621 38264 81633 38267
rect 71648 38236 81633 38264
rect 71648 38224 71654 38236
rect 81621 38233 81633 38236
rect 81667 38264 81679 38267
rect 83182 38264 83188 38276
rect 81667 38236 83188 38264
rect 81667 38233 81679 38236
rect 81621 38227 81679 38233
rect 83182 38224 83188 38236
rect 83240 38224 83246 38276
rect 84657 38267 84715 38273
rect 84657 38233 84669 38267
rect 84703 38264 84715 38267
rect 85393 38267 85451 38273
rect 85393 38264 85405 38267
rect 84703 38236 85405 38264
rect 84703 38233 84715 38236
rect 84657 38227 84715 38233
rect 85393 38233 85405 38236
rect 85439 38233 85451 38267
rect 85393 38227 85451 38233
rect 72694 38196 72700 38208
rect 67560 38168 72700 38196
rect 72694 38156 72700 38168
rect 72752 38156 72758 38208
rect 74166 38196 74172 38208
rect 74127 38168 74172 38196
rect 74166 38156 74172 38168
rect 74224 38156 74230 38208
rect 77478 38196 77484 38208
rect 77439 38168 77484 38196
rect 77478 38156 77484 38168
rect 77536 38196 77542 38208
rect 81526 38196 81532 38208
rect 77536 38168 81532 38196
rect 77536 38156 77542 38168
rect 81526 38156 81532 38168
rect 81584 38156 81590 38208
rect 81710 38156 81716 38208
rect 81768 38196 81774 38208
rect 82449 38199 82507 38205
rect 82449 38196 82461 38199
rect 81768 38168 82461 38196
rect 81768 38156 81774 38168
rect 82449 38165 82461 38168
rect 82495 38196 82507 38199
rect 82633 38199 82691 38205
rect 82633 38196 82645 38199
rect 82495 38168 82645 38196
rect 82495 38165 82507 38168
rect 82449 38159 82507 38165
rect 82633 38165 82645 38168
rect 82679 38165 82691 38199
rect 83090 38196 83096 38208
rect 83051 38168 83096 38196
rect 82633 38159 82691 38165
rect 83090 38156 83096 38168
rect 83148 38156 83154 38208
rect 83200 38196 83228 38224
rect 84933 38199 84991 38205
rect 84933 38196 84945 38199
rect 83200 38168 84945 38196
rect 84933 38165 84945 38168
rect 84979 38196 84991 38199
rect 85500 38196 85528 38295
rect 88518 38292 88524 38344
rect 88576 38341 88582 38344
rect 88576 38335 88634 38341
rect 88576 38301 88588 38335
rect 88622 38332 88634 38335
rect 88797 38335 88855 38341
rect 88622 38301 88656 38332
rect 88576 38295 88656 38301
rect 88797 38301 88809 38335
rect 88843 38332 88855 38335
rect 88843 38304 89668 38332
rect 88843 38301 88855 38304
rect 88797 38295 88855 38301
rect 88576 38292 88582 38295
rect 88628 38264 88656 38295
rect 89441 38267 89499 38273
rect 89441 38264 89453 38267
rect 88628 38236 89453 38264
rect 89441 38233 89453 38236
rect 89487 38233 89499 38267
rect 89441 38227 89499 38233
rect 89640 38208 89668 38304
rect 90082 38292 90088 38344
rect 90140 38332 90146 38344
rect 90910 38332 90916 38344
rect 90140 38304 90916 38332
rect 90140 38292 90146 38304
rect 90910 38292 90916 38304
rect 90968 38332 90974 38344
rect 91005 38335 91063 38341
rect 91005 38332 91017 38335
rect 90968 38304 91017 38332
rect 90968 38292 90974 38304
rect 91005 38301 91017 38304
rect 91051 38301 91063 38335
rect 91005 38295 91063 38301
rect 91480 38264 91508 38363
rect 91557 38335 91615 38341
rect 91557 38301 91569 38335
rect 91603 38301 91615 38335
rect 91557 38295 91615 38301
rect 94317 38335 94375 38341
rect 94317 38301 94329 38335
rect 94363 38301 94375 38335
rect 94590 38332 94596 38344
rect 94551 38304 94596 38332
rect 94317 38295 94375 38301
rect 90284 38236 91508 38264
rect 88702 38196 88708 38208
rect 84979 38168 85528 38196
rect 88663 38168 88708 38196
rect 84979 38165 84991 38168
rect 84933 38159 84991 38165
rect 88702 38156 88708 38168
rect 88760 38156 88766 38208
rect 89622 38196 89628 38208
rect 89583 38168 89628 38196
rect 89622 38156 89628 38168
rect 89680 38156 89686 38208
rect 89714 38156 89720 38208
rect 89772 38196 89778 38208
rect 90284 38205 90312 38236
rect 90269 38199 90327 38205
rect 90269 38196 90281 38199
rect 89772 38168 90281 38196
rect 89772 38156 89778 38168
rect 90269 38165 90281 38168
rect 90315 38165 90327 38199
rect 90269 38159 90327 38165
rect 91002 38156 91008 38208
rect 91060 38196 91066 38208
rect 91572 38196 91600 38295
rect 91060 38168 91600 38196
rect 94225 38199 94283 38205
rect 91060 38156 91066 38168
rect 94225 38165 94237 38199
rect 94271 38196 94283 38199
rect 94332 38196 94360 38295
rect 94590 38292 94596 38304
rect 94648 38292 94654 38344
rect 94498 38196 94504 38208
rect 94271 38168 94504 38196
rect 94271 38165 94283 38168
rect 94225 38159 94283 38165
rect 94498 38156 94504 38168
rect 94556 38156 94562 38208
rect 1104 38106 105616 38128
rect 1104 38054 4246 38106
rect 4298 38054 4310 38106
rect 4362 38054 4374 38106
rect 4426 38054 4438 38106
rect 4490 38054 34966 38106
rect 35018 38054 35030 38106
rect 35082 38054 35094 38106
rect 35146 38054 35158 38106
rect 35210 38054 65686 38106
rect 65738 38054 65750 38106
rect 65802 38054 65814 38106
rect 65866 38054 65878 38106
rect 65930 38054 96406 38106
rect 96458 38054 96470 38106
rect 96522 38054 96534 38106
rect 96586 38054 96598 38106
rect 96650 38054 105616 38106
rect 1104 38032 105616 38054
rect 4798 37952 4804 38004
rect 4856 37992 4862 38004
rect 5169 37995 5227 38001
rect 5169 37992 5181 37995
rect 4856 37964 5181 37992
rect 4856 37952 4862 37964
rect 5169 37961 5181 37964
rect 5215 37961 5227 37995
rect 5169 37955 5227 37961
rect 10594 37952 10600 38004
rect 10652 37992 10658 38004
rect 49786 37992 49792 38004
rect 10652 37964 49792 37992
rect 10652 37952 10658 37964
rect 49786 37952 49792 37964
rect 49844 37952 49850 38004
rect 49878 37952 49884 38004
rect 49936 37992 49942 38004
rect 51166 37992 51172 38004
rect 49936 37964 51172 37992
rect 49936 37952 49942 37964
rect 51166 37952 51172 37964
rect 51224 37952 51230 38004
rect 51258 37952 51264 38004
rect 51316 37992 51322 38004
rect 58986 37992 58992 38004
rect 51316 37964 58572 37992
rect 58947 37964 58992 37992
rect 51316 37952 51322 37964
rect 26326 37924 26332 37936
rect 23492 37896 26332 37924
rect 2774 37816 2780 37868
rect 2832 37856 2838 37868
rect 8297 37859 8355 37865
rect 2832 37828 2877 37856
rect 2832 37816 2838 37828
rect 8297 37825 8309 37859
rect 8343 37856 8355 37859
rect 10778 37856 10784 37868
rect 8343 37828 10784 37856
rect 8343 37825 8355 37828
rect 8297 37819 8355 37825
rect 10778 37816 10784 37828
rect 10836 37816 10842 37868
rect 12710 37856 12716 37868
rect 12671 37828 12716 37856
rect 12710 37816 12716 37828
rect 12768 37816 12774 37868
rect 18509 37859 18567 37865
rect 18509 37856 18521 37859
rect 18156 37828 18521 37856
rect 18156 37800 18184 37828
rect 18509 37825 18521 37828
rect 18555 37825 18567 37859
rect 18509 37819 18567 37825
rect 19245 37859 19303 37865
rect 19245 37825 19257 37859
rect 19291 37856 19303 37859
rect 21085 37859 21143 37865
rect 21085 37856 21097 37859
rect 19291 37828 21097 37856
rect 19291 37825 19303 37828
rect 19245 37819 19303 37825
rect 21085 37825 21097 37828
rect 21131 37856 21143 37859
rect 21174 37856 21180 37868
rect 21131 37828 21180 37856
rect 21131 37825 21143 37828
rect 21085 37819 21143 37825
rect 21174 37816 21180 37828
rect 21232 37816 21238 37868
rect 23492 37856 23520 37896
rect 26326 37884 26332 37896
rect 26384 37884 26390 37936
rect 26418 37884 26424 37936
rect 26476 37924 26482 37936
rect 26605 37927 26663 37933
rect 26605 37924 26617 37927
rect 26476 37896 26617 37924
rect 26476 37884 26482 37896
rect 26605 37893 26617 37896
rect 26651 37893 26663 37927
rect 26605 37887 26663 37893
rect 27065 37927 27123 37933
rect 27065 37893 27077 37927
rect 27111 37924 27123 37927
rect 27154 37924 27160 37936
rect 27111 37896 27160 37924
rect 27111 37893 27123 37896
rect 27065 37887 27123 37893
rect 27154 37884 27160 37896
rect 27212 37884 27218 37936
rect 31478 37924 31484 37936
rect 31439 37896 31484 37924
rect 31478 37884 31484 37896
rect 31536 37924 31542 37936
rect 31665 37927 31723 37933
rect 31665 37924 31677 37927
rect 31536 37896 31677 37924
rect 31536 37884 31542 37896
rect 31665 37893 31677 37896
rect 31711 37924 31723 37927
rect 31938 37924 31944 37936
rect 31711 37896 31944 37924
rect 31711 37893 31723 37896
rect 31665 37887 31723 37893
rect 31938 37884 31944 37896
rect 31996 37884 32002 37936
rect 39022 37884 39028 37936
rect 39080 37924 39086 37936
rect 40773 37927 40831 37933
rect 40773 37924 40785 37927
rect 39080 37896 40785 37924
rect 39080 37884 39086 37896
rect 40773 37893 40785 37896
rect 40819 37893 40831 37927
rect 45370 37924 45376 37936
rect 45331 37896 45376 37924
rect 40773 37887 40831 37893
rect 45370 37884 45376 37896
rect 45428 37884 45434 37936
rect 56318 37924 56324 37936
rect 45480 37896 55904 37924
rect 56279 37896 56324 37924
rect 21836 37828 23520 37856
rect 25654 37828 25912 37856
rect 2501 37791 2559 37797
rect 2501 37757 2513 37791
rect 2547 37788 2559 37791
rect 4985 37791 5043 37797
rect 2547 37760 4292 37788
rect 2547 37757 2559 37760
rect 2501 37751 2559 37757
rect 4264 37664 4292 37760
rect 4985 37757 4997 37791
rect 5031 37788 5043 37791
rect 5442 37788 5448 37800
rect 5031 37760 5448 37788
rect 5031 37757 5043 37760
rect 4985 37751 5043 37757
rect 5442 37748 5448 37760
rect 5500 37748 5506 37800
rect 8202 37788 8208 37800
rect 8163 37760 8208 37788
rect 8202 37748 8208 37760
rect 8260 37748 8266 37800
rect 8478 37748 8484 37800
rect 8536 37788 8542 37800
rect 8573 37791 8631 37797
rect 8573 37788 8585 37791
rect 8536 37760 8585 37788
rect 8536 37748 8542 37760
rect 8573 37757 8585 37760
rect 8619 37757 8631 37791
rect 8573 37751 8631 37757
rect 8757 37791 8815 37797
rect 8757 37757 8769 37791
rect 8803 37788 8815 37791
rect 12158 37788 12164 37800
rect 8803 37760 12164 37788
rect 8803 37757 8815 37760
rect 8757 37751 8815 37757
rect 12158 37748 12164 37760
rect 12216 37748 12222 37800
rect 12437 37791 12495 37797
rect 12437 37757 12449 37791
rect 12483 37788 12495 37791
rect 18138 37788 18144 37800
rect 12483 37760 13768 37788
rect 18099 37760 18144 37788
rect 12483 37757 12495 37760
rect 12437 37751 12495 37757
rect 6546 37680 6552 37732
rect 6604 37720 6610 37732
rect 7561 37723 7619 37729
rect 7561 37720 7573 37723
rect 6604 37692 7573 37720
rect 6604 37680 6610 37692
rect 7561 37689 7573 37692
rect 7607 37689 7619 37723
rect 7561 37683 7619 37689
rect 13740 37664 13768 37760
rect 18138 37748 18144 37760
rect 18196 37748 18202 37800
rect 18322 37748 18328 37800
rect 18380 37788 18386 37800
rect 19150 37788 19156 37800
rect 18380 37760 19156 37788
rect 18380 37748 18386 37760
rect 19150 37748 19156 37760
rect 19208 37748 19214 37800
rect 19521 37791 19579 37797
rect 19521 37757 19533 37791
rect 19567 37788 19579 37791
rect 20806 37788 20812 37800
rect 19567 37760 20812 37788
rect 19567 37757 19579 37760
rect 19521 37751 19579 37757
rect 20806 37748 20812 37760
rect 20864 37748 20870 37800
rect 20901 37791 20959 37797
rect 20901 37757 20913 37791
rect 20947 37788 20959 37791
rect 21729 37791 21787 37797
rect 21729 37788 21741 37791
rect 20947 37760 21741 37788
rect 20947 37757 20959 37760
rect 20901 37751 20959 37757
rect 21729 37757 21741 37760
rect 21775 37757 21787 37791
rect 21729 37751 21787 37757
rect 14090 37720 14096 37732
rect 14003 37692 14096 37720
rect 14090 37680 14096 37692
rect 14148 37720 14154 37732
rect 21836 37720 21864 37828
rect 23382 37748 23388 37800
rect 23440 37788 23446 37800
rect 25654 37797 25682 37828
rect 25639 37791 25697 37797
rect 25639 37788 25651 37791
rect 23440 37760 25651 37788
rect 23440 37748 23446 37760
rect 25639 37757 25651 37760
rect 25685 37757 25697 37791
rect 25774 37788 25780 37800
rect 25735 37760 25780 37788
rect 25639 37751 25697 37757
rect 25774 37748 25780 37760
rect 25832 37748 25838 37800
rect 14148 37692 18460 37720
rect 14148 37680 14154 37692
rect 3418 37612 3424 37664
rect 3476 37652 3482 37664
rect 3881 37655 3939 37661
rect 3881 37652 3893 37655
rect 3476 37624 3893 37652
rect 3476 37612 3482 37624
rect 3881 37621 3893 37624
rect 3927 37621 3939 37655
rect 4246 37652 4252 37664
rect 4207 37624 4252 37652
rect 3881 37615 3939 37621
rect 4246 37612 4252 37624
rect 4304 37612 4310 37664
rect 13722 37612 13728 37664
rect 13780 37652 13786 37664
rect 14185 37655 14243 37661
rect 14185 37652 14197 37655
rect 13780 37624 14197 37652
rect 13780 37612 13786 37624
rect 14185 37621 14197 37624
rect 14231 37621 14243 37655
rect 18322 37652 18328 37664
rect 18283 37624 18328 37652
rect 14185 37615 14243 37621
rect 18322 37612 18328 37624
rect 18380 37612 18386 37664
rect 18432 37652 18460 37692
rect 20272 37692 21864 37720
rect 25409 37723 25467 37729
rect 20272 37652 20300 37692
rect 25409 37689 25421 37723
rect 25455 37720 25467 37723
rect 25792 37720 25820 37748
rect 25455 37692 25820 37720
rect 25884 37720 25912 37828
rect 28902 37816 28908 37868
rect 28960 37856 28966 37868
rect 32217 37859 32275 37865
rect 32217 37856 32229 37859
rect 28960 37828 32229 37856
rect 28960 37816 28966 37828
rect 32217 37825 32229 37828
rect 32263 37825 32275 37859
rect 32217 37819 32275 37825
rect 36998 37816 37004 37868
rect 37056 37856 37062 37868
rect 38105 37859 38163 37865
rect 38105 37856 38117 37859
rect 37056 37828 38117 37856
rect 37056 37816 37062 37828
rect 38105 37825 38117 37828
rect 38151 37825 38163 37859
rect 38105 37819 38163 37825
rect 39298 37816 39304 37868
rect 39356 37856 39362 37868
rect 39485 37859 39543 37865
rect 39485 37856 39497 37859
rect 39356 37828 39497 37856
rect 39356 37816 39362 37828
rect 39485 37825 39497 37828
rect 39531 37856 39543 37859
rect 39942 37856 39948 37868
rect 39531 37828 39948 37856
rect 39531 37825 39543 37828
rect 39485 37819 39543 37825
rect 39942 37816 39948 37828
rect 40000 37816 40006 37868
rect 40126 37816 40132 37868
rect 40184 37856 40190 37868
rect 40644 37859 40702 37865
rect 40644 37856 40656 37859
rect 40184 37828 40656 37856
rect 40184 37816 40190 37828
rect 40644 37825 40656 37828
rect 40690 37825 40702 37859
rect 40862 37856 40868 37868
rect 40823 37828 40868 37856
rect 40644 37819 40702 37825
rect 40862 37816 40868 37828
rect 40920 37816 40926 37868
rect 41230 37856 41236 37868
rect 41191 37828 41236 37856
rect 41230 37816 41236 37828
rect 41288 37816 41294 37868
rect 26142 37788 26148 37800
rect 26103 37760 26148 37788
rect 26142 37748 26148 37760
rect 26200 37748 26206 37800
rect 26237 37791 26295 37797
rect 26237 37757 26249 37791
rect 26283 37788 26295 37791
rect 27890 37788 27896 37800
rect 26283 37760 27896 37788
rect 26283 37757 26295 37760
rect 26237 37751 26295 37757
rect 26252 37720 26280 37751
rect 27890 37748 27896 37760
rect 27948 37748 27954 37800
rect 31846 37788 31852 37800
rect 31807 37760 31852 37788
rect 31846 37748 31852 37760
rect 31904 37748 31910 37800
rect 31938 37748 31944 37800
rect 31996 37788 32002 37800
rect 33594 37788 33600 37800
rect 31996 37760 32041 37788
rect 33555 37760 33600 37788
rect 31996 37748 32002 37760
rect 33594 37748 33600 37760
rect 33652 37748 33658 37800
rect 37550 37748 37556 37800
rect 37608 37788 37614 37800
rect 37829 37791 37887 37797
rect 37829 37788 37841 37791
rect 37608 37760 37841 37788
rect 37608 37748 37614 37760
rect 37829 37757 37841 37760
rect 37875 37757 37887 37791
rect 40402 37788 40408 37800
rect 37829 37751 37887 37757
rect 37936 37760 40408 37788
rect 25884 37692 26280 37720
rect 25455 37689 25467 37692
rect 25409 37683 25467 37689
rect 35986 37680 35992 37732
rect 36044 37720 36050 37732
rect 37936 37720 37964 37760
rect 40402 37748 40408 37760
rect 40460 37748 40466 37800
rect 40497 37791 40555 37797
rect 40497 37757 40509 37791
rect 40543 37788 40555 37791
rect 41138 37788 41144 37800
rect 40543 37760 41144 37788
rect 40543 37757 40555 37760
rect 40497 37751 40555 37757
rect 41138 37748 41144 37760
rect 41196 37748 41202 37800
rect 43809 37791 43867 37797
rect 43809 37788 43821 37791
rect 41248 37760 43821 37788
rect 36044 37692 37964 37720
rect 36044 37680 36050 37692
rect 39390 37680 39396 37732
rect 39448 37720 39454 37732
rect 41248 37720 41276 37760
rect 43809 37757 43821 37760
rect 43855 37757 43867 37791
rect 43809 37751 43867 37757
rect 43993 37791 44051 37797
rect 43993 37757 44005 37791
rect 44039 37788 44051 37791
rect 44082 37788 44088 37800
rect 44039 37760 44088 37788
rect 44039 37757 44051 37760
rect 43993 37751 44051 37757
rect 44082 37748 44088 37760
rect 44140 37748 44146 37800
rect 44450 37788 44456 37800
rect 44411 37760 44456 37788
rect 44450 37748 44456 37760
rect 44508 37748 44514 37800
rect 44545 37791 44603 37797
rect 44545 37757 44557 37791
rect 44591 37788 44603 37791
rect 45388 37788 45416 37884
rect 44591 37760 45416 37788
rect 44591 37757 44603 37760
rect 44545 37751 44603 37757
rect 39448 37692 41276 37720
rect 39448 37680 39454 37692
rect 42886 37680 42892 37732
rect 42944 37720 42950 37732
rect 45480 37720 45508 37896
rect 45554 37816 45560 37868
rect 45612 37856 45618 37868
rect 45612 37828 45657 37856
rect 45612 37816 45618 37828
rect 46658 37816 46664 37868
rect 46716 37856 46722 37868
rect 49602 37856 49608 37868
rect 46716 37828 49608 37856
rect 46716 37816 46722 37828
rect 49602 37816 49608 37828
rect 49660 37816 49666 37868
rect 51261 37859 51319 37865
rect 51261 37825 51273 37859
rect 51307 37856 51319 37859
rect 51350 37856 51356 37868
rect 51307 37828 51356 37856
rect 51307 37825 51319 37828
rect 51261 37819 51319 37825
rect 51350 37816 51356 37828
rect 51408 37856 51414 37868
rect 51721 37859 51779 37865
rect 51721 37856 51733 37859
rect 51408 37828 51733 37856
rect 51408 37816 51414 37828
rect 51721 37825 51733 37828
rect 51767 37825 51779 37859
rect 53374 37856 53380 37868
rect 51721 37819 51779 37825
rect 52840 37828 53380 37856
rect 46198 37748 46204 37800
rect 46256 37788 46262 37800
rect 50706 37788 50712 37800
rect 46256 37760 50712 37788
rect 46256 37748 46262 37760
rect 50706 37748 50712 37760
rect 50764 37748 50770 37800
rect 51445 37791 51503 37797
rect 51445 37757 51457 37791
rect 51491 37788 51503 37791
rect 51534 37788 51540 37800
rect 51491 37760 51540 37788
rect 51491 37757 51503 37760
rect 51445 37751 51503 37757
rect 51534 37748 51540 37760
rect 51592 37748 51598 37800
rect 51810 37748 51816 37800
rect 51868 37788 51874 37800
rect 51905 37791 51963 37797
rect 51905 37788 51917 37791
rect 51868 37760 51917 37788
rect 51868 37748 51874 37760
rect 51905 37757 51917 37760
rect 51951 37757 51963 37791
rect 52362 37788 52368 37800
rect 52323 37760 52368 37788
rect 51905 37751 51963 37757
rect 52362 37748 52368 37760
rect 52420 37748 52426 37800
rect 52454 37748 52460 37800
rect 52512 37788 52518 37800
rect 52840 37788 52868 37828
rect 53374 37816 53380 37828
rect 53432 37816 53438 37868
rect 55876 37856 55904 37896
rect 56318 37884 56324 37896
rect 56376 37884 56382 37936
rect 58544 37924 58572 37964
rect 58986 37952 58992 37964
rect 59044 37952 59050 38004
rect 60258 37995 60316 38001
rect 60258 37961 60270 37995
rect 60304 37992 60316 37995
rect 60642 37992 60648 38004
rect 60304 37964 60648 37992
rect 60304 37961 60316 37964
rect 60258 37955 60316 37961
rect 60642 37952 60648 37964
rect 60700 37952 60706 38004
rect 62114 37952 62120 38004
rect 62172 37992 62178 38004
rect 62850 37992 62856 38004
rect 62172 37964 62856 37992
rect 62172 37952 62178 37964
rect 62850 37952 62856 37964
rect 62908 37952 62914 38004
rect 64432 37964 82860 37992
rect 64432 37924 64460 37964
rect 58544 37896 64460 37924
rect 65426 37884 65432 37936
rect 65484 37924 65490 37936
rect 77478 37924 77484 37936
rect 65484 37896 70348 37924
rect 65484 37884 65490 37896
rect 59722 37856 59728 37868
rect 55876 37828 59728 37856
rect 59722 37816 59728 37828
rect 59780 37816 59786 37868
rect 59906 37856 59912 37868
rect 59867 37828 59912 37856
rect 59906 37816 59912 37828
rect 59964 37816 59970 37868
rect 60458 37856 60464 37868
rect 60419 37828 60464 37856
rect 60458 37816 60464 37828
rect 60516 37816 60522 37868
rect 64230 37816 64236 37868
rect 64288 37856 64294 37868
rect 64417 37859 64475 37865
rect 64417 37856 64429 37859
rect 64288 37828 64429 37856
rect 64288 37816 64294 37828
rect 64417 37825 64429 37828
rect 64463 37825 64475 37859
rect 64690 37856 64696 37868
rect 64651 37828 64696 37856
rect 64417 37819 64475 37825
rect 64690 37816 64696 37828
rect 64748 37816 64754 37868
rect 68741 37859 68799 37865
rect 68741 37825 68753 37859
rect 68787 37856 68799 37859
rect 70213 37859 70271 37865
rect 70213 37856 70225 37859
rect 68787 37828 70225 37856
rect 68787 37825 68799 37828
rect 68741 37819 68799 37825
rect 70213 37825 70225 37828
rect 70259 37825 70271 37859
rect 70213 37819 70271 37825
rect 52512 37760 52868 37788
rect 52512 37748 52518 37760
rect 56226 37748 56232 37800
rect 56284 37788 56290 37800
rect 57333 37791 57391 37797
rect 56284 37760 56329 37788
rect 56284 37748 56290 37760
rect 57333 37757 57345 37791
rect 57379 37788 57391 37791
rect 57422 37788 57428 37800
rect 57379 37760 57428 37788
rect 57379 37757 57391 37760
rect 57333 37751 57391 37757
rect 57422 37748 57428 37760
rect 57480 37788 57486 37800
rect 57609 37791 57667 37797
rect 57609 37788 57621 37791
rect 57480 37760 57621 37788
rect 57480 37748 57486 37760
rect 57609 37757 57621 37760
rect 57655 37757 57667 37791
rect 57609 37751 57667 37757
rect 57885 37791 57943 37797
rect 57885 37757 57897 37791
rect 57931 37788 57943 37791
rect 58250 37788 58256 37800
rect 57931 37760 58256 37788
rect 57931 37757 57943 37760
rect 57885 37751 57943 37757
rect 58250 37748 58256 37760
rect 58308 37748 58314 37800
rect 59924 37788 59952 37816
rect 60323 37791 60381 37797
rect 60323 37788 60335 37791
rect 59924 37760 60335 37788
rect 60323 37757 60335 37760
rect 60369 37757 60381 37791
rect 60323 37751 60381 37757
rect 60829 37791 60887 37797
rect 60829 37757 60841 37791
rect 60875 37788 60887 37791
rect 64322 37788 64328 37800
rect 60875 37760 64328 37788
rect 60875 37757 60887 37760
rect 60829 37751 60887 37757
rect 64322 37748 64328 37760
rect 64380 37748 64386 37800
rect 68557 37791 68615 37797
rect 68557 37757 68569 37791
rect 68603 37788 68615 37791
rect 68649 37791 68707 37797
rect 68649 37788 68661 37791
rect 68603 37760 68661 37788
rect 68603 37757 68615 37760
rect 68557 37751 68615 37757
rect 68649 37757 68661 37760
rect 68695 37757 68707 37791
rect 68922 37788 68928 37800
rect 68883 37760 68928 37788
rect 68649 37751 68707 37757
rect 68922 37748 68928 37760
rect 68980 37748 68986 37800
rect 70320 37788 70348 37896
rect 70412 37896 77484 37924
rect 70412 37788 70440 37896
rect 77478 37884 77484 37896
rect 77536 37884 77542 37936
rect 82832 37924 82860 37964
rect 82906 37952 82912 38004
rect 82964 37992 82970 38004
rect 84105 37995 84163 38001
rect 84105 37992 84117 37995
rect 82964 37964 84117 37992
rect 82964 37952 82970 37964
rect 84105 37961 84117 37964
rect 84151 37961 84163 37995
rect 84105 37955 84163 37961
rect 85853 37927 85911 37933
rect 85853 37924 85865 37927
rect 82832 37896 85865 37924
rect 85853 37893 85865 37896
rect 85899 37924 85911 37927
rect 89165 37927 89223 37933
rect 89165 37924 89177 37927
rect 85899 37896 89177 37924
rect 85899 37893 85911 37896
rect 85853 37887 85911 37893
rect 89165 37893 89177 37896
rect 89211 37893 89223 37927
rect 89438 37924 89444 37936
rect 89399 37896 89444 37924
rect 89165 37887 89223 37893
rect 71590 37856 71596 37868
rect 71551 37828 71596 37856
rect 71590 37816 71596 37828
rect 71648 37816 71654 37868
rect 72694 37856 72700 37868
rect 72655 37828 72700 37856
rect 72694 37816 72700 37828
rect 72752 37816 72758 37868
rect 76742 37856 76748 37868
rect 76703 37828 76748 37856
rect 76742 37816 76748 37828
rect 76800 37856 76806 37868
rect 81621 37859 81679 37865
rect 76800 37828 76880 37856
rect 76800 37816 76806 37828
rect 70320 37760 70440 37788
rect 70486 37748 70492 37800
rect 70544 37788 70550 37800
rect 70673 37791 70731 37797
rect 70673 37788 70685 37791
rect 70544 37760 70685 37788
rect 70544 37748 70550 37760
rect 70673 37757 70685 37760
rect 70719 37757 70731 37791
rect 70673 37751 70731 37757
rect 70762 37748 70768 37800
rect 70820 37788 70826 37800
rect 70857 37791 70915 37797
rect 70857 37788 70869 37791
rect 70820 37760 70869 37788
rect 70820 37748 70826 37760
rect 70857 37757 70869 37760
rect 70903 37788 70915 37791
rect 71038 37788 71044 37800
rect 70903 37760 71044 37788
rect 70903 37757 70915 37760
rect 70857 37751 70915 37757
rect 71038 37748 71044 37760
rect 71096 37748 71102 37800
rect 71222 37788 71228 37800
rect 71183 37760 71228 37788
rect 71222 37748 71228 37760
rect 71280 37748 71286 37800
rect 71314 37748 71320 37800
rect 71372 37788 71378 37800
rect 72234 37788 72240 37800
rect 71372 37760 71417 37788
rect 72195 37760 72240 37788
rect 71372 37748 71378 37760
rect 72234 37748 72240 37760
rect 72292 37748 72298 37800
rect 72329 37791 72387 37797
rect 72329 37757 72341 37791
rect 72375 37757 72387 37791
rect 72329 37751 72387 37757
rect 42944 37692 45508 37720
rect 42944 37680 42950 37692
rect 45554 37680 45560 37732
rect 45612 37720 45618 37732
rect 48314 37720 48320 37732
rect 45612 37692 48320 37720
rect 45612 37680 45618 37692
rect 48314 37680 48320 37692
rect 48372 37680 48378 37732
rect 48406 37680 48412 37732
rect 48464 37720 48470 37732
rect 59725 37723 59783 37729
rect 59725 37720 59737 37723
rect 48464 37692 57560 37720
rect 48464 37680 48470 37692
rect 18432 37624 20300 37652
rect 20346 37612 20352 37664
rect 20404 37652 20410 37664
rect 21634 37652 21640 37664
rect 20404 37624 21640 37652
rect 20404 37612 20410 37624
rect 21634 37612 21640 37624
rect 21692 37612 21698 37664
rect 21818 37652 21824 37664
rect 21779 37624 21824 37652
rect 21818 37612 21824 37624
rect 21876 37612 21882 37664
rect 32030 37612 32036 37664
rect 32088 37652 32094 37664
rect 37550 37652 37556 37664
rect 32088 37624 37556 37652
rect 32088 37612 32094 37624
rect 37550 37612 37556 37624
rect 37608 37652 37614 37664
rect 37645 37655 37703 37661
rect 37645 37652 37657 37655
rect 37608 37624 37657 37652
rect 37608 37612 37614 37624
rect 37645 37621 37657 37624
rect 37691 37621 37703 37655
rect 37645 37615 37703 37621
rect 37734 37612 37740 37664
rect 37792 37652 37798 37664
rect 38930 37652 38936 37664
rect 37792 37624 38936 37652
rect 37792 37612 37798 37624
rect 38930 37612 38936 37624
rect 38988 37612 38994 37664
rect 40126 37612 40132 37664
rect 40184 37652 40190 37664
rect 40221 37655 40279 37661
rect 40221 37652 40233 37655
rect 40184 37624 40233 37652
rect 40184 37612 40190 37624
rect 40221 37621 40233 37624
rect 40267 37621 40279 37655
rect 40221 37615 40279 37621
rect 42794 37612 42800 37664
rect 42852 37652 42858 37664
rect 44082 37652 44088 37664
rect 42852 37624 44088 37652
rect 42852 37612 42858 37624
rect 44082 37612 44088 37624
rect 44140 37612 44146 37664
rect 45005 37655 45063 37661
rect 45005 37621 45017 37655
rect 45051 37652 45063 37655
rect 46658 37652 46664 37664
rect 45051 37624 46664 37652
rect 45051 37621 45063 37624
rect 45005 37615 45063 37621
rect 46658 37612 46664 37624
rect 46716 37612 46722 37664
rect 47854 37612 47860 37664
rect 47912 37652 47918 37664
rect 52454 37652 52460 37664
rect 47912 37624 52460 37652
rect 47912 37612 47918 37624
rect 52454 37612 52460 37624
rect 52512 37612 52518 37664
rect 52914 37652 52920 37664
rect 52875 37624 52920 37652
rect 52914 37612 52920 37624
rect 52972 37612 52978 37664
rect 53285 37655 53343 37661
rect 53285 37621 53297 37655
rect 53331 37652 53343 37655
rect 53374 37652 53380 37664
rect 53331 37624 53380 37652
rect 53331 37621 53343 37624
rect 53285 37615 53343 37621
rect 53374 37612 53380 37624
rect 53432 37612 53438 37664
rect 54202 37612 54208 37664
rect 54260 37652 54266 37664
rect 57333 37655 57391 37661
rect 57333 37652 57345 37655
rect 54260 37624 57345 37652
rect 54260 37612 54266 37624
rect 57333 37621 57345 37624
rect 57379 37652 57391 37655
rect 57425 37655 57483 37661
rect 57425 37652 57437 37655
rect 57379 37624 57437 37652
rect 57379 37621 57391 37624
rect 57333 37615 57391 37621
rect 57425 37621 57437 37624
rect 57471 37621 57483 37655
rect 57532 37652 57560 37692
rect 58544 37692 59737 37720
rect 58544 37652 58572 37692
rect 59725 37689 59737 37692
rect 59771 37720 59783 37723
rect 60093 37723 60151 37729
rect 60093 37720 60105 37723
rect 59771 37692 60105 37720
rect 59771 37689 59783 37692
rect 59725 37683 59783 37689
rect 60093 37689 60105 37692
rect 60139 37689 60151 37723
rect 60093 37683 60151 37689
rect 66073 37723 66131 37729
rect 66073 37689 66085 37723
rect 66119 37720 66131 37723
rect 69290 37720 69296 37732
rect 66119 37692 69296 37720
rect 66119 37689 66131 37692
rect 66073 37683 66131 37689
rect 69290 37680 69296 37692
rect 69348 37680 69354 37732
rect 69566 37680 69572 37732
rect 69624 37720 69630 37732
rect 72344 37720 72372 37751
rect 72418 37748 72424 37800
rect 72476 37788 72482 37800
rect 76852 37797 76880 37828
rect 81621 37825 81633 37859
rect 81667 37856 81679 37859
rect 83090 37856 83096 37868
rect 81667 37828 83096 37856
rect 81667 37825 81679 37828
rect 81621 37819 81679 37825
rect 83090 37816 83096 37828
rect 83148 37816 83154 37868
rect 89180 37856 89208 37887
rect 89438 37884 89444 37896
rect 89496 37924 89502 37936
rect 90177 37927 90235 37933
rect 90177 37924 90189 37927
rect 89496 37896 90189 37924
rect 89496 37884 89502 37896
rect 90177 37893 90189 37896
rect 90223 37924 90235 37927
rect 91278 37924 91284 37936
rect 90223 37896 91284 37924
rect 90223 37893 90235 37896
rect 90177 37887 90235 37893
rect 91278 37884 91284 37896
rect 91336 37884 91342 37936
rect 89898 37856 89904 37868
rect 89180 37828 89760 37856
rect 89859 37828 89904 37856
rect 72513 37791 72571 37797
rect 72513 37788 72525 37791
rect 72476 37760 72525 37788
rect 72476 37748 72482 37760
rect 72513 37757 72525 37760
rect 72559 37757 72571 37791
rect 72513 37751 72571 37757
rect 76837 37791 76895 37797
rect 76837 37757 76849 37791
rect 76883 37757 76895 37791
rect 77478 37788 77484 37800
rect 77439 37760 77484 37788
rect 76837 37751 76895 37757
rect 77478 37748 77484 37760
rect 77536 37748 77542 37800
rect 77662 37788 77668 37800
rect 77623 37760 77668 37788
rect 77662 37748 77668 37760
rect 77720 37748 77726 37800
rect 81253 37791 81311 37797
rect 81253 37757 81265 37791
rect 81299 37788 81311 37791
rect 81345 37791 81403 37797
rect 81345 37788 81357 37791
rect 81299 37760 81357 37788
rect 81299 37757 81311 37760
rect 81253 37751 81311 37757
rect 81345 37757 81357 37760
rect 81391 37788 81403 37791
rect 82538 37788 82544 37800
rect 81391 37760 82544 37788
rect 81391 37757 81403 37760
rect 81345 37751 81403 37757
rect 82538 37748 82544 37760
rect 82596 37748 82602 37800
rect 83826 37788 83832 37800
rect 83787 37760 83832 37788
rect 83826 37748 83832 37760
rect 83884 37748 83890 37800
rect 84013 37791 84071 37797
rect 84013 37757 84025 37791
rect 84059 37757 84071 37791
rect 85666 37788 85672 37800
rect 85627 37760 85672 37788
rect 84013 37751 84071 37757
rect 81434 37720 81440 37732
rect 69624 37692 72372 37720
rect 72804 37692 81440 37720
rect 69624 37680 69630 37692
rect 64230 37652 64236 37664
rect 57532 37624 58572 37652
rect 64191 37624 64236 37652
rect 57425 37615 57483 37621
rect 64230 37612 64236 37624
rect 64288 37652 64294 37664
rect 64414 37652 64420 37664
rect 64288 37624 64420 37652
rect 64288 37612 64294 37624
rect 64414 37612 64420 37624
rect 64472 37652 64478 37664
rect 65334 37652 65340 37664
rect 64472 37624 65340 37652
rect 64472 37612 64478 37624
rect 65334 37612 65340 37624
rect 65392 37612 65398 37664
rect 68557 37655 68615 37661
rect 68557 37621 68569 37655
rect 68603 37652 68615 37655
rect 68922 37652 68928 37664
rect 68603 37624 68928 37652
rect 68603 37621 68615 37624
rect 68557 37615 68615 37621
rect 68922 37612 68928 37624
rect 68980 37612 68986 37664
rect 69106 37652 69112 37664
rect 69067 37624 69112 37652
rect 69106 37612 69112 37624
rect 69164 37612 69170 37664
rect 71222 37612 71228 37664
rect 71280 37652 71286 37664
rect 71777 37655 71835 37661
rect 71777 37652 71789 37655
rect 71280 37624 71789 37652
rect 71280 37612 71286 37624
rect 71777 37621 71789 37624
rect 71823 37652 71835 37655
rect 72804 37652 72832 37692
rect 81434 37680 81440 37692
rect 81492 37680 81498 37732
rect 84028 37720 84056 37751
rect 85666 37748 85672 37760
rect 85724 37748 85730 37800
rect 89640 37797 89668 37828
rect 89732 37800 89760 37828
rect 89898 37816 89904 37828
rect 89956 37816 89962 37868
rect 91554 37856 91560 37868
rect 91515 37828 91560 37856
rect 91554 37816 91560 37828
rect 91612 37816 91618 37868
rect 94041 37859 94099 37865
rect 94041 37825 94053 37859
rect 94087 37856 94099 37859
rect 94590 37856 94596 37868
rect 94087 37828 94596 37856
rect 94087 37825 94099 37828
rect 94041 37819 94099 37825
rect 94590 37816 94596 37828
rect 94648 37816 94654 37868
rect 89349 37791 89407 37797
rect 89349 37757 89361 37791
rect 89395 37757 89407 37791
rect 89349 37751 89407 37757
rect 89595 37791 89668 37797
rect 89595 37757 89607 37791
rect 89641 37760 89668 37791
rect 89641 37757 89653 37760
rect 89595 37751 89653 37757
rect 83660 37692 84056 37720
rect 89364 37720 89392 37751
rect 89714 37748 89720 37800
rect 89772 37788 89778 37800
rect 91189 37791 91247 37797
rect 91189 37788 91201 37791
rect 89772 37760 91201 37788
rect 89772 37748 89778 37760
rect 91189 37757 91201 37760
rect 91235 37788 91247 37791
rect 91649 37791 91707 37797
rect 91649 37788 91661 37791
rect 91235 37760 91661 37788
rect 91235 37757 91247 37760
rect 91189 37751 91247 37757
rect 91649 37757 91661 37760
rect 91695 37757 91707 37791
rect 93305 37791 93363 37797
rect 93305 37788 93317 37791
rect 91649 37751 91707 37757
rect 93136 37760 93317 37788
rect 91002 37720 91008 37732
rect 89364 37692 91008 37720
rect 71823 37624 72832 37652
rect 76929 37655 76987 37661
rect 71823 37621 71835 37624
rect 71777 37615 71835 37621
rect 76929 37621 76941 37655
rect 76975 37652 76987 37655
rect 77294 37652 77300 37664
rect 76975 37624 77300 37652
rect 76975 37621 76987 37624
rect 76929 37615 76987 37621
rect 77294 37612 77300 37624
rect 77352 37612 77358 37664
rect 81452 37652 81480 37680
rect 83660 37661 83688 37692
rect 91002 37680 91008 37692
rect 91060 37680 91066 37732
rect 82725 37655 82783 37661
rect 82725 37652 82737 37655
rect 81452 37624 82737 37652
rect 82725 37621 82737 37624
rect 82771 37652 82783 37655
rect 83645 37655 83703 37661
rect 83645 37652 83657 37655
rect 82771 37624 83657 37652
rect 82771 37621 82783 37624
rect 82725 37615 82783 37621
rect 83645 37621 83657 37624
rect 83691 37621 83703 37655
rect 83645 37615 83703 37621
rect 90726 37612 90732 37664
rect 90784 37652 90790 37664
rect 93136 37661 93164 37760
rect 93305 37757 93317 37760
rect 93351 37757 93363 37791
rect 93486 37788 93492 37800
rect 93447 37760 93492 37788
rect 93305 37751 93363 37757
rect 93486 37748 93492 37760
rect 93544 37748 93550 37800
rect 93578 37748 93584 37800
rect 93636 37788 93642 37800
rect 94961 37791 95019 37797
rect 94961 37788 94973 37791
rect 93636 37760 93681 37788
rect 94792 37760 94973 37788
rect 93636 37748 93642 37760
rect 94792 37661 94820 37760
rect 94961 37757 94973 37760
rect 95007 37757 95019 37791
rect 95234 37788 95240 37800
rect 95195 37760 95240 37788
rect 94961 37751 95019 37757
rect 95234 37748 95240 37760
rect 95292 37748 95298 37800
rect 96617 37791 96675 37797
rect 96617 37757 96629 37791
rect 96663 37788 96675 37791
rect 97074 37788 97080 37800
rect 96663 37760 97080 37788
rect 96663 37757 96675 37760
rect 96617 37751 96675 37757
rect 97074 37748 97080 37760
rect 97132 37748 97138 37800
rect 95145 37723 95203 37729
rect 95145 37689 95157 37723
rect 95191 37720 95203 37723
rect 95326 37720 95332 37732
rect 95191 37692 95332 37720
rect 95191 37689 95203 37692
rect 95145 37683 95203 37689
rect 95326 37680 95332 37692
rect 95384 37680 95390 37732
rect 95694 37720 95700 37732
rect 95655 37692 95700 37720
rect 95694 37680 95700 37692
rect 95752 37680 95758 37732
rect 93121 37655 93179 37661
rect 93121 37652 93133 37655
rect 90784 37624 93133 37652
rect 90784 37612 90790 37624
rect 93121 37621 93133 37624
rect 93167 37652 93179 37655
rect 94777 37655 94835 37661
rect 94777 37652 94789 37655
rect 93167 37624 94789 37652
rect 93167 37621 93179 37624
rect 93121 37615 93179 37621
rect 94777 37621 94789 37624
rect 94823 37621 94835 37655
rect 96706 37652 96712 37664
rect 96667 37624 96712 37652
rect 94777 37615 94835 37621
rect 96706 37612 96712 37624
rect 96764 37612 96770 37664
rect 1104 37562 105616 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 50326 37562
rect 50378 37510 50390 37562
rect 50442 37510 50454 37562
rect 50506 37510 50518 37562
rect 50570 37510 81046 37562
rect 81098 37510 81110 37562
rect 81162 37510 81174 37562
rect 81226 37510 81238 37562
rect 81290 37510 105616 37562
rect 1104 37488 105616 37510
rect 8941 37451 8999 37457
rect 8941 37417 8953 37451
rect 8987 37448 8999 37451
rect 16022 37448 16028 37460
rect 8987 37420 16028 37448
rect 8987 37417 8999 37420
rect 8941 37411 8999 37417
rect 8205 37383 8263 37389
rect 8205 37349 8217 37383
rect 8251 37380 8263 37383
rect 8570 37380 8576 37392
rect 8251 37352 8576 37380
rect 8251 37349 8263 37352
rect 8205 37343 8263 37349
rect 8570 37340 8576 37352
rect 8628 37340 8634 37392
rect 4341 37315 4399 37321
rect 4341 37281 4353 37315
rect 4387 37312 4399 37315
rect 4614 37312 4620 37324
rect 4387 37284 4620 37312
rect 4387 37281 4399 37284
rect 4341 37275 4399 37281
rect 4614 37272 4620 37284
rect 4672 37272 4678 37324
rect 8389 37315 8447 37321
rect 8389 37281 8401 37315
rect 8435 37312 8447 37315
rect 8956 37312 8984 37411
rect 16022 37408 16028 37420
rect 16080 37408 16086 37460
rect 19426 37448 19432 37460
rect 19387 37420 19432 37448
rect 19426 37408 19432 37420
rect 19484 37408 19490 37460
rect 19797 37451 19855 37457
rect 19797 37417 19809 37451
rect 19843 37448 19855 37451
rect 19978 37448 19984 37460
rect 19843 37420 19984 37448
rect 19843 37417 19855 37420
rect 19797 37411 19855 37417
rect 19978 37408 19984 37420
rect 20036 37448 20042 37460
rect 20714 37448 20720 37460
rect 20036 37420 20720 37448
rect 20036 37408 20042 37420
rect 20714 37408 20720 37420
rect 20772 37408 20778 37460
rect 20806 37408 20812 37460
rect 20864 37448 20870 37460
rect 22097 37451 22155 37457
rect 22097 37448 22109 37451
rect 20864 37420 22109 37448
rect 20864 37408 20870 37420
rect 22097 37417 22109 37420
rect 22143 37417 22155 37451
rect 23382 37448 23388 37460
rect 23343 37420 23388 37448
rect 22097 37411 22155 37417
rect 23382 37408 23388 37420
rect 23440 37408 23446 37460
rect 24486 37448 24492 37460
rect 24447 37420 24492 37448
rect 24486 37408 24492 37420
rect 24544 37408 24550 37460
rect 25777 37451 25835 37457
rect 25777 37417 25789 37451
rect 25823 37448 25835 37451
rect 26234 37448 26240 37460
rect 25823 37420 26240 37448
rect 25823 37417 25835 37420
rect 25777 37411 25835 37417
rect 26234 37408 26240 37420
rect 26292 37408 26298 37460
rect 28810 37408 28816 37460
rect 28868 37448 28874 37460
rect 28997 37451 29055 37457
rect 28997 37448 29009 37451
rect 28868 37420 29009 37448
rect 28868 37408 28874 37420
rect 28997 37417 29009 37420
rect 29043 37417 29055 37451
rect 28997 37411 29055 37417
rect 31846 37408 31852 37460
rect 31904 37448 31910 37460
rect 34425 37451 34483 37457
rect 34425 37448 34437 37451
rect 31904 37420 34437 37448
rect 31904 37408 31910 37420
rect 34425 37417 34437 37420
rect 34471 37417 34483 37451
rect 40037 37451 40095 37457
rect 40037 37448 40049 37451
rect 34425 37411 34483 37417
rect 34532 37420 40049 37448
rect 13262 37340 13268 37392
rect 13320 37380 13326 37392
rect 34532 37380 34560 37420
rect 40037 37417 40049 37420
rect 40083 37448 40095 37451
rect 40310 37448 40316 37460
rect 40083 37420 40316 37448
rect 40083 37417 40095 37420
rect 40037 37411 40095 37417
rect 40310 37408 40316 37420
rect 40368 37408 40374 37460
rect 40862 37448 40868 37460
rect 40823 37420 40868 37448
rect 40862 37408 40868 37420
rect 40920 37408 40926 37460
rect 41414 37408 41420 37460
rect 41472 37448 41478 37460
rect 47946 37448 47952 37460
rect 41472 37420 47952 37448
rect 41472 37408 41478 37420
rect 47946 37408 47952 37420
rect 48004 37408 48010 37460
rect 51166 37408 51172 37460
rect 51224 37448 51230 37460
rect 57974 37448 57980 37460
rect 51224 37420 57560 37448
rect 57935 37420 57980 37448
rect 51224 37408 51230 37420
rect 37734 37380 37740 37392
rect 13320 37352 34560 37380
rect 36372 37352 37740 37380
rect 13320 37340 13326 37352
rect 8435 37284 8984 37312
rect 8435 37281 8447 37284
rect 8389 37275 8447 37281
rect 12158 37272 12164 37324
rect 12216 37312 12222 37324
rect 12437 37315 12495 37321
rect 12437 37312 12449 37315
rect 12216 37284 12449 37312
rect 12216 37272 12222 37284
rect 12437 37281 12449 37284
rect 12483 37281 12495 37315
rect 12437 37275 12495 37281
rect 12529 37315 12587 37321
rect 12529 37281 12541 37315
rect 12575 37312 12587 37315
rect 13173 37315 13231 37321
rect 13173 37312 13185 37315
rect 12575 37284 13185 37312
rect 12575 37281 12587 37284
rect 12529 37275 12587 37281
rect 13173 37281 13185 37284
rect 13219 37312 13231 37315
rect 13909 37315 13967 37321
rect 13909 37312 13921 37315
rect 13219 37284 13921 37312
rect 13219 37281 13231 37284
rect 13173 37275 13231 37281
rect 13909 37281 13921 37284
rect 13955 37312 13967 37315
rect 14550 37312 14556 37324
rect 13955 37284 14556 37312
rect 13955 37281 13967 37284
rect 13909 37275 13967 37281
rect 14550 37272 14556 37284
rect 14608 37272 14614 37324
rect 18141 37315 18199 37321
rect 18141 37281 18153 37315
rect 18187 37312 18199 37315
rect 18230 37312 18236 37324
rect 18187 37284 18236 37312
rect 18187 37281 18199 37284
rect 18141 37275 18199 37281
rect 18230 37272 18236 37284
rect 18288 37272 18294 37324
rect 18414 37312 18420 37324
rect 18327 37284 18420 37312
rect 18414 37272 18420 37284
rect 18472 37312 18478 37324
rect 18782 37312 18788 37324
rect 18472 37284 18788 37312
rect 18472 37272 18478 37284
rect 18782 37272 18788 37284
rect 18840 37312 18846 37324
rect 18969 37315 19027 37321
rect 18969 37312 18981 37315
rect 18840 37284 18981 37312
rect 18840 37272 18846 37284
rect 18969 37281 18981 37284
rect 19015 37281 19027 37315
rect 18969 37275 19027 37281
rect 19153 37315 19211 37321
rect 19153 37281 19165 37315
rect 19199 37312 19211 37315
rect 19199 37284 19748 37312
rect 19199 37281 19211 37284
rect 19153 37275 19211 37281
rect 4065 37247 4123 37253
rect 4065 37213 4077 37247
rect 4111 37244 4123 37247
rect 4246 37244 4252 37256
rect 4111 37216 4252 37244
rect 4111 37213 4123 37216
rect 4065 37207 4123 37213
rect 4246 37204 4252 37216
rect 4304 37244 4310 37256
rect 4798 37244 4804 37256
rect 4304 37216 4804 37244
rect 4304 37204 4310 37216
rect 4798 37204 4804 37216
rect 4856 37244 4862 37256
rect 5813 37247 5871 37253
rect 5813 37244 5825 37247
rect 4856 37216 5825 37244
rect 4856 37204 4862 37216
rect 5813 37213 5825 37216
rect 5859 37213 5871 37247
rect 5813 37207 5871 37213
rect 8938 37204 8944 37256
rect 8996 37244 9002 37256
rect 8996 37216 13768 37244
rect 8996 37204 9002 37216
rect 10042 37136 10048 37188
rect 10100 37176 10106 37188
rect 13630 37176 13636 37188
rect 10100 37148 13636 37176
rect 10100 37136 10106 37148
rect 13630 37136 13636 37148
rect 13688 37136 13694 37188
rect 13740 37176 13768 37216
rect 13814 37204 13820 37256
rect 13872 37244 13878 37256
rect 19720 37244 19748 37284
rect 19794 37272 19800 37324
rect 19852 37312 19858 37324
rect 21082 37312 21088 37324
rect 19852 37284 21088 37312
rect 19852 37272 19858 37284
rect 21082 37272 21088 37284
rect 21140 37312 21146 37324
rect 21637 37315 21695 37321
rect 21637 37312 21649 37315
rect 21140 37284 21649 37312
rect 21140 37272 21146 37284
rect 21637 37281 21649 37284
rect 21683 37281 21695 37315
rect 21818 37312 21824 37324
rect 21779 37284 21824 37312
rect 21637 37275 21695 37281
rect 21818 37272 21824 37284
rect 21876 37312 21882 37324
rect 22925 37315 22983 37321
rect 21876 37284 22232 37312
rect 21876 37272 21882 37284
rect 19978 37244 19984 37256
rect 13872 37216 13917 37244
rect 19720 37216 19984 37244
rect 13872 37204 13878 37216
rect 19978 37204 19984 37216
rect 20036 37204 20042 37256
rect 20898 37244 20904 37256
rect 20859 37216 20904 37244
rect 20898 37204 20904 37216
rect 20956 37204 20962 37256
rect 22204 37244 22232 37284
rect 22925 37281 22937 37315
rect 22971 37312 22983 37315
rect 23201 37315 23259 37321
rect 23201 37312 23213 37315
rect 22971 37284 23213 37312
rect 22971 37281 22983 37284
rect 22925 37275 22983 37281
rect 23201 37281 23213 37284
rect 23247 37312 23259 37315
rect 24762 37312 24768 37324
rect 23247 37284 24768 37312
rect 23247 37281 23259 37284
rect 23201 37275 23259 37281
rect 24762 37272 24768 37284
rect 24820 37272 24826 37324
rect 25038 37312 25044 37324
rect 24999 37284 25044 37312
rect 25038 37272 25044 37284
rect 25096 37272 25102 37324
rect 25406 37312 25412 37324
rect 25367 37284 25412 37312
rect 25406 37272 25412 37284
rect 25464 37272 25470 37324
rect 25593 37315 25651 37321
rect 25593 37281 25605 37315
rect 25639 37312 25651 37315
rect 26234 37312 26240 37324
rect 25639 37284 26240 37312
rect 25639 37281 25651 37284
rect 25593 37275 25651 37281
rect 26234 37272 26240 37284
rect 26292 37272 26298 37324
rect 27338 37312 27344 37324
rect 27299 37284 27344 37312
rect 27338 37272 27344 37284
rect 27396 37312 27402 37324
rect 27525 37315 27583 37321
rect 27525 37312 27537 37315
rect 27396 37284 27537 37312
rect 27396 37272 27402 37284
rect 27525 37281 27537 37284
rect 27571 37281 27583 37315
rect 27525 37275 27583 37281
rect 27709 37315 27767 37321
rect 27709 37281 27721 37315
rect 27755 37312 27767 37315
rect 27798 37312 27804 37324
rect 27755 37284 27804 37312
rect 27755 37281 27767 37284
rect 27709 37275 27767 37281
rect 27798 37272 27804 37284
rect 27856 37312 27862 37324
rect 28261 37315 28319 37321
rect 28261 37312 28273 37315
rect 27856 37284 28273 37312
rect 27856 37272 27862 37284
rect 28261 37281 28273 37284
rect 28307 37281 28319 37315
rect 28261 37275 28319 37281
rect 28445 37315 28503 37321
rect 28445 37281 28457 37315
rect 28491 37312 28503 37315
rect 28718 37312 28724 37324
rect 28491 37284 28724 37312
rect 28491 37281 28503 37284
rect 28445 37275 28503 37281
rect 28718 37272 28724 37284
rect 28776 37272 28782 37324
rect 32493 37315 32551 37321
rect 32493 37281 32505 37315
rect 32539 37312 32551 37315
rect 32677 37315 32735 37321
rect 32677 37312 32689 37315
rect 32539 37284 32689 37312
rect 32539 37281 32551 37284
rect 32493 37275 32551 37281
rect 32677 37281 32689 37284
rect 32723 37312 32735 37315
rect 32766 37312 32772 37324
rect 32723 37284 32772 37312
rect 32723 37281 32735 37284
rect 32677 37275 32735 37281
rect 32766 37272 32772 37284
rect 32824 37272 32830 37324
rect 34609 37315 34667 37321
rect 34609 37281 34621 37315
rect 34655 37312 34667 37315
rect 34698 37312 34704 37324
rect 34655 37284 34704 37312
rect 34655 37281 34667 37284
rect 34609 37275 34667 37281
rect 34698 37272 34704 37284
rect 34756 37272 34762 37324
rect 34790 37272 34796 37324
rect 34848 37312 34854 37324
rect 35161 37315 35219 37321
rect 35161 37312 35173 37315
rect 34848 37284 35173 37312
rect 34848 37272 34854 37284
rect 35161 37281 35173 37284
rect 35207 37312 35219 37315
rect 35621 37315 35679 37321
rect 35621 37312 35633 37315
rect 35207 37284 35633 37312
rect 35207 37281 35219 37284
rect 35161 37275 35219 37281
rect 35621 37281 35633 37284
rect 35667 37312 35679 37315
rect 35710 37312 35716 37324
rect 35667 37284 35716 37312
rect 35667 37281 35679 37284
rect 35621 37275 35679 37281
rect 35710 37272 35716 37284
rect 35768 37272 35774 37324
rect 36170 37312 36176 37324
rect 36131 37284 36176 37312
rect 36170 37272 36176 37284
rect 36228 37272 36234 37324
rect 36372 37321 36400 37352
rect 37734 37340 37740 37352
rect 37792 37340 37798 37392
rect 39390 37380 39396 37392
rect 39351 37352 39396 37380
rect 39390 37340 39396 37352
rect 39448 37340 39454 37392
rect 40218 37380 40224 37392
rect 40179 37352 40224 37380
rect 40218 37340 40224 37352
rect 40276 37340 40282 37392
rect 44637 37383 44695 37389
rect 44637 37380 44649 37383
rect 43640 37352 44649 37380
rect 36357 37315 36415 37321
rect 36357 37281 36369 37315
rect 36403 37281 36415 37315
rect 38013 37315 38071 37321
rect 38013 37312 38025 37315
rect 36357 37275 36415 37281
rect 36740 37284 38025 37312
rect 22465 37247 22523 37253
rect 22465 37244 22477 37247
rect 22204 37216 22477 37244
rect 22465 37213 22477 37216
rect 22511 37244 22523 37247
rect 24946 37244 24952 37256
rect 22511 37216 24952 37244
rect 22511 37213 22523 37216
rect 22465 37207 22523 37213
rect 24946 37204 24952 37216
rect 25004 37204 25010 37256
rect 25133 37247 25191 37253
rect 25133 37213 25145 37247
rect 25179 37244 25191 37247
rect 25961 37247 26019 37253
rect 25961 37244 25973 37247
rect 25179 37216 25973 37244
rect 25179 37213 25191 37216
rect 25133 37207 25191 37213
rect 25961 37213 25973 37216
rect 26007 37244 26019 37247
rect 26050 37244 26056 37256
rect 26007 37216 26056 37244
rect 26007 37213 26019 37216
rect 25961 37207 26019 37213
rect 26050 37204 26056 37216
rect 26108 37204 26114 37256
rect 28810 37204 28816 37256
rect 28868 37244 28874 37256
rect 35253 37247 35311 37253
rect 35253 37244 35265 37247
rect 28868 37216 35265 37244
rect 28868 37204 28874 37216
rect 35253 37213 35265 37216
rect 35299 37244 35311 37247
rect 35434 37244 35440 37256
rect 35299 37216 35440 37244
rect 35299 37213 35311 37216
rect 35253 37207 35311 37213
rect 35434 37204 35440 37216
rect 35492 37204 35498 37256
rect 36740 37253 36768 37284
rect 38013 37281 38025 37284
rect 38059 37281 38071 37315
rect 43640 37312 43668 37352
rect 44637 37349 44649 37352
rect 44683 37380 44695 37383
rect 44683 37352 44864 37380
rect 44683 37349 44695 37352
rect 44637 37343 44695 37349
rect 38013 37275 38071 37281
rect 38120 37284 39988 37312
rect 36725 37247 36783 37253
rect 36725 37213 36737 37247
rect 36771 37213 36783 37247
rect 37550 37244 37556 37256
rect 37511 37216 37556 37244
rect 36725 37207 36783 37213
rect 37550 37204 37556 37216
rect 37608 37204 37614 37256
rect 37734 37244 37740 37256
rect 37695 37216 37740 37244
rect 37734 37204 37740 37216
rect 37792 37244 37798 37256
rect 38120 37244 38148 37284
rect 37792 37216 38148 37244
rect 39960 37244 39988 37284
rect 40420 37284 43668 37312
rect 43809 37315 43867 37321
rect 40420 37244 40448 37284
rect 43809 37281 43821 37315
rect 43855 37312 43867 37315
rect 44726 37312 44732 37324
rect 43855 37284 44732 37312
rect 43855 37281 43867 37284
rect 43809 37275 43867 37281
rect 44726 37272 44732 37284
rect 44784 37272 44790 37324
rect 44836 37321 44864 37352
rect 45830 37340 45836 37392
rect 45888 37380 45894 37392
rect 48958 37380 48964 37392
rect 45888 37352 48964 37380
rect 45888 37340 45894 37352
rect 48958 37340 48964 37352
rect 49016 37340 49022 37392
rect 49068 37352 50936 37380
rect 44821 37315 44879 37321
rect 44821 37281 44833 37315
rect 44867 37281 44879 37315
rect 45097 37315 45155 37321
rect 45097 37312 45109 37315
rect 44821 37275 44879 37281
rect 44928 37284 45109 37312
rect 40586 37244 40592 37256
rect 39960 37216 40448 37244
rect 40547 37216 40592 37244
rect 37792 37204 37798 37216
rect 40586 37204 40592 37216
rect 40644 37204 40650 37256
rect 43901 37247 43959 37253
rect 43901 37213 43913 37247
rect 43947 37244 43959 37247
rect 43990 37244 43996 37256
rect 43947 37216 43996 37244
rect 43947 37213 43959 37216
rect 43901 37207 43959 37213
rect 43990 37204 43996 37216
rect 44048 37204 44054 37256
rect 44082 37204 44088 37256
rect 44140 37244 44146 37256
rect 44928 37244 44956 37284
rect 45097 37281 45109 37284
rect 45143 37281 45155 37315
rect 45097 37275 45155 37281
rect 46477 37315 46535 37321
rect 46477 37281 46489 37315
rect 46523 37312 46535 37315
rect 47854 37312 47860 37324
rect 46523 37284 47860 37312
rect 46523 37281 46535 37284
rect 46477 37275 46535 37281
rect 47854 37272 47860 37284
rect 47912 37272 47918 37324
rect 47946 37272 47952 37324
rect 48004 37312 48010 37324
rect 48590 37312 48596 37324
rect 48004 37284 48596 37312
rect 48004 37272 48010 37284
rect 48590 37272 48596 37284
rect 48648 37272 48654 37324
rect 48682 37272 48688 37324
rect 48740 37312 48746 37324
rect 49068 37321 49096 37352
rect 49053 37315 49111 37321
rect 49053 37312 49065 37315
rect 48740 37284 49065 37312
rect 48740 37272 48746 37284
rect 49053 37281 49065 37284
rect 49099 37281 49111 37315
rect 50062 37312 50068 37324
rect 50023 37284 50068 37312
rect 49053 37275 49111 37281
rect 50062 37272 50068 37284
rect 50120 37312 50126 37324
rect 50249 37315 50307 37321
rect 50249 37312 50261 37315
rect 50120 37284 50261 37312
rect 50120 37272 50126 37284
rect 50249 37281 50261 37284
rect 50295 37281 50307 37315
rect 50249 37275 50307 37281
rect 50433 37315 50491 37321
rect 50433 37281 50445 37315
rect 50479 37312 50491 37315
rect 50798 37312 50804 37324
rect 50479 37284 50804 37312
rect 50479 37281 50491 37284
rect 50433 37275 50491 37281
rect 50798 37272 50804 37284
rect 50856 37272 50862 37324
rect 50908 37321 50936 37352
rect 51534 37340 51540 37392
rect 51592 37380 51598 37392
rect 52362 37380 52368 37392
rect 51592 37352 52368 37380
rect 51592 37340 51598 37352
rect 52362 37340 52368 37352
rect 52420 37340 52426 37392
rect 52914 37340 52920 37392
rect 52972 37380 52978 37392
rect 54573 37383 54631 37389
rect 54573 37380 54585 37383
rect 52972 37352 54585 37380
rect 52972 37340 52978 37352
rect 54573 37349 54585 37352
rect 54619 37349 54631 37383
rect 55309 37383 55367 37389
rect 55309 37380 55321 37383
rect 54573 37343 54631 37349
rect 54680 37352 55321 37380
rect 50893 37315 50951 37321
rect 50893 37281 50905 37315
rect 50939 37281 50951 37315
rect 50893 37275 50951 37281
rect 50985 37315 51043 37321
rect 50985 37281 50997 37315
rect 51031 37312 51043 37315
rect 51997 37315 52055 37321
rect 51997 37312 52009 37315
rect 51031 37284 52009 37312
rect 51031 37281 51043 37284
rect 50985 37275 51043 37281
rect 51997 37281 52009 37284
rect 52043 37312 52055 37315
rect 52043 37284 52500 37312
rect 52043 37281 52055 37284
rect 51997 37275 52055 37281
rect 44140 37216 44956 37244
rect 52472 37244 52500 37284
rect 52546 37272 52552 37324
rect 52604 37312 52610 37324
rect 54680 37312 54708 37352
rect 55309 37349 55321 37352
rect 55355 37349 55367 37383
rect 55309 37343 55367 37349
rect 56318 37340 56324 37392
rect 56376 37380 56382 37392
rect 57532 37380 57560 37420
rect 57974 37408 57980 37420
rect 58032 37408 58038 37460
rect 60458 37408 60464 37460
rect 60516 37448 60522 37460
rect 69106 37448 69112 37460
rect 60516 37420 69112 37448
rect 60516 37408 60522 37420
rect 69106 37408 69112 37420
rect 69164 37408 69170 37460
rect 69566 37448 69572 37460
rect 69527 37420 69572 37448
rect 69566 37408 69572 37420
rect 69624 37408 69630 37460
rect 70673 37451 70731 37457
rect 70673 37448 70685 37451
rect 69952 37420 70685 37448
rect 65426 37380 65432 37392
rect 56376 37352 57468 37380
rect 57532 37352 65432 37380
rect 56376 37340 56382 37352
rect 55122 37312 55128 37324
rect 52604 37284 54708 37312
rect 54772 37284 55128 37312
rect 52604 37272 52610 37284
rect 53834 37244 53840 37256
rect 52472 37216 53840 37244
rect 44140 37204 44146 37216
rect 53834 37204 53840 37216
rect 53892 37204 53898 37256
rect 54772 37253 54800 37284
rect 55122 37272 55128 37284
rect 55180 37272 55186 37324
rect 56965 37315 57023 37321
rect 56965 37312 56977 37315
rect 56428 37284 56977 37312
rect 54720 37247 54800 37253
rect 54720 37213 54732 37247
rect 54766 37216 54800 37247
rect 54938 37244 54944 37256
rect 54899 37216 54944 37244
rect 54766 37213 54778 37216
rect 54720 37207 54778 37213
rect 54938 37204 54944 37216
rect 54996 37204 55002 37256
rect 56226 37244 56232 37256
rect 56187 37216 56232 37244
rect 56226 37204 56232 37216
rect 56284 37244 56290 37256
rect 56428 37253 56456 37284
rect 56965 37281 56977 37284
rect 57011 37312 57023 37315
rect 57330 37312 57336 37324
rect 57011 37284 57336 37312
rect 57011 37281 57023 37284
rect 56965 37275 57023 37281
rect 57330 37272 57336 37284
rect 57388 37272 57394 37324
rect 57440 37321 57468 37352
rect 65426 37340 65432 37352
rect 65484 37340 65490 37392
rect 57425 37315 57483 37321
rect 57425 37281 57437 37315
rect 57471 37281 57483 37315
rect 57425 37275 57483 37281
rect 57514 37272 57520 37324
rect 57572 37312 57578 37324
rect 62209 37315 62267 37321
rect 62209 37312 62221 37315
rect 57572 37284 62221 37312
rect 57572 37272 57578 37284
rect 62209 37281 62221 37284
rect 62255 37312 62267 37315
rect 62393 37315 62451 37321
rect 62393 37312 62405 37315
rect 62255 37284 62405 37312
rect 62255 37281 62267 37284
rect 62209 37275 62267 37281
rect 62393 37281 62405 37284
rect 62439 37312 62451 37315
rect 62945 37315 63003 37321
rect 62945 37312 62957 37315
rect 62439 37284 62957 37312
rect 62439 37281 62451 37284
rect 62393 37275 62451 37281
rect 62945 37281 62957 37284
rect 62991 37312 63003 37315
rect 63497 37315 63555 37321
rect 63497 37312 63509 37315
rect 62991 37284 63509 37312
rect 62991 37281 63003 37284
rect 62945 37275 63003 37281
rect 63497 37281 63509 37284
rect 63543 37281 63555 37315
rect 63497 37275 63555 37281
rect 63681 37315 63739 37321
rect 63681 37281 63693 37315
rect 63727 37312 63739 37315
rect 63862 37312 63868 37324
rect 63727 37284 63868 37312
rect 63727 37281 63739 37284
rect 63681 37275 63739 37281
rect 63862 37272 63868 37284
rect 63920 37312 63926 37324
rect 69952 37321 69980 37420
rect 70673 37417 70685 37420
rect 70719 37448 70731 37451
rect 70762 37448 70768 37460
rect 70719 37420 70768 37448
rect 70719 37417 70731 37420
rect 70673 37411 70731 37417
rect 70762 37408 70768 37420
rect 70820 37408 70826 37460
rect 70857 37451 70915 37457
rect 70857 37417 70869 37451
rect 70903 37448 70915 37451
rect 71222 37448 71228 37460
rect 70903 37420 71228 37448
rect 70903 37417 70915 37420
rect 70857 37411 70915 37417
rect 69937 37315 69995 37321
rect 63920 37284 64828 37312
rect 63920 37272 63926 37284
rect 56413 37247 56471 37253
rect 56413 37244 56425 37247
rect 56284 37216 56425 37244
rect 56284 37204 56290 37216
rect 56413 37213 56425 37216
rect 56459 37213 56471 37247
rect 56413 37207 56471 37213
rect 56594 37204 56600 37256
rect 56652 37244 56658 37256
rect 56781 37247 56839 37253
rect 56781 37244 56793 37247
rect 56652 37216 56793 37244
rect 56652 37204 56658 37216
rect 56781 37213 56793 37216
rect 56827 37213 56839 37247
rect 56781 37207 56839 37213
rect 62574 37204 62580 37256
rect 62632 37244 62638 37256
rect 62761 37247 62819 37253
rect 62761 37244 62773 37247
rect 62632 37216 62773 37244
rect 62632 37204 62638 37216
rect 62761 37213 62773 37216
rect 62807 37213 62819 37247
rect 64800 37244 64828 37284
rect 69937 37281 69949 37315
rect 69983 37281 69995 37315
rect 69937 37275 69995 37281
rect 70305 37315 70363 37321
rect 70305 37281 70317 37315
rect 70351 37312 70363 37315
rect 70872 37312 70900 37411
rect 71222 37408 71228 37420
rect 71280 37408 71286 37460
rect 71685 37451 71743 37457
rect 71685 37417 71697 37451
rect 71731 37448 71743 37451
rect 72234 37448 72240 37460
rect 71731 37420 72240 37448
rect 71731 37417 71743 37420
rect 71685 37411 71743 37417
rect 72234 37408 72240 37420
rect 72292 37408 72298 37460
rect 72786 37448 72792 37460
rect 72747 37420 72792 37448
rect 72786 37408 72792 37420
rect 72844 37408 72850 37460
rect 73154 37408 73160 37460
rect 73212 37448 73218 37460
rect 75365 37451 75423 37457
rect 75365 37448 75377 37451
rect 73212 37420 75377 37448
rect 73212 37408 73218 37420
rect 75365 37417 75377 37420
rect 75411 37417 75423 37451
rect 75365 37411 75423 37417
rect 82814 37408 82820 37460
rect 82872 37448 82878 37460
rect 83185 37451 83243 37457
rect 83185 37448 83197 37451
rect 82872 37420 83197 37448
rect 82872 37408 82878 37420
rect 83185 37417 83197 37420
rect 83231 37417 83243 37451
rect 83185 37411 83243 37417
rect 88702 37408 88708 37460
rect 88760 37448 88766 37460
rect 96706 37448 96712 37460
rect 88760 37420 96712 37448
rect 88760 37408 88766 37420
rect 71774 37340 71780 37392
rect 71832 37380 71838 37392
rect 72804 37380 72832 37408
rect 71832 37352 72832 37380
rect 82909 37383 82967 37389
rect 71832 37340 71838 37352
rect 70351 37284 70900 37312
rect 70351 37281 70363 37284
rect 70305 37275 70363 37281
rect 71498 37272 71504 37324
rect 71556 37312 71562 37324
rect 72068 37321 72096 37352
rect 82909 37349 82921 37383
rect 82955 37380 82967 37383
rect 82998 37380 83004 37392
rect 82955 37352 83004 37380
rect 82955 37349 82967 37352
rect 82909 37343 82967 37349
rect 82998 37340 83004 37352
rect 83056 37340 83062 37392
rect 85574 37380 85580 37392
rect 85040 37352 85580 37380
rect 71869 37315 71927 37321
rect 71869 37312 71881 37315
rect 71556 37284 71881 37312
rect 71556 37272 71562 37284
rect 71869 37281 71881 37284
rect 71915 37281 71927 37315
rect 71869 37275 71927 37281
rect 72053 37315 72111 37321
rect 72053 37281 72065 37315
rect 72099 37281 72111 37315
rect 72053 37275 72111 37281
rect 72421 37315 72479 37321
rect 72421 37281 72433 37315
rect 72467 37312 72479 37315
rect 72970 37312 72976 37324
rect 72467 37284 72976 37312
rect 72467 37281 72479 37284
rect 72421 37275 72479 37281
rect 72970 37272 72976 37284
rect 73028 37272 73034 37324
rect 75181 37315 75239 37321
rect 75181 37281 75193 37315
rect 75227 37312 75239 37315
rect 75914 37312 75920 37324
rect 75227 37284 75920 37312
rect 75227 37281 75239 37284
rect 75181 37275 75239 37281
rect 75914 37272 75920 37284
rect 75972 37272 75978 37324
rect 82817 37315 82875 37321
rect 82817 37281 82829 37315
rect 82863 37312 82875 37315
rect 83093 37315 83151 37321
rect 83093 37312 83105 37315
rect 82863 37284 83105 37312
rect 82863 37281 82875 37284
rect 82817 37275 82875 37281
rect 83093 37281 83105 37284
rect 83139 37312 83151 37315
rect 83182 37312 83188 37324
rect 83139 37284 83188 37312
rect 83139 37281 83151 37284
rect 83093 37275 83151 37281
rect 83182 37272 83188 37284
rect 83240 37272 83246 37324
rect 85040 37321 85068 37352
rect 85574 37340 85580 37352
rect 85632 37340 85638 37392
rect 85025 37315 85083 37321
rect 85025 37281 85037 37315
rect 85071 37281 85083 37315
rect 85025 37275 85083 37281
rect 85301 37315 85359 37321
rect 85301 37281 85313 37315
rect 85347 37312 85359 37315
rect 86218 37312 86224 37324
rect 85347 37284 86224 37312
rect 85347 37281 85359 37284
rect 85301 37275 85359 37281
rect 86218 37272 86224 37284
rect 86276 37272 86282 37324
rect 86862 37272 86868 37324
rect 86920 37312 86926 37324
rect 89441 37315 89499 37321
rect 89441 37312 89453 37315
rect 86920 37284 89453 37312
rect 86920 37272 86926 37284
rect 89441 37281 89453 37284
rect 89487 37281 89499 37315
rect 89441 37275 89499 37281
rect 69750 37244 69756 37256
rect 64800 37216 67588 37244
rect 69711 37216 69756 37244
rect 62761 37207 62819 37213
rect 20806 37176 20812 37188
rect 13740 37148 20812 37176
rect 20806 37136 20812 37148
rect 20864 37136 20870 37188
rect 22278 37136 22284 37188
rect 22336 37176 22342 37188
rect 22925 37179 22983 37185
rect 22925 37176 22937 37179
rect 22336 37148 22937 37176
rect 22336 37136 22342 37148
rect 22925 37145 22937 37148
rect 22971 37176 22983 37179
rect 23017 37179 23075 37185
rect 23017 37176 23029 37179
rect 22971 37148 23029 37176
rect 22971 37145 22983 37148
rect 22925 37139 22983 37145
rect 23017 37145 23029 37148
rect 23063 37145 23075 37179
rect 23017 37139 23075 37145
rect 28721 37179 28779 37185
rect 28721 37145 28733 37179
rect 28767 37176 28779 37179
rect 67450 37176 67456 37188
rect 28767 37148 37596 37176
rect 28767 37145 28779 37148
rect 28721 37139 28779 37145
rect 4062 37068 4068 37120
rect 4120 37108 4126 37120
rect 5445 37111 5503 37117
rect 5445 37108 5457 37111
rect 4120 37080 5457 37108
rect 4120 37068 4126 37080
rect 5445 37077 5457 37080
rect 5491 37077 5503 37111
rect 5445 37071 5503 37077
rect 7650 37068 7656 37120
rect 7708 37108 7714 37120
rect 8481 37111 8539 37117
rect 8481 37108 8493 37111
rect 7708 37080 8493 37108
rect 7708 37068 7714 37080
rect 8481 37077 8493 37080
rect 8527 37077 8539 37111
rect 8481 37071 8539 37077
rect 12526 37068 12532 37120
rect 12584 37108 12590 37120
rect 12713 37111 12771 37117
rect 12713 37108 12725 37111
rect 12584 37080 12725 37108
rect 12584 37068 12590 37080
rect 12713 37077 12725 37080
rect 12759 37077 12771 37111
rect 12713 37071 12771 37077
rect 12894 37068 12900 37120
rect 12952 37108 12958 37120
rect 14093 37111 14151 37117
rect 14093 37108 14105 37111
rect 12952 37080 14105 37108
rect 12952 37068 12958 37080
rect 14093 37077 14105 37080
rect 14139 37077 14151 37111
rect 14093 37071 14151 37077
rect 18230 37068 18236 37120
rect 18288 37108 18294 37120
rect 20625 37111 20683 37117
rect 20625 37108 20637 37111
rect 18288 37080 20637 37108
rect 18288 37068 18294 37080
rect 20625 37077 20637 37080
rect 20671 37108 20683 37111
rect 20898 37108 20904 37120
rect 20671 37080 20904 37108
rect 20671 37077 20683 37080
rect 20625 37071 20683 37077
rect 20898 37068 20904 37080
rect 20956 37068 20962 37120
rect 20990 37068 20996 37120
rect 21048 37108 21054 37120
rect 31754 37108 31760 37120
rect 21048 37080 31760 37108
rect 21048 37068 21054 37080
rect 31754 37068 31760 37080
rect 31812 37068 31818 37120
rect 31938 37068 31944 37120
rect 31996 37108 32002 37120
rect 32674 37108 32680 37120
rect 31996 37080 32680 37108
rect 31996 37068 32002 37080
rect 32674 37068 32680 37080
rect 32732 37068 32738 37120
rect 32861 37111 32919 37117
rect 32861 37077 32873 37111
rect 32907 37108 32919 37111
rect 35986 37108 35992 37120
rect 32907 37080 35992 37108
rect 32907 37077 32919 37080
rect 32861 37071 32919 37077
rect 35986 37068 35992 37080
rect 36044 37068 36050 37120
rect 37568 37108 37596 37148
rect 38672 37148 44864 37176
rect 38672 37108 38700 37148
rect 37568 37080 38700 37108
rect 40310 37068 40316 37120
rect 40368 37117 40374 37120
rect 40368 37111 40417 37117
rect 40368 37077 40371 37111
rect 40405 37077 40417 37111
rect 40494 37108 40500 37120
rect 40455 37080 40500 37108
rect 40368 37071 40417 37077
rect 40368 37068 40374 37071
rect 40494 37068 40500 37080
rect 40552 37068 40558 37120
rect 44836 37108 44864 37148
rect 45756 37148 67456 37176
rect 45756 37108 45784 37148
rect 67450 37136 67456 37148
rect 67508 37136 67514 37188
rect 44836 37080 45784 37108
rect 48498 37068 48504 37120
rect 48556 37108 48562 37120
rect 49142 37108 49148 37120
rect 48556 37080 49148 37108
rect 48556 37068 48562 37080
rect 49142 37068 49148 37080
rect 49200 37068 49206 37120
rect 49234 37068 49240 37120
rect 49292 37108 49298 37120
rect 49329 37111 49387 37117
rect 49329 37108 49341 37111
rect 49292 37080 49341 37108
rect 49292 37068 49298 37080
rect 49329 37077 49341 37080
rect 49375 37077 49387 37111
rect 49329 37071 49387 37077
rect 50798 37068 50804 37120
rect 50856 37108 50862 37120
rect 51445 37111 51503 37117
rect 51445 37108 51457 37111
rect 50856 37080 51457 37108
rect 50856 37068 50862 37080
rect 51445 37077 51457 37080
rect 51491 37077 51503 37111
rect 51445 37071 51503 37077
rect 51626 37068 51632 37120
rect 51684 37108 51690 37120
rect 51721 37111 51779 37117
rect 51721 37108 51733 37111
rect 51684 37080 51733 37108
rect 51684 37068 51690 37080
rect 51721 37077 51733 37080
rect 51767 37077 51779 37111
rect 54846 37108 54852 37120
rect 54807 37080 54852 37108
rect 51721 37071 51779 37077
rect 54846 37068 54852 37080
rect 54904 37068 54910 37120
rect 56594 37108 56600 37120
rect 56555 37080 56600 37108
rect 56594 37068 56600 37080
rect 56652 37068 56658 37120
rect 62574 37108 62580 37120
rect 62535 37080 62580 37108
rect 62574 37068 62580 37080
rect 62632 37068 62638 37120
rect 63957 37111 64015 37117
rect 63957 37077 63969 37111
rect 64003 37108 64015 37111
rect 64782 37108 64788 37120
rect 64003 37080 64788 37108
rect 64003 37077 64015 37080
rect 63957 37071 64015 37077
rect 64782 37068 64788 37080
rect 64840 37068 64846 37120
rect 67560 37108 67588 37216
rect 69750 37204 69756 37216
rect 69808 37204 69814 37256
rect 70213 37247 70271 37253
rect 70213 37213 70225 37247
rect 70259 37213 70271 37247
rect 72326 37244 72332 37256
rect 72287 37216 72332 37244
rect 70213 37207 70271 37213
rect 69290 37136 69296 37188
rect 69348 37176 69354 37188
rect 70228 37176 70256 37207
rect 72326 37204 72332 37216
rect 72384 37204 72390 37256
rect 77021 37247 77079 37253
rect 77021 37244 77033 37247
rect 76760 37216 77033 37244
rect 69348 37148 70256 37176
rect 69348 37136 69354 37148
rect 76760 37120 76788 37216
rect 77021 37213 77033 37216
rect 77067 37213 77079 37247
rect 77021 37207 77079 37213
rect 77297 37247 77355 37253
rect 77297 37213 77309 37247
rect 77343 37244 77355 37247
rect 77386 37244 77392 37256
rect 77343 37216 77392 37244
rect 77343 37213 77355 37216
rect 77297 37207 77355 37213
rect 77386 37204 77392 37216
rect 77444 37204 77450 37256
rect 84470 37244 84476 37256
rect 84431 37216 84476 37244
rect 84470 37204 84476 37216
rect 84528 37204 84534 37256
rect 85485 37247 85543 37253
rect 85485 37213 85497 37247
rect 85531 37213 85543 37247
rect 85485 37207 85543 37213
rect 85500 37120 85528 37207
rect 89456 37176 89484 37275
rect 89548 37253 89576 37420
rect 90177 37383 90235 37389
rect 90177 37349 90189 37383
rect 90223 37380 90235 37383
rect 91002 37380 91008 37392
rect 90223 37352 91008 37380
rect 90223 37349 90235 37352
rect 90177 37343 90235 37349
rect 91002 37340 91008 37352
rect 91060 37340 91066 37392
rect 91278 37380 91284 37392
rect 91239 37352 91284 37380
rect 91278 37340 91284 37352
rect 91336 37340 91342 37392
rect 91465 37383 91523 37389
rect 91465 37349 91477 37383
rect 91511 37380 91523 37383
rect 91554 37380 91560 37392
rect 91511 37352 91560 37380
rect 91511 37349 91523 37352
rect 91465 37343 91523 37349
rect 91554 37340 91560 37352
rect 91612 37340 91618 37392
rect 89714 37272 89720 37324
rect 89772 37312 89778 37324
rect 91296 37312 91324 37340
rect 94240 37321 94268 37420
rect 96706 37408 96712 37420
rect 96764 37408 96770 37460
rect 94590 37340 94596 37392
rect 94648 37380 94654 37392
rect 95237 37383 95295 37389
rect 95237 37380 95249 37383
rect 94648 37352 95249 37380
rect 94648 37340 94654 37352
rect 95237 37349 95249 37352
rect 95283 37349 95295 37383
rect 95237 37343 95295 37349
rect 91649 37315 91707 37321
rect 91649 37312 91661 37315
rect 89772 37284 89817 37312
rect 91296 37284 91661 37312
rect 89772 37272 89778 37284
rect 91649 37281 91661 37284
rect 91695 37281 91707 37315
rect 91649 37275 91707 37281
rect 94041 37315 94099 37321
rect 94041 37281 94053 37315
rect 94087 37312 94099 37315
rect 94225 37315 94283 37321
rect 94087 37284 94176 37312
rect 94087 37281 94099 37284
rect 94041 37275 94099 37281
rect 89533 37247 89591 37253
rect 89533 37213 89545 37247
rect 89579 37213 89591 37247
rect 89533 37207 89591 37213
rect 92017 37247 92075 37253
rect 92017 37213 92029 37247
rect 92063 37244 92075 37247
rect 93578 37244 93584 37256
rect 92063 37216 93584 37244
rect 92063 37213 92075 37216
rect 92017 37207 92075 37213
rect 93578 37204 93584 37216
rect 93636 37204 93642 37256
rect 94148 37176 94176 37284
rect 94225 37281 94237 37315
rect 94271 37281 94283 37315
rect 95252 37312 95280 37343
rect 95421 37315 95479 37321
rect 95421 37312 95433 37315
rect 95252 37284 95433 37312
rect 94225 37275 94283 37281
rect 95421 37281 95433 37284
rect 95467 37281 95479 37315
rect 95694 37312 95700 37324
rect 95655 37284 95700 37312
rect 95421 37275 95479 37281
rect 95694 37272 95700 37284
rect 95752 37272 95758 37324
rect 94593 37247 94651 37253
rect 94593 37213 94605 37247
rect 94639 37244 94651 37247
rect 95234 37244 95240 37256
rect 94639 37216 95240 37244
rect 94639 37213 94651 37216
rect 94593 37207 94651 37213
rect 95234 37204 95240 37216
rect 95292 37204 95298 37256
rect 95142 37176 95148 37188
rect 89456 37148 94084 37176
rect 94148 37148 95148 37176
rect 70486 37108 70492 37120
rect 67560 37080 70492 37108
rect 70486 37068 70492 37080
rect 70544 37068 70550 37120
rect 72970 37108 72976 37120
rect 72931 37080 72976 37108
rect 72970 37068 72976 37080
rect 73028 37068 73034 37120
rect 76742 37108 76748 37120
rect 76703 37080 76748 37108
rect 76742 37068 76748 37080
rect 76800 37068 76806 37120
rect 78398 37108 78404 37120
rect 78359 37080 78404 37108
rect 78398 37068 78404 37080
rect 78456 37068 78462 37120
rect 84286 37108 84292 37120
rect 84247 37080 84292 37108
rect 84286 37068 84292 37080
rect 84344 37108 84350 37120
rect 85482 37108 85488 37120
rect 84344 37080 85488 37108
rect 84344 37068 84350 37080
rect 85482 37068 85488 37080
rect 85540 37068 85546 37120
rect 87414 37068 87420 37120
rect 87472 37108 87478 37120
rect 89714 37108 89720 37120
rect 87472 37080 89720 37108
rect 87472 37068 87478 37080
rect 89714 37068 89720 37080
rect 89772 37108 89778 37120
rect 90361 37111 90419 37117
rect 90361 37108 90373 37111
rect 89772 37080 90373 37108
rect 89772 37068 89778 37080
rect 90361 37077 90373 37080
rect 90407 37108 90419 37111
rect 93670 37108 93676 37120
rect 90407 37080 93676 37108
rect 90407 37077 90419 37080
rect 90361 37071 90419 37077
rect 93670 37068 93676 37080
rect 93728 37068 93734 37120
rect 94056 37108 94084 37148
rect 95142 37136 95148 37148
rect 95200 37136 95206 37188
rect 95050 37108 95056 37120
rect 94056 37080 95056 37108
rect 95050 37068 95056 37080
rect 95108 37068 95114 37120
rect 96985 37111 97043 37117
rect 96985 37077 96997 37111
rect 97031 37108 97043 37111
rect 97074 37108 97080 37120
rect 97031 37080 97080 37108
rect 97031 37077 97043 37080
rect 96985 37071 97043 37077
rect 97074 37068 97080 37080
rect 97132 37068 97138 37120
rect 1104 37018 105616 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 65686 37018
rect 65738 36966 65750 37018
rect 65802 36966 65814 37018
rect 65866 36966 65878 37018
rect 65930 36966 96406 37018
rect 96458 36966 96470 37018
rect 96522 36966 96534 37018
rect 96586 36966 96598 37018
rect 96650 36966 105616 37018
rect 1104 36944 105616 36966
rect 3234 36864 3240 36916
rect 3292 36904 3298 36916
rect 3881 36907 3939 36913
rect 3881 36904 3893 36907
rect 3292 36876 3893 36904
rect 3292 36864 3298 36876
rect 3881 36873 3893 36876
rect 3927 36873 3939 36907
rect 3881 36867 3939 36873
rect 3988 36876 12664 36904
rect 3694 36796 3700 36848
rect 3752 36836 3758 36848
rect 3988 36836 4016 36876
rect 9766 36836 9772 36848
rect 3752 36808 4016 36836
rect 5368 36808 9772 36836
rect 3752 36796 3758 36808
rect 2498 36768 2504 36780
rect 2411 36740 2504 36768
rect 2498 36728 2504 36740
rect 2556 36768 2562 36780
rect 4614 36768 4620 36780
rect 2556 36740 4620 36768
rect 2556 36728 2562 36740
rect 4614 36728 4620 36740
rect 4672 36728 4678 36780
rect 2777 36703 2835 36709
rect 2777 36669 2789 36703
rect 2823 36700 2835 36703
rect 4249 36703 4307 36709
rect 4249 36700 4261 36703
rect 2823 36672 4261 36700
rect 2823 36669 2835 36672
rect 2777 36663 2835 36669
rect 4249 36669 4261 36672
rect 4295 36700 4307 36703
rect 5368 36700 5396 36808
rect 9766 36796 9772 36808
rect 9824 36796 9830 36848
rect 10042 36836 10048 36848
rect 9876 36808 10048 36836
rect 8754 36728 8760 36780
rect 8812 36768 8818 36780
rect 9876 36777 9904 36808
rect 10042 36796 10048 36808
rect 10100 36796 10106 36848
rect 12636 36836 12664 36876
rect 12710 36864 12716 36916
rect 12768 36904 12774 36916
rect 28810 36904 28816 36916
rect 12768 36876 12813 36904
rect 12912 36876 28816 36904
rect 12768 36864 12774 36876
rect 12912 36836 12940 36876
rect 28810 36864 28816 36876
rect 28868 36864 28874 36916
rect 34790 36904 34796 36916
rect 28920 36876 34796 36904
rect 12636 36808 12940 36836
rect 13538 36796 13544 36848
rect 13596 36836 13602 36848
rect 14185 36839 14243 36845
rect 14185 36836 14197 36839
rect 13596 36808 14197 36836
rect 13596 36796 13602 36808
rect 14185 36805 14197 36808
rect 14231 36805 14243 36839
rect 14185 36799 14243 36805
rect 17037 36839 17095 36845
rect 17037 36805 17049 36839
rect 17083 36836 17095 36839
rect 18414 36836 18420 36848
rect 17083 36808 18420 36836
rect 17083 36805 17095 36808
rect 17037 36799 17095 36805
rect 18414 36796 18420 36808
rect 18472 36796 18478 36848
rect 22649 36839 22707 36845
rect 22649 36805 22661 36839
rect 22695 36836 22707 36839
rect 28920 36836 28948 36876
rect 34790 36864 34796 36876
rect 34848 36864 34854 36916
rect 35434 36864 35440 36916
rect 35492 36904 35498 36916
rect 35621 36907 35679 36913
rect 35621 36904 35633 36907
rect 35492 36876 35633 36904
rect 35492 36864 35498 36876
rect 35621 36873 35633 36876
rect 35667 36873 35679 36907
rect 36998 36904 37004 36916
rect 36959 36876 37004 36904
rect 35621 36867 35679 36873
rect 32030 36836 32036 36848
rect 22695 36808 28948 36836
rect 31404 36808 32036 36836
rect 22695 36805 22707 36808
rect 22649 36799 22707 36805
rect 9401 36771 9459 36777
rect 9401 36768 9413 36771
rect 8812 36740 9413 36768
rect 8812 36728 8818 36740
rect 9401 36737 9413 36740
rect 9447 36768 9459 36771
rect 9861 36771 9919 36777
rect 9447 36740 9812 36768
rect 9447 36737 9459 36740
rect 9401 36731 9459 36737
rect 4295 36672 5396 36700
rect 4295 36669 4307 36672
rect 4249 36663 4307 36669
rect 5442 36660 5448 36712
rect 5500 36700 5506 36712
rect 6917 36703 6975 36709
rect 6917 36700 6929 36703
rect 5500 36672 6929 36700
rect 5500 36660 5506 36672
rect 6917 36669 6929 36672
rect 6963 36700 6975 36703
rect 7098 36700 7104 36712
rect 6963 36672 7104 36700
rect 6963 36669 6975 36672
rect 6917 36663 6975 36669
rect 7098 36660 7104 36672
rect 7156 36660 7162 36712
rect 7650 36700 7656 36712
rect 7611 36672 7656 36700
rect 7650 36660 7656 36672
rect 7708 36660 7714 36712
rect 7929 36703 7987 36709
rect 7929 36669 7941 36703
rect 7975 36700 7987 36703
rect 8849 36703 8907 36709
rect 8849 36700 8861 36703
rect 7975 36672 8861 36700
rect 7975 36669 7987 36672
rect 7929 36663 7987 36669
rect 8849 36669 8861 36672
rect 8895 36669 8907 36703
rect 8849 36663 8907 36669
rect 9582 36660 9588 36712
rect 9640 36700 9646 36712
rect 9677 36703 9735 36709
rect 9677 36700 9689 36703
rect 9640 36672 9689 36700
rect 9640 36660 9646 36672
rect 9677 36669 9689 36672
rect 9723 36669 9735 36703
rect 9784 36700 9812 36740
rect 9861 36737 9873 36771
rect 9907 36737 9919 36771
rect 9861 36731 9919 36737
rect 10226 36728 10232 36780
rect 10284 36768 10290 36780
rect 12805 36771 12863 36777
rect 12805 36768 12817 36771
rect 10284 36740 12817 36768
rect 10284 36728 10290 36740
rect 12805 36737 12817 36740
rect 12851 36737 12863 36771
rect 12805 36731 12863 36737
rect 13173 36771 13231 36777
rect 13173 36737 13185 36771
rect 13219 36768 13231 36771
rect 13262 36768 13268 36780
rect 13219 36740 13268 36768
rect 13219 36737 13231 36740
rect 13173 36731 13231 36737
rect 13262 36728 13268 36740
rect 13320 36728 13326 36780
rect 20809 36771 20867 36777
rect 20809 36768 20821 36771
rect 19076 36740 20821 36768
rect 19076 36712 19104 36740
rect 20809 36737 20821 36740
rect 20855 36737 20867 36771
rect 20809 36731 20867 36737
rect 24121 36771 24179 36777
rect 24121 36737 24133 36771
rect 24167 36768 24179 36771
rect 24946 36768 24952 36780
rect 24167 36740 24952 36768
rect 24167 36737 24179 36740
rect 24121 36731 24179 36737
rect 24946 36728 24952 36740
rect 25004 36728 25010 36780
rect 26786 36728 26792 36780
rect 26844 36768 26850 36780
rect 27801 36771 27859 36777
rect 27801 36768 27813 36771
rect 26844 36740 27108 36768
rect 26844 36728 26850 36740
rect 10137 36703 10195 36709
rect 10137 36700 10149 36703
rect 9784 36672 10149 36700
rect 9677 36663 9735 36669
rect 10137 36669 10149 36672
rect 10183 36669 10195 36703
rect 10137 36663 10195 36669
rect 11422 36660 11428 36712
rect 11480 36700 11486 36712
rect 12342 36700 12348 36712
rect 11480 36672 12348 36700
rect 11480 36660 11486 36672
rect 12342 36660 12348 36672
rect 12400 36660 12406 36712
rect 12584 36703 12642 36709
rect 12584 36669 12596 36703
rect 12630 36700 12642 36703
rect 12894 36700 12900 36712
rect 12630 36672 12900 36700
rect 12630 36669 12642 36672
rect 12584 36663 12642 36669
rect 12894 36660 12900 36672
rect 12952 36660 12958 36712
rect 13998 36700 14004 36712
rect 13959 36672 14004 36700
rect 13998 36660 14004 36672
rect 14056 36660 14062 36712
rect 14090 36660 14096 36712
rect 14148 36700 14154 36712
rect 16669 36703 16727 36709
rect 16669 36700 16681 36703
rect 14148 36672 16681 36700
rect 14148 36660 14154 36672
rect 16669 36669 16681 36672
rect 16715 36700 16727 36703
rect 16853 36703 16911 36709
rect 16853 36700 16865 36703
rect 16715 36672 16865 36700
rect 16715 36669 16727 36672
rect 16669 36663 16727 36669
rect 16853 36669 16865 36672
rect 16899 36700 16911 36703
rect 18874 36700 18880 36712
rect 16899 36672 18880 36700
rect 16899 36669 16911 36672
rect 16853 36663 16911 36669
rect 18874 36660 18880 36672
rect 18932 36660 18938 36712
rect 19058 36700 19064 36712
rect 19019 36672 19064 36700
rect 19058 36660 19064 36672
rect 19116 36660 19122 36712
rect 19334 36660 19340 36712
rect 19392 36700 19398 36712
rect 22278 36700 22284 36712
rect 19392 36672 19437 36700
rect 19996 36672 22284 36700
rect 19392 36660 19398 36672
rect 3970 36592 3976 36644
rect 4028 36632 4034 36644
rect 12250 36632 12256 36644
rect 4028 36604 12256 36632
rect 4028 36592 4034 36604
rect 12250 36592 12256 36604
rect 12308 36592 12314 36644
rect 12437 36635 12495 36641
rect 12437 36601 12449 36635
rect 12483 36632 12495 36635
rect 12802 36632 12808 36644
rect 12483 36604 12808 36632
rect 12483 36601 12495 36604
rect 12437 36595 12495 36601
rect 12802 36592 12808 36604
rect 12860 36592 12866 36644
rect 13630 36592 13636 36644
rect 13688 36632 13694 36644
rect 18966 36632 18972 36644
rect 13688 36604 18972 36632
rect 13688 36592 13694 36604
rect 18966 36592 18972 36604
rect 19024 36592 19030 36644
rect 4525 36567 4583 36573
rect 4525 36533 4537 36567
rect 4571 36564 4583 36567
rect 4614 36564 4620 36576
rect 4571 36536 4620 36564
rect 4571 36533 4583 36536
rect 4525 36527 4583 36533
rect 4614 36524 4620 36536
rect 4672 36524 4678 36576
rect 4890 36524 4896 36576
rect 4948 36564 4954 36576
rect 7009 36567 7067 36573
rect 7009 36564 7021 36567
rect 4948 36536 7021 36564
rect 4948 36524 4954 36536
rect 7009 36533 7021 36536
rect 7055 36533 7067 36567
rect 7009 36527 7067 36533
rect 8570 36524 8576 36576
rect 8628 36564 8634 36576
rect 14182 36564 14188 36576
rect 8628 36536 14188 36564
rect 8628 36524 8634 36536
rect 14182 36524 14188 36536
rect 14240 36524 14246 36576
rect 14274 36524 14280 36576
rect 14332 36564 14338 36576
rect 14461 36567 14519 36573
rect 14461 36564 14473 36567
rect 14332 36536 14473 36564
rect 14332 36524 14338 36536
rect 14461 36533 14473 36536
rect 14507 36564 14519 36567
rect 19996 36564 20024 36672
rect 22278 36660 22284 36672
rect 22336 36660 22342 36712
rect 22373 36703 22431 36709
rect 22373 36669 22385 36703
rect 22419 36700 22431 36703
rect 22465 36703 22523 36709
rect 22465 36700 22477 36703
rect 22419 36672 22477 36700
rect 22419 36669 22431 36672
rect 22373 36663 22431 36669
rect 22465 36669 22477 36672
rect 22511 36669 22523 36703
rect 24302 36700 24308 36712
rect 24263 36672 24308 36700
rect 22465 36663 22523 36669
rect 20070 36592 20076 36644
rect 20128 36632 20134 36644
rect 22388 36632 22416 36663
rect 24302 36660 24308 36672
rect 24360 36660 24366 36712
rect 25038 36700 25044 36712
rect 24999 36672 25044 36700
rect 25038 36660 25044 36672
rect 25096 36660 25102 36712
rect 25406 36700 25412 36712
rect 25367 36672 25412 36700
rect 25406 36660 25412 36672
rect 25464 36660 25470 36712
rect 27080 36709 27108 36740
rect 27632 36740 27813 36768
rect 25501 36703 25559 36709
rect 25501 36669 25513 36703
rect 25547 36669 25559 36703
rect 25501 36663 25559 36669
rect 26881 36703 26939 36709
rect 26881 36669 26893 36703
rect 26927 36669 26939 36703
rect 26881 36663 26939 36669
rect 27065 36703 27123 36709
rect 27065 36669 27077 36703
rect 27111 36669 27123 36703
rect 27065 36663 27123 36669
rect 20128 36604 22416 36632
rect 24320 36632 24348 36660
rect 25516 36632 25544 36663
rect 26418 36632 26424 36644
rect 24320 36604 25544 36632
rect 26379 36604 26424 36632
rect 20128 36592 20134 36604
rect 26418 36592 26424 36604
rect 26476 36592 26482 36644
rect 26896 36632 26924 36663
rect 27154 36660 27160 36712
rect 27212 36700 27218 36712
rect 27632 36709 27660 36740
rect 27801 36737 27813 36740
rect 27847 36768 27859 36771
rect 28626 36768 28632 36780
rect 27847 36740 28632 36768
rect 27847 36737 27859 36740
rect 27801 36731 27859 36737
rect 28626 36728 28632 36740
rect 28684 36728 28690 36780
rect 30285 36771 30343 36777
rect 30285 36737 30297 36771
rect 30331 36768 30343 36771
rect 31404 36768 31432 36808
rect 32030 36796 32036 36808
rect 32088 36796 32094 36848
rect 30331 36740 31432 36768
rect 31941 36771 31999 36777
rect 30331 36737 30343 36740
rect 30285 36731 30343 36737
rect 31941 36737 31953 36771
rect 31987 36768 31999 36771
rect 32122 36768 32128 36780
rect 31987 36740 32128 36768
rect 31987 36737 31999 36740
rect 31941 36731 31999 36737
rect 32122 36728 32128 36740
rect 32180 36768 32186 36780
rect 34701 36771 34759 36777
rect 34701 36768 34713 36771
rect 32180 36740 34713 36768
rect 32180 36728 32186 36740
rect 34701 36737 34713 36740
rect 34747 36737 34759 36771
rect 35636 36768 35664 36867
rect 36998 36864 37004 36876
rect 37056 36864 37062 36916
rect 39117 36907 39175 36913
rect 39117 36873 39129 36907
rect 39163 36904 39175 36907
rect 39393 36907 39451 36913
rect 39393 36904 39405 36907
rect 39163 36876 39405 36904
rect 39163 36873 39175 36876
rect 39117 36867 39175 36873
rect 39393 36873 39405 36876
rect 39439 36904 39451 36907
rect 39482 36904 39488 36916
rect 39439 36876 39488 36904
rect 39439 36873 39451 36876
rect 39393 36867 39451 36873
rect 39482 36864 39488 36876
rect 39540 36864 39546 36916
rect 49786 36864 49792 36916
rect 49844 36904 49850 36916
rect 53745 36907 53803 36913
rect 49844 36876 53696 36904
rect 49844 36864 49850 36876
rect 35710 36796 35716 36848
rect 35768 36836 35774 36848
rect 43162 36836 43168 36848
rect 35768 36808 43168 36836
rect 35768 36796 35774 36808
rect 43162 36796 43168 36808
rect 43220 36796 43226 36848
rect 44174 36836 44180 36848
rect 44135 36808 44180 36836
rect 44174 36796 44180 36808
rect 44232 36796 44238 36848
rect 48038 36796 48044 36848
rect 48096 36836 48102 36848
rect 50430 36836 50436 36848
rect 48096 36808 50436 36836
rect 48096 36796 48102 36808
rect 50430 36796 50436 36808
rect 50488 36796 50494 36848
rect 50706 36836 50712 36848
rect 50667 36808 50712 36836
rect 50706 36796 50712 36808
rect 50764 36796 50770 36848
rect 53668 36836 53696 36876
rect 53745 36873 53757 36907
rect 53791 36904 53803 36907
rect 54938 36904 54944 36916
rect 53791 36876 54944 36904
rect 53791 36873 53803 36876
rect 53745 36867 53803 36873
rect 54938 36864 54944 36876
rect 54996 36864 55002 36916
rect 60734 36904 60740 36916
rect 55876 36876 60740 36904
rect 54849 36839 54907 36845
rect 54849 36836 54861 36839
rect 53668 36808 54861 36836
rect 54849 36805 54861 36808
rect 54895 36836 54907 36839
rect 55876 36836 55904 36876
rect 60734 36864 60740 36876
rect 60792 36864 60798 36916
rect 91002 36904 91008 36916
rect 60844 36876 91008 36904
rect 54895 36808 55904 36836
rect 54895 36805 54907 36808
rect 54849 36799 54907 36805
rect 35805 36771 35863 36777
rect 35805 36768 35817 36771
rect 35636 36740 35817 36768
rect 34701 36731 34759 36737
rect 35805 36737 35817 36740
rect 35851 36737 35863 36771
rect 35805 36731 35863 36737
rect 38102 36728 38108 36780
rect 38160 36768 38166 36780
rect 48498 36768 48504 36780
rect 38160 36740 48504 36768
rect 38160 36728 38166 36740
rect 48498 36728 48504 36740
rect 48556 36728 48562 36780
rect 48682 36768 48688 36780
rect 48643 36740 48688 36768
rect 48682 36728 48688 36740
rect 48740 36728 48746 36780
rect 50249 36771 50307 36777
rect 50249 36737 50261 36771
rect 50295 36768 50307 36771
rect 50580 36771 50638 36777
rect 50580 36768 50592 36771
rect 50295 36740 50592 36768
rect 50295 36737 50307 36740
rect 50249 36731 50307 36737
rect 50580 36737 50592 36740
rect 50626 36737 50638 36771
rect 50798 36768 50804 36780
rect 50759 36740 50804 36768
rect 50580 36731 50638 36737
rect 50798 36728 50804 36740
rect 50856 36728 50862 36780
rect 51166 36768 51172 36780
rect 51127 36740 51172 36768
rect 51166 36728 51172 36740
rect 51224 36728 51230 36780
rect 52454 36728 52460 36780
rect 52512 36768 52518 36780
rect 54297 36771 54355 36777
rect 52512 36740 52960 36768
rect 52512 36728 52518 36740
rect 27433 36703 27491 36709
rect 27433 36700 27445 36703
rect 27212 36672 27445 36700
rect 27212 36660 27218 36672
rect 27433 36669 27445 36672
rect 27479 36669 27491 36703
rect 27433 36663 27491 36669
rect 27617 36703 27675 36709
rect 27617 36669 27629 36703
rect 27663 36669 27675 36703
rect 27617 36663 27675 36669
rect 27985 36703 28043 36709
rect 27985 36669 27997 36703
rect 28031 36700 28043 36703
rect 28718 36700 28724 36712
rect 28031 36672 28724 36700
rect 28031 36669 28043 36672
rect 27985 36663 28043 36669
rect 28000 36632 28028 36663
rect 28718 36660 28724 36672
rect 28776 36660 28782 36712
rect 30374 36660 30380 36712
rect 30432 36700 30438 36712
rect 30561 36703 30619 36709
rect 30561 36700 30573 36703
rect 30432 36672 30573 36700
rect 30432 36660 30438 36672
rect 30561 36669 30573 36672
rect 30607 36669 30619 36703
rect 30561 36663 30619 36669
rect 31846 36660 31852 36712
rect 31904 36700 31910 36712
rect 32953 36703 33011 36709
rect 32953 36700 32965 36703
rect 31904 36672 32965 36700
rect 31904 36660 31910 36672
rect 32953 36669 32965 36672
rect 32999 36669 33011 36703
rect 32953 36663 33011 36669
rect 35529 36703 35587 36709
rect 35529 36669 35541 36703
rect 35575 36700 35587 36703
rect 35986 36700 35992 36712
rect 35575 36672 35992 36700
rect 35575 36669 35587 36672
rect 35529 36663 35587 36669
rect 35986 36660 35992 36672
rect 36044 36660 36050 36712
rect 36446 36660 36452 36712
rect 36504 36700 36510 36712
rect 36541 36703 36599 36709
rect 36541 36700 36553 36703
rect 36504 36672 36553 36700
rect 36504 36660 36510 36672
rect 36541 36669 36553 36672
rect 36587 36669 36599 36703
rect 36541 36663 36599 36669
rect 36722 36660 36728 36712
rect 36780 36700 36786 36712
rect 39117 36703 39175 36709
rect 39117 36700 39129 36703
rect 36780 36672 39129 36700
rect 36780 36660 36786 36672
rect 39117 36669 39129 36672
rect 39163 36669 39175 36703
rect 39298 36700 39304 36712
rect 39259 36672 39304 36700
rect 39117 36663 39175 36669
rect 39298 36660 39304 36672
rect 39356 36660 39362 36712
rect 44085 36703 44143 36709
rect 44085 36669 44097 36703
rect 44131 36700 44143 36703
rect 44450 36700 44456 36712
rect 44131 36672 44456 36700
rect 44131 36669 44143 36672
rect 44085 36663 44143 36669
rect 44450 36660 44456 36672
rect 44508 36660 44514 36712
rect 46937 36703 46995 36709
rect 46937 36669 46949 36703
rect 46983 36700 46995 36703
rect 47029 36703 47087 36709
rect 47029 36700 47041 36703
rect 46983 36672 47041 36700
rect 46983 36669 46995 36672
rect 46937 36663 46995 36669
rect 47029 36669 47041 36672
rect 47075 36669 47087 36703
rect 47302 36700 47308 36712
rect 47263 36672 47308 36700
rect 47029 36663 47087 36669
rect 38562 36632 38568 36644
rect 26896 36604 28028 36632
rect 32600 36604 38568 36632
rect 20622 36564 20628 36576
rect 14507 36536 20024 36564
rect 20583 36536 20628 36564
rect 14507 36533 14519 36536
rect 14461 36527 14519 36533
rect 20622 36524 20628 36536
rect 20680 36524 20686 36576
rect 24486 36564 24492 36576
rect 24447 36536 24492 36564
rect 24486 36524 24492 36536
rect 24544 36524 24550 36576
rect 25130 36524 25136 36576
rect 25188 36564 25194 36576
rect 32600 36564 32628 36604
rect 38562 36592 38568 36604
rect 38620 36592 38626 36644
rect 43346 36592 43352 36644
rect 43404 36632 43410 36644
rect 46952 36632 46980 36663
rect 47302 36660 47308 36672
rect 47360 36660 47366 36712
rect 48961 36703 49019 36709
rect 48961 36700 48973 36703
rect 48424 36672 48973 36700
rect 43404 36604 46980 36632
rect 43404 36592 43410 36604
rect 32766 36564 32772 36576
rect 25188 36536 32628 36564
rect 32727 36536 32772 36564
rect 25188 36524 25194 36536
rect 32766 36524 32772 36536
rect 32824 36524 32830 36576
rect 34701 36567 34759 36573
rect 34701 36533 34713 36567
rect 34747 36564 34759 36567
rect 37826 36564 37832 36576
rect 34747 36536 37832 36564
rect 34747 36533 34759 36536
rect 34701 36527 34759 36533
rect 37826 36524 37832 36536
rect 37884 36524 37890 36576
rect 38654 36524 38660 36576
rect 38712 36564 38718 36576
rect 43254 36564 43260 36576
rect 38712 36536 43260 36564
rect 38712 36524 38718 36536
rect 43254 36524 43260 36536
rect 43312 36524 43318 36576
rect 48314 36524 48320 36576
rect 48372 36564 48378 36576
rect 48424 36564 48452 36672
rect 48961 36669 48973 36672
rect 49007 36669 49019 36703
rect 48961 36663 49019 36669
rect 49145 36703 49203 36709
rect 49145 36669 49157 36703
rect 49191 36669 49203 36703
rect 49145 36663 49203 36669
rect 49160 36576 49188 36663
rect 49234 36660 49240 36712
rect 49292 36700 49298 36712
rect 49605 36703 49663 36709
rect 49605 36700 49617 36703
rect 49292 36672 49617 36700
rect 49292 36660 49298 36672
rect 49605 36669 49617 36672
rect 49651 36669 49663 36703
rect 49605 36663 49663 36669
rect 49697 36703 49755 36709
rect 49697 36669 49709 36703
rect 49743 36669 49755 36703
rect 49697 36663 49755 36669
rect 50433 36703 50491 36709
rect 50433 36669 50445 36703
rect 50479 36700 50491 36703
rect 51442 36700 51448 36712
rect 50479 36672 51448 36700
rect 50479 36669 50491 36672
rect 50433 36663 50491 36669
rect 49712 36632 49740 36663
rect 51442 36660 51448 36672
rect 51500 36660 51506 36712
rect 52730 36700 52736 36712
rect 52691 36672 52736 36700
rect 52730 36660 52736 36672
rect 52788 36660 52794 36712
rect 52825 36703 52883 36709
rect 52825 36669 52837 36703
rect 52871 36669 52883 36703
rect 52932 36700 52960 36740
rect 54297 36737 54309 36771
rect 54343 36768 54355 36771
rect 55030 36768 55036 36780
rect 54343 36740 55036 36768
rect 54343 36737 54355 36740
rect 54297 36731 54355 36737
rect 53193 36703 53251 36709
rect 53193 36700 53205 36703
rect 52932 36672 53205 36700
rect 52825 36663 52883 36669
rect 53193 36669 53205 36672
rect 53239 36669 53251 36703
rect 53193 36663 53251 36669
rect 53285 36703 53343 36709
rect 53285 36669 53297 36703
rect 53331 36700 53343 36703
rect 53834 36700 53840 36712
rect 53331 36672 53840 36700
rect 53331 36669 53343 36672
rect 53285 36663 53343 36669
rect 50890 36632 50896 36644
rect 49712 36604 50896 36632
rect 50890 36592 50896 36604
rect 50948 36632 50954 36644
rect 51261 36635 51319 36641
rect 51261 36632 51273 36635
rect 50948 36604 51273 36632
rect 50948 36592 50954 36604
rect 51261 36601 51273 36604
rect 51307 36601 51319 36635
rect 52454 36632 52460 36644
rect 52367 36604 52460 36632
rect 51261 36595 51319 36601
rect 52454 36592 52460 36604
rect 52512 36632 52518 36644
rect 52840 36632 52868 36663
rect 53834 36660 53840 36672
rect 53892 36700 53898 36712
rect 54312 36700 54340 36731
rect 55030 36728 55036 36740
rect 55088 36728 55094 36780
rect 55306 36768 55312 36780
rect 55267 36740 55312 36768
rect 55306 36728 55312 36740
rect 55364 36728 55370 36780
rect 55876 36709 55904 36808
rect 56042 36796 56048 36848
rect 56100 36836 56106 36848
rect 56594 36836 56600 36848
rect 56100 36808 56600 36836
rect 56100 36796 56106 36808
rect 56594 36796 56600 36808
rect 56652 36836 56658 36848
rect 57149 36839 57207 36845
rect 57149 36836 57161 36839
rect 56652 36808 57161 36836
rect 56652 36796 56658 36808
rect 57149 36805 57161 36808
rect 57195 36805 57207 36839
rect 57149 36799 57207 36805
rect 58250 36796 58256 36848
rect 58308 36836 58314 36848
rect 58437 36839 58495 36845
rect 58437 36836 58449 36839
rect 58308 36808 58449 36836
rect 58308 36796 58314 36808
rect 58437 36805 58449 36808
rect 58483 36805 58495 36839
rect 58437 36799 58495 36805
rect 58526 36796 58532 36848
rect 58584 36836 58590 36848
rect 60844 36836 60872 36876
rect 91002 36864 91008 36876
rect 91060 36864 91066 36916
rect 91097 36907 91155 36913
rect 91097 36873 91109 36907
rect 91143 36904 91155 36907
rect 91278 36904 91284 36916
rect 91143 36876 91284 36904
rect 91143 36873 91155 36876
rect 91097 36867 91155 36873
rect 91278 36864 91284 36876
rect 91336 36864 91342 36916
rect 91373 36907 91431 36913
rect 91373 36873 91385 36907
rect 91419 36904 91431 36907
rect 93394 36904 93400 36916
rect 91419 36876 93400 36904
rect 91419 36873 91431 36876
rect 91373 36867 91431 36873
rect 64414 36836 64420 36848
rect 58584 36808 60872 36836
rect 64375 36808 64420 36836
rect 58584 36796 58590 36808
rect 64414 36796 64420 36808
rect 64472 36836 64478 36848
rect 71685 36839 71743 36845
rect 71685 36836 71697 36839
rect 64472 36808 64552 36836
rect 64472 36796 64478 36808
rect 55953 36771 56011 36777
rect 55953 36737 55965 36771
rect 55999 36768 56011 36771
rect 56686 36768 56692 36780
rect 55999 36740 56692 36768
rect 55999 36737 56011 36740
rect 55953 36731 56011 36737
rect 56686 36728 56692 36740
rect 56744 36768 56750 36780
rect 64524 36777 64552 36808
rect 71240 36808 71697 36836
rect 64509 36771 64567 36777
rect 56744 36740 57652 36768
rect 56744 36728 56750 36740
rect 53892 36672 54340 36700
rect 55861 36703 55919 36709
rect 53892 36660 53898 36672
rect 55861 36669 55873 36703
rect 55907 36669 55919 36703
rect 55861 36663 55919 36669
rect 56229 36703 56287 36709
rect 56229 36669 56241 36703
rect 56275 36669 56287 36703
rect 56229 36663 56287 36669
rect 53742 36632 53748 36644
rect 52512 36604 53748 36632
rect 52512 36592 52518 36604
rect 53742 36592 53748 36604
rect 53800 36592 53806 36644
rect 53944 36604 54892 36632
rect 48777 36567 48835 36573
rect 48777 36564 48789 36567
rect 48372 36536 48789 36564
rect 48372 36524 48378 36536
rect 48777 36533 48789 36536
rect 48823 36533 48835 36567
rect 49142 36564 49148 36576
rect 49055 36536 49148 36564
rect 48777 36527 48835 36533
rect 49142 36524 49148 36536
rect 49200 36564 49206 36576
rect 51537 36567 51595 36573
rect 51537 36564 51549 36567
rect 49200 36536 51549 36564
rect 49200 36524 49206 36536
rect 51537 36533 51549 36536
rect 51583 36564 51595 36567
rect 51718 36564 51724 36576
rect 51583 36536 51724 36564
rect 51583 36533 51595 36536
rect 51537 36527 51595 36533
rect 51718 36524 51724 36536
rect 51776 36524 51782 36576
rect 51902 36524 51908 36576
rect 51960 36564 51966 36576
rect 53944 36564 53972 36604
rect 54110 36564 54116 36576
rect 51960 36536 53972 36564
rect 54071 36536 54116 36564
rect 51960 36524 51966 36536
rect 54110 36524 54116 36536
rect 54168 36524 54174 36576
rect 54864 36564 54892 36604
rect 55033 36567 55091 36573
rect 55033 36564 55045 36567
rect 54864 36536 55045 36564
rect 55033 36533 55045 36536
rect 55079 36564 55091 36567
rect 56244 36564 56272 36663
rect 56318 36660 56324 36712
rect 56376 36700 56382 36712
rect 56778 36700 56784 36712
rect 56376 36672 56421 36700
rect 56739 36672 56784 36700
rect 56376 36660 56382 36672
rect 56778 36660 56784 36672
rect 56836 36700 56842 36712
rect 56965 36703 57023 36709
rect 56965 36700 56977 36703
rect 56836 36672 56977 36700
rect 56836 36660 56842 36672
rect 56965 36669 56977 36672
rect 57011 36669 57023 36703
rect 56965 36663 57023 36669
rect 57149 36703 57207 36709
rect 57149 36669 57161 36703
rect 57195 36700 57207 36703
rect 57333 36703 57391 36709
rect 57333 36700 57345 36703
rect 57195 36672 57345 36700
rect 57195 36669 57207 36672
rect 57149 36663 57207 36669
rect 57333 36669 57345 36672
rect 57379 36669 57391 36703
rect 57333 36663 57391 36669
rect 57517 36703 57575 36709
rect 57517 36669 57529 36703
rect 57563 36669 57575 36703
rect 57624 36700 57652 36740
rect 64509 36737 64521 36771
rect 64555 36737 64567 36771
rect 64782 36768 64788 36780
rect 64743 36740 64788 36768
rect 64509 36731 64567 36737
rect 64782 36728 64788 36740
rect 64840 36728 64846 36780
rect 69014 36728 69020 36780
rect 69072 36768 69078 36780
rect 70305 36771 70363 36777
rect 70305 36768 70317 36771
rect 69072 36740 70317 36768
rect 69072 36728 69078 36740
rect 70305 36737 70317 36740
rect 70351 36737 70363 36771
rect 71038 36768 71044 36780
rect 70999 36740 71044 36768
rect 70305 36731 70363 36737
rect 71038 36728 71044 36740
rect 71096 36728 71102 36780
rect 57977 36703 58035 36709
rect 57977 36700 57989 36703
rect 57624 36672 57989 36700
rect 57517 36663 57575 36669
rect 57977 36669 57989 36672
rect 58023 36669 58035 36703
rect 57977 36663 58035 36669
rect 58069 36703 58127 36709
rect 58069 36669 58081 36703
rect 58115 36669 58127 36703
rect 69290 36700 69296 36712
rect 58069 36663 58127 36669
rect 64616 36672 66484 36700
rect 69251 36672 69296 36700
rect 57532 36632 57560 36663
rect 57882 36632 57888 36644
rect 57532 36604 57888 36632
rect 57882 36592 57888 36604
rect 57940 36632 57946 36644
rect 58084 36632 58112 36663
rect 62114 36632 62120 36644
rect 57940 36604 62120 36632
rect 57940 36592 57946 36604
rect 62114 36592 62120 36604
rect 62172 36592 62178 36644
rect 63126 36592 63132 36644
rect 63184 36632 63190 36644
rect 64616 36632 64644 36672
rect 63184 36604 64644 36632
rect 66456 36632 66484 36672
rect 69290 36660 69296 36672
rect 69348 36660 69354 36712
rect 70949 36703 71007 36709
rect 70949 36669 70961 36703
rect 70995 36700 71007 36703
rect 71240 36700 71268 36808
rect 71685 36805 71697 36808
rect 71731 36836 71743 36839
rect 71774 36836 71780 36848
rect 71731 36808 71780 36836
rect 71731 36805 71743 36808
rect 71685 36799 71743 36805
rect 71774 36796 71780 36808
rect 71832 36796 71838 36848
rect 71869 36839 71927 36845
rect 71869 36805 71881 36839
rect 71915 36836 71927 36839
rect 72970 36836 72976 36848
rect 71915 36808 72976 36836
rect 71915 36805 71927 36808
rect 71869 36799 71927 36805
rect 71884 36768 71912 36799
rect 72970 36796 72976 36808
rect 73028 36836 73034 36848
rect 85117 36839 85175 36845
rect 73028 36808 84976 36836
rect 73028 36796 73034 36808
rect 77294 36768 77300 36780
rect 71332 36740 71912 36768
rect 77255 36740 77300 36768
rect 71332 36709 71360 36740
rect 77294 36728 77300 36740
rect 77352 36728 77358 36780
rect 77478 36728 77484 36780
rect 77536 36768 77542 36780
rect 77757 36771 77815 36777
rect 77757 36768 77769 36771
rect 77536 36740 77769 36768
rect 77536 36728 77542 36740
rect 77757 36737 77769 36740
rect 77803 36768 77815 36771
rect 78677 36771 78735 36777
rect 78677 36768 78689 36771
rect 77803 36740 78689 36768
rect 77803 36737 77815 36740
rect 77757 36731 77815 36737
rect 78677 36737 78689 36740
rect 78723 36737 78735 36771
rect 78677 36731 78735 36737
rect 79226 36728 79232 36780
rect 79284 36768 79290 36780
rect 79284 36740 81572 36768
rect 79284 36728 79290 36740
rect 70995 36672 71268 36700
rect 71317 36703 71375 36709
rect 70995 36669 71007 36672
rect 70949 36663 71007 36669
rect 71317 36669 71329 36703
rect 71363 36669 71375 36703
rect 71317 36663 71375 36669
rect 71406 36660 71412 36712
rect 71464 36700 71470 36712
rect 76745 36703 76803 36709
rect 71464 36672 71509 36700
rect 71464 36660 71470 36672
rect 76745 36669 76757 36703
rect 76791 36700 76803 36703
rect 77386 36700 77392 36712
rect 76791 36672 77392 36700
rect 76791 36669 76803 36672
rect 76745 36663 76803 36669
rect 77386 36660 77392 36672
rect 77444 36660 77450 36712
rect 77573 36703 77631 36709
rect 77573 36669 77585 36703
rect 77619 36700 77631 36703
rect 77662 36700 77668 36712
rect 77619 36672 77668 36700
rect 77619 36669 77631 36672
rect 77573 36663 77631 36669
rect 77662 36660 77668 36672
rect 77720 36660 77726 36712
rect 78398 36700 78404 36712
rect 78311 36672 78404 36700
rect 78398 36660 78404 36672
rect 78456 36700 78462 36712
rect 78585 36703 78643 36709
rect 78585 36700 78597 36703
rect 78456 36672 78597 36700
rect 78456 36660 78462 36672
rect 78585 36669 78597 36672
rect 78631 36669 78643 36703
rect 78585 36663 78643 36669
rect 78766 36660 78772 36712
rect 78824 36700 78830 36712
rect 81544 36709 81572 36740
rect 79965 36703 80023 36709
rect 79965 36700 79977 36703
rect 78824 36672 79977 36700
rect 78824 36660 78830 36672
rect 79965 36669 79977 36672
rect 80011 36700 80023 36703
rect 80425 36703 80483 36709
rect 80425 36700 80437 36703
rect 80011 36672 80437 36700
rect 80011 36669 80023 36672
rect 79965 36663 80023 36669
rect 80425 36669 80437 36672
rect 80471 36669 80483 36703
rect 80425 36663 80483 36669
rect 81529 36703 81587 36709
rect 81529 36669 81541 36703
rect 81575 36669 81587 36703
rect 81529 36663 81587 36669
rect 69385 36635 69443 36641
rect 69385 36632 69397 36635
rect 66456 36604 69397 36632
rect 63184 36592 63190 36604
rect 69385 36601 69397 36604
rect 69431 36632 69443 36635
rect 69750 36632 69756 36644
rect 69431 36604 69756 36632
rect 69431 36601 69443 36604
rect 69385 36595 69443 36601
rect 69750 36592 69756 36604
rect 69808 36592 69814 36644
rect 58618 36564 58624 36576
rect 55079 36536 58624 36564
rect 55079 36533 55091 36536
rect 55033 36527 55091 36533
rect 58618 36524 58624 36536
rect 58676 36524 58682 36576
rect 66070 36564 66076 36576
rect 66031 36536 66076 36564
rect 66070 36524 66076 36536
rect 66128 36524 66134 36576
rect 77294 36524 77300 36576
rect 77352 36564 77358 36576
rect 78416 36573 78444 36660
rect 79778 36632 79784 36644
rect 79739 36604 79784 36632
rect 79778 36592 79784 36604
rect 79836 36592 79842 36644
rect 78401 36567 78459 36573
rect 78401 36564 78413 36567
rect 77352 36536 78413 36564
rect 77352 36524 77358 36536
rect 78401 36533 78413 36536
rect 78447 36533 78459 36567
rect 78401 36527 78459 36533
rect 80054 36524 80060 36576
rect 80112 36564 80118 36576
rect 81710 36564 81716 36576
rect 80112 36536 80157 36564
rect 81671 36536 81716 36564
rect 80112 36524 80118 36536
rect 81710 36524 81716 36536
rect 81768 36524 81774 36576
rect 84286 36524 84292 36576
rect 84344 36564 84350 36576
rect 84841 36567 84899 36573
rect 84841 36564 84853 36567
rect 84344 36536 84853 36564
rect 84344 36524 84350 36536
rect 84841 36533 84853 36536
rect 84887 36533 84899 36567
rect 84948 36564 84976 36808
rect 85117 36805 85129 36839
rect 85163 36836 85175 36839
rect 85206 36836 85212 36848
rect 85163 36808 85212 36836
rect 85163 36805 85175 36808
rect 85117 36799 85175 36805
rect 85206 36796 85212 36808
rect 85264 36796 85270 36848
rect 85574 36836 85580 36848
rect 85535 36808 85580 36836
rect 85574 36796 85580 36808
rect 85632 36796 85638 36848
rect 85224 36700 85252 36796
rect 86218 36768 86224 36780
rect 86179 36740 86224 36768
rect 86218 36728 86224 36740
rect 86276 36768 86282 36780
rect 88426 36768 88432 36780
rect 86276 36740 88432 36768
rect 86276 36728 86282 36740
rect 88426 36728 88432 36740
rect 88484 36728 88490 36780
rect 90085 36771 90143 36777
rect 90085 36737 90097 36771
rect 90131 36768 90143 36771
rect 91278 36768 91284 36780
rect 90131 36740 91284 36768
rect 90131 36737 90143 36740
rect 90085 36731 90143 36737
rect 91278 36728 91284 36740
rect 91336 36728 91342 36780
rect 85393 36703 85451 36709
rect 85393 36700 85405 36703
rect 85224 36672 85405 36700
rect 85393 36669 85405 36672
rect 85439 36669 85451 36703
rect 85393 36663 85451 36669
rect 85482 36660 85488 36712
rect 85540 36700 85546 36712
rect 85945 36703 86003 36709
rect 85945 36700 85957 36703
rect 85540 36672 85957 36700
rect 85540 36660 85546 36672
rect 85945 36669 85957 36672
rect 85991 36669 86003 36703
rect 85945 36663 86003 36669
rect 89717 36703 89775 36709
rect 89717 36669 89729 36703
rect 89763 36669 89775 36703
rect 91005 36703 91063 36709
rect 91005 36700 91017 36703
rect 89717 36663 89775 36669
rect 90284 36672 91017 36700
rect 89162 36592 89168 36644
rect 89220 36632 89226 36644
rect 89533 36635 89591 36641
rect 89533 36632 89545 36635
rect 89220 36604 89545 36632
rect 89220 36592 89226 36604
rect 89533 36601 89545 36604
rect 89579 36601 89591 36635
rect 89732 36632 89760 36663
rect 90174 36632 90180 36644
rect 89732 36604 90180 36632
rect 89533 36595 89591 36601
rect 90174 36592 90180 36604
rect 90232 36592 90238 36644
rect 90284 36564 90312 36672
rect 91005 36669 91017 36672
rect 91051 36700 91063 36703
rect 91480 36700 91508 36876
rect 93394 36864 93400 36876
rect 93452 36864 93458 36916
rect 93857 36907 93915 36913
rect 93857 36873 93869 36907
rect 93903 36904 93915 36907
rect 94038 36904 94044 36916
rect 93903 36876 94044 36904
rect 93903 36873 93915 36876
rect 93857 36867 93915 36873
rect 94038 36864 94044 36876
rect 94096 36864 94102 36916
rect 95326 36864 95332 36916
rect 95384 36904 95390 36916
rect 96893 36907 96951 36913
rect 96893 36904 96905 36907
rect 95384 36876 96905 36904
rect 95384 36864 95390 36876
rect 96893 36873 96905 36876
rect 96939 36873 96951 36907
rect 96893 36867 96951 36873
rect 95234 36768 95240 36780
rect 92952 36740 95240 36768
rect 92952 36709 92980 36740
rect 95234 36728 95240 36740
rect 95292 36728 95298 36780
rect 91051 36672 91508 36700
rect 92937 36703 92995 36709
rect 91051 36669 91063 36672
rect 91005 36663 91063 36669
rect 92937 36669 92949 36703
rect 92983 36669 92995 36703
rect 92937 36663 92995 36669
rect 93029 36703 93087 36709
rect 93029 36669 93041 36703
rect 93075 36700 93087 36703
rect 94593 36703 94651 36709
rect 94593 36700 94605 36703
rect 93075 36672 94605 36700
rect 93075 36669 93087 36672
rect 93029 36663 93087 36669
rect 94593 36669 94605 36672
rect 94639 36669 94651 36703
rect 94593 36663 94651 36669
rect 92750 36592 92756 36644
rect 92808 36632 92814 36644
rect 93949 36635 94007 36641
rect 93949 36632 93961 36635
rect 92808 36604 93961 36632
rect 92808 36592 92814 36604
rect 93949 36601 93961 36604
rect 93995 36601 94007 36635
rect 94608 36632 94636 36663
rect 94682 36660 94688 36712
rect 94740 36700 94746 36712
rect 94958 36700 94964 36712
rect 94740 36672 94785 36700
rect 94919 36672 94964 36700
rect 94740 36660 94746 36672
rect 94958 36660 94964 36672
rect 95016 36660 95022 36712
rect 95050 36660 95056 36712
rect 95108 36700 95114 36712
rect 95108 36672 95153 36700
rect 95108 36660 95114 36672
rect 95326 36660 95332 36712
rect 95384 36700 95390 36712
rect 96801 36703 96859 36709
rect 96801 36700 96813 36703
rect 95384 36672 96813 36700
rect 95384 36660 95390 36672
rect 96801 36669 96813 36672
rect 96847 36700 96859 36703
rect 97258 36700 97264 36712
rect 96847 36672 97264 36700
rect 96847 36669 96859 36672
rect 96801 36663 96859 36669
rect 97258 36660 97264 36672
rect 97316 36660 97322 36712
rect 96617 36635 96675 36641
rect 96617 36632 96629 36635
rect 94608 36604 96629 36632
rect 93949 36595 94007 36601
rect 96617 36601 96629 36604
rect 96663 36601 96675 36635
rect 96617 36595 96675 36601
rect 84948 36536 90312 36564
rect 84841 36527 84899 36533
rect 90910 36524 90916 36576
rect 90968 36564 90974 36576
rect 93581 36567 93639 36573
rect 93581 36564 93593 36567
rect 90968 36536 93593 36564
rect 90968 36524 90974 36536
rect 93581 36533 93593 36536
rect 93627 36564 93639 36567
rect 94682 36564 94688 36576
rect 93627 36536 94688 36564
rect 93627 36533 93639 36536
rect 93581 36527 93639 36533
rect 94682 36524 94688 36536
rect 94740 36524 94746 36576
rect 1104 36474 105616 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 50326 36474
rect 50378 36422 50390 36474
rect 50442 36422 50454 36474
rect 50506 36422 50518 36474
rect 50570 36422 81046 36474
rect 81098 36422 81110 36474
rect 81162 36422 81174 36474
rect 81226 36422 81238 36474
rect 81290 36422 105616 36474
rect 1104 36400 105616 36422
rect 8938 36360 8944 36372
rect 8899 36332 8944 36360
rect 8938 36320 8944 36332
rect 8996 36320 9002 36372
rect 11790 36360 11796 36372
rect 11751 36332 11796 36360
rect 11790 36320 11796 36332
rect 11848 36320 11854 36372
rect 24486 36360 24492 36372
rect 11900 36332 24492 36360
rect 5074 36252 5080 36304
rect 5132 36292 5138 36304
rect 11900 36292 11928 36332
rect 24486 36320 24492 36332
rect 24544 36320 24550 36372
rect 24762 36320 24768 36372
rect 24820 36360 24826 36372
rect 26234 36360 26240 36372
rect 24820 36332 26240 36360
rect 24820 36320 24826 36332
rect 26234 36320 26240 36332
rect 26292 36360 26298 36372
rect 26789 36363 26847 36369
rect 26789 36360 26801 36363
rect 26292 36332 26801 36360
rect 26292 36320 26298 36332
rect 26789 36329 26801 36332
rect 26835 36360 26847 36363
rect 26970 36360 26976 36372
rect 26835 36332 26976 36360
rect 26835 36329 26847 36332
rect 26789 36323 26847 36329
rect 26970 36320 26976 36332
rect 27028 36320 27034 36372
rect 27157 36363 27215 36369
rect 27157 36329 27169 36363
rect 27203 36360 27215 36363
rect 27203 36332 29040 36360
rect 27203 36329 27215 36332
rect 27157 36323 27215 36329
rect 5132 36264 11928 36292
rect 12437 36295 12495 36301
rect 5132 36252 5138 36264
rect 12437 36261 12449 36295
rect 12483 36292 12495 36295
rect 12894 36292 12900 36304
rect 12483 36264 12900 36292
rect 12483 36261 12495 36264
rect 12437 36255 12495 36261
rect 12894 36252 12900 36264
rect 12952 36252 12958 36304
rect 24305 36295 24363 36301
rect 24305 36292 24317 36295
rect 13740 36264 24317 36292
rect 8570 36224 8576 36236
rect 8531 36196 8576 36224
rect 8570 36184 8576 36196
rect 8628 36184 8634 36236
rect 8757 36227 8815 36233
rect 8757 36193 8769 36227
rect 8803 36224 8815 36227
rect 8938 36224 8944 36236
rect 8803 36196 8944 36224
rect 8803 36193 8815 36196
rect 8757 36187 8815 36193
rect 8938 36184 8944 36196
rect 8996 36184 9002 36236
rect 11333 36227 11391 36233
rect 11333 36193 11345 36227
rect 11379 36224 11391 36227
rect 11790 36224 11796 36236
rect 11379 36196 11796 36224
rect 11379 36193 11391 36196
rect 11333 36187 11391 36193
rect 11790 36184 11796 36196
rect 11848 36184 11854 36236
rect 12776 36227 12834 36233
rect 12776 36193 12788 36227
rect 12822 36224 12834 36227
rect 12986 36224 12992 36236
rect 12822 36196 12992 36224
rect 12822 36193 12834 36196
rect 12776 36187 12834 36193
rect 12986 36184 12992 36196
rect 13044 36184 13050 36236
rect 7742 36156 7748 36168
rect 7703 36128 7748 36156
rect 7742 36116 7748 36128
rect 7800 36116 7806 36168
rect 8297 36159 8355 36165
rect 8297 36125 8309 36159
rect 8343 36156 8355 36159
rect 8662 36156 8668 36168
rect 8343 36128 8668 36156
rect 8343 36125 8355 36128
rect 8297 36119 8355 36125
rect 8662 36116 8668 36128
rect 8720 36116 8726 36168
rect 13170 36156 13176 36168
rect 13131 36128 13176 36156
rect 13170 36116 13176 36128
rect 13228 36116 13234 36168
rect 5994 36048 6000 36100
rect 6052 36088 6058 36100
rect 11517 36091 11575 36097
rect 6052 36060 9168 36088
rect 6052 36048 6058 36060
rect 8754 35980 8760 36032
rect 8812 36020 8818 36032
rect 9033 36023 9091 36029
rect 9033 36020 9045 36023
rect 8812 35992 9045 36020
rect 8812 35980 8818 35992
rect 9033 35989 9045 35992
rect 9079 35989 9091 36023
rect 9140 36020 9168 36060
rect 11517 36057 11529 36091
rect 11563 36088 11575 36091
rect 12342 36088 12348 36100
rect 11563 36060 12348 36088
rect 11563 36057 11575 36060
rect 11517 36051 11575 36057
rect 12342 36048 12348 36060
rect 12400 36048 12406 36100
rect 12526 36048 12532 36100
rect 12584 36097 12590 36100
rect 12584 36091 12633 36097
rect 12584 36057 12587 36091
rect 12621 36057 12633 36091
rect 12710 36088 12716 36100
rect 12671 36060 12716 36088
rect 12584 36051 12633 36057
rect 12584 36048 12590 36051
rect 12710 36048 12716 36060
rect 12768 36048 12774 36100
rect 13740 36020 13768 36264
rect 24305 36261 24317 36264
rect 24351 36261 24363 36295
rect 24305 36255 24363 36261
rect 24394 36252 24400 36304
rect 24452 36292 24458 36304
rect 24452 36264 28948 36292
rect 24452 36252 24458 36264
rect 13906 36184 13912 36236
rect 13964 36224 13970 36236
rect 14001 36227 14059 36233
rect 14001 36224 14013 36227
rect 13964 36196 14013 36224
rect 13964 36184 13970 36196
rect 14001 36193 14013 36196
rect 14047 36193 14059 36227
rect 14001 36187 14059 36193
rect 17865 36227 17923 36233
rect 17865 36193 17877 36227
rect 17911 36224 17923 36227
rect 18414 36224 18420 36236
rect 17911 36196 18420 36224
rect 17911 36193 17923 36196
rect 17865 36187 17923 36193
rect 18414 36184 18420 36196
rect 18472 36184 18478 36236
rect 18601 36227 18659 36233
rect 18601 36193 18613 36227
rect 18647 36224 18659 36227
rect 19153 36227 19211 36233
rect 19153 36224 19165 36227
rect 18647 36196 19165 36224
rect 18647 36193 18659 36196
rect 18601 36187 18659 36193
rect 19153 36193 19165 36196
rect 19199 36193 19211 36227
rect 20898 36224 20904 36236
rect 20859 36196 20904 36224
rect 19153 36187 19211 36193
rect 17681 36159 17739 36165
rect 17681 36156 17693 36159
rect 17512 36128 17693 36156
rect 14182 36088 14188 36100
rect 14095 36060 14188 36088
rect 14182 36048 14188 36060
rect 14240 36088 14246 36100
rect 15562 36088 15568 36100
rect 14240 36060 15568 36088
rect 14240 36048 14246 36060
rect 15562 36048 15568 36060
rect 15620 36048 15626 36100
rect 13906 36020 13912 36032
rect 9140 35992 13768 36020
rect 13867 35992 13912 36020
rect 9033 35983 9091 35989
rect 13906 35980 13912 35992
rect 13964 35980 13970 36032
rect 17310 35980 17316 36032
rect 17368 36020 17374 36032
rect 17512 36029 17540 36128
rect 17681 36125 17693 36128
rect 17727 36125 17739 36159
rect 19168 36156 19196 36187
rect 20898 36184 20904 36196
rect 20956 36184 20962 36236
rect 24118 36224 24124 36236
rect 24079 36196 24124 36224
rect 24118 36184 24124 36196
rect 24176 36184 24182 36236
rect 24949 36227 25007 36233
rect 24949 36193 24961 36227
rect 24995 36224 25007 36227
rect 25038 36224 25044 36236
rect 24995 36196 25044 36224
rect 24995 36193 25007 36196
rect 24949 36187 25007 36193
rect 25038 36184 25044 36196
rect 25096 36184 25102 36236
rect 25317 36227 25375 36233
rect 25317 36193 25329 36227
rect 25363 36224 25375 36227
rect 25406 36224 25412 36236
rect 25363 36196 25412 36224
rect 25363 36193 25375 36196
rect 25317 36187 25375 36193
rect 25406 36184 25412 36196
rect 25464 36184 25470 36236
rect 25516 36233 25544 36264
rect 25501 36227 25559 36233
rect 25501 36193 25513 36227
rect 25547 36193 25559 36227
rect 26970 36224 26976 36236
rect 26931 36196 26976 36224
rect 25501 36187 25559 36193
rect 26970 36184 26976 36196
rect 27028 36184 27034 36236
rect 19168 36128 20300 36156
rect 17681 36119 17739 36125
rect 18782 36088 18788 36100
rect 18743 36060 18788 36088
rect 18782 36048 18788 36060
rect 18840 36048 18846 36100
rect 18874 36048 18880 36100
rect 18932 36088 18938 36100
rect 20162 36088 20168 36100
rect 18932 36060 20168 36088
rect 18932 36048 18938 36060
rect 20162 36048 20168 36060
rect 20220 36048 20226 36100
rect 17497 36023 17555 36029
rect 17497 36020 17509 36023
rect 17368 35992 17509 36020
rect 17368 35980 17374 35992
rect 17497 35989 17509 35992
rect 17543 35989 17555 36023
rect 17497 35983 17555 35989
rect 18138 35980 18144 36032
rect 18196 36020 18202 36032
rect 19242 36020 19248 36032
rect 18196 35992 19248 36020
rect 18196 35980 18202 35992
rect 19242 35980 19248 35992
rect 19300 36020 19306 36032
rect 20070 36020 20076 36032
rect 19300 35992 20076 36020
rect 19300 35980 19306 35992
rect 20070 35980 20076 35992
rect 20128 35980 20134 36032
rect 20272 36020 20300 36128
rect 20714 36116 20720 36168
rect 20772 36156 20778 36168
rect 24029 36159 24087 36165
rect 24029 36156 24041 36159
rect 20772 36128 24041 36156
rect 20772 36116 20778 36128
rect 24029 36125 24041 36128
rect 24075 36156 24087 36159
rect 24857 36159 24915 36165
rect 24857 36156 24869 36159
rect 24075 36128 24869 36156
rect 24075 36125 24087 36128
rect 24029 36119 24087 36125
rect 24857 36125 24869 36128
rect 24903 36156 24915 36159
rect 25130 36156 25136 36168
rect 24903 36128 25136 36156
rect 24903 36125 24915 36128
rect 24857 36119 24915 36125
rect 25130 36116 25136 36128
rect 25188 36116 25194 36168
rect 28813 36159 28871 36165
rect 28813 36125 28825 36159
rect 28859 36125 28871 36159
rect 28813 36119 28871 36125
rect 23842 36088 23848 36100
rect 22204 36060 23848 36088
rect 20993 36023 21051 36029
rect 20993 36020 21005 36023
rect 20272 35992 21005 36020
rect 20993 35989 21005 35992
rect 21039 36020 21051 36023
rect 22204 36020 22232 36060
rect 23842 36048 23848 36060
rect 23900 36048 23906 36100
rect 25406 36048 25412 36100
rect 25464 36088 25470 36100
rect 27154 36088 27160 36100
rect 25464 36060 27160 36088
rect 25464 36048 25470 36060
rect 27154 36048 27160 36060
rect 27212 36048 27218 36100
rect 21039 35992 22232 36020
rect 21039 35989 21051 35992
rect 20993 35983 21051 35989
rect 28442 35980 28448 36032
rect 28500 36020 28506 36032
rect 28629 36023 28687 36029
rect 28629 36020 28641 36023
rect 28500 35992 28641 36020
rect 28500 35980 28506 35992
rect 28629 35989 28641 35992
rect 28675 36020 28687 36023
rect 28828 36020 28856 36119
rect 28920 36088 28948 36264
rect 29012 36233 29040 36332
rect 29086 36320 29092 36372
rect 29144 36360 29150 36372
rect 29144 36332 29592 36360
rect 29144 36320 29150 36332
rect 29564 36292 29592 36332
rect 29638 36320 29644 36372
rect 29696 36360 29702 36372
rect 36633 36363 36691 36369
rect 29696 36332 36584 36360
rect 29696 36320 29702 36332
rect 31113 36295 31171 36301
rect 31113 36292 31125 36295
rect 29564 36264 31125 36292
rect 28997 36227 29055 36233
rect 28997 36193 29009 36227
rect 29043 36224 29055 36227
rect 29362 36224 29368 36236
rect 29043 36196 29368 36224
rect 29043 36193 29055 36196
rect 28997 36187 29055 36193
rect 29362 36184 29368 36196
rect 29420 36184 29426 36236
rect 29546 36184 29552 36236
rect 29604 36224 29610 36236
rect 29748 36233 29776 36264
rect 31113 36261 31125 36264
rect 31159 36261 31171 36295
rect 36446 36292 36452 36304
rect 31113 36255 31171 36261
rect 36188 36264 36452 36292
rect 29733 36227 29791 36233
rect 29604 36196 29649 36224
rect 29604 36184 29610 36196
rect 29733 36193 29745 36227
rect 29779 36193 29791 36227
rect 29733 36187 29791 36193
rect 31021 36227 31079 36233
rect 31021 36193 31033 36227
rect 31067 36224 31079 36227
rect 31938 36224 31944 36236
rect 31067 36196 31944 36224
rect 31067 36193 31079 36196
rect 31021 36187 31079 36193
rect 31938 36184 31944 36196
rect 31996 36184 32002 36236
rect 32122 36224 32128 36236
rect 32083 36196 32128 36224
rect 32122 36184 32128 36196
rect 32180 36184 32186 36236
rect 35618 36224 35624 36236
rect 35531 36196 35624 36224
rect 35618 36184 35624 36196
rect 35676 36224 35682 36236
rect 36188 36233 36216 36264
rect 36446 36252 36452 36264
rect 36504 36252 36510 36304
rect 36556 36292 36584 36332
rect 36633 36329 36645 36363
rect 36679 36360 36691 36363
rect 47302 36360 47308 36372
rect 36679 36332 47308 36360
rect 36679 36329 36691 36332
rect 36633 36323 36691 36329
rect 47302 36320 47308 36332
rect 47360 36320 47366 36372
rect 50985 36363 51043 36369
rect 50985 36360 50997 36363
rect 50172 36332 50997 36360
rect 43438 36292 43444 36304
rect 36556 36264 43444 36292
rect 43438 36252 43444 36264
rect 43496 36252 43502 36304
rect 44910 36252 44916 36304
rect 44968 36292 44974 36304
rect 45005 36295 45063 36301
rect 45005 36292 45017 36295
rect 44968 36264 45017 36292
rect 44968 36252 44974 36264
rect 45005 36261 45017 36264
rect 45051 36261 45063 36295
rect 45005 36255 45063 36261
rect 50172 36236 50200 36332
rect 50985 36329 50997 36332
rect 51031 36360 51043 36363
rect 51810 36360 51816 36372
rect 51031 36332 51816 36360
rect 51031 36329 51043 36332
rect 50985 36323 51043 36329
rect 51810 36320 51816 36332
rect 51868 36320 51874 36372
rect 54846 36320 54852 36372
rect 54904 36360 54910 36372
rect 57517 36363 57575 36369
rect 57517 36360 57529 36363
rect 54904 36332 57529 36360
rect 54904 36320 54910 36332
rect 57517 36329 57529 36332
rect 57563 36329 57575 36363
rect 57517 36323 57575 36329
rect 59173 36363 59231 36369
rect 59173 36329 59185 36363
rect 59219 36360 59231 36363
rect 60734 36360 60740 36372
rect 59219 36332 60740 36360
rect 59219 36329 59231 36332
rect 59173 36323 59231 36329
rect 60734 36320 60740 36332
rect 60792 36320 60798 36372
rect 60826 36320 60832 36372
rect 60884 36360 60890 36372
rect 62301 36363 62359 36369
rect 62301 36360 62313 36363
rect 60884 36332 62313 36360
rect 60884 36320 60890 36332
rect 62301 36329 62313 36332
rect 62347 36360 62359 36363
rect 63310 36360 63316 36372
rect 62347 36332 63316 36360
rect 62347 36329 62359 36332
rect 62301 36323 62359 36329
rect 63310 36320 63316 36332
rect 63368 36320 63374 36372
rect 71498 36360 71504 36372
rect 71459 36332 71504 36360
rect 71498 36320 71504 36332
rect 71556 36320 71562 36372
rect 72881 36363 72939 36369
rect 72881 36329 72893 36363
rect 72927 36360 72939 36363
rect 83734 36360 83740 36372
rect 72927 36332 83740 36360
rect 72927 36329 72939 36332
rect 72881 36323 72939 36329
rect 83734 36320 83740 36332
rect 83792 36320 83798 36372
rect 88797 36363 88855 36369
rect 88797 36360 88809 36363
rect 84304 36332 88809 36360
rect 50706 36292 50712 36304
rect 50667 36264 50712 36292
rect 50706 36252 50712 36264
rect 50764 36252 50770 36304
rect 51074 36252 51080 36304
rect 51132 36292 51138 36304
rect 51132 36264 51672 36292
rect 51132 36252 51138 36264
rect 51644 36236 51672 36264
rect 53374 36252 53380 36304
rect 53432 36292 53438 36304
rect 53432 36264 75868 36292
rect 53432 36252 53438 36264
rect 36173 36227 36231 36233
rect 36173 36224 36185 36227
rect 35676 36196 36185 36224
rect 35676 36184 35682 36196
rect 36173 36193 36185 36196
rect 36219 36193 36231 36227
rect 36173 36187 36231 36193
rect 36357 36227 36415 36233
rect 36357 36193 36369 36227
rect 36403 36224 36415 36227
rect 36909 36227 36967 36233
rect 36909 36224 36921 36227
rect 36403 36196 36921 36224
rect 36403 36193 36415 36196
rect 36357 36187 36415 36193
rect 31754 36116 31760 36168
rect 31812 36156 31818 36168
rect 31812 36128 34560 36156
rect 31812 36116 31818 36128
rect 29638 36088 29644 36100
rect 28920 36060 29644 36088
rect 29638 36048 29644 36060
rect 29696 36048 29702 36100
rect 30098 36048 30104 36100
rect 30156 36088 30162 36100
rect 32217 36091 32275 36097
rect 32217 36088 32229 36091
rect 30156 36060 32229 36088
rect 30156 36048 30162 36060
rect 32217 36057 32229 36060
rect 32263 36057 32275 36091
rect 34532 36088 34560 36128
rect 35342 36116 35348 36168
rect 35400 36156 35406 36168
rect 35437 36159 35495 36165
rect 35437 36156 35449 36159
rect 35400 36128 35449 36156
rect 35400 36116 35406 36128
rect 35437 36125 35449 36128
rect 35483 36125 35495 36159
rect 35437 36119 35495 36125
rect 36556 36088 36584 36196
rect 36909 36193 36921 36196
rect 36955 36224 36967 36227
rect 38102 36224 38108 36236
rect 36955 36196 38108 36224
rect 36955 36193 36967 36196
rect 36909 36187 36967 36193
rect 38102 36184 38108 36196
rect 38160 36184 38166 36236
rect 39025 36227 39083 36233
rect 39025 36193 39037 36227
rect 39071 36224 39083 36227
rect 39390 36224 39396 36236
rect 39071 36196 39396 36224
rect 39071 36193 39083 36196
rect 39025 36187 39083 36193
rect 39390 36184 39396 36196
rect 39448 36184 39454 36236
rect 42794 36184 42800 36236
rect 42852 36224 42858 36236
rect 43165 36227 43223 36233
rect 43165 36224 43177 36227
rect 42852 36196 43177 36224
rect 42852 36184 42858 36196
rect 43165 36193 43177 36196
rect 43211 36224 43223 36227
rect 43346 36224 43352 36236
rect 43211 36196 43352 36224
rect 43211 36193 43223 36196
rect 43165 36187 43223 36193
rect 43346 36184 43352 36196
rect 43404 36184 43410 36236
rect 49605 36227 49663 36233
rect 49605 36193 49617 36227
rect 49651 36224 49663 36227
rect 49970 36224 49976 36236
rect 49651 36196 49976 36224
rect 49651 36193 49663 36196
rect 49605 36187 49663 36193
rect 49970 36184 49976 36196
rect 50028 36184 50034 36236
rect 50154 36224 50160 36236
rect 50067 36196 50160 36224
rect 50154 36184 50160 36196
rect 50212 36184 50218 36236
rect 50338 36224 50344 36236
rect 50299 36196 50344 36224
rect 50338 36184 50344 36196
rect 50396 36184 50402 36236
rect 51626 36184 51632 36236
rect 51684 36224 51690 36236
rect 52730 36224 52736 36236
rect 51684 36196 52736 36224
rect 51684 36184 51690 36196
rect 52730 36184 52736 36196
rect 52788 36224 52794 36236
rect 54110 36224 54116 36236
rect 52788 36196 54116 36224
rect 52788 36184 52794 36196
rect 54110 36184 54116 36196
rect 54168 36224 54174 36236
rect 56505 36227 56563 36233
rect 54168 36196 56456 36224
rect 54168 36184 54174 36196
rect 38930 36116 38936 36168
rect 38988 36156 38994 36168
rect 39117 36159 39175 36165
rect 39117 36156 39129 36159
rect 38988 36128 39129 36156
rect 38988 36116 38994 36128
rect 39117 36125 39129 36128
rect 39163 36125 39175 36159
rect 43622 36156 43628 36168
rect 43583 36128 43628 36156
rect 39117 36119 39175 36125
rect 43622 36116 43628 36128
rect 43680 36116 43686 36168
rect 49421 36159 49479 36165
rect 49421 36156 49433 36159
rect 49068 36128 49433 36156
rect 34532 36060 36584 36088
rect 32217 36051 32275 36057
rect 28675 35992 28856 36020
rect 30009 36023 30067 36029
rect 28675 35989 28687 35992
rect 28629 35983 28687 35989
rect 30009 35989 30021 36023
rect 30055 36020 30067 36023
rect 30558 36020 30564 36032
rect 30055 35992 30564 36020
rect 30055 35989 30067 35992
rect 30009 35983 30067 35989
rect 30558 35980 30564 35992
rect 30616 35980 30622 36032
rect 35342 36020 35348 36032
rect 35303 35992 35348 36020
rect 35342 35980 35348 35992
rect 35400 35980 35406 36032
rect 48774 35980 48780 36032
rect 48832 36020 48838 36032
rect 49068 36029 49096 36128
rect 49421 36125 49433 36128
rect 49467 36125 49479 36159
rect 56321 36159 56379 36165
rect 56321 36156 56333 36159
rect 49421 36119 49479 36125
rect 55968 36128 56333 36156
rect 55968 36032 55996 36128
rect 56321 36125 56333 36128
rect 56367 36125 56379 36159
rect 56321 36119 56379 36125
rect 49053 36023 49111 36029
rect 49053 36020 49065 36023
rect 48832 35992 49065 36020
rect 48832 35980 48838 35992
rect 49053 35989 49065 35992
rect 49099 35989 49111 36023
rect 49053 35983 49111 35989
rect 49329 36023 49387 36029
rect 49329 35989 49341 36023
rect 49375 36020 49387 36023
rect 49510 36020 49516 36032
rect 49375 35992 49516 36020
rect 49375 35989 49387 35992
rect 49329 35983 49387 35989
rect 49510 35980 49516 35992
rect 49568 36020 49574 36032
rect 50338 36020 50344 36032
rect 49568 35992 50344 36020
rect 49568 35980 49574 35992
rect 50338 35980 50344 35992
rect 50396 35980 50402 36032
rect 51166 36020 51172 36032
rect 51127 35992 51172 36020
rect 51166 35980 51172 35992
rect 51224 35980 51230 36032
rect 55950 36020 55956 36032
rect 55911 35992 55956 36020
rect 55950 35980 55956 35992
rect 56008 35980 56014 36032
rect 56226 36020 56232 36032
rect 56187 35992 56232 36020
rect 56226 35980 56232 35992
rect 56284 35980 56290 36032
rect 56428 36020 56456 36196
rect 56505 36193 56517 36227
rect 56551 36193 56563 36227
rect 56505 36187 56563 36193
rect 56520 36088 56548 36187
rect 56594 36184 56600 36236
rect 56652 36224 56658 36236
rect 56965 36227 57023 36233
rect 56965 36224 56977 36227
rect 56652 36196 56977 36224
rect 56652 36184 56658 36196
rect 56965 36193 56977 36196
rect 57011 36193 57023 36227
rect 56965 36187 57023 36193
rect 57057 36227 57115 36233
rect 57057 36193 57069 36227
rect 57103 36224 57115 36227
rect 58526 36224 58532 36236
rect 57103 36196 57836 36224
rect 58487 36196 58532 36224
rect 57103 36193 57115 36196
rect 57057 36187 57115 36193
rect 57808 36168 57836 36196
rect 58526 36184 58532 36196
rect 58584 36184 58590 36236
rect 58618 36184 58624 36236
rect 58676 36224 58682 36236
rect 62485 36227 62543 36233
rect 62485 36224 62497 36227
rect 58676 36196 62497 36224
rect 58676 36184 58682 36196
rect 62485 36193 62497 36196
rect 62531 36224 62543 36227
rect 62531 36196 63264 36224
rect 62531 36193 62543 36196
rect 62485 36187 62543 36193
rect 57790 36156 57796 36168
rect 57751 36128 57796 36156
rect 57790 36116 57796 36128
rect 57848 36116 57854 36168
rect 58897 36159 58955 36165
rect 58897 36125 58909 36159
rect 58943 36156 58955 36159
rect 59814 36156 59820 36168
rect 58943 36128 59820 36156
rect 58943 36125 58955 36128
rect 58897 36119 58955 36125
rect 59814 36116 59820 36128
rect 59872 36116 59878 36168
rect 62666 36156 62672 36168
rect 62627 36128 62672 36156
rect 62666 36116 62672 36128
rect 62724 36116 62730 36168
rect 63126 36156 63132 36168
rect 63087 36128 63132 36156
rect 63126 36116 63132 36128
rect 63184 36116 63190 36168
rect 63236 36156 63264 36196
rect 63310 36184 63316 36236
rect 63368 36224 63374 36236
rect 63681 36227 63739 36233
rect 63368 36196 63413 36224
rect 63368 36184 63374 36196
rect 63681 36193 63693 36227
rect 63727 36193 63739 36227
rect 63862 36224 63868 36236
rect 63823 36196 63868 36224
rect 63681 36187 63739 36193
rect 63494 36156 63500 36168
rect 63236 36128 63500 36156
rect 63494 36116 63500 36128
rect 63552 36156 63558 36168
rect 63696 36156 63724 36187
rect 63862 36184 63868 36196
rect 63920 36184 63926 36236
rect 66070 36184 66076 36236
rect 66128 36224 66134 36236
rect 69845 36227 69903 36233
rect 69845 36224 69857 36227
rect 66128 36196 69857 36224
rect 66128 36184 66134 36196
rect 69845 36193 69857 36196
rect 69891 36224 69903 36227
rect 71314 36224 71320 36236
rect 69891 36196 71320 36224
rect 69891 36193 69903 36196
rect 69845 36187 69903 36193
rect 71314 36184 71320 36196
rect 71372 36184 71378 36236
rect 71409 36227 71467 36233
rect 71409 36193 71421 36227
rect 71455 36224 71467 36227
rect 71774 36224 71780 36236
rect 71455 36196 71780 36224
rect 71455 36193 71467 36196
rect 71409 36187 71467 36193
rect 71774 36184 71780 36196
rect 71832 36224 71838 36236
rect 72326 36224 72332 36236
rect 71832 36196 72332 36224
rect 71832 36184 71838 36196
rect 72326 36184 72332 36196
rect 72384 36184 72390 36236
rect 73062 36224 73068 36236
rect 73023 36196 73068 36224
rect 73062 36184 73068 36196
rect 73120 36224 73126 36236
rect 73617 36227 73675 36233
rect 73617 36224 73629 36227
rect 73120 36196 73629 36224
rect 73120 36184 73126 36196
rect 73617 36193 73629 36196
rect 73663 36193 73675 36227
rect 73617 36187 73675 36193
rect 64414 36156 64420 36168
rect 63552 36128 64420 36156
rect 63552 36116 63558 36128
rect 64414 36116 64420 36128
rect 64472 36116 64478 36168
rect 69937 36159 69995 36165
rect 69937 36125 69949 36159
rect 69983 36156 69995 36159
rect 70486 36156 70492 36168
rect 69983 36128 70492 36156
rect 69983 36125 69995 36128
rect 69937 36119 69995 36125
rect 70486 36116 70492 36128
rect 70544 36116 70550 36168
rect 72973 36159 73031 36165
rect 72973 36125 72985 36159
rect 73019 36156 73031 36159
rect 73154 36156 73160 36168
rect 73019 36128 73160 36156
rect 73019 36125 73031 36128
rect 72973 36119 73031 36125
rect 73154 36116 73160 36128
rect 73212 36156 73218 36168
rect 73801 36159 73859 36165
rect 73801 36156 73813 36159
rect 73212 36128 73813 36156
rect 73212 36116 73218 36128
rect 73801 36125 73813 36128
rect 73847 36125 73859 36159
rect 73801 36119 73859 36125
rect 58069 36091 58127 36097
rect 58069 36088 58081 36091
rect 56520 36060 58081 36088
rect 58069 36057 58081 36060
rect 58115 36088 58127 36091
rect 72881 36091 72939 36097
rect 72881 36088 72893 36091
rect 58115 36060 72893 36088
rect 58115 36057 58127 36060
rect 58069 36051 58127 36057
rect 72881 36057 72893 36060
rect 72927 36057 72939 36091
rect 72881 36051 72939 36057
rect 58434 36020 58440 36032
rect 56428 35992 58440 36020
rect 58434 35980 58440 35992
rect 58492 35980 58498 36032
rect 58618 35980 58624 36032
rect 58676 36029 58682 36032
rect 58676 36023 58725 36029
rect 58676 35989 58679 36023
rect 58713 35989 58725 36023
rect 58802 36020 58808 36032
rect 58763 35992 58808 36020
rect 58676 35983 58725 35989
rect 58676 35980 58682 35983
rect 58802 35980 58808 35992
rect 58860 35980 58866 36032
rect 70210 35980 70216 36032
rect 70268 36020 70274 36032
rect 71498 36020 71504 36032
rect 70268 35992 71504 36020
rect 70268 35980 70274 35992
rect 71498 35980 71504 35992
rect 71556 35980 71562 36032
rect 73246 36020 73252 36032
rect 73207 35992 73252 36020
rect 73246 35980 73252 35992
rect 73304 35980 73310 36032
rect 75840 36020 75868 36264
rect 77662 36252 77668 36304
rect 77720 36292 77726 36304
rect 79321 36295 79379 36301
rect 79321 36292 79333 36295
rect 77720 36264 79333 36292
rect 77720 36252 77726 36264
rect 79321 36261 79333 36264
rect 79367 36292 79379 36295
rect 80054 36292 80060 36304
rect 79367 36264 80060 36292
rect 79367 36261 79379 36264
rect 79321 36255 79379 36261
rect 80054 36252 80060 36264
rect 80112 36252 80118 36304
rect 81710 36252 81716 36304
rect 81768 36292 81774 36304
rect 84304 36292 84332 36332
rect 81768 36264 84332 36292
rect 81768 36252 81774 36264
rect 77570 36224 77576 36236
rect 77531 36196 77576 36224
rect 77570 36184 77576 36196
rect 77628 36184 77634 36236
rect 78217 36227 78275 36233
rect 78217 36193 78229 36227
rect 78263 36224 78275 36227
rect 78493 36227 78551 36233
rect 78493 36224 78505 36227
rect 78263 36196 78505 36224
rect 78263 36193 78275 36196
rect 78217 36187 78275 36193
rect 78493 36193 78505 36196
rect 78539 36224 78551 36227
rect 78766 36224 78772 36236
rect 78539 36196 78772 36224
rect 78539 36193 78551 36196
rect 78493 36187 78551 36193
rect 75914 36116 75920 36168
rect 75972 36156 75978 36168
rect 77846 36156 77852 36168
rect 75972 36128 77852 36156
rect 75972 36116 75978 36128
rect 77846 36116 77852 36128
rect 77904 36116 77910 36168
rect 77941 36159 77999 36165
rect 77941 36125 77953 36159
rect 77987 36156 77999 36159
rect 78030 36156 78036 36168
rect 77987 36128 78036 36156
rect 77987 36125 77999 36128
rect 77941 36119 77999 36125
rect 78030 36116 78036 36128
rect 78088 36116 78094 36168
rect 77938 36020 77944 36032
rect 75840 35992 77944 36020
rect 77938 35980 77944 35992
rect 77996 36020 78002 36032
rect 78232 36020 78260 36187
rect 78766 36184 78772 36196
rect 78824 36184 78830 36236
rect 79226 36224 79232 36236
rect 79187 36196 79232 36224
rect 79226 36184 79232 36196
rect 79284 36184 79290 36236
rect 79413 36227 79471 36233
rect 79413 36193 79425 36227
rect 79459 36193 79471 36227
rect 84470 36224 84476 36236
rect 84431 36196 84476 36224
rect 79413 36187 79471 36193
rect 78306 36116 78312 36168
rect 78364 36156 78370 36168
rect 79428 36156 79456 36187
rect 84470 36184 84476 36196
rect 84528 36184 84534 36236
rect 85853 36227 85911 36233
rect 85853 36193 85865 36227
rect 85899 36224 85911 36227
rect 86681 36227 86739 36233
rect 86681 36224 86693 36227
rect 85899 36196 86693 36224
rect 85899 36193 85911 36196
rect 85853 36187 85911 36193
rect 86681 36193 86693 36196
rect 86727 36193 86739 36227
rect 88352 36224 88380 36332
rect 88797 36329 88809 36332
rect 88843 36329 88855 36363
rect 97258 36360 97264 36372
rect 97219 36332 97264 36360
rect 88797 36323 88855 36329
rect 97258 36320 97264 36332
rect 97316 36320 97322 36372
rect 88426 36252 88432 36304
rect 88484 36292 88490 36304
rect 89165 36295 89223 36301
rect 89165 36292 89177 36295
rect 88484 36264 89177 36292
rect 88484 36252 88490 36264
rect 89165 36261 89177 36264
rect 89211 36261 89223 36295
rect 89165 36255 89223 36261
rect 88981 36227 89039 36233
rect 88981 36224 88993 36227
rect 88352 36196 88993 36224
rect 86681 36187 86739 36193
rect 88981 36193 88993 36196
rect 89027 36193 89039 36227
rect 88981 36187 89039 36193
rect 89257 36227 89315 36233
rect 89257 36193 89269 36227
rect 89303 36224 89315 36227
rect 89714 36224 89720 36236
rect 89303 36196 89720 36224
rect 89303 36193 89315 36196
rect 89257 36187 89315 36193
rect 84197 36159 84255 36165
rect 84197 36156 84209 36159
rect 78364 36128 79456 36156
rect 84028 36128 84209 36156
rect 78364 36116 78370 36128
rect 79594 36020 79600 36032
rect 77996 35992 78260 36020
rect 79555 35992 79600 36020
rect 77996 35980 78002 35992
rect 79594 35980 79600 35992
rect 79652 35980 79658 36032
rect 82538 35980 82544 36032
rect 82596 36020 82602 36032
rect 84028 36029 84056 36128
rect 84197 36125 84209 36128
rect 84243 36156 84255 36159
rect 86218 36156 86224 36168
rect 84243 36128 86224 36156
rect 84243 36125 84255 36128
rect 84197 36119 84255 36125
rect 86218 36116 86224 36128
rect 86276 36116 86282 36168
rect 88996 36156 89024 36187
rect 89714 36184 89720 36196
rect 89772 36184 89778 36236
rect 90545 36227 90603 36233
rect 90545 36193 90557 36227
rect 90591 36224 90603 36227
rect 91738 36224 91744 36236
rect 90591 36196 91744 36224
rect 90591 36193 90603 36196
rect 90545 36187 90603 36193
rect 91738 36184 91744 36196
rect 91796 36184 91802 36236
rect 92750 36224 92756 36236
rect 92711 36196 92756 36224
rect 92750 36184 92756 36196
rect 92808 36184 92814 36236
rect 92845 36227 92903 36233
rect 92845 36193 92857 36227
rect 92891 36224 92903 36227
rect 94869 36227 94927 36233
rect 94869 36224 94881 36227
rect 92891 36196 94881 36224
rect 92891 36193 92903 36196
rect 92845 36187 92903 36193
rect 94869 36193 94881 36196
rect 94915 36193 94927 36227
rect 97074 36224 97080 36236
rect 97035 36196 97080 36224
rect 94869 36187 94927 36193
rect 97074 36184 97080 36196
rect 97132 36184 97138 36236
rect 90726 36156 90732 36168
rect 88996 36128 90732 36156
rect 90726 36116 90732 36128
rect 90784 36116 90790 36168
rect 94590 36156 94596 36168
rect 94424 36128 94596 36156
rect 84013 36023 84071 36029
rect 84013 36020 84025 36023
rect 82596 35992 84025 36020
rect 82596 35980 82602 35992
rect 84013 35989 84025 35992
rect 84059 35989 84071 36023
rect 86770 36020 86776 36032
rect 86731 35992 86776 36020
rect 84013 35983 84071 35989
rect 86770 35980 86776 35992
rect 86828 35980 86834 36032
rect 89441 36023 89499 36029
rect 89441 35989 89453 36023
rect 89487 36020 89499 36023
rect 89530 36020 89536 36032
rect 89487 35992 89536 36020
rect 89487 35989 89499 35992
rect 89441 35983 89499 35989
rect 89530 35980 89536 35992
rect 89588 35980 89594 36032
rect 90634 36020 90640 36032
rect 90595 35992 90640 36020
rect 90634 35980 90640 35992
rect 90692 35980 90698 36032
rect 93946 35980 93952 36032
rect 94004 36020 94010 36032
rect 94424 36029 94452 36128
rect 94590 36116 94596 36128
rect 94648 36116 94654 36168
rect 94409 36023 94467 36029
rect 94409 36020 94421 36023
rect 94004 35992 94421 36020
rect 94004 35980 94010 35992
rect 94409 35989 94421 35992
rect 94455 35989 94467 36023
rect 94409 35983 94467 35989
rect 96157 36023 96215 36029
rect 96157 35989 96169 36023
rect 96203 36020 96215 36023
rect 96706 36020 96712 36032
rect 96203 35992 96712 36020
rect 96203 35989 96215 35992
rect 96157 35983 96215 35989
rect 96706 35980 96712 35992
rect 96764 35980 96770 36032
rect 1104 35930 105616 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 65686 35930
rect 65738 35878 65750 35930
rect 65802 35878 65814 35930
rect 65866 35878 65878 35930
rect 65930 35878 96406 35930
rect 96458 35878 96470 35930
rect 96522 35878 96534 35930
rect 96586 35878 96598 35930
rect 96650 35878 105616 35930
rect 1104 35856 105616 35878
rect 9769 35819 9827 35825
rect 9769 35785 9781 35819
rect 9815 35816 9827 35819
rect 19613 35819 19671 35825
rect 9815 35788 19012 35816
rect 9815 35785 9827 35788
rect 9769 35779 9827 35785
rect 5166 35708 5172 35760
rect 5224 35748 5230 35760
rect 7193 35751 7251 35757
rect 7193 35748 7205 35751
rect 5224 35720 7205 35748
rect 5224 35708 5230 35720
rect 7193 35717 7205 35720
rect 7239 35717 7251 35751
rect 7193 35711 7251 35717
rect 2777 35683 2835 35689
rect 2777 35649 2789 35683
rect 2823 35680 2835 35683
rect 2866 35680 2872 35692
rect 2823 35652 2872 35680
rect 2823 35649 2835 35652
rect 2777 35643 2835 35649
rect 2866 35640 2872 35652
rect 2924 35640 2930 35692
rect 7742 35640 7748 35692
rect 7800 35680 7806 35692
rect 7929 35683 7987 35689
rect 7929 35680 7941 35683
rect 7800 35652 7941 35680
rect 7800 35640 7806 35652
rect 7929 35649 7941 35652
rect 7975 35649 7987 35683
rect 9493 35683 9551 35689
rect 9493 35680 9505 35683
rect 7929 35643 7987 35649
rect 8496 35652 9505 35680
rect 2501 35615 2559 35621
rect 2501 35581 2513 35615
rect 2547 35612 2559 35615
rect 4154 35612 4160 35624
rect 2547 35584 4160 35612
rect 2547 35581 2559 35584
rect 2501 35575 2559 35581
rect 4154 35572 4160 35584
rect 4212 35572 4218 35624
rect 5445 35615 5503 35621
rect 5445 35581 5457 35615
rect 5491 35612 5503 35615
rect 5534 35612 5540 35624
rect 5491 35584 5540 35612
rect 5491 35581 5503 35584
rect 5445 35575 5503 35581
rect 5534 35572 5540 35584
rect 5592 35572 5598 35624
rect 5718 35612 5724 35624
rect 5679 35584 5724 35612
rect 5718 35572 5724 35584
rect 5776 35572 5782 35624
rect 7098 35612 7104 35624
rect 7059 35584 7104 35612
rect 7098 35572 7104 35584
rect 7156 35572 7162 35624
rect 7837 35615 7895 35621
rect 7837 35581 7849 35615
rect 7883 35612 7895 35615
rect 8496 35612 8524 35652
rect 9493 35649 9505 35652
rect 9539 35649 9551 35683
rect 9493 35643 9551 35649
rect 7883 35584 8524 35612
rect 9217 35615 9275 35621
rect 7883 35581 7895 35584
rect 7837 35575 7895 35581
rect 9217 35581 9229 35615
rect 9263 35612 9275 35615
rect 9784 35612 9812 35779
rect 15194 35748 15200 35760
rect 11164 35720 15200 35748
rect 9263 35584 9812 35612
rect 9263 35581 9275 35584
rect 9217 35575 9275 35581
rect 10870 35572 10876 35624
rect 10928 35612 10934 35624
rect 10965 35615 11023 35621
rect 10965 35612 10977 35615
rect 10928 35584 10977 35612
rect 10928 35572 10934 35584
rect 10965 35581 10977 35584
rect 11011 35581 11023 35615
rect 10965 35575 11023 35581
rect 3970 35504 3976 35556
rect 4028 35544 4034 35556
rect 9033 35547 9091 35553
rect 4028 35516 5304 35544
rect 4028 35504 4034 35516
rect 3234 35436 3240 35488
rect 3292 35476 3298 35488
rect 3881 35479 3939 35485
rect 3881 35476 3893 35479
rect 3292 35448 3893 35476
rect 3292 35436 3298 35448
rect 3881 35445 3893 35448
rect 3927 35445 3939 35479
rect 3881 35439 3939 35445
rect 4154 35436 4160 35488
rect 4212 35476 4218 35488
rect 4341 35479 4399 35485
rect 4341 35476 4353 35479
rect 4212 35448 4353 35476
rect 4212 35436 4218 35448
rect 4341 35445 4353 35448
rect 4387 35476 4399 35479
rect 4706 35476 4712 35488
rect 4387 35448 4712 35476
rect 4387 35445 4399 35448
rect 4341 35439 4399 35445
rect 4706 35436 4712 35448
rect 4764 35436 4770 35488
rect 5276 35485 5304 35516
rect 9033 35513 9045 35547
rect 9079 35544 9091 35547
rect 9582 35544 9588 35556
rect 9079 35516 9588 35544
rect 9079 35513 9091 35516
rect 9033 35507 9091 35513
rect 9582 35504 9588 35516
rect 9640 35544 9646 35556
rect 11164 35544 11192 35720
rect 15194 35708 15200 35720
rect 15252 35708 15258 35760
rect 12802 35680 12808 35692
rect 12763 35652 12808 35680
rect 12802 35640 12808 35652
rect 12860 35640 12866 35692
rect 13998 35680 14004 35692
rect 13556 35652 14004 35680
rect 11422 35572 11428 35624
rect 11480 35612 11486 35624
rect 13556 35621 13584 35652
rect 13998 35640 14004 35652
rect 14056 35640 14062 35692
rect 15289 35683 15347 35689
rect 15289 35649 15301 35683
rect 15335 35680 15347 35683
rect 16025 35683 16083 35689
rect 16025 35680 16037 35683
rect 15335 35652 16037 35680
rect 15335 35649 15347 35652
rect 15289 35643 15347 35649
rect 16025 35649 16037 35652
rect 16071 35680 16083 35683
rect 17954 35680 17960 35692
rect 16071 35652 17960 35680
rect 16071 35649 16083 35652
rect 16025 35643 16083 35649
rect 17954 35640 17960 35652
rect 18012 35640 18018 35692
rect 18325 35683 18383 35689
rect 18325 35649 18337 35683
rect 18371 35680 18383 35683
rect 18782 35680 18788 35692
rect 18371 35652 18788 35680
rect 18371 35649 18383 35652
rect 18325 35643 18383 35649
rect 18782 35640 18788 35652
rect 18840 35640 18846 35692
rect 18984 35680 19012 35788
rect 19613 35785 19625 35819
rect 19659 35816 19671 35819
rect 20898 35816 20904 35828
rect 19659 35788 20904 35816
rect 19659 35785 19671 35788
rect 19613 35779 19671 35785
rect 20898 35776 20904 35788
rect 20956 35776 20962 35828
rect 25225 35819 25283 35825
rect 25225 35785 25237 35819
rect 25271 35816 25283 35819
rect 25406 35816 25412 35828
rect 25271 35788 25412 35816
rect 25271 35785 25283 35788
rect 25225 35779 25283 35785
rect 25406 35776 25412 35788
rect 25464 35776 25470 35828
rect 25498 35776 25504 35828
rect 25556 35816 25562 35828
rect 57882 35816 57888 35828
rect 25556 35788 57888 35816
rect 25556 35776 25562 35788
rect 57882 35776 57888 35788
rect 57940 35776 57946 35828
rect 70486 35776 70492 35828
rect 70544 35816 70550 35828
rect 71038 35816 71044 35828
rect 70544 35788 71044 35816
rect 70544 35776 70550 35788
rect 71038 35776 71044 35788
rect 71096 35816 71102 35828
rect 71409 35819 71467 35825
rect 71409 35816 71421 35819
rect 71096 35788 71421 35816
rect 71096 35776 71102 35788
rect 71409 35785 71421 35788
rect 71455 35785 71467 35819
rect 71409 35779 71467 35785
rect 73062 35776 73068 35828
rect 73120 35816 73126 35828
rect 74261 35819 74319 35825
rect 74261 35816 74273 35819
rect 73120 35788 74273 35816
rect 73120 35776 73126 35788
rect 74261 35785 74273 35788
rect 74307 35816 74319 35819
rect 77662 35816 77668 35828
rect 74307 35788 77668 35816
rect 74307 35785 74319 35788
rect 74261 35779 74319 35785
rect 77662 35776 77668 35788
rect 77720 35776 77726 35828
rect 77938 35825 77944 35828
rect 77922 35819 77944 35825
rect 77922 35785 77934 35819
rect 77922 35779 77944 35785
rect 77938 35776 77944 35779
rect 77996 35776 78002 35828
rect 78033 35819 78091 35825
rect 78033 35785 78045 35819
rect 78079 35816 78091 35819
rect 79597 35819 79655 35825
rect 79597 35816 79609 35819
rect 78079 35788 79609 35816
rect 78079 35785 78091 35788
rect 78033 35779 78091 35785
rect 79597 35785 79609 35788
rect 79643 35785 79655 35819
rect 79597 35779 79655 35785
rect 79778 35776 79784 35828
rect 79836 35816 79842 35828
rect 80057 35819 80115 35825
rect 80057 35816 80069 35819
rect 79836 35788 80069 35816
rect 79836 35776 79842 35788
rect 80057 35785 80069 35788
rect 80103 35785 80115 35819
rect 80057 35779 80115 35785
rect 86037 35819 86095 35825
rect 86037 35785 86049 35819
rect 86083 35816 86095 35819
rect 86862 35816 86868 35828
rect 86083 35788 86868 35816
rect 86083 35785 86095 35788
rect 86037 35779 86095 35785
rect 86862 35776 86868 35788
rect 86920 35776 86926 35828
rect 94133 35819 94191 35825
rect 94133 35785 94145 35819
rect 94179 35816 94191 35819
rect 96709 35819 96767 35825
rect 96709 35816 96721 35819
rect 94179 35788 96721 35816
rect 94179 35785 94191 35788
rect 94133 35779 94191 35785
rect 96709 35785 96721 35788
rect 96755 35785 96767 35819
rect 96709 35779 96767 35785
rect 20714 35748 20720 35760
rect 20675 35720 20720 35748
rect 20714 35708 20720 35720
rect 20772 35708 20778 35760
rect 25130 35708 25136 35760
rect 25188 35748 25194 35760
rect 30282 35748 30288 35760
rect 25188 35720 30288 35748
rect 25188 35708 25194 35720
rect 30282 35708 30288 35720
rect 30340 35708 30346 35760
rect 32122 35708 32128 35760
rect 32180 35748 32186 35760
rect 32766 35748 32772 35760
rect 32180 35720 32772 35748
rect 32180 35708 32186 35720
rect 32766 35708 32772 35720
rect 32824 35748 32830 35760
rect 42794 35748 42800 35760
rect 32824 35720 42800 35748
rect 32824 35708 32830 35720
rect 42794 35708 42800 35720
rect 42852 35708 42858 35760
rect 42886 35708 42892 35760
rect 42944 35708 42950 35760
rect 44450 35748 44456 35760
rect 44411 35720 44456 35748
rect 44450 35708 44456 35720
rect 44508 35708 44514 35760
rect 49786 35748 49792 35760
rect 44560 35720 49792 35748
rect 24118 35680 24124 35692
rect 18984 35652 24124 35680
rect 24118 35640 24124 35652
rect 24176 35640 24182 35692
rect 26881 35683 26939 35689
rect 26881 35649 26893 35683
rect 26927 35649 26939 35683
rect 26881 35643 26939 35649
rect 12989 35615 13047 35621
rect 12989 35612 13001 35615
rect 11480 35584 13001 35612
rect 11480 35572 11486 35584
rect 12989 35581 13001 35584
rect 13035 35581 13047 35615
rect 12989 35575 13047 35581
rect 13173 35615 13231 35621
rect 13173 35581 13185 35615
rect 13219 35581 13231 35615
rect 13173 35575 13231 35581
rect 13541 35615 13599 35621
rect 13541 35581 13553 35615
rect 13587 35581 13599 35615
rect 13541 35575 13599 35581
rect 9640 35516 11192 35544
rect 9640 35504 9646 35516
rect 5261 35479 5319 35485
rect 5261 35445 5273 35479
rect 5307 35445 5319 35479
rect 10870 35476 10876 35488
rect 10831 35448 10876 35476
rect 5261 35439 5319 35445
rect 10870 35436 10876 35448
rect 10928 35436 10934 35488
rect 11164 35485 11192 35516
rect 11149 35479 11207 35485
rect 11149 35445 11161 35479
rect 11195 35445 11207 35479
rect 13188 35476 13216 35575
rect 13630 35572 13636 35624
rect 13688 35612 13694 35624
rect 15194 35612 15200 35624
rect 13688 35584 13733 35612
rect 15155 35584 15200 35612
rect 13688 35572 13694 35584
rect 15194 35572 15200 35584
rect 15252 35572 15258 35624
rect 15562 35612 15568 35624
rect 15523 35584 15568 35612
rect 15562 35572 15568 35584
rect 15620 35572 15626 35624
rect 15749 35615 15807 35621
rect 15749 35581 15761 35615
rect 15795 35612 15807 35615
rect 15841 35615 15899 35621
rect 15841 35612 15853 35615
rect 15795 35584 15853 35612
rect 15795 35581 15807 35584
rect 15749 35575 15807 35581
rect 15841 35581 15853 35584
rect 15887 35581 15899 35615
rect 15841 35575 15899 35581
rect 18049 35615 18107 35621
rect 18049 35581 18061 35615
rect 18095 35612 18107 35615
rect 19058 35612 19064 35624
rect 18095 35584 19064 35612
rect 18095 35581 18107 35584
rect 18049 35575 18107 35581
rect 13446 35504 13452 35556
rect 13504 35544 13510 35556
rect 14553 35547 14611 35553
rect 14553 35544 14565 35547
rect 13504 35516 14565 35544
rect 13504 35504 13510 35516
rect 14553 35513 14565 35516
rect 14599 35513 14611 35547
rect 14553 35507 14611 35513
rect 13814 35476 13820 35488
rect 13188 35448 13820 35476
rect 11149 35439 11207 35445
rect 13814 35436 13820 35448
rect 13872 35436 13878 35488
rect 13998 35476 14004 35488
rect 13959 35448 14004 35476
rect 13998 35436 14004 35448
rect 14056 35436 14062 35488
rect 15856 35476 15884 35575
rect 19058 35572 19064 35584
rect 19116 35612 19122 35624
rect 19978 35612 19984 35624
rect 19116 35584 19984 35612
rect 19116 35572 19122 35584
rect 19978 35572 19984 35584
rect 20036 35572 20042 35624
rect 20622 35612 20628 35624
rect 20583 35584 20628 35612
rect 20622 35572 20628 35584
rect 20680 35572 20686 35624
rect 25041 35615 25099 35621
rect 25041 35581 25053 35615
rect 25087 35612 25099 35615
rect 25130 35612 25136 35624
rect 25087 35584 25136 35612
rect 25087 35581 25099 35584
rect 25041 35575 25099 35581
rect 19150 35504 19156 35556
rect 19208 35544 19214 35556
rect 24857 35547 24915 35553
rect 24857 35544 24869 35547
rect 19208 35516 24869 35544
rect 19208 35504 19214 35516
rect 24857 35513 24869 35516
rect 24903 35544 24915 35547
rect 25056 35544 25084 35575
rect 25130 35572 25136 35584
rect 25188 35572 25194 35624
rect 26786 35612 26792 35624
rect 25792 35584 26792 35612
rect 24903 35516 25084 35544
rect 24903 35513 24915 35516
rect 24857 35507 24915 35513
rect 19426 35476 19432 35488
rect 15856 35448 19432 35476
rect 19426 35436 19432 35448
rect 19484 35436 19490 35488
rect 19889 35479 19947 35485
rect 19889 35445 19901 35479
rect 19935 35476 19947 35479
rect 19978 35476 19984 35488
rect 19935 35448 19984 35476
rect 19935 35445 19947 35448
rect 19889 35439 19947 35445
rect 19978 35436 19984 35448
rect 20036 35476 20042 35488
rect 21818 35476 21824 35488
rect 20036 35448 21824 35476
rect 20036 35436 20042 35448
rect 21818 35436 21824 35448
rect 21876 35436 21882 35488
rect 25038 35436 25044 35488
rect 25096 35476 25102 35488
rect 25792 35476 25820 35584
rect 26786 35572 26792 35584
rect 26844 35572 26850 35624
rect 26896 35544 26924 35643
rect 26970 35640 26976 35692
rect 27028 35680 27034 35692
rect 30558 35680 30564 35692
rect 27028 35652 30420 35680
rect 30519 35652 30564 35680
rect 27028 35640 27034 35652
rect 27154 35612 27160 35624
rect 27115 35584 27160 35612
rect 27154 35572 27160 35584
rect 27212 35572 27218 35624
rect 27341 35615 27399 35621
rect 27341 35581 27353 35615
rect 27387 35612 27399 35615
rect 28902 35612 28908 35624
rect 27387 35584 28908 35612
rect 27387 35581 27399 35584
rect 27341 35575 27399 35581
rect 28902 35572 28908 35584
rect 28960 35572 28966 35624
rect 29086 35572 29092 35624
rect 29144 35612 29150 35624
rect 30285 35615 30343 35621
rect 30285 35612 30297 35615
rect 29144 35584 30297 35612
rect 29144 35572 29150 35584
rect 30285 35581 30297 35584
rect 30331 35581 30343 35615
rect 30392 35612 30420 35652
rect 30558 35640 30564 35652
rect 30616 35640 30622 35692
rect 35342 35680 35348 35692
rect 35303 35652 35348 35680
rect 35342 35640 35348 35652
rect 35400 35640 35406 35692
rect 36633 35683 36691 35689
rect 35544 35652 35756 35680
rect 30392 35584 31248 35612
rect 30285 35575 30343 35581
rect 30098 35544 30104 35556
rect 26896 35516 30104 35544
rect 30098 35504 30104 35516
rect 30156 35504 30162 35556
rect 25096 35448 25820 35476
rect 26421 35479 26479 35485
rect 25096 35436 25102 35448
rect 26421 35445 26433 35479
rect 26467 35476 26479 35479
rect 26510 35476 26516 35488
rect 26467 35448 26516 35476
rect 26467 35445 26479 35448
rect 26421 35439 26479 35445
rect 26510 35436 26516 35448
rect 26568 35436 26574 35488
rect 26602 35436 26608 35488
rect 26660 35476 26666 35488
rect 30190 35476 30196 35488
rect 26660 35448 30196 35476
rect 26660 35436 26666 35448
rect 30190 35436 30196 35448
rect 30248 35436 30254 35488
rect 30300 35476 30328 35575
rect 31220 35544 31248 35584
rect 31294 35572 31300 35624
rect 31352 35612 31358 35624
rect 35544 35621 35572 35652
rect 35529 35615 35587 35621
rect 35529 35612 35541 35615
rect 31352 35584 35541 35612
rect 31352 35572 31358 35584
rect 35529 35581 35541 35584
rect 35575 35581 35587 35615
rect 35728 35612 35756 35652
rect 36633 35649 36645 35683
rect 36679 35680 36691 35683
rect 42610 35680 42616 35692
rect 36679 35652 42616 35680
rect 36679 35649 36691 35652
rect 36633 35643 36691 35649
rect 42610 35640 42616 35652
rect 42668 35640 42674 35692
rect 42904 35680 42932 35708
rect 43165 35683 43223 35689
rect 43165 35680 43177 35683
rect 42904 35652 43177 35680
rect 43165 35649 43177 35652
rect 43211 35649 43223 35683
rect 43165 35643 43223 35649
rect 44082 35640 44088 35692
rect 44140 35680 44146 35692
rect 44560 35680 44588 35720
rect 49786 35708 49792 35720
rect 49844 35708 49850 35760
rect 51350 35708 51356 35760
rect 51408 35748 51414 35760
rect 51997 35751 52055 35757
rect 51997 35748 52009 35751
rect 51408 35720 52009 35748
rect 51408 35708 51414 35720
rect 51997 35717 52009 35720
rect 52043 35717 52055 35751
rect 51997 35711 52055 35717
rect 54570 35708 54576 35760
rect 54628 35748 54634 35760
rect 54628 35720 55076 35748
rect 54628 35708 54634 35720
rect 44140 35652 44588 35680
rect 44140 35640 44146 35652
rect 48774 35640 48780 35692
rect 48832 35680 48838 35692
rect 50433 35683 50491 35689
rect 48832 35652 49556 35680
rect 48832 35640 48838 35652
rect 36081 35615 36139 35621
rect 36081 35612 36093 35615
rect 35728 35584 36093 35612
rect 35529 35575 35587 35581
rect 36081 35581 36093 35584
rect 36127 35612 36139 35615
rect 36170 35612 36176 35624
rect 36127 35584 36176 35612
rect 36127 35581 36139 35584
rect 36081 35575 36139 35581
rect 36170 35572 36176 35584
rect 36228 35572 36234 35624
rect 36265 35615 36323 35621
rect 36265 35581 36277 35615
rect 36311 35581 36323 35615
rect 36265 35575 36323 35581
rect 36280 35544 36308 35575
rect 36446 35572 36452 35624
rect 36504 35612 36510 35624
rect 39666 35612 39672 35624
rect 36504 35584 39672 35612
rect 36504 35572 36510 35584
rect 39666 35572 39672 35584
rect 39724 35572 39730 35624
rect 42794 35572 42800 35624
rect 42852 35612 42858 35624
rect 42889 35615 42947 35621
rect 42889 35612 42901 35615
rect 42852 35584 42901 35612
rect 42852 35572 42858 35584
rect 42889 35581 42901 35584
rect 42935 35581 42947 35615
rect 49145 35615 49203 35621
rect 49145 35612 49157 35615
rect 42889 35575 42947 35581
rect 42996 35584 43852 35612
rect 36909 35547 36967 35553
rect 36909 35544 36921 35547
rect 31220 35516 36921 35544
rect 36909 35513 36921 35516
rect 36955 35544 36967 35547
rect 41230 35544 41236 35556
rect 36955 35516 41236 35544
rect 36955 35513 36967 35516
rect 36909 35507 36967 35513
rect 41230 35504 41236 35516
rect 41288 35504 41294 35556
rect 42058 35504 42064 35556
rect 42116 35544 42122 35556
rect 42996 35544 43024 35584
rect 42116 35516 43024 35544
rect 43824 35544 43852 35584
rect 48976 35584 49157 35612
rect 48866 35544 48872 35556
rect 43824 35516 48872 35544
rect 42116 35504 42122 35516
rect 48866 35504 48872 35516
rect 48924 35504 48930 35556
rect 48976 35488 49004 35584
rect 49145 35581 49157 35584
rect 49191 35612 49203 35615
rect 49234 35612 49240 35624
rect 49191 35584 49240 35612
rect 49191 35581 49203 35584
rect 49145 35575 49203 35581
rect 49234 35572 49240 35584
rect 49292 35572 49298 35624
rect 49329 35615 49387 35621
rect 49329 35581 49341 35615
rect 49375 35581 49387 35615
rect 49528 35612 49556 35652
rect 50433 35649 50445 35683
rect 50479 35680 50491 35683
rect 51868 35683 51926 35689
rect 51868 35680 51880 35683
rect 50479 35652 51880 35680
rect 50479 35649 50491 35652
rect 50433 35643 50491 35649
rect 51868 35649 51880 35652
rect 51914 35649 51926 35683
rect 51868 35643 51926 35649
rect 52089 35683 52147 35689
rect 52089 35649 52101 35683
rect 52135 35680 52147 35683
rect 54938 35680 54944 35692
rect 52135 35652 54944 35680
rect 52135 35649 52147 35652
rect 52089 35643 52147 35649
rect 54938 35640 54944 35652
rect 54996 35640 55002 35692
rect 55048 35689 55076 35720
rect 55122 35708 55128 35760
rect 55180 35748 55186 35760
rect 56137 35751 56195 35757
rect 56137 35748 56149 35751
rect 55180 35720 56149 35748
rect 55180 35708 55186 35720
rect 56137 35717 56149 35720
rect 56183 35717 56195 35751
rect 57514 35748 57520 35760
rect 56137 35711 56195 35717
rect 56704 35720 57520 35748
rect 55033 35683 55091 35689
rect 55033 35649 55045 35683
rect 55079 35649 55091 35683
rect 55033 35643 55091 35649
rect 56594 35640 56600 35692
rect 56652 35680 56658 35692
rect 56704 35689 56732 35720
rect 57514 35708 57520 35720
rect 57572 35748 57578 35760
rect 63313 35751 63371 35757
rect 57572 35720 59124 35748
rect 57572 35708 57578 35720
rect 56689 35683 56747 35689
rect 56689 35680 56701 35683
rect 56652 35652 56701 35680
rect 56652 35640 56658 35652
rect 56689 35649 56701 35652
rect 56735 35649 56747 35683
rect 56962 35680 56968 35692
rect 56923 35652 56968 35680
rect 56689 35643 56747 35649
rect 56962 35640 56968 35652
rect 57020 35680 57026 35692
rect 58618 35680 58624 35692
rect 57020 35652 57652 35680
rect 58579 35652 58624 35680
rect 57020 35640 57026 35652
rect 49789 35615 49847 35621
rect 49789 35612 49801 35615
rect 49528 35584 49801 35612
rect 49329 35575 49387 35581
rect 49789 35581 49801 35584
rect 49835 35581 49847 35615
rect 49789 35575 49847 35581
rect 49881 35615 49939 35621
rect 49881 35581 49893 35615
rect 49927 35612 49939 35615
rect 49970 35612 49976 35624
rect 49927 35584 49976 35612
rect 49927 35581 49939 35584
rect 49881 35575 49939 35581
rect 49344 35544 49372 35575
rect 49970 35572 49976 35584
rect 50028 35612 50034 35624
rect 50706 35612 50712 35624
rect 50028 35584 50712 35612
rect 50028 35572 50034 35584
rect 50706 35572 50712 35584
rect 50764 35572 50770 35624
rect 55214 35572 55220 35624
rect 55272 35612 55278 35624
rect 55677 35615 55735 35621
rect 55272 35584 55317 35612
rect 55272 35572 55278 35584
rect 55677 35581 55689 35615
rect 55723 35581 55735 35615
rect 55677 35575 55735 35581
rect 50890 35544 50896 35556
rect 49344 35516 50896 35544
rect 50890 35504 50896 35516
rect 50948 35504 50954 35556
rect 51718 35504 51724 35556
rect 51776 35544 51782 35556
rect 51776 35516 51820 35544
rect 51776 35504 51782 35516
rect 54478 35504 54484 35556
rect 54536 35544 54542 35556
rect 54849 35547 54907 35553
rect 54849 35544 54861 35547
rect 54536 35516 54861 35544
rect 54536 35504 54542 35516
rect 54849 35513 54861 35516
rect 54895 35544 54907 35547
rect 55692 35544 55720 35575
rect 55766 35572 55772 35624
rect 55824 35612 55830 35624
rect 57333 35615 57391 35621
rect 57333 35612 57345 35615
rect 55824 35584 55869 35612
rect 56060 35584 57345 35612
rect 55824 35572 55830 35584
rect 54895 35516 55720 35544
rect 54895 35513 54907 35516
rect 54849 35507 54907 35513
rect 31754 35476 31760 35488
rect 30300 35448 31760 35476
rect 31754 35436 31760 35448
rect 31812 35436 31818 35488
rect 31849 35479 31907 35485
rect 31849 35445 31861 35479
rect 31895 35476 31907 35479
rect 31938 35476 31944 35488
rect 31895 35448 31944 35476
rect 31895 35445 31907 35448
rect 31849 35439 31907 35445
rect 31938 35436 31944 35448
rect 31996 35436 32002 35488
rect 34606 35436 34612 35488
rect 34664 35476 34670 35488
rect 35161 35479 35219 35485
rect 35161 35476 35173 35479
rect 34664 35448 35173 35476
rect 34664 35436 34670 35448
rect 35161 35445 35173 35448
rect 35207 35476 35219 35479
rect 35342 35476 35348 35488
rect 35207 35448 35348 35476
rect 35207 35445 35219 35448
rect 35161 35439 35219 35445
rect 35342 35436 35348 35448
rect 35400 35436 35406 35488
rect 36262 35436 36268 35488
rect 36320 35476 36326 35488
rect 42978 35476 42984 35488
rect 36320 35448 42984 35476
rect 36320 35436 36326 35448
rect 42978 35436 42984 35448
rect 43036 35436 43042 35488
rect 48774 35476 48780 35488
rect 48735 35448 48780 35476
rect 48774 35436 48780 35448
rect 48832 35436 48838 35488
rect 48958 35476 48964 35488
rect 48919 35448 48964 35476
rect 48958 35436 48964 35448
rect 49016 35436 49022 35488
rect 50706 35476 50712 35488
rect 50619 35448 50712 35476
rect 50706 35436 50712 35448
rect 50764 35476 50770 35488
rect 51166 35476 51172 35488
rect 50764 35448 51172 35476
rect 50764 35436 50770 35448
rect 51166 35436 51172 35448
rect 51224 35476 51230 35488
rect 51994 35476 52000 35488
rect 51224 35448 52000 35476
rect 51224 35436 51230 35448
rect 51994 35436 52000 35448
rect 52052 35436 52058 35488
rect 52362 35476 52368 35488
rect 52323 35448 52368 35476
rect 52362 35436 52368 35448
rect 52420 35436 52426 35488
rect 54570 35436 54576 35488
rect 54628 35476 54634 35488
rect 54665 35479 54723 35485
rect 54665 35476 54677 35479
rect 54628 35448 54677 35476
rect 54628 35436 54634 35448
rect 54665 35445 54677 35448
rect 54711 35445 54723 35479
rect 55692 35476 55720 35516
rect 56060 35476 56088 35584
rect 57333 35581 57345 35584
rect 57379 35581 57391 35615
rect 57514 35612 57520 35624
rect 57475 35584 57520 35612
rect 57333 35575 57391 35581
rect 57514 35572 57520 35584
rect 57572 35572 57578 35624
rect 57624 35612 57652 35652
rect 58618 35640 58624 35652
rect 58676 35640 58682 35692
rect 59096 35624 59124 35720
rect 63313 35717 63325 35751
rect 63359 35748 63371 35751
rect 63494 35748 63500 35760
rect 63359 35720 63500 35748
rect 63359 35717 63371 35720
rect 63313 35711 63371 35717
rect 63494 35708 63500 35720
rect 63552 35708 63558 35760
rect 63678 35748 63684 35760
rect 63639 35720 63684 35748
rect 63678 35708 63684 35720
rect 63736 35708 63742 35760
rect 67453 35751 67511 35757
rect 64156 35720 67404 35748
rect 64156 35689 64184 35720
rect 64141 35683 64199 35689
rect 64141 35649 64153 35683
rect 64187 35649 64199 35683
rect 64141 35643 64199 35649
rect 66254 35640 66260 35692
rect 66312 35680 66318 35692
rect 67376 35680 67404 35720
rect 67453 35717 67465 35751
rect 67499 35748 67511 35751
rect 68738 35748 68744 35760
rect 67499 35720 68744 35748
rect 67499 35717 67511 35720
rect 67453 35711 67511 35717
rect 68738 35708 68744 35720
rect 68796 35708 68802 35760
rect 76101 35751 76159 35757
rect 76101 35717 76113 35751
rect 76147 35748 76159 35751
rect 77570 35748 77576 35760
rect 76147 35720 77576 35748
rect 76147 35717 76159 35720
rect 76101 35711 76159 35717
rect 77570 35708 77576 35720
rect 77628 35708 77634 35760
rect 78401 35751 78459 35757
rect 78401 35717 78413 35751
rect 78447 35748 78459 35751
rect 84470 35748 84476 35760
rect 78447 35720 84476 35748
rect 78447 35717 78459 35720
rect 78401 35711 78459 35717
rect 84470 35708 84476 35720
rect 84528 35708 84534 35760
rect 85669 35751 85727 35757
rect 85669 35748 85681 35751
rect 84948 35720 85681 35748
rect 70210 35680 70216 35692
rect 66312 35652 66357 35680
rect 67376 35652 70216 35680
rect 66312 35640 66318 35652
rect 57977 35615 58035 35621
rect 57977 35612 57989 35615
rect 57624 35584 57989 35612
rect 57977 35581 57989 35584
rect 58023 35581 58035 35615
rect 57977 35575 58035 35581
rect 58069 35615 58127 35621
rect 58069 35581 58081 35615
rect 58115 35612 58127 35615
rect 59078 35612 59084 35624
rect 58115 35584 58940 35612
rect 59039 35584 59084 35612
rect 58115 35581 58127 35584
rect 58069 35575 58127 35581
rect 56134 35504 56140 35556
rect 56192 35544 56198 35556
rect 58084 35544 58112 35575
rect 56192 35516 58112 35544
rect 56192 35504 56198 35516
rect 58912 35488 58940 35584
rect 59078 35572 59084 35584
rect 59136 35572 59142 35624
rect 63129 35615 63187 35621
rect 63129 35581 63141 35615
rect 63175 35612 63187 35615
rect 63310 35612 63316 35624
rect 63175 35584 63316 35612
rect 63175 35581 63187 35584
rect 63129 35575 63187 35581
rect 63310 35572 63316 35584
rect 63368 35612 63374 35624
rect 64049 35615 64107 35621
rect 64049 35612 64061 35615
rect 63368 35584 64061 35612
rect 63368 35572 63374 35584
rect 64049 35581 64061 35584
rect 64095 35581 64107 35615
rect 64414 35612 64420 35624
rect 64375 35584 64420 35612
rect 64049 35575 64107 35581
rect 64414 35572 64420 35584
rect 64472 35572 64478 35624
rect 64598 35612 64604 35624
rect 64559 35584 64604 35612
rect 64598 35572 64604 35584
rect 64656 35572 64662 35624
rect 66441 35615 66499 35621
rect 66441 35612 66453 35615
rect 65904 35584 66453 35612
rect 56505 35479 56563 35485
rect 56505 35476 56517 35479
rect 55692 35448 56517 35476
rect 54665 35439 54723 35445
rect 56505 35445 56517 35448
rect 56551 35445 56563 35479
rect 58894 35476 58900 35488
rect 58855 35448 58900 35476
rect 56505 35439 56563 35445
rect 58894 35436 58900 35448
rect 58952 35436 58958 35488
rect 62022 35436 62028 35488
rect 62080 35476 62086 35488
rect 65904 35485 65932 35584
rect 66441 35581 66453 35584
rect 66487 35612 66499 35615
rect 66993 35615 67051 35621
rect 66993 35612 67005 35615
rect 66487 35584 67005 35612
rect 66487 35581 66499 35584
rect 66441 35575 66499 35581
rect 66993 35581 67005 35584
rect 67039 35581 67051 35615
rect 66993 35575 67051 35581
rect 67177 35615 67235 35621
rect 67177 35581 67189 35615
rect 67223 35612 67235 35615
rect 67376 35612 67404 35652
rect 70210 35640 70216 35652
rect 70268 35640 70274 35692
rect 77478 35640 77484 35692
rect 77536 35680 77542 35692
rect 77536 35652 77708 35680
rect 77536 35640 77542 35652
rect 67223 35584 67404 35612
rect 67223 35581 67235 35584
rect 67177 35575 67235 35581
rect 68554 35572 68560 35624
rect 68612 35612 68618 35624
rect 69106 35621 69112 35624
rect 68833 35615 68891 35621
rect 68833 35612 68845 35615
rect 68612 35584 68845 35612
rect 68612 35572 68618 35584
rect 68833 35581 68845 35584
rect 68879 35581 68891 35615
rect 68833 35575 68891 35581
rect 69103 35575 69112 35621
rect 69164 35612 69170 35624
rect 70489 35615 70547 35621
rect 69164 35584 69203 35612
rect 69106 35572 69112 35575
rect 69164 35572 69170 35584
rect 70489 35581 70501 35615
rect 70535 35612 70547 35615
rect 71317 35615 71375 35621
rect 71317 35612 71329 35615
rect 70535 35584 71329 35612
rect 70535 35581 70547 35584
rect 70489 35575 70547 35581
rect 71317 35581 71329 35584
rect 71363 35612 71375 35615
rect 71406 35612 71412 35624
rect 71363 35584 71412 35612
rect 71363 35581 71375 35584
rect 71317 35575 71375 35581
rect 71406 35572 71412 35584
rect 71464 35572 71470 35624
rect 74169 35615 74227 35621
rect 74169 35581 74181 35615
rect 74215 35612 74227 35615
rect 74258 35612 74264 35624
rect 74215 35584 74264 35612
rect 74215 35581 74227 35584
rect 74169 35575 74227 35581
rect 74258 35572 74264 35584
rect 74316 35612 74322 35624
rect 74445 35615 74503 35621
rect 74445 35612 74457 35615
rect 74316 35584 74457 35612
rect 74316 35572 74322 35584
rect 74445 35581 74457 35584
rect 74491 35581 74503 35615
rect 74445 35575 74503 35581
rect 75914 35572 75920 35624
rect 75972 35612 75978 35624
rect 76193 35615 76251 35621
rect 76193 35612 76205 35615
rect 75972 35584 76205 35612
rect 75972 35572 75978 35584
rect 76193 35581 76205 35584
rect 76239 35581 76251 35615
rect 76193 35575 76251 35581
rect 76282 35572 76288 35624
rect 76340 35612 76346 35624
rect 76469 35615 76527 35621
rect 76469 35612 76481 35615
rect 76340 35584 76481 35612
rect 76340 35572 76346 35584
rect 76469 35581 76481 35584
rect 76515 35581 76527 35615
rect 76469 35575 76527 35581
rect 76650 35572 76656 35624
rect 76708 35612 76714 35624
rect 77386 35612 77392 35624
rect 76708 35584 77392 35612
rect 76708 35572 76714 35584
rect 77386 35572 77392 35584
rect 77444 35572 77450 35624
rect 77680 35612 77708 35652
rect 77757 35615 77815 35621
rect 77757 35612 77769 35615
rect 77680 35584 77769 35612
rect 77757 35581 77769 35584
rect 77803 35581 77815 35615
rect 77757 35575 77815 35581
rect 77938 35572 77944 35624
rect 77996 35612 78002 35624
rect 78096 35615 78154 35621
rect 78096 35612 78108 35615
rect 77996 35584 78108 35612
rect 77996 35572 78002 35584
rect 78096 35581 78108 35584
rect 78142 35612 78154 35615
rect 79965 35615 80023 35621
rect 79965 35612 79977 35615
rect 78142 35584 79977 35612
rect 78142 35581 78154 35584
rect 78096 35575 78154 35581
rect 79965 35581 79977 35584
rect 80011 35612 80023 35615
rect 80425 35615 80483 35621
rect 80425 35612 80437 35615
rect 80011 35584 80437 35612
rect 80011 35581 80023 35584
rect 79965 35575 80023 35581
rect 80425 35581 80437 35584
rect 80471 35581 80483 35615
rect 83734 35612 83740 35624
rect 83695 35584 83740 35612
rect 80425 35575 80483 35581
rect 83734 35572 83740 35584
rect 83792 35612 83798 35624
rect 84105 35615 84163 35621
rect 84105 35612 84117 35615
rect 83792 35584 84117 35612
rect 83792 35572 83798 35584
rect 84105 35581 84117 35584
rect 84151 35612 84163 35615
rect 84948 35612 84976 35720
rect 85669 35717 85681 35720
rect 85715 35717 85727 35751
rect 85669 35711 85727 35717
rect 85540 35683 85598 35689
rect 85540 35649 85552 35683
rect 85586 35680 85598 35683
rect 85586 35649 85620 35680
rect 85540 35643 85620 35649
rect 84151 35584 84976 35612
rect 84151 35581 84163 35584
rect 84105 35575 84163 35581
rect 65978 35504 65984 35556
rect 66036 35544 66042 35556
rect 68646 35544 68652 35556
rect 66036 35516 68652 35544
rect 66036 35504 66042 35516
rect 68646 35504 68652 35516
rect 68704 35504 68710 35556
rect 76101 35547 76159 35553
rect 69768 35516 70808 35544
rect 65705 35479 65763 35485
rect 65705 35476 65717 35479
rect 62080 35448 65717 35476
rect 62080 35436 62086 35448
rect 65705 35445 65717 35448
rect 65751 35476 65763 35479
rect 65889 35479 65947 35485
rect 65889 35476 65901 35479
rect 65751 35448 65901 35476
rect 65751 35445 65763 35448
rect 65705 35439 65763 35445
rect 65889 35445 65901 35448
rect 65935 35445 65947 35479
rect 66070 35476 66076 35488
rect 66031 35448 66076 35476
rect 65889 35439 65947 35445
rect 66070 35436 66076 35448
rect 66128 35436 66134 35488
rect 66162 35436 66168 35488
rect 66220 35476 66226 35488
rect 69768 35476 69796 35516
rect 66220 35448 69796 35476
rect 66220 35436 66226 35448
rect 69842 35436 69848 35488
rect 69900 35476 69906 35488
rect 70486 35476 70492 35488
rect 69900 35448 70492 35476
rect 69900 35436 69906 35448
rect 70486 35436 70492 35448
rect 70544 35436 70550 35488
rect 70578 35436 70584 35488
rect 70636 35476 70642 35488
rect 70780 35476 70808 35516
rect 76101 35513 76113 35547
rect 76147 35544 76159 35547
rect 76377 35547 76435 35553
rect 76377 35544 76389 35547
rect 76147 35516 76389 35544
rect 76147 35513 76159 35516
rect 76101 35507 76159 35513
rect 76377 35513 76389 35516
rect 76423 35513 76435 35547
rect 76377 35507 76435 35513
rect 76558 35504 76564 35556
rect 76616 35544 76622 35556
rect 76929 35547 76987 35553
rect 76929 35544 76941 35547
rect 76616 35516 76941 35544
rect 76616 35504 76622 35516
rect 76929 35513 76941 35516
rect 76975 35513 76987 35547
rect 77662 35544 77668 35556
rect 77623 35516 77668 35544
rect 76929 35507 76987 35513
rect 77662 35504 77668 35516
rect 77720 35504 77726 35556
rect 78677 35547 78735 35553
rect 78677 35513 78689 35547
rect 78723 35544 78735 35547
rect 78766 35544 78772 35556
rect 78723 35516 78772 35544
rect 78723 35513 78735 35516
rect 78677 35507 78735 35513
rect 78766 35504 78772 35516
rect 78824 35504 78830 35556
rect 79597 35547 79655 35553
rect 79597 35513 79609 35547
rect 79643 35544 79655 35547
rect 79778 35544 79784 35556
rect 79643 35516 79784 35544
rect 79643 35513 79655 35516
rect 79597 35507 79655 35513
rect 79778 35504 79784 35516
rect 79836 35504 79842 35556
rect 85390 35544 85396 35556
rect 85351 35516 85396 35544
rect 85390 35504 85396 35516
rect 85448 35504 85454 35556
rect 85592 35544 85620 35643
rect 85684 35612 85712 35711
rect 85850 35708 85856 35760
rect 85908 35748 85914 35760
rect 93857 35751 93915 35757
rect 93857 35748 93869 35751
rect 85908 35720 93869 35748
rect 85908 35708 85914 35720
rect 93857 35717 93869 35720
rect 93903 35748 93915 35751
rect 94038 35748 94044 35760
rect 93903 35720 94044 35748
rect 93903 35717 93915 35720
rect 93857 35711 93915 35717
rect 94038 35708 94044 35720
rect 94096 35708 94102 35760
rect 85758 35640 85764 35692
rect 85816 35680 85822 35692
rect 86405 35683 86463 35689
rect 86405 35680 86417 35683
rect 85816 35652 86417 35680
rect 85816 35640 85822 35652
rect 86405 35649 86417 35652
rect 86451 35649 86463 35683
rect 88426 35680 88432 35692
rect 88387 35652 88432 35680
rect 86405 35643 86463 35649
rect 88426 35640 88432 35652
rect 88484 35640 88490 35692
rect 89180 35652 89668 35680
rect 86221 35615 86279 35621
rect 86221 35612 86233 35615
rect 85684 35584 86233 35612
rect 86221 35581 86233 35584
rect 86267 35612 86279 35615
rect 86770 35612 86776 35624
rect 86267 35584 86776 35612
rect 86267 35581 86279 35584
rect 86221 35575 86279 35581
rect 86770 35572 86776 35584
rect 86828 35572 86834 35624
rect 88150 35612 88156 35624
rect 87708 35584 88156 35612
rect 87708 35544 87736 35584
rect 88150 35572 88156 35584
rect 88208 35572 88214 35624
rect 88242 35572 88248 35624
rect 88300 35572 88306 35624
rect 85592 35516 87736 35544
rect 87969 35547 88027 35553
rect 87969 35513 87981 35547
rect 88015 35544 88027 35547
rect 88260 35544 88288 35572
rect 88015 35516 88288 35544
rect 88015 35513 88027 35516
rect 87969 35507 88027 35513
rect 79502 35476 79508 35488
rect 70636 35448 70681 35476
rect 70780 35448 79508 35476
rect 70636 35436 70642 35448
rect 79502 35436 79508 35448
rect 79560 35436 79566 35488
rect 80146 35436 80152 35488
rect 80204 35476 80210 35488
rect 83921 35479 83979 35485
rect 83921 35476 83933 35479
rect 80204 35448 83933 35476
rect 80204 35436 80210 35448
rect 83921 35445 83933 35448
rect 83967 35476 83979 35479
rect 84286 35476 84292 35488
rect 83967 35448 84292 35476
rect 83967 35445 83979 35448
rect 83921 35439 83979 35445
rect 84286 35436 84292 35448
rect 84344 35436 84350 35488
rect 88978 35436 88984 35488
rect 89036 35476 89042 35488
rect 89180 35485 89208 35652
rect 89533 35615 89591 35621
rect 89533 35581 89545 35615
rect 89579 35581 89591 35615
rect 89640 35612 89668 35652
rect 89714 35640 89720 35692
rect 89772 35680 89778 35692
rect 90726 35680 90732 35692
rect 89772 35652 89817 35680
rect 90687 35652 90732 35680
rect 89772 35640 89778 35652
rect 90726 35640 90732 35652
rect 90784 35680 90790 35692
rect 91005 35683 91063 35689
rect 91005 35680 91017 35683
rect 90784 35652 91017 35680
rect 90784 35640 90790 35652
rect 91005 35649 91017 35652
rect 91051 35649 91063 35683
rect 91005 35643 91063 35649
rect 89901 35615 89959 35621
rect 89640 35584 89760 35612
rect 89533 35575 89591 35581
rect 89165 35479 89223 35485
rect 89165 35476 89177 35479
rect 89036 35448 89177 35476
rect 89036 35436 89042 35448
rect 89165 35445 89177 35448
rect 89211 35445 89223 35479
rect 89548 35476 89576 35575
rect 89732 35544 89760 35584
rect 89901 35581 89913 35615
rect 89947 35581 89959 35615
rect 91278 35612 91284 35624
rect 91239 35584 91284 35612
rect 89901 35575 89959 35581
rect 89916 35544 89944 35575
rect 91278 35572 91284 35584
rect 91336 35572 91342 35624
rect 93670 35612 93676 35624
rect 93583 35584 93676 35612
rect 93670 35572 93676 35584
rect 93728 35612 93734 35624
rect 94148 35612 94176 35779
rect 95234 35680 95240 35692
rect 95195 35652 95240 35680
rect 95234 35640 95240 35652
rect 95292 35640 95298 35692
rect 94958 35612 94964 35624
rect 93728 35584 94176 35612
rect 94608 35584 94964 35612
rect 93728 35572 93734 35584
rect 89732 35516 89944 35544
rect 91189 35547 91247 35553
rect 91189 35513 91201 35547
rect 91235 35513 91247 35547
rect 91189 35507 91247 35513
rect 91741 35547 91799 35553
rect 91741 35513 91753 35547
rect 91787 35544 91799 35547
rect 94130 35544 94136 35556
rect 91787 35516 94136 35544
rect 91787 35513 91799 35516
rect 91741 35507 91799 35513
rect 91204 35476 91232 35507
rect 94130 35504 94136 35516
rect 94188 35504 94194 35556
rect 91278 35476 91284 35488
rect 89548 35448 91284 35476
rect 89165 35439 89223 35445
rect 91278 35436 91284 35448
rect 91336 35436 91342 35488
rect 94038 35436 94044 35488
rect 94096 35476 94102 35488
rect 94608 35485 94636 35584
rect 94958 35572 94964 35584
rect 95016 35572 95022 35624
rect 96617 35615 96675 35621
rect 96617 35581 96629 35615
rect 96663 35612 96675 35615
rect 96706 35612 96712 35624
rect 96663 35584 96712 35612
rect 96663 35581 96675 35584
rect 96617 35575 96675 35581
rect 96706 35572 96712 35584
rect 96764 35572 96770 35624
rect 94777 35547 94835 35553
rect 94777 35513 94789 35547
rect 94823 35544 94835 35547
rect 95050 35544 95056 35556
rect 94823 35516 95056 35544
rect 94823 35513 94835 35516
rect 94777 35507 94835 35513
rect 95050 35504 95056 35516
rect 95108 35504 95114 35556
rect 94593 35479 94651 35485
rect 94593 35476 94605 35479
rect 94096 35448 94605 35476
rect 94096 35436 94102 35448
rect 94593 35445 94605 35448
rect 94639 35445 94651 35479
rect 94593 35439 94651 35445
rect 1104 35386 105616 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 50326 35386
rect 50378 35334 50390 35386
rect 50442 35334 50454 35386
rect 50506 35334 50518 35386
rect 50570 35334 81046 35386
rect 81098 35334 81110 35386
rect 81162 35334 81174 35386
rect 81226 35334 81238 35386
rect 81290 35334 105616 35386
rect 1104 35312 105616 35334
rect 5810 35272 5816 35284
rect 5771 35244 5816 35272
rect 5810 35232 5816 35244
rect 5868 35232 5874 35284
rect 7374 35272 7380 35284
rect 7335 35244 7380 35272
rect 7374 35232 7380 35244
rect 7432 35232 7438 35284
rect 13906 35232 13912 35284
rect 13964 35272 13970 35284
rect 15010 35272 15016 35284
rect 13964 35244 15016 35272
rect 13964 35232 13970 35244
rect 15010 35232 15016 35244
rect 15068 35272 15074 35284
rect 19150 35272 19156 35284
rect 15068 35244 19156 35272
rect 15068 35232 15074 35244
rect 19150 35232 19156 35244
rect 19208 35232 19214 35284
rect 19334 35232 19340 35284
rect 19392 35272 19398 35284
rect 19429 35275 19487 35281
rect 19429 35272 19441 35275
rect 19392 35244 19441 35272
rect 19392 35232 19398 35244
rect 19429 35241 19441 35244
rect 19475 35241 19487 35275
rect 19429 35235 19487 35241
rect 19797 35275 19855 35281
rect 19797 35241 19809 35275
rect 19843 35272 19855 35275
rect 20714 35272 20720 35284
rect 19843 35244 20720 35272
rect 19843 35241 19855 35244
rect 19797 35235 19855 35241
rect 3878 35164 3884 35216
rect 3936 35204 3942 35216
rect 9950 35204 9956 35216
rect 3936 35176 9956 35204
rect 3936 35164 3942 35176
rect 9950 35164 9956 35176
rect 10008 35164 10014 35216
rect 12894 35204 12900 35216
rect 12855 35176 12900 35204
rect 12894 35164 12900 35176
rect 12952 35164 12958 35216
rect 13814 35204 13820 35216
rect 13556 35176 13820 35204
rect 5534 35096 5540 35148
rect 5592 35136 5598 35148
rect 5721 35139 5779 35145
rect 5721 35136 5733 35139
rect 5592 35108 5733 35136
rect 5592 35096 5598 35108
rect 5721 35105 5733 35108
rect 5767 35105 5779 35139
rect 6270 35136 6276 35148
rect 6231 35108 6276 35136
rect 5721 35099 5779 35105
rect 6270 35096 6276 35108
rect 6328 35096 6334 35148
rect 7098 35096 7104 35148
rect 7156 35136 7162 35148
rect 7285 35139 7343 35145
rect 7285 35136 7297 35139
rect 7156 35108 7297 35136
rect 7156 35096 7162 35108
rect 7285 35105 7297 35108
rect 7331 35105 7343 35139
rect 7285 35099 7343 35105
rect 7837 35139 7895 35145
rect 7837 35105 7849 35139
rect 7883 35136 7895 35139
rect 13446 35136 13452 35148
rect 7883 35108 13452 35136
rect 7883 35105 7895 35108
rect 7837 35099 7895 35105
rect 13446 35096 13452 35108
rect 13504 35096 13510 35148
rect 13556 35145 13584 35176
rect 13814 35164 13820 35176
rect 13872 35204 13878 35216
rect 14369 35207 14427 35213
rect 14369 35204 14381 35207
rect 13872 35176 14381 35204
rect 13872 35164 13878 35176
rect 14369 35173 14381 35176
rect 14415 35204 14427 35207
rect 19702 35204 19708 35216
rect 14415 35176 19708 35204
rect 14415 35173 14427 35176
rect 14369 35167 14427 35173
rect 19702 35164 19708 35176
rect 19760 35164 19766 35216
rect 13541 35139 13599 35145
rect 13541 35105 13553 35139
rect 13587 35105 13599 35139
rect 13541 35099 13599 35105
rect 13909 35139 13967 35145
rect 13909 35105 13921 35139
rect 13955 35136 13967 35139
rect 13998 35136 14004 35148
rect 13955 35108 14004 35136
rect 13955 35105 13967 35108
rect 13909 35099 13967 35105
rect 13998 35096 14004 35108
rect 14056 35096 14062 35148
rect 14093 35139 14151 35145
rect 14093 35105 14105 35139
rect 14139 35136 14151 35139
rect 14458 35136 14464 35148
rect 14139 35108 14464 35136
rect 14139 35105 14151 35108
rect 14093 35099 14151 35105
rect 14458 35096 14464 35108
rect 14516 35096 14522 35148
rect 18322 35096 18328 35148
rect 18380 35136 18386 35148
rect 18417 35139 18475 35145
rect 18417 35136 18429 35139
rect 18380 35108 18429 35136
rect 18380 35096 18386 35108
rect 18417 35105 18429 35108
rect 18463 35136 18475 35139
rect 18969 35139 19027 35145
rect 18969 35136 18981 35139
rect 18463 35108 18981 35136
rect 18463 35105 18475 35108
rect 18417 35099 18475 35105
rect 18969 35105 18981 35108
rect 19015 35105 19027 35139
rect 18969 35099 19027 35105
rect 19153 35139 19211 35145
rect 19153 35105 19165 35139
rect 19199 35136 19211 35139
rect 19812 35136 19840 35235
rect 20714 35232 20720 35244
rect 20772 35232 20778 35284
rect 22186 35232 22192 35284
rect 22244 35272 22250 35284
rect 25133 35275 25191 35281
rect 25133 35272 25145 35275
rect 22244 35244 25145 35272
rect 22244 35232 22250 35244
rect 25133 35241 25145 35244
rect 25179 35272 25191 35275
rect 25314 35272 25320 35284
rect 25179 35244 25320 35272
rect 25179 35241 25191 35244
rect 25133 35235 25191 35241
rect 25314 35232 25320 35244
rect 25372 35232 25378 35284
rect 28261 35275 28319 35281
rect 28261 35241 28273 35275
rect 28307 35272 28319 35275
rect 30374 35272 30380 35284
rect 28307 35244 29408 35272
rect 30335 35244 30380 35272
rect 28307 35241 28319 35244
rect 28261 35235 28319 35241
rect 24397 35207 24455 35213
rect 24397 35204 24409 35207
rect 22756 35176 24409 35204
rect 21818 35136 21824 35148
rect 19199 35108 19840 35136
rect 21779 35108 21824 35136
rect 19199 35105 19211 35108
rect 19153 35099 19211 35105
rect 21818 35096 21824 35108
rect 21876 35096 21882 35148
rect 22370 35136 22376 35148
rect 21928 35108 22376 35136
rect 3602 35028 3608 35080
rect 3660 35068 3666 35080
rect 9398 35068 9404 35080
rect 3660 35040 9404 35068
rect 3660 35028 3666 35040
rect 9398 35028 9404 35040
rect 9456 35028 9462 35080
rect 13633 35071 13691 35077
rect 13633 35037 13645 35071
rect 13679 35068 13691 35071
rect 14016 35068 14044 35096
rect 14642 35068 14648 35080
rect 13679 35040 13952 35068
rect 14016 35040 14648 35068
rect 13679 35037 13691 35040
rect 13633 35031 13691 35037
rect 13924 35012 13952 35040
rect 14642 35028 14648 35040
rect 14700 35028 14706 35080
rect 18233 35071 18291 35077
rect 18233 35068 18245 35071
rect 18064 35040 18245 35068
rect 3418 34960 3424 35012
rect 3476 35000 3482 35012
rect 3786 35000 3792 35012
rect 3476 34972 3792 35000
rect 3476 34960 3482 34972
rect 3786 34960 3792 34972
rect 3844 34960 3850 35012
rect 13906 34960 13912 35012
rect 13964 35000 13970 35012
rect 14185 35003 14243 35009
rect 14185 35000 14197 35003
rect 13964 34972 14197 35000
rect 13964 34960 13970 34972
rect 14185 34969 14197 34972
rect 14231 34969 14243 35003
rect 14185 34963 14243 34969
rect 4062 34892 4068 34944
rect 4120 34932 4126 34944
rect 15654 34932 15660 34944
rect 4120 34904 15660 34932
rect 4120 34892 4126 34904
rect 15654 34892 15660 34904
rect 15712 34892 15718 34944
rect 17310 34892 17316 34944
rect 17368 34932 17374 34944
rect 18064 34941 18092 35040
rect 18233 35037 18245 35040
rect 18279 35037 18291 35071
rect 21928 35068 21956 35108
rect 22370 35096 22376 35108
rect 22428 35136 22434 35148
rect 22756 35136 22784 35176
rect 24397 35173 24409 35176
rect 24443 35204 24455 35207
rect 24443 35176 29316 35204
rect 24443 35173 24455 35176
rect 24397 35167 24455 35173
rect 24302 35136 24308 35148
rect 22428 35108 22784 35136
rect 24263 35108 24308 35136
rect 22428 35096 22434 35108
rect 24302 35096 24308 35108
rect 24360 35096 24366 35148
rect 25314 35136 25320 35148
rect 25275 35108 25320 35136
rect 25314 35096 25320 35108
rect 25372 35096 25378 35148
rect 28074 35136 28080 35148
rect 28035 35108 28080 35136
rect 28074 35096 28080 35108
rect 28132 35096 28138 35148
rect 28442 35096 28448 35148
rect 28500 35136 28506 35148
rect 29181 35139 29239 35145
rect 29181 35136 29193 35139
rect 28500 35108 29193 35136
rect 28500 35096 28506 35108
rect 29181 35105 29193 35108
rect 29227 35105 29239 35139
rect 29181 35099 29239 35105
rect 18233 35031 18291 35037
rect 21836 35040 21956 35068
rect 18138 34960 18144 35012
rect 18196 35000 18202 35012
rect 21836 35000 21864 35040
rect 22094 35028 22100 35080
rect 22152 35068 22158 35080
rect 22152 35040 22197 35068
rect 22152 35028 22158 35040
rect 22278 35028 22284 35080
rect 22336 35068 22342 35080
rect 22830 35068 22836 35080
rect 22336 35040 22836 35068
rect 22336 35028 22342 35040
rect 22830 35028 22836 35040
rect 22888 35028 22894 35080
rect 22922 35028 22928 35080
rect 22980 35068 22986 35080
rect 22980 35040 29224 35068
rect 22980 35028 22986 35040
rect 18196 34972 21864 35000
rect 18196 34960 18202 34972
rect 25038 34960 25044 35012
rect 25096 35000 25102 35012
rect 25501 35003 25559 35009
rect 25501 35000 25513 35003
rect 25096 34972 25513 35000
rect 25096 34960 25102 34972
rect 25501 34969 25513 34972
rect 25547 34969 25559 35003
rect 29086 35000 29092 35012
rect 25501 34963 25559 34969
rect 25608 34972 29092 35000
rect 18049 34935 18107 34941
rect 18049 34932 18061 34935
rect 17368 34904 18061 34932
rect 17368 34892 17374 34904
rect 18049 34901 18061 34904
rect 18095 34901 18107 34935
rect 18049 34895 18107 34901
rect 18782 34892 18788 34944
rect 18840 34932 18846 34944
rect 22278 34932 22284 34944
rect 18840 34904 22284 34932
rect 18840 34892 18846 34904
rect 22278 34892 22284 34904
rect 22336 34892 22342 34944
rect 23382 34932 23388 34944
rect 23343 34904 23388 34932
rect 23382 34892 23388 34904
rect 23440 34892 23446 34944
rect 23658 34932 23664 34944
rect 23571 34904 23664 34932
rect 23658 34892 23664 34904
rect 23716 34932 23722 34944
rect 25608 34932 25636 34972
rect 29086 34960 29092 34972
rect 29144 34960 29150 35012
rect 23716 34904 25636 34932
rect 23716 34892 23722 34904
rect 26050 34892 26056 34944
rect 26108 34932 26114 34944
rect 27614 34932 27620 34944
rect 26108 34904 27620 34932
rect 26108 34892 26114 34904
rect 27614 34892 27620 34904
rect 27672 34932 27678 34944
rect 27893 34935 27951 34941
rect 27893 34932 27905 34935
rect 27672 34904 27905 34932
rect 27672 34892 27678 34904
rect 27893 34901 27905 34904
rect 27939 34932 27951 34935
rect 28074 34932 28080 34944
rect 27939 34904 28080 34932
rect 27939 34901 27951 34904
rect 27893 34895 27951 34901
rect 28074 34892 28080 34904
rect 28132 34892 28138 34944
rect 28442 34892 28448 34944
rect 28500 34932 28506 34944
rect 28997 34935 29055 34941
rect 28997 34932 29009 34935
rect 28500 34904 29009 34932
rect 28500 34892 28506 34904
rect 28997 34901 29009 34904
rect 29043 34901 29055 34935
rect 29196 34932 29224 35040
rect 29288 35000 29316 35176
rect 29380 35145 29408 35244
rect 30374 35232 30380 35244
rect 30432 35232 30438 35284
rect 30466 35232 30472 35284
rect 30524 35272 30530 35284
rect 34333 35275 34391 35281
rect 34333 35272 34345 35275
rect 30524 35244 34345 35272
rect 30524 35232 30530 35244
rect 34333 35241 34345 35244
rect 34379 35272 34391 35275
rect 34701 35275 34759 35281
rect 34379 35244 34560 35272
rect 34379 35241 34391 35244
rect 34333 35235 34391 35241
rect 31294 35204 31300 35216
rect 29932 35176 31300 35204
rect 29932 35145 29960 35176
rect 31294 35164 31300 35176
rect 31352 35164 31358 35216
rect 32876 35176 33916 35204
rect 32876 35148 32904 35176
rect 29365 35139 29423 35145
rect 29365 35105 29377 35139
rect 29411 35136 29423 35139
rect 29917 35139 29975 35145
rect 29917 35136 29929 35139
rect 29411 35108 29929 35136
rect 29411 35105 29423 35108
rect 29365 35099 29423 35105
rect 29917 35105 29929 35108
rect 29963 35105 29975 35139
rect 30098 35136 30104 35148
rect 30059 35108 30104 35136
rect 29917 35099 29975 35105
rect 30098 35096 30104 35108
rect 30156 35096 30162 35148
rect 30282 35096 30288 35148
rect 30340 35096 30346 35148
rect 32306 35145 32312 35148
rect 31481 35139 31539 35145
rect 31481 35105 31493 35139
rect 31527 35136 31539 35139
rect 32294 35139 32312 35145
rect 31527 35108 32260 35136
rect 31527 35105 31539 35108
rect 31481 35099 31539 35105
rect 30300 35068 30328 35096
rect 31662 35068 31668 35080
rect 30300 35040 31668 35068
rect 31662 35028 31668 35040
rect 31720 35028 31726 35080
rect 31754 35028 31760 35080
rect 31812 35068 31818 35080
rect 32125 35071 32183 35077
rect 32125 35068 32137 35071
rect 31812 35040 32137 35068
rect 31812 35028 31818 35040
rect 32125 35037 32137 35040
rect 32171 35037 32183 35071
rect 32232 35068 32260 35108
rect 32294 35105 32306 35139
rect 32294 35099 32312 35105
rect 32306 35096 32312 35099
rect 32364 35096 32370 35148
rect 32769 35139 32827 35145
rect 32769 35136 32781 35139
rect 32508 35108 32781 35136
rect 32508 35068 32536 35108
rect 32769 35105 32781 35108
rect 32815 35105 32827 35139
rect 32769 35099 32827 35105
rect 32858 35096 32864 35148
rect 32916 35136 32922 35148
rect 32916 35108 33009 35136
rect 32916 35096 32922 35108
rect 33318 35096 33324 35148
rect 33376 35136 33382 35148
rect 33376 35108 33456 35136
rect 33376 35096 33382 35108
rect 33428 35077 33456 35108
rect 33888 35080 33916 35176
rect 34532 35145 34560 35244
rect 34701 35241 34713 35275
rect 34747 35272 34759 35275
rect 38930 35272 38936 35284
rect 34747 35244 35572 35272
rect 34747 35241 34759 35244
rect 34701 35235 34759 35241
rect 35544 35145 35572 35244
rect 36464 35244 38936 35272
rect 34517 35139 34575 35145
rect 34517 35105 34529 35139
rect 34563 35105 34575 35139
rect 34517 35099 34575 35105
rect 35529 35139 35587 35145
rect 35529 35105 35541 35139
rect 35575 35136 35587 35139
rect 36262 35136 36268 35148
rect 35575 35108 36268 35136
rect 35575 35105 35587 35108
rect 35529 35099 35587 35105
rect 36262 35096 36268 35108
rect 36320 35096 36326 35148
rect 32232 35040 32536 35068
rect 33413 35071 33471 35077
rect 32125 35031 32183 35037
rect 33413 35037 33425 35071
rect 33459 35037 33471 35071
rect 33870 35068 33876 35080
rect 33831 35040 33876 35068
rect 33413 35031 33471 35037
rect 33870 35028 33876 35040
rect 33928 35028 33934 35080
rect 35618 35068 35624 35080
rect 35579 35040 35624 35068
rect 35618 35028 35624 35040
rect 35676 35028 35682 35080
rect 36357 35071 36415 35077
rect 36357 35037 36369 35071
rect 36403 35068 36415 35071
rect 36464 35068 36492 35244
rect 38930 35232 38936 35244
rect 38988 35232 38994 35284
rect 39025 35275 39083 35281
rect 39025 35241 39037 35275
rect 39071 35272 39083 35275
rect 40494 35272 40500 35284
rect 39071 35244 40500 35272
rect 39071 35241 39083 35244
rect 39025 35235 39083 35241
rect 40494 35232 40500 35244
rect 40552 35232 40558 35284
rect 42245 35275 42303 35281
rect 42245 35241 42257 35275
rect 42291 35272 42303 35275
rect 42886 35272 42892 35284
rect 42291 35244 42892 35272
rect 42291 35241 42303 35244
rect 42245 35235 42303 35241
rect 42886 35232 42892 35244
rect 42944 35232 42950 35284
rect 43990 35232 43996 35284
rect 44048 35272 44054 35284
rect 48038 35272 48044 35284
rect 44048 35244 44496 35272
rect 44048 35232 44054 35244
rect 36814 35164 36820 35216
rect 36872 35204 36878 35216
rect 41690 35204 41696 35216
rect 36872 35176 41696 35204
rect 36872 35164 36878 35176
rect 41690 35164 41696 35176
rect 41748 35164 41754 35216
rect 42978 35164 42984 35216
rect 43036 35204 43042 35216
rect 43073 35207 43131 35213
rect 43073 35204 43085 35207
rect 43036 35176 43085 35204
rect 43036 35164 43042 35176
rect 43073 35173 43085 35176
rect 43119 35204 43131 35207
rect 44082 35204 44088 35216
rect 43119 35176 44088 35204
rect 43119 35173 43131 35176
rect 43073 35167 43131 35173
rect 36630 35145 36636 35148
rect 36604 35139 36636 35145
rect 36604 35105 36616 35139
rect 36604 35099 36636 35105
rect 36630 35096 36636 35099
rect 36688 35096 36694 35148
rect 36722 35096 36728 35148
rect 36780 35136 36786 35148
rect 36780 35108 36825 35136
rect 36780 35096 36786 35108
rect 37274 35096 37280 35148
rect 37332 35136 37338 35148
rect 37829 35139 37887 35145
rect 37829 35136 37841 35139
rect 37332 35108 37841 35136
rect 37332 35096 37338 35108
rect 37829 35105 37841 35108
rect 37875 35105 37887 35139
rect 38010 35136 38016 35148
rect 37971 35108 38016 35136
rect 37829 35099 37887 35105
rect 36998 35068 37004 35080
rect 36403 35040 36492 35068
rect 36911 35040 37004 35068
rect 36403 35037 36415 35040
rect 36357 35031 36415 35037
rect 36998 35028 37004 35040
rect 37056 35068 37062 35080
rect 37737 35071 37795 35077
rect 37737 35068 37749 35071
rect 37056 35040 37749 35068
rect 37056 35028 37062 35040
rect 37737 35037 37749 35040
rect 37783 35037 37795 35071
rect 37844 35068 37872 35099
rect 38010 35096 38016 35108
rect 38068 35096 38074 35148
rect 38473 35139 38531 35145
rect 38473 35136 38485 35139
rect 38120 35108 38485 35136
rect 38120 35068 38148 35108
rect 38473 35105 38485 35108
rect 38519 35105 38531 35139
rect 38473 35099 38531 35105
rect 38565 35139 38623 35145
rect 38565 35105 38577 35139
rect 38611 35136 38623 35139
rect 38654 35136 38660 35148
rect 38611 35108 38660 35136
rect 38611 35105 38623 35108
rect 38565 35099 38623 35105
rect 38654 35096 38660 35108
rect 38712 35136 38718 35148
rect 39393 35139 39451 35145
rect 39393 35136 39405 35139
rect 38712 35108 39405 35136
rect 38712 35096 38718 35108
rect 39393 35105 39405 35108
rect 39439 35136 39451 35139
rect 39574 35136 39580 35148
rect 39439 35108 39580 35136
rect 39439 35105 39451 35108
rect 39393 35099 39451 35105
rect 39574 35096 39580 35108
rect 39632 35096 39638 35148
rect 40586 35136 40592 35148
rect 40499 35108 40592 35136
rect 40586 35096 40592 35108
rect 40644 35136 40650 35148
rect 40773 35139 40831 35145
rect 40773 35136 40785 35139
rect 40644 35108 40785 35136
rect 40644 35096 40650 35108
rect 40773 35105 40785 35108
rect 40819 35136 40831 35139
rect 41233 35139 41291 35145
rect 41233 35136 41245 35139
rect 40819 35108 41245 35136
rect 40819 35105 40831 35108
rect 40773 35099 40831 35105
rect 41233 35105 41245 35108
rect 41279 35136 41291 35139
rect 41782 35136 41788 35148
rect 41279 35108 41788 35136
rect 41279 35105 41291 35108
rect 41233 35099 41291 35105
rect 41782 35096 41788 35108
rect 41840 35096 41846 35148
rect 44008 35145 44036 35176
rect 44082 35164 44088 35176
rect 44140 35164 44146 35216
rect 41969 35139 42027 35145
rect 41969 35105 41981 35139
rect 42015 35136 42027 35139
rect 43993 35139 44051 35145
rect 42015 35108 43576 35136
rect 42015 35105 42027 35108
rect 41969 35099 42027 35105
rect 37844 35040 38148 35068
rect 39040 35040 40908 35068
rect 37737 35031 37795 35037
rect 38746 35000 38752 35012
rect 29288 34972 38752 35000
rect 38746 34960 38752 34972
rect 38804 34960 38810 35012
rect 31481 34935 31539 34941
rect 31481 34932 31493 34935
rect 29196 34904 31493 34932
rect 28997 34895 29055 34901
rect 31481 34901 31493 34904
rect 31527 34932 31539 34935
rect 31573 34935 31631 34941
rect 31573 34932 31585 34935
rect 31527 34904 31585 34932
rect 31527 34901 31539 34904
rect 31481 34895 31539 34901
rect 31573 34901 31585 34904
rect 31619 34901 31631 34935
rect 31573 34895 31631 34901
rect 31662 34892 31668 34944
rect 31720 34932 31726 34944
rect 33502 34932 33508 34944
rect 31720 34904 33508 34932
rect 31720 34892 31726 34904
rect 33502 34892 33508 34904
rect 33560 34892 33566 34944
rect 33594 34892 33600 34944
rect 33652 34932 33658 34944
rect 33689 34935 33747 34941
rect 33689 34932 33701 34935
rect 33652 34904 33701 34932
rect 33652 34892 33658 34904
rect 33689 34901 33701 34904
rect 33735 34932 33747 34935
rect 37090 34932 37096 34944
rect 33735 34904 37096 34932
rect 33735 34901 33747 34904
rect 33689 34895 33747 34901
rect 37090 34892 37096 34904
rect 37148 34892 37154 34944
rect 37274 34932 37280 34944
rect 37235 34904 37280 34932
rect 37274 34892 37280 34904
rect 37332 34932 37338 34944
rect 37461 34935 37519 34941
rect 37461 34932 37473 34935
rect 37332 34904 37473 34932
rect 37332 34892 37338 34904
rect 37461 34901 37473 34904
rect 37507 34901 37519 34935
rect 37461 34895 37519 34901
rect 37737 34935 37795 34941
rect 37737 34901 37749 34935
rect 37783 34932 37795 34935
rect 39040 34932 39068 35040
rect 40880 35000 40908 35040
rect 40954 35028 40960 35080
rect 41012 35068 41018 35080
rect 41141 35071 41199 35077
rect 41141 35068 41153 35071
rect 41012 35040 41153 35068
rect 41012 35028 41018 35040
rect 41141 35037 41153 35040
rect 41187 35037 41199 35071
rect 43438 35068 43444 35080
rect 43399 35040 43444 35068
rect 41141 35031 41199 35037
rect 43438 35028 43444 35040
rect 43496 35028 43502 35080
rect 43548 35068 43576 35108
rect 43993 35105 44005 35139
rect 44039 35105 44051 35139
rect 44358 35136 44364 35148
rect 44319 35108 44364 35136
rect 43993 35099 44051 35105
rect 44358 35096 44364 35108
rect 44416 35096 44422 35148
rect 44468 35145 44496 35244
rect 47504 35244 48044 35272
rect 46566 35164 46572 35216
rect 46624 35204 46630 35216
rect 46624 35176 47256 35204
rect 46624 35164 46630 35176
rect 44453 35139 44511 35145
rect 44453 35105 44465 35139
rect 44499 35105 44511 35139
rect 44453 35099 44511 35105
rect 47121 35139 47179 35145
rect 47121 35105 47133 35139
rect 47167 35105 47179 35139
rect 47228 35136 47256 35176
rect 47504 35136 47532 35244
rect 48038 35232 48044 35244
rect 48096 35232 48102 35284
rect 48133 35275 48191 35281
rect 48133 35241 48145 35275
rect 48179 35272 48191 35275
rect 49878 35272 49884 35284
rect 48179 35244 49884 35272
rect 48179 35241 48191 35244
rect 48133 35235 48191 35241
rect 49878 35232 49884 35244
rect 49936 35232 49942 35284
rect 49970 35232 49976 35284
rect 50028 35272 50034 35284
rect 51626 35272 51632 35284
rect 50028 35244 50752 35272
rect 50028 35232 50034 35244
rect 47762 35164 47768 35216
rect 47820 35204 47826 35216
rect 47820 35176 50200 35204
rect 47820 35164 47826 35176
rect 47581 35139 47639 35145
rect 47581 35136 47593 35139
rect 47228 35108 47593 35136
rect 47121 35099 47179 35105
rect 47581 35105 47593 35108
rect 47627 35105 47639 35139
rect 47581 35099 47639 35105
rect 47673 35139 47731 35145
rect 47673 35105 47685 35139
rect 47719 35136 47731 35139
rect 48501 35139 48559 35145
rect 48501 35136 48513 35139
rect 47719 35108 48513 35136
rect 47719 35105 47731 35108
rect 47673 35099 47731 35105
rect 48501 35105 48513 35108
rect 48547 35136 48559 35139
rect 49142 35136 49148 35148
rect 48547 35108 49148 35136
rect 48547 35105 48559 35108
rect 48501 35099 48559 35105
rect 44085 35071 44143 35077
rect 44085 35068 44097 35071
rect 43548 35040 44097 35068
rect 44085 35037 44097 35040
rect 44131 35068 44143 35071
rect 44174 35068 44180 35080
rect 44131 35040 44180 35068
rect 44131 35037 44143 35040
rect 44085 35031 44143 35037
rect 44174 35028 44180 35040
rect 44232 35028 44238 35080
rect 46750 35028 46756 35080
rect 46808 35068 46814 35080
rect 46937 35071 46995 35077
rect 46937 35068 46949 35071
rect 46808 35040 46949 35068
rect 46808 35028 46814 35040
rect 46937 35037 46949 35040
rect 46983 35037 46995 35071
rect 46937 35031 46995 35037
rect 42889 35003 42947 35009
rect 40880 34972 42564 35000
rect 37783 34904 39068 34932
rect 42536 34932 42564 34972
rect 42889 34969 42901 35003
rect 42935 35000 42947 35003
rect 44266 35000 44272 35012
rect 42935 34972 44272 35000
rect 42935 34969 42947 34972
rect 42889 34963 42947 34969
rect 42904 34932 42932 34963
rect 44266 34960 44272 34972
rect 44324 34960 44330 35012
rect 47136 35000 47164 35099
rect 49142 35096 49148 35108
rect 49200 35096 49206 35148
rect 49602 35096 49608 35148
rect 49660 35136 49666 35148
rect 50065 35139 50123 35145
rect 50065 35136 50077 35139
rect 49660 35108 50077 35136
rect 49660 35096 49666 35108
rect 50065 35105 50077 35108
rect 50111 35105 50123 35139
rect 50065 35099 50123 35105
rect 48866 35028 48872 35080
rect 48924 35068 48930 35080
rect 49881 35071 49939 35077
rect 49881 35068 49893 35071
rect 48924 35040 49893 35068
rect 48924 35028 48930 35040
rect 49881 35037 49893 35040
rect 49927 35068 49939 35071
rect 49970 35068 49976 35080
rect 49927 35040 49976 35068
rect 49927 35037 49939 35040
rect 49881 35031 49939 35037
rect 49970 35028 49976 35040
rect 50028 35028 50034 35080
rect 48685 35003 48743 35009
rect 48685 35000 48697 35003
rect 47136 34972 48697 35000
rect 48685 34969 48697 34972
rect 48731 35000 48743 35003
rect 50172 35000 50200 35176
rect 50246 35096 50252 35148
rect 50304 35136 50310 35148
rect 50724 35145 50752 35244
rect 50816 35244 51632 35272
rect 50816 35145 50844 35244
rect 51626 35232 51632 35244
rect 51684 35232 51690 35284
rect 51994 35232 52000 35284
rect 52052 35272 52058 35284
rect 56134 35272 56140 35284
rect 52052 35244 56140 35272
rect 52052 35232 52058 35244
rect 56134 35232 56140 35244
rect 56192 35232 56198 35284
rect 56318 35272 56324 35284
rect 56279 35244 56324 35272
rect 56318 35232 56324 35244
rect 56376 35232 56382 35284
rect 56502 35232 56508 35284
rect 56560 35272 56566 35284
rect 56560 35244 58940 35272
rect 56560 35232 56566 35244
rect 52362 35164 52368 35216
rect 52420 35204 52426 35216
rect 57974 35204 57980 35216
rect 52420 35176 57980 35204
rect 52420 35164 52426 35176
rect 57974 35164 57980 35176
rect 58032 35164 58038 35216
rect 58069 35207 58127 35213
rect 58069 35173 58081 35207
rect 58115 35204 58127 35207
rect 58802 35204 58808 35216
rect 58115 35176 58808 35204
rect 58115 35173 58127 35176
rect 58069 35167 58127 35173
rect 58802 35164 58808 35176
rect 58860 35164 58866 35216
rect 58912 35204 58940 35244
rect 59814 35232 59820 35284
rect 59872 35272 59878 35284
rect 63313 35275 63371 35281
rect 63313 35272 63325 35275
rect 59872 35244 63325 35272
rect 59872 35232 59878 35244
rect 63313 35241 63325 35244
rect 63359 35241 63371 35275
rect 65797 35275 65855 35281
rect 65797 35272 65809 35275
rect 63313 35235 63371 35241
rect 64524 35244 65809 35272
rect 64524 35204 64552 35244
rect 65797 35241 65809 35244
rect 65843 35272 65855 35275
rect 65889 35275 65947 35281
rect 65889 35272 65901 35275
rect 65843 35244 65901 35272
rect 65843 35241 65855 35244
rect 65797 35235 65855 35241
rect 65889 35241 65901 35244
rect 65935 35272 65947 35275
rect 66073 35275 66131 35281
rect 66073 35272 66085 35275
rect 65935 35244 66085 35272
rect 65935 35241 65947 35244
rect 65889 35235 65947 35241
rect 66073 35241 66085 35244
rect 66119 35272 66131 35275
rect 66119 35244 67220 35272
rect 66119 35241 66131 35244
rect 66073 35235 66131 35241
rect 58912 35176 64552 35204
rect 64598 35164 64604 35216
rect 64656 35204 64662 35216
rect 64656 35176 67128 35204
rect 64656 35164 64662 35176
rect 67100 35148 67128 35176
rect 50709 35139 50767 35145
rect 50304 35108 50349 35136
rect 50304 35096 50310 35108
rect 50709 35105 50721 35139
rect 50755 35105 50767 35139
rect 50709 35099 50767 35105
rect 50801 35139 50859 35145
rect 50801 35105 50813 35139
rect 50847 35105 50859 35139
rect 53282 35136 53288 35148
rect 53243 35108 53288 35136
rect 50801 35099 50859 35105
rect 53282 35096 53288 35108
rect 53340 35096 53346 35148
rect 53834 35096 53840 35148
rect 53892 35136 53898 35148
rect 54573 35139 54631 35145
rect 54573 35136 54585 35139
rect 53892 35108 54585 35136
rect 53892 35096 53898 35108
rect 54573 35105 54585 35108
rect 54619 35105 54631 35139
rect 54573 35099 54631 35105
rect 55766 35096 55772 35148
rect 55824 35136 55830 35148
rect 56689 35139 56747 35145
rect 56689 35136 56701 35139
rect 55824 35108 56701 35136
rect 55824 35096 55830 35108
rect 56689 35105 56701 35108
rect 56735 35136 56747 35139
rect 56735 35108 56916 35136
rect 56735 35105 56747 35108
rect 56689 35099 56747 35105
rect 51350 35068 51356 35080
rect 51311 35040 51356 35068
rect 51350 35028 51356 35040
rect 51408 35028 51414 35080
rect 51810 35068 51816 35080
rect 51771 35040 51816 35068
rect 51810 35028 51816 35040
rect 51868 35028 51874 35080
rect 51994 35028 52000 35080
rect 52052 35068 52058 35080
rect 56134 35068 56140 35080
rect 52052 35040 56140 35068
rect 52052 35028 52058 35040
rect 56134 35028 56140 35040
rect 56192 35028 56198 35080
rect 56410 35028 56416 35080
rect 56468 35068 56474 35080
rect 56781 35071 56839 35077
rect 56781 35068 56793 35071
rect 56468 35040 56793 35068
rect 56468 35028 56474 35040
rect 56781 35037 56793 35040
rect 56827 35037 56839 35071
rect 56888 35068 56916 35108
rect 56962 35096 56968 35148
rect 57020 35136 57026 35148
rect 57425 35139 57483 35145
rect 57425 35136 57437 35139
rect 57020 35108 57065 35136
rect 57164 35108 57437 35136
rect 57020 35096 57026 35108
rect 57164 35068 57192 35108
rect 57425 35105 57437 35108
rect 57471 35105 57483 35139
rect 57425 35099 57483 35105
rect 57517 35139 57575 35145
rect 57517 35105 57529 35139
rect 57563 35136 57575 35139
rect 58345 35139 58403 35145
rect 58345 35136 58357 35139
rect 57563 35108 58357 35136
rect 57563 35105 57575 35108
rect 57517 35099 57575 35105
rect 58345 35105 58357 35108
rect 58391 35136 58403 35139
rect 58434 35136 58440 35148
rect 58391 35108 58440 35136
rect 58391 35105 58403 35108
rect 58345 35099 58403 35105
rect 58434 35096 58440 35108
rect 58492 35096 58498 35148
rect 58529 35139 58587 35145
rect 58529 35105 58541 35139
rect 58575 35136 58587 35139
rect 58618 35136 58624 35148
rect 58575 35108 58624 35136
rect 58575 35105 58587 35108
rect 58529 35099 58587 35105
rect 58618 35096 58624 35108
rect 58676 35096 58682 35148
rect 62301 35139 62359 35145
rect 62301 35105 62313 35139
rect 62347 35105 62359 35139
rect 62758 35136 62764 35148
rect 62719 35108 62764 35136
rect 62301 35099 62359 35105
rect 56888 35040 57192 35068
rect 56781 35031 56839 35037
rect 57974 35028 57980 35080
rect 58032 35068 58038 35080
rect 61194 35068 61200 35080
rect 58032 35040 61200 35068
rect 58032 35028 58038 35040
rect 61194 35028 61200 35040
rect 61252 35028 61258 35080
rect 62117 35071 62175 35077
rect 62117 35037 62129 35071
rect 62163 35037 62175 35071
rect 62117 35031 62175 35037
rect 62022 35000 62028 35012
rect 48731 34972 50108 35000
rect 50172 34972 62028 35000
rect 48731 34969 48743 34972
rect 48685 34963 48743 34969
rect 46566 34932 46572 34944
rect 42536 34904 42932 34932
rect 46527 34904 46572 34932
rect 37783 34901 37795 34904
rect 37737 34895 37795 34901
rect 46566 34892 46572 34904
rect 46624 34892 46630 34944
rect 46750 34932 46756 34944
rect 46711 34904 46756 34932
rect 46750 34892 46756 34904
rect 46808 34892 46814 34944
rect 46842 34892 46848 34944
rect 46900 34932 46906 34944
rect 49418 34932 49424 34944
rect 46900 34904 49424 34932
rect 46900 34892 46906 34904
rect 49418 34892 49424 34904
rect 49476 34892 49482 34944
rect 49602 34892 49608 34944
rect 49660 34932 49666 34944
rect 49697 34935 49755 34941
rect 49697 34932 49709 34935
rect 49660 34904 49709 34932
rect 49660 34892 49666 34904
rect 49697 34901 49709 34904
rect 49743 34901 49755 34935
rect 50080 34932 50108 34972
rect 62022 34960 62028 34972
rect 62080 34960 62086 35012
rect 51994 34932 52000 34944
rect 50080 34904 52000 34932
rect 49697 34895 49755 34901
rect 51994 34892 52000 34904
rect 52052 34892 52058 34944
rect 53006 34892 53012 34944
rect 53064 34932 53070 34944
rect 53377 34935 53435 34941
rect 53377 34932 53389 34935
rect 53064 34904 53389 34932
rect 53064 34892 53070 34904
rect 53377 34901 53389 34904
rect 53423 34901 53435 34935
rect 54018 34932 54024 34944
rect 53979 34904 54024 34932
rect 53377 34895 53435 34901
rect 54018 34892 54024 34904
rect 54076 34892 54082 34944
rect 54202 34932 54208 34944
rect 54163 34904 54208 34932
rect 54202 34892 54208 34904
rect 54260 34892 54266 34944
rect 54754 34932 54760 34944
rect 54715 34904 54760 34932
rect 54754 34892 54760 34904
rect 54812 34892 54818 34944
rect 54846 34892 54852 34944
rect 54904 34932 54910 34944
rect 54941 34935 54999 34941
rect 54941 34932 54953 34935
rect 54904 34904 54953 34932
rect 54904 34892 54910 34904
rect 54941 34901 54953 34904
rect 54987 34901 54999 34935
rect 56410 34932 56416 34944
rect 56371 34904 56416 34932
rect 54941 34895 54999 34901
rect 56410 34892 56416 34904
rect 56468 34892 56474 34944
rect 56962 34892 56968 34944
rect 57020 34932 57026 34944
rect 57790 34932 57796 34944
rect 57020 34904 57796 34932
rect 57020 34892 57026 34904
rect 57790 34892 57796 34904
rect 57848 34932 57854 34944
rect 58618 34932 58624 34944
rect 57848 34904 58624 34932
rect 57848 34892 57854 34904
rect 58618 34892 58624 34904
rect 58676 34892 58682 34944
rect 61746 34932 61752 34944
rect 61707 34904 61752 34932
rect 61746 34892 61752 34904
rect 61804 34932 61810 34944
rect 61933 34935 61991 34941
rect 61933 34932 61945 34935
rect 61804 34904 61945 34932
rect 61804 34892 61810 34904
rect 61933 34901 61945 34904
rect 61979 34932 61991 34935
rect 62132 34932 62160 35031
rect 62316 35000 62344 35099
rect 62758 35096 62764 35108
rect 62816 35096 62822 35148
rect 62853 35139 62911 35145
rect 62853 35105 62865 35139
rect 62899 35136 62911 35139
rect 63034 35136 63040 35148
rect 62899 35108 63040 35136
rect 62899 35105 62911 35108
rect 62853 35099 62911 35105
rect 63034 35096 63040 35108
rect 63092 35096 63098 35148
rect 64322 35096 64328 35148
rect 64380 35136 64386 35148
rect 64693 35139 64751 35145
rect 64693 35136 64705 35139
rect 64380 35108 64705 35136
rect 64380 35096 64386 35108
rect 64693 35105 64705 35108
rect 64739 35105 64751 35139
rect 64693 35099 64751 35105
rect 65797 35139 65855 35145
rect 65797 35105 65809 35139
rect 65843 35136 65855 35139
rect 66625 35139 66683 35145
rect 66625 35136 66637 35139
rect 65843 35108 66637 35136
rect 65843 35105 65855 35108
rect 65797 35099 65855 35105
rect 66625 35105 66637 35108
rect 66671 35105 66683 35139
rect 66625 35099 66683 35105
rect 66714 35096 66720 35148
rect 66772 35136 66778 35148
rect 67082 35136 67088 35148
rect 66772 35108 66817 35136
rect 66995 35108 67088 35136
rect 66772 35096 66778 35108
rect 67082 35096 67088 35108
rect 67140 35096 67146 35148
rect 67192 35145 67220 35244
rect 69198 35232 69204 35284
rect 69256 35272 69262 35284
rect 87414 35272 87420 35284
rect 69256 35244 87420 35272
rect 69256 35232 69262 35244
rect 87414 35232 87420 35244
rect 87472 35232 87478 35284
rect 88426 35232 88432 35284
rect 88484 35272 88490 35284
rect 90637 35275 90695 35281
rect 90637 35272 90649 35275
rect 88484 35244 90649 35272
rect 88484 35232 88490 35244
rect 90637 35241 90649 35244
rect 90683 35241 90695 35275
rect 90637 35235 90695 35241
rect 67266 35164 67272 35216
rect 67324 35204 67330 35216
rect 68922 35204 68928 35216
rect 67324 35176 68928 35204
rect 67324 35164 67330 35176
rect 68922 35164 68928 35176
rect 68980 35164 68986 35216
rect 70489 35207 70547 35213
rect 70489 35173 70501 35207
rect 70535 35204 70547 35207
rect 71774 35204 71780 35216
rect 70535 35176 71780 35204
rect 70535 35173 70547 35176
rect 70489 35167 70547 35173
rect 71774 35164 71780 35176
rect 71832 35164 71838 35216
rect 75917 35207 75975 35213
rect 75196 35176 75592 35204
rect 67177 35139 67235 35145
rect 67177 35105 67189 35139
rect 67223 35105 67235 35139
rect 67177 35099 67235 35105
rect 68738 35096 68744 35148
rect 68796 35136 68802 35148
rect 69109 35139 69167 35145
rect 69109 35136 69121 35139
rect 68796 35108 69121 35136
rect 68796 35096 68802 35108
rect 69109 35105 69121 35108
rect 69155 35105 69167 35139
rect 69109 35099 69167 35105
rect 73157 35139 73215 35145
rect 73157 35105 73169 35139
rect 73203 35136 73215 35139
rect 73246 35136 73252 35148
rect 73203 35108 73252 35136
rect 73203 35105 73215 35108
rect 73157 35099 73215 35105
rect 73246 35096 73252 35108
rect 73304 35096 73310 35148
rect 74166 35136 74172 35148
rect 73632 35108 74172 35136
rect 64785 35071 64843 35077
rect 64785 35037 64797 35071
rect 64831 35068 64843 35071
rect 66346 35068 66352 35080
rect 64831 35040 66352 35068
rect 64831 35037 64843 35040
rect 64785 35031 64843 35037
rect 66346 35028 66352 35040
rect 66404 35028 66410 35080
rect 68554 35028 68560 35080
rect 68612 35068 68618 35080
rect 68833 35071 68891 35077
rect 68833 35068 68845 35071
rect 68612 35040 68845 35068
rect 68612 35028 68618 35040
rect 68833 35037 68845 35040
rect 68879 35068 68891 35071
rect 70578 35068 70584 35080
rect 68879 35040 70584 35068
rect 68879 35037 68891 35040
rect 68833 35031 68891 35037
rect 70578 35028 70584 35040
rect 70636 35068 70642 35080
rect 72881 35071 72939 35077
rect 72881 35068 72893 35071
rect 70636 35040 72893 35068
rect 70636 35028 70642 35040
rect 72881 35037 72893 35040
rect 72927 35068 72939 35071
rect 73632 35068 73660 35108
rect 74166 35096 74172 35108
rect 74224 35136 74230 35148
rect 74626 35136 74632 35148
rect 74224 35108 74632 35136
rect 74224 35096 74230 35108
rect 74626 35096 74632 35108
rect 74684 35096 74690 35148
rect 74258 35068 74264 35080
rect 72927 35040 73660 35068
rect 74219 35040 74264 35068
rect 72927 35037 72939 35040
rect 72881 35031 72939 35037
rect 74258 35028 74264 35040
rect 74316 35068 74322 35080
rect 75196 35077 75224 35176
rect 75362 35136 75368 35148
rect 75323 35108 75368 35136
rect 75362 35096 75368 35108
rect 75420 35096 75426 35148
rect 75564 35145 75592 35176
rect 75917 35173 75929 35207
rect 75963 35204 75975 35207
rect 76282 35204 76288 35216
rect 75963 35176 76288 35204
rect 75963 35173 75975 35176
rect 75917 35167 75975 35173
rect 76282 35164 76288 35176
rect 76340 35164 76346 35216
rect 78306 35204 78312 35216
rect 76392 35176 78312 35204
rect 75549 35139 75607 35145
rect 75549 35105 75561 35139
rect 75595 35105 75607 35139
rect 75549 35099 75607 35105
rect 75638 35096 75644 35148
rect 75696 35136 75702 35148
rect 76392 35136 76420 35176
rect 78306 35164 78312 35176
rect 78364 35164 78370 35216
rect 84470 35164 84476 35216
rect 84528 35204 84534 35216
rect 84528 35176 84608 35204
rect 84528 35164 84534 35176
rect 75696 35108 76420 35136
rect 77021 35139 77079 35145
rect 75696 35096 75702 35108
rect 77021 35105 77033 35139
rect 77067 35136 77079 35139
rect 77110 35136 77116 35148
rect 77067 35108 77116 35136
rect 77067 35105 77079 35108
rect 77021 35099 77079 35105
rect 77110 35096 77116 35108
rect 77168 35096 77174 35148
rect 78493 35139 78551 35145
rect 78493 35105 78505 35139
rect 78539 35136 78551 35139
rect 79594 35136 79600 35148
rect 78539 35108 79600 35136
rect 78539 35105 78551 35108
rect 78493 35099 78551 35105
rect 79594 35096 79600 35108
rect 79652 35096 79658 35148
rect 81342 35096 81348 35148
rect 81400 35136 81406 35148
rect 83274 35136 83280 35148
rect 81400 35108 83136 35136
rect 83235 35108 83280 35136
rect 81400 35096 81406 35108
rect 75181 35071 75239 35077
rect 75181 35068 75193 35071
rect 74316 35040 75193 35068
rect 74316 35028 74322 35040
rect 75181 35037 75193 35040
rect 75227 35037 75239 35071
rect 75380 35068 75408 35096
rect 76009 35071 76067 35077
rect 76009 35068 76021 35071
rect 75380 35040 76021 35068
rect 75181 35031 75239 35037
rect 76009 35037 76021 35040
rect 76055 35068 76067 35071
rect 78217 35071 78275 35077
rect 78217 35068 78229 35071
rect 76055 35040 77248 35068
rect 76055 35037 76067 35040
rect 76009 35031 76067 35037
rect 63681 35003 63739 35009
rect 63681 35000 63693 35003
rect 62316 34972 63693 35000
rect 63681 34969 63693 34972
rect 63727 35000 63739 35003
rect 67266 35000 67272 35012
rect 63727 34972 67272 35000
rect 63727 34969 63739 34972
rect 63681 34963 63739 34969
rect 67266 34960 67272 34972
rect 67324 34960 67330 35012
rect 67637 35003 67695 35009
rect 67637 34969 67649 35003
rect 67683 35000 67695 35003
rect 68738 35000 68744 35012
rect 67683 34972 68744 35000
rect 67683 34969 67695 34972
rect 67637 34963 67695 34969
rect 68738 34960 68744 34972
rect 68796 34960 68802 35012
rect 77018 35000 77024 35012
rect 74644 34972 77024 35000
rect 62758 34932 62764 34944
rect 61979 34904 62764 34932
rect 61979 34901 61991 34904
rect 61933 34895 61991 34901
rect 62758 34892 62764 34904
rect 62816 34892 62822 34944
rect 63126 34892 63132 34944
rect 63184 34932 63190 34944
rect 63862 34932 63868 34944
rect 63184 34904 63868 34932
rect 63184 34892 63190 34904
rect 63862 34892 63868 34904
rect 63920 34932 63926 34944
rect 64506 34932 64512 34944
rect 63920 34904 64512 34932
rect 63920 34892 63926 34904
rect 64506 34892 64512 34904
rect 64564 34892 64570 34944
rect 66162 34892 66168 34944
rect 66220 34932 66226 34944
rect 66257 34935 66315 34941
rect 66257 34932 66269 34935
rect 66220 34904 66269 34932
rect 66220 34892 66226 34904
rect 66257 34901 66269 34904
rect 66303 34932 66315 34935
rect 66714 34932 66720 34944
rect 66303 34904 66720 34932
rect 66303 34901 66315 34904
rect 66257 34895 66315 34901
rect 66714 34892 66720 34904
rect 66772 34892 66778 34944
rect 67082 34892 67088 34944
rect 67140 34932 67146 34944
rect 69842 34932 69848 34944
rect 67140 34904 69848 34932
rect 67140 34892 67146 34904
rect 69842 34892 69848 34904
rect 69900 34892 69906 34944
rect 69934 34892 69940 34944
rect 69992 34932 69998 34944
rect 74644 34932 74672 34972
rect 77018 34960 77024 34972
rect 77076 34960 77082 35012
rect 77220 35009 77248 35040
rect 78048 35040 78229 35068
rect 77205 35003 77263 35009
rect 77205 34969 77217 35003
rect 77251 34969 77263 35003
rect 77205 34963 77263 34969
rect 78048 34944 78076 35040
rect 78217 35037 78229 35040
rect 78263 35068 78275 35071
rect 82081 35071 82139 35077
rect 78263 35040 82032 35068
rect 78263 35037 78275 35040
rect 78217 35031 78275 35037
rect 82004 35000 82032 35040
rect 82081 35037 82093 35071
rect 82127 35068 82139 35071
rect 82262 35068 82268 35080
rect 82127 35040 82268 35068
rect 82127 35037 82139 35040
rect 82081 35031 82139 35037
rect 82262 35028 82268 35040
rect 82320 35028 82326 35080
rect 82538 35000 82544 35012
rect 82004 34972 82544 35000
rect 82538 34960 82544 34972
rect 82596 34960 82602 35012
rect 69992 34904 74672 34932
rect 69992 34892 69998 34904
rect 75086 34892 75092 34944
rect 75144 34932 75150 34944
rect 77294 34932 77300 34944
rect 75144 34904 77300 34932
rect 75144 34892 75150 34904
rect 77294 34892 77300 34904
rect 77352 34892 77358 34944
rect 78030 34932 78036 34944
rect 77991 34904 78036 34932
rect 78030 34892 78036 34904
rect 78088 34892 78094 34944
rect 78950 34892 78956 34944
rect 79008 34932 79014 34944
rect 79597 34935 79655 34941
rect 79597 34932 79609 34935
rect 79008 34904 79609 34932
rect 79008 34892 79014 34904
rect 79597 34901 79609 34904
rect 79643 34901 79655 34935
rect 81802 34932 81808 34944
rect 81763 34904 81808 34932
rect 79597 34895 79655 34901
rect 81802 34892 81808 34904
rect 81860 34892 81866 34944
rect 82078 34892 82084 34944
rect 82136 34932 82142 34944
rect 82173 34935 82231 34941
rect 82173 34932 82185 34935
rect 82136 34904 82185 34932
rect 82136 34892 82142 34904
rect 82173 34901 82185 34904
rect 82219 34901 82231 34935
rect 83108 34932 83136 35108
rect 83274 35096 83280 35108
rect 83332 35136 83338 35148
rect 84013 35139 84071 35145
rect 83332 35108 83964 35136
rect 83332 35096 83338 35108
rect 83936 35077 83964 35108
rect 84013 35105 84025 35139
rect 84059 35136 84071 35139
rect 84059 35108 84332 35136
rect 84059 35105 84071 35108
rect 84013 35099 84071 35105
rect 83921 35071 83979 35077
rect 83921 35037 83933 35071
rect 83967 35037 83979 35071
rect 84304 35068 84332 35108
rect 84378 35096 84384 35148
rect 84436 35136 84442 35148
rect 84580 35145 84608 35176
rect 84746 35164 84752 35216
rect 84804 35204 84810 35216
rect 84804 35176 84849 35204
rect 84804 35164 84810 35176
rect 86034 35164 86040 35216
rect 86092 35204 86098 35216
rect 86092 35176 86137 35204
rect 86092 35164 86098 35176
rect 86218 35164 86224 35216
rect 86276 35204 86282 35216
rect 86276 35176 89116 35204
rect 86276 35164 86282 35176
rect 84565 35139 84623 35145
rect 84436 35108 84481 35136
rect 84436 35096 84442 35108
rect 84565 35105 84577 35139
rect 84611 35136 84623 35139
rect 85390 35136 85396 35148
rect 84611 35108 85396 35136
rect 84611 35105 84623 35108
rect 84565 35099 84623 35105
rect 85390 35096 85396 35108
rect 85448 35096 85454 35148
rect 85574 35136 85580 35148
rect 85535 35108 85580 35136
rect 85574 35096 85580 35108
rect 85632 35096 85638 35148
rect 85945 35139 86003 35145
rect 85945 35105 85957 35139
rect 85991 35136 86003 35139
rect 88242 35136 88248 35148
rect 85991 35108 88248 35136
rect 85991 35105 86003 35108
rect 85945 35099 86003 35105
rect 88242 35096 88248 35108
rect 88300 35096 88306 35148
rect 89088 35145 89116 35176
rect 89073 35139 89131 35145
rect 89073 35105 89085 35139
rect 89119 35136 89131 35139
rect 89530 35136 89536 35148
rect 89119 35108 89300 35136
rect 89491 35108 89536 35136
rect 89119 35105 89131 35108
rect 89073 35099 89131 35105
rect 88337 35071 88395 35077
rect 88337 35068 88349 35071
rect 84304 35040 88349 35068
rect 83921 35031 83979 35037
rect 88337 35037 88349 35040
rect 88383 35068 88395 35071
rect 89162 35068 89168 35080
rect 88383 35040 89168 35068
rect 88383 35037 88395 35040
rect 88337 35031 88395 35037
rect 89162 35028 89168 35040
rect 89220 35028 89226 35080
rect 89272 35077 89300 35108
rect 89530 35096 89536 35108
rect 89588 35096 89594 35148
rect 91738 35136 91744 35148
rect 91651 35108 91744 35136
rect 91738 35096 91744 35108
rect 91796 35136 91802 35148
rect 94130 35136 94136 35148
rect 91796 35108 93992 35136
rect 94091 35108 94136 35136
rect 91796 35096 91802 35108
rect 89257 35071 89315 35077
rect 89257 35037 89269 35071
rect 89303 35068 89315 35071
rect 93581 35071 93639 35077
rect 93581 35068 93593 35071
rect 89303 35040 93593 35068
rect 89303 35037 89315 35040
rect 89257 35031 89315 35037
rect 93581 35037 93593 35040
rect 93627 35068 93639 35071
rect 93854 35068 93860 35080
rect 93627 35040 93860 35068
rect 93627 35037 93639 35040
rect 93581 35031 93639 35037
rect 93854 35028 93860 35040
rect 93912 35028 93918 35080
rect 93964 35068 93992 35108
rect 94130 35096 94136 35108
rect 94188 35096 94194 35148
rect 95237 35071 95295 35077
rect 95237 35068 95249 35071
rect 93964 35040 95249 35068
rect 95237 35037 95249 35040
rect 95283 35037 95295 35071
rect 95237 35031 95295 35037
rect 83458 35000 83464 35012
rect 83419 34972 83464 35000
rect 83458 34960 83464 34972
rect 83516 34960 83522 35012
rect 83550 34960 83556 35012
rect 83608 35000 83614 35012
rect 83608 34972 88472 35000
rect 83608 34960 83614 34972
rect 88334 34932 88340 34944
rect 83108 34904 88340 34932
rect 82173 34895 82231 34901
rect 88334 34892 88340 34904
rect 88392 34892 88398 34944
rect 88444 34932 88472 34972
rect 90174 34932 90180 34944
rect 88444 34904 90180 34932
rect 90174 34892 90180 34904
rect 90232 34932 90238 34944
rect 91925 34935 91983 34941
rect 91925 34932 91937 34935
rect 90232 34904 91937 34932
rect 90232 34892 90238 34904
rect 91925 34901 91937 34904
rect 91971 34901 91983 34935
rect 91925 34895 91983 34901
rect 1104 34842 105616 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 65686 34842
rect 65738 34790 65750 34842
rect 65802 34790 65814 34842
rect 65866 34790 65878 34842
rect 65930 34790 96406 34842
rect 96458 34790 96470 34842
rect 96522 34790 96534 34842
rect 96586 34790 96598 34842
rect 96650 34790 105616 34842
rect 1104 34768 105616 34790
rect 4341 34731 4399 34737
rect 4341 34697 4353 34731
rect 4387 34728 4399 34731
rect 4614 34728 4620 34740
rect 4387 34700 4620 34728
rect 4387 34697 4399 34700
rect 4341 34691 4399 34697
rect 4614 34688 4620 34700
rect 4672 34688 4678 34740
rect 11422 34728 11428 34740
rect 11383 34700 11428 34728
rect 11422 34688 11428 34700
rect 11480 34688 11486 34740
rect 13078 34688 13084 34740
rect 13136 34728 13142 34740
rect 13722 34728 13728 34740
rect 13136 34700 13728 34728
rect 13136 34688 13142 34700
rect 13722 34688 13728 34700
rect 13780 34728 13786 34740
rect 14458 34728 14464 34740
rect 13780 34700 14044 34728
rect 14419 34700 14464 34728
rect 13780 34688 13786 34700
rect 14016 34660 14044 34700
rect 14458 34688 14464 34700
rect 14516 34728 14522 34740
rect 15286 34728 15292 34740
rect 14516 34700 15292 34728
rect 14516 34688 14522 34700
rect 15286 34688 15292 34700
rect 15344 34688 15350 34740
rect 18782 34728 18788 34740
rect 18743 34700 18788 34728
rect 18782 34688 18788 34700
rect 18840 34688 18846 34740
rect 19426 34688 19432 34740
rect 19484 34728 19490 34740
rect 21174 34728 21180 34740
rect 19484 34700 21180 34728
rect 19484 34688 19490 34700
rect 21174 34688 21180 34700
rect 21232 34688 21238 34740
rect 21729 34731 21787 34737
rect 21729 34697 21741 34731
rect 21775 34728 21787 34731
rect 22094 34728 22100 34740
rect 21775 34700 22100 34728
rect 21775 34697 21787 34700
rect 21729 34691 21787 34697
rect 22094 34688 22100 34700
rect 22152 34688 22158 34740
rect 22278 34728 22284 34740
rect 22239 34700 22284 34728
rect 22278 34688 22284 34700
rect 22336 34688 22342 34740
rect 24857 34731 24915 34737
rect 24857 34697 24869 34731
rect 24903 34728 24915 34731
rect 35989 34731 36047 34737
rect 24903 34700 35940 34728
rect 24903 34697 24915 34700
rect 24857 34691 24915 34697
rect 14366 34660 14372 34672
rect 14016 34632 14372 34660
rect 14366 34620 14372 34632
rect 14424 34620 14430 34672
rect 22186 34660 22192 34672
rect 14476 34632 22192 34660
rect 2498 34592 2504 34604
rect 2459 34564 2504 34592
rect 2498 34552 2504 34564
rect 2556 34552 2562 34604
rect 2777 34595 2835 34601
rect 2777 34561 2789 34595
rect 2823 34592 2835 34595
rect 3142 34592 3148 34604
rect 2823 34564 3148 34592
rect 2823 34561 2835 34564
rect 2777 34555 2835 34561
rect 3142 34552 3148 34564
rect 3200 34552 3206 34604
rect 10870 34552 10876 34604
rect 10928 34592 10934 34604
rect 14476 34592 14504 34632
rect 22186 34620 22192 34632
rect 22244 34620 22250 34672
rect 23477 34663 23535 34669
rect 23477 34629 23489 34663
rect 23523 34660 23535 34663
rect 24872 34660 24900 34691
rect 23523 34632 24900 34660
rect 23523 34629 23535 34632
rect 23477 34623 23535 34629
rect 25314 34620 25320 34672
rect 25372 34660 25378 34672
rect 30466 34660 30472 34672
rect 25372 34632 30472 34660
rect 25372 34620 25378 34632
rect 30466 34620 30472 34632
rect 30524 34620 30530 34672
rect 30668 34632 33364 34660
rect 10928 34564 14504 34592
rect 10928 34552 10934 34564
rect 17770 34552 17776 34604
rect 17828 34592 17834 34604
rect 20070 34592 20076 34604
rect 17828 34564 20076 34592
rect 17828 34552 17834 34564
rect 20070 34552 20076 34564
rect 20128 34552 20134 34604
rect 20272 34564 20760 34592
rect 5445 34527 5503 34533
rect 5445 34493 5457 34527
rect 5491 34493 5503 34527
rect 5445 34487 5503 34493
rect 5721 34527 5779 34533
rect 5721 34493 5733 34527
rect 5767 34524 5779 34527
rect 5902 34524 5908 34536
rect 5767 34496 5908 34524
rect 5767 34493 5779 34496
rect 5721 34487 5779 34493
rect 4062 34416 4068 34468
rect 4120 34456 4126 34468
rect 5460 34456 5488 34487
rect 5902 34484 5908 34496
rect 5960 34484 5966 34536
rect 6270 34484 6276 34536
rect 6328 34524 6334 34536
rect 6825 34527 6883 34533
rect 6825 34524 6837 34527
rect 6328 34496 6837 34524
rect 6328 34484 6334 34496
rect 6825 34493 6837 34496
rect 6871 34493 6883 34527
rect 7282 34524 7288 34536
rect 7243 34496 7288 34524
rect 6825 34487 6883 34493
rect 7282 34484 7288 34496
rect 7340 34484 7346 34536
rect 11333 34527 11391 34533
rect 11333 34493 11345 34527
rect 11379 34524 11391 34527
rect 11379 34496 13032 34524
rect 11379 34493 11391 34496
rect 11333 34487 11391 34493
rect 5534 34456 5540 34468
rect 4120 34428 5396 34456
rect 5447 34428 5540 34456
rect 4120 34416 4126 34428
rect 3878 34388 3884 34400
rect 3839 34360 3884 34388
rect 3878 34348 3884 34360
rect 3936 34348 3942 34400
rect 5258 34388 5264 34400
rect 5219 34360 5264 34388
rect 5258 34348 5264 34360
rect 5316 34348 5322 34400
rect 5368 34388 5396 34428
rect 5534 34416 5540 34428
rect 5592 34456 5598 34468
rect 6288 34456 6316 34484
rect 12618 34456 12624 34468
rect 5592 34428 6316 34456
rect 6380 34428 12624 34456
rect 5592 34416 5598 34428
rect 6380 34388 6408 34428
rect 12618 34416 12624 34428
rect 12676 34416 12682 34468
rect 6914 34388 6920 34400
rect 5368 34360 6408 34388
rect 6875 34360 6920 34388
rect 6914 34348 6920 34360
rect 6972 34348 6978 34400
rect 13004 34388 13032 34496
rect 13078 34484 13084 34536
rect 13136 34524 13142 34536
rect 13357 34527 13415 34533
rect 13136 34496 13181 34524
rect 13136 34484 13142 34496
rect 13357 34493 13369 34527
rect 13403 34524 13415 34527
rect 13722 34524 13728 34536
rect 13403 34496 13728 34524
rect 13403 34493 13415 34496
rect 13357 34487 13415 34493
rect 13722 34484 13728 34496
rect 13780 34484 13786 34536
rect 14366 34484 14372 34536
rect 14424 34524 14430 34536
rect 14829 34527 14887 34533
rect 14829 34524 14841 34527
rect 14424 34496 14841 34524
rect 14424 34484 14430 34496
rect 14829 34493 14841 34496
rect 14875 34493 14887 34527
rect 14829 34487 14887 34493
rect 16574 34484 16580 34536
rect 16632 34524 16638 34536
rect 16632 34496 17908 34524
rect 16632 34484 16638 34496
rect 17880 34456 17908 34496
rect 17954 34484 17960 34536
rect 18012 34524 18018 34536
rect 18601 34527 18659 34533
rect 18601 34524 18613 34527
rect 18012 34496 18613 34524
rect 18012 34484 18018 34496
rect 18601 34493 18613 34496
rect 18647 34493 18659 34527
rect 18601 34487 18659 34493
rect 18708 34496 19932 34524
rect 18708 34456 18736 34496
rect 17880 34428 18736 34456
rect 19904 34456 19932 34496
rect 19978 34484 19984 34536
rect 20036 34524 20042 34536
rect 20272 34524 20300 34564
rect 20036 34496 20300 34524
rect 20036 34484 20042 34496
rect 20346 34484 20352 34536
rect 20404 34524 20410 34536
rect 20732 34533 20760 34564
rect 23382 34552 23388 34604
rect 23440 34592 23446 34604
rect 26145 34595 26203 34601
rect 23440 34564 24072 34592
rect 23440 34552 23446 34564
rect 20533 34527 20591 34533
rect 20533 34524 20545 34527
rect 20404 34496 20545 34524
rect 20404 34484 20410 34496
rect 20533 34493 20545 34496
rect 20579 34493 20591 34527
rect 20533 34487 20591 34493
rect 20717 34527 20775 34533
rect 20717 34493 20729 34527
rect 20763 34493 20775 34527
rect 21174 34524 21180 34536
rect 21135 34496 21180 34524
rect 20717 34487 20775 34493
rect 21174 34484 21180 34496
rect 21232 34484 21238 34536
rect 21266 34484 21272 34536
rect 21324 34524 21330 34536
rect 23661 34527 23719 34533
rect 23661 34524 23673 34527
rect 21324 34496 21369 34524
rect 23584 34496 23673 34524
rect 21324 34484 21330 34496
rect 23584 34456 23612 34496
rect 23661 34493 23673 34496
rect 23707 34524 23719 34527
rect 24044 34524 24072 34564
rect 26145 34561 26157 34595
rect 26191 34592 26203 34595
rect 30668 34592 30696 34632
rect 32214 34592 32220 34604
rect 26191 34564 30696 34592
rect 30760 34564 31248 34592
rect 32175 34564 32220 34592
rect 26191 34561 26203 34564
rect 26145 34555 26203 34561
rect 30760 34536 30788 34564
rect 24765 34527 24823 34533
rect 24765 34524 24777 34527
rect 23707 34496 23980 34524
rect 24044 34496 24777 34524
rect 23707 34493 23719 34496
rect 23661 34487 23719 34493
rect 19904 34428 23612 34456
rect 23952 34456 23980 34496
rect 24765 34493 24777 34496
rect 24811 34493 24823 34527
rect 24765 34487 24823 34493
rect 26421 34527 26479 34533
rect 26421 34493 26433 34527
rect 26467 34493 26479 34527
rect 26421 34487 26479 34493
rect 24029 34459 24087 34465
rect 24029 34456 24041 34459
rect 23952 34428 24041 34456
rect 24029 34425 24041 34428
rect 24075 34456 24087 34459
rect 26050 34456 26056 34468
rect 24075 34428 26056 34456
rect 24075 34425 24087 34428
rect 24029 34419 24087 34425
rect 26050 34416 26056 34428
rect 26108 34416 26114 34468
rect 26234 34456 26240 34468
rect 26195 34428 26240 34456
rect 26234 34416 26240 34428
rect 26292 34456 26298 34468
rect 26436 34456 26464 34487
rect 26694 34484 26700 34536
rect 26752 34524 26758 34536
rect 30558 34524 30564 34536
rect 26752 34496 30564 34524
rect 26752 34484 26758 34496
rect 30558 34484 30564 34496
rect 30616 34484 30622 34536
rect 30742 34524 30748 34536
rect 30703 34496 30748 34524
rect 30742 34484 30748 34496
rect 30800 34484 30806 34536
rect 30926 34524 30932 34536
rect 30887 34496 30932 34524
rect 30926 34484 30932 34496
rect 30984 34484 30990 34536
rect 31113 34527 31171 34533
rect 31113 34493 31125 34527
rect 31159 34493 31171 34527
rect 31220 34524 31248 34564
rect 32214 34552 32220 34564
rect 32272 34552 32278 34604
rect 32677 34595 32735 34601
rect 32677 34592 32689 34595
rect 32416 34564 32689 34592
rect 31573 34527 31631 34533
rect 31573 34524 31585 34527
rect 31220 34496 31585 34524
rect 31113 34487 31171 34493
rect 31573 34493 31585 34496
rect 31619 34493 31631 34527
rect 31573 34487 31631 34493
rect 31665 34527 31723 34533
rect 31665 34493 31677 34527
rect 31711 34524 31723 34527
rect 32416 34524 32444 34564
rect 32677 34561 32689 34564
rect 32723 34592 32735 34595
rect 32858 34592 32864 34604
rect 32723 34564 32864 34592
rect 32723 34561 32735 34564
rect 32677 34555 32735 34561
rect 32858 34552 32864 34564
rect 32916 34552 32922 34604
rect 33336 34592 33364 34632
rect 33502 34620 33508 34672
rect 33560 34660 33566 34672
rect 35621 34663 35679 34669
rect 35621 34660 35633 34663
rect 33560 34632 35633 34660
rect 33560 34620 33566 34632
rect 35621 34629 35633 34632
rect 35667 34660 35679 34663
rect 35912 34660 35940 34700
rect 35989 34697 36001 34731
rect 36035 34728 36047 34731
rect 36630 34728 36636 34740
rect 36035 34700 36636 34728
rect 36035 34697 36047 34700
rect 35989 34691 36047 34697
rect 36630 34688 36636 34700
rect 36688 34728 36694 34740
rect 36998 34728 37004 34740
rect 36688 34700 37004 34728
rect 36688 34688 36694 34700
rect 36998 34688 37004 34700
rect 37056 34688 37062 34740
rect 37277 34731 37335 34737
rect 37277 34697 37289 34731
rect 37323 34728 37335 34731
rect 38838 34728 38844 34740
rect 37323 34700 38844 34728
rect 37323 34697 37335 34700
rect 37277 34691 37335 34697
rect 38838 34688 38844 34700
rect 38896 34688 38902 34740
rect 39022 34728 39028 34740
rect 38983 34700 39028 34728
rect 39022 34688 39028 34700
rect 39080 34688 39086 34740
rect 39393 34731 39451 34737
rect 39393 34697 39405 34731
rect 39439 34728 39451 34731
rect 39574 34728 39580 34740
rect 39439 34700 39580 34728
rect 39439 34697 39451 34700
rect 39393 34691 39451 34697
rect 39574 34688 39580 34700
rect 39632 34688 39638 34740
rect 39666 34688 39672 34740
rect 39724 34728 39730 34740
rect 41233 34731 41291 34737
rect 41233 34728 41245 34731
rect 39724 34700 41245 34728
rect 39724 34688 39730 34700
rect 41233 34697 41245 34700
rect 41279 34728 41291 34731
rect 41506 34728 41512 34740
rect 41279 34700 41512 34728
rect 41279 34697 41291 34700
rect 41233 34691 41291 34697
rect 41506 34688 41512 34700
rect 41564 34688 41570 34740
rect 41690 34688 41696 34740
rect 41748 34728 41754 34740
rect 42886 34728 42892 34740
rect 41748 34700 42892 34728
rect 41748 34688 41754 34700
rect 42886 34688 42892 34700
rect 42944 34688 42950 34740
rect 42981 34731 43039 34737
rect 42981 34697 42993 34731
rect 43027 34728 43039 34731
rect 43622 34728 43628 34740
rect 43027 34700 43628 34728
rect 43027 34697 43039 34700
rect 42981 34691 43039 34697
rect 43622 34688 43628 34700
rect 43680 34688 43686 34740
rect 81342 34728 81348 34740
rect 43732 34700 81348 34728
rect 42058 34660 42064 34672
rect 35667 34632 35848 34660
rect 35912 34632 42064 34660
rect 35667 34629 35679 34632
rect 35621 34623 35679 34629
rect 33336 34564 33824 34592
rect 31711 34496 32444 34524
rect 32493 34527 32551 34533
rect 31711 34493 31723 34496
rect 31665 34487 31723 34493
rect 32493 34493 32505 34527
rect 32539 34524 32551 34527
rect 33318 34524 33324 34536
rect 32539 34496 33324 34524
rect 32539 34493 32551 34496
rect 32493 34487 32551 34493
rect 26292 34428 26464 34456
rect 26292 34416 26298 34428
rect 13630 34388 13636 34400
rect 13004 34360 13636 34388
rect 13630 34348 13636 34360
rect 13688 34348 13694 34400
rect 19978 34348 19984 34400
rect 20036 34388 20042 34400
rect 20165 34391 20223 34397
rect 20165 34388 20177 34391
rect 20036 34360 20177 34388
rect 20036 34348 20042 34360
rect 20165 34357 20177 34360
rect 20211 34357 20223 34391
rect 20346 34388 20352 34400
rect 20307 34360 20352 34388
rect 20165 34351 20223 34357
rect 20346 34348 20352 34360
rect 20404 34348 20410 34400
rect 21174 34348 21180 34400
rect 21232 34388 21238 34400
rect 22097 34391 22155 34397
rect 22097 34388 22109 34391
rect 21232 34360 22109 34388
rect 21232 34348 21238 34360
rect 22097 34357 22109 34360
rect 22143 34388 22155 34391
rect 23477 34391 23535 34397
rect 23477 34388 23489 34391
rect 22143 34360 23489 34388
rect 22143 34357 22155 34360
rect 22097 34351 22155 34357
rect 23477 34357 23489 34360
rect 23523 34357 23535 34391
rect 23842 34388 23848 34400
rect 23755 34360 23848 34388
rect 23477 34351 23535 34357
rect 23842 34348 23848 34360
rect 23900 34388 23906 34400
rect 26145 34391 26203 34397
rect 26145 34388 26157 34391
rect 23900 34360 26157 34388
rect 23900 34348 23906 34360
rect 26145 34357 26157 34360
rect 26191 34357 26203 34391
rect 26602 34388 26608 34400
rect 26563 34360 26608 34388
rect 26145 34351 26203 34357
rect 26602 34348 26608 34360
rect 26660 34348 26666 34400
rect 31128 34388 31156 34487
rect 32306 34388 32312 34400
rect 31128 34360 32312 34388
rect 32306 34348 32312 34360
rect 32364 34388 32370 34400
rect 32508 34388 32536 34487
rect 33318 34484 33324 34496
rect 33376 34484 33382 34536
rect 33796 34456 33824 34564
rect 35820 34533 35848 34632
rect 42058 34620 42064 34632
rect 42116 34620 42122 34672
rect 43732 34660 43760 34700
rect 81342 34688 81348 34700
rect 81400 34688 81406 34740
rect 81434 34688 81440 34740
rect 81492 34728 81498 34740
rect 81492 34700 88012 34728
rect 81492 34688 81498 34700
rect 49881 34663 49939 34669
rect 49881 34660 49893 34663
rect 42168 34632 43760 34660
rect 44468 34632 49893 34660
rect 42168 34592 42196 34632
rect 37844 34564 38148 34592
rect 35805 34527 35863 34533
rect 35805 34493 35817 34527
rect 35851 34493 35863 34527
rect 37458 34524 37464 34536
rect 37419 34496 37464 34524
rect 35805 34487 35863 34493
rect 37458 34484 37464 34496
rect 37516 34524 37522 34536
rect 37844 34533 37872 34564
rect 37645 34527 37703 34533
rect 37645 34524 37657 34527
rect 37516 34496 37657 34524
rect 37516 34484 37522 34496
rect 37645 34493 37657 34496
rect 37691 34524 37703 34527
rect 37829 34527 37887 34533
rect 37829 34524 37841 34527
rect 37691 34496 37841 34524
rect 37691 34493 37703 34496
rect 37645 34487 37703 34493
rect 37829 34493 37841 34496
rect 37875 34493 37887 34527
rect 38010 34524 38016 34536
rect 37923 34496 38016 34524
rect 37829 34487 37887 34493
rect 38010 34484 38016 34496
rect 38068 34484 38074 34536
rect 38120 34524 38148 34564
rect 38948 34564 42196 34592
rect 38473 34527 38531 34533
rect 38473 34524 38485 34527
rect 38120 34496 38485 34524
rect 38473 34493 38485 34496
rect 38519 34493 38531 34527
rect 38473 34487 38531 34493
rect 38565 34527 38623 34533
rect 38565 34493 38577 34527
rect 38611 34524 38623 34527
rect 38654 34524 38660 34536
rect 38611 34496 38660 34524
rect 38611 34493 38623 34496
rect 38565 34487 38623 34493
rect 37277 34459 37335 34465
rect 37277 34456 37289 34459
rect 33796 34428 37289 34456
rect 37277 34425 37289 34428
rect 37323 34425 37335 34459
rect 38028 34456 38056 34484
rect 38580 34456 38608 34487
rect 38654 34484 38660 34496
rect 38712 34484 38718 34536
rect 38948 34524 38976 34564
rect 42978 34552 42984 34604
rect 43036 34592 43042 34604
rect 44468 34592 44496 34632
rect 49881 34629 49893 34632
rect 49927 34660 49939 34663
rect 52273 34663 52331 34669
rect 52273 34660 52285 34663
rect 49927 34632 52285 34660
rect 49927 34629 49939 34632
rect 49881 34623 49939 34629
rect 52273 34629 52285 34632
rect 52319 34629 52331 34663
rect 52273 34623 52331 34629
rect 52457 34663 52515 34669
rect 52457 34629 52469 34663
rect 52503 34660 52515 34663
rect 52638 34660 52644 34672
rect 52503 34632 52644 34660
rect 52503 34629 52515 34632
rect 52457 34623 52515 34629
rect 43036 34564 44496 34592
rect 43036 34552 43042 34564
rect 44542 34552 44548 34604
rect 44600 34592 44606 34604
rect 51902 34592 51908 34604
rect 44600 34564 51908 34592
rect 44600 34552 44606 34564
rect 51902 34552 51908 34564
rect 51960 34552 51966 34604
rect 38764 34496 38976 34524
rect 38028 34428 38608 34456
rect 37277 34419 37335 34425
rect 32364 34360 32536 34388
rect 32364 34348 32370 34360
rect 37090 34348 37096 34400
rect 37148 34388 37154 34400
rect 38764 34388 38792 34496
rect 40034 34484 40040 34536
rect 40092 34524 40098 34536
rect 40954 34524 40960 34536
rect 40092 34496 40960 34524
rect 40092 34484 40098 34496
rect 40954 34484 40960 34496
rect 41012 34524 41018 34536
rect 41601 34527 41659 34533
rect 41601 34524 41613 34527
rect 41012 34496 41613 34524
rect 41012 34484 41018 34496
rect 41601 34493 41613 34496
rect 41647 34524 41659 34527
rect 41785 34527 41843 34533
rect 41785 34524 41797 34527
rect 41647 34496 41797 34524
rect 41647 34493 41659 34496
rect 41601 34487 41659 34493
rect 41785 34493 41797 34496
rect 41831 34493 41843 34527
rect 41969 34527 42027 34533
rect 41969 34524 41981 34527
rect 41785 34487 41843 34493
rect 41892 34496 41981 34524
rect 41506 34456 41512 34468
rect 41419 34428 41512 34456
rect 41506 34416 41512 34428
rect 41564 34456 41570 34468
rect 41892 34456 41920 34496
rect 41969 34493 41981 34496
rect 42015 34524 42027 34527
rect 42521 34527 42579 34533
rect 42521 34524 42533 34527
rect 42015 34496 42533 34524
rect 42015 34493 42027 34496
rect 41969 34487 42027 34493
rect 42521 34493 42533 34496
rect 42567 34524 42579 34527
rect 42705 34527 42763 34533
rect 42567 34496 42656 34524
rect 42567 34493 42579 34496
rect 42521 34487 42579 34493
rect 41564 34428 41920 34456
rect 42628 34456 42656 34496
rect 42705 34493 42717 34527
rect 42751 34524 42763 34527
rect 43990 34524 43996 34536
rect 42751 34496 43996 34524
rect 42751 34493 42763 34496
rect 42705 34487 42763 34493
rect 43990 34484 43996 34496
rect 44048 34484 44054 34536
rect 51810 34524 51816 34536
rect 44100 34496 51816 34524
rect 44100 34456 44128 34496
rect 51810 34484 51816 34496
rect 51868 34484 51874 34536
rect 52288 34524 52316 34623
rect 52638 34620 52644 34632
rect 52696 34620 52702 34672
rect 59078 34660 59084 34672
rect 56060 34632 59084 34660
rect 53006 34592 53012 34604
rect 52967 34564 53012 34592
rect 53006 34552 53012 34564
rect 53064 34552 53070 34604
rect 53926 34552 53932 34604
rect 53984 34592 53990 34604
rect 55033 34595 55091 34601
rect 55033 34592 55045 34595
rect 53984 34564 55045 34592
rect 53984 34552 53990 34564
rect 55033 34561 55045 34564
rect 55079 34561 55091 34595
rect 56060 34592 56088 34632
rect 59078 34620 59084 34632
rect 59136 34620 59142 34672
rect 59832 34632 64092 34660
rect 55033 34555 55091 34561
rect 55252 34564 56088 34592
rect 52641 34527 52699 34533
rect 52641 34524 52653 34527
rect 52288 34496 52653 34524
rect 52641 34493 52653 34496
rect 52687 34493 52699 34527
rect 52641 34487 52699 34493
rect 52733 34527 52791 34533
rect 52733 34493 52745 34527
rect 52779 34493 52791 34527
rect 54110 34524 54116 34536
rect 52733 34487 52791 34493
rect 53760 34496 54116 34524
rect 42628 34428 44128 34456
rect 48501 34459 48559 34465
rect 41564 34416 41570 34428
rect 48501 34425 48513 34459
rect 48547 34456 48559 34459
rect 48593 34459 48651 34465
rect 48593 34456 48605 34459
rect 48547 34428 48605 34456
rect 48547 34425 48559 34428
rect 48501 34419 48559 34425
rect 48593 34425 48605 34428
rect 48639 34456 48651 34459
rect 52546 34456 52552 34468
rect 48639 34428 52552 34456
rect 48639 34425 48651 34428
rect 48593 34419 48651 34425
rect 52546 34416 52552 34428
rect 52604 34416 52610 34468
rect 37148 34360 38792 34388
rect 37148 34348 37154 34360
rect 49970 34348 49976 34400
rect 50028 34388 50034 34400
rect 52362 34388 52368 34400
rect 50028 34360 52368 34388
rect 50028 34348 50034 34360
rect 52362 34348 52368 34360
rect 52420 34348 52426 34400
rect 52748 34388 52776 34487
rect 53760 34388 53788 34496
rect 54110 34484 54116 34496
rect 54168 34484 54174 34536
rect 54294 34484 54300 34536
rect 54352 34524 54358 34536
rect 54481 34527 54539 34533
rect 54481 34524 54493 34527
rect 54352 34496 54493 34524
rect 54352 34484 54358 34496
rect 54481 34493 54493 34496
rect 54527 34493 54539 34527
rect 54665 34527 54723 34533
rect 54665 34524 54677 34527
rect 54481 34487 54539 34493
rect 54588 34496 54677 34524
rect 54386 34456 54392 34468
rect 54299 34428 54392 34456
rect 54386 34416 54392 34428
rect 54444 34456 54450 34468
rect 54588 34456 54616 34496
rect 54665 34493 54677 34496
rect 54711 34493 54723 34527
rect 54846 34524 54852 34536
rect 54807 34496 54852 34524
rect 54665 34487 54723 34493
rect 54846 34484 54852 34496
rect 54904 34484 54910 34536
rect 54938 34484 54944 34536
rect 54996 34524 55002 34536
rect 55252 34524 55280 34564
rect 56134 34552 56140 34604
rect 56192 34592 56198 34604
rect 56689 34595 56747 34601
rect 56689 34592 56701 34595
rect 56192 34564 56701 34592
rect 56192 34552 56198 34564
rect 56689 34561 56701 34564
rect 56735 34561 56747 34595
rect 56689 34555 56747 34561
rect 56965 34595 57023 34601
rect 56965 34561 56977 34595
rect 57011 34592 57023 34595
rect 58986 34592 58992 34604
rect 57011 34564 57652 34592
rect 58899 34564 58992 34592
rect 57011 34561 57023 34564
rect 56965 34555 57023 34561
rect 55398 34524 55404 34536
rect 54996 34496 55280 34524
rect 55359 34496 55404 34524
rect 54996 34484 55002 34496
rect 55398 34484 55404 34496
rect 55456 34484 55462 34536
rect 56980 34524 57008 34555
rect 56612 34496 57008 34524
rect 57333 34527 57391 34533
rect 55214 34456 55220 34468
rect 54444 34428 54616 34456
rect 55175 34428 55220 34456
rect 54444 34416 54450 34428
rect 55214 34416 55220 34428
rect 55272 34416 55278 34468
rect 52748 34360 53788 34388
rect 54570 34348 54576 34400
rect 54628 34388 54634 34400
rect 56612 34388 56640 34496
rect 57333 34493 57345 34527
rect 57379 34493 57391 34527
rect 57514 34524 57520 34536
rect 57475 34496 57520 34524
rect 57333 34487 57391 34493
rect 56778 34456 56784 34468
rect 56739 34428 56784 34456
rect 56778 34416 56784 34428
rect 56836 34456 56842 34468
rect 57348 34456 57376 34487
rect 57514 34484 57520 34496
rect 57572 34484 57578 34536
rect 57624 34524 57652 34564
rect 58986 34552 58992 34564
rect 59044 34592 59050 34604
rect 59832 34592 59860 34632
rect 59044 34564 59860 34592
rect 59044 34552 59050 34564
rect 57882 34524 57888 34536
rect 57624 34496 57888 34524
rect 57882 34484 57888 34496
rect 57940 34524 57946 34536
rect 57974 34524 57980 34536
rect 57940 34496 57980 34524
rect 57940 34484 57946 34496
rect 57974 34484 57980 34496
rect 58032 34484 58038 34536
rect 58069 34527 58127 34533
rect 58069 34493 58081 34527
rect 58115 34493 58127 34527
rect 58894 34524 58900 34536
rect 58855 34496 58900 34524
rect 58069 34487 58127 34493
rect 56836 34428 57376 34456
rect 56836 34416 56842 34428
rect 54628 34360 56640 34388
rect 56689 34391 56747 34397
rect 54628 34348 54634 34360
rect 56689 34357 56701 34391
rect 56735 34388 56747 34391
rect 57514 34388 57520 34400
rect 56735 34360 57520 34388
rect 56735 34357 56747 34360
rect 56689 34351 56747 34357
rect 57514 34348 57520 34360
rect 57572 34348 57578 34400
rect 58082 34388 58110 34487
rect 58894 34484 58900 34496
rect 58952 34484 58958 34536
rect 59078 34484 59084 34536
rect 59136 34524 59142 34536
rect 62945 34527 63003 34533
rect 62945 34524 62957 34527
rect 59136 34496 62436 34524
rect 59136 34484 59142 34496
rect 58158 34388 58164 34400
rect 58082 34360 58164 34388
rect 58158 34348 58164 34360
rect 58216 34348 58222 34400
rect 58526 34388 58532 34400
rect 58487 34360 58532 34388
rect 58526 34348 58532 34360
rect 58584 34348 58590 34400
rect 62408 34388 62436 34496
rect 62684 34496 62957 34524
rect 62482 34416 62488 34468
rect 62540 34456 62546 34468
rect 62684 34465 62712 34496
rect 62945 34493 62957 34496
rect 62991 34493 63003 34527
rect 63126 34524 63132 34536
rect 63087 34496 63132 34524
rect 62945 34487 63003 34493
rect 62669 34459 62727 34465
rect 62669 34456 62681 34459
rect 62540 34428 62681 34456
rect 62540 34416 62546 34428
rect 62669 34425 62681 34428
rect 62715 34425 62727 34459
rect 62960 34456 62988 34487
rect 63126 34484 63132 34496
rect 63184 34484 63190 34536
rect 63589 34527 63647 34533
rect 63589 34493 63601 34527
rect 63635 34493 63647 34527
rect 63589 34487 63647 34493
rect 63681 34527 63739 34533
rect 63681 34493 63693 34527
rect 63727 34524 63739 34527
rect 63862 34524 63868 34536
rect 63727 34496 63868 34524
rect 63727 34493 63739 34496
rect 63681 34487 63739 34493
rect 63604 34456 63632 34487
rect 63862 34484 63868 34496
rect 63920 34484 63926 34536
rect 62960 34428 63632 34456
rect 64064 34456 64092 34632
rect 65334 34620 65340 34672
rect 65392 34660 65398 34672
rect 65797 34663 65855 34669
rect 65797 34660 65809 34663
rect 65392 34632 65809 34660
rect 65392 34620 65398 34632
rect 65797 34629 65809 34632
rect 65843 34660 65855 34663
rect 65843 34632 65932 34660
rect 65843 34629 65855 34632
rect 65797 34623 65855 34629
rect 65904 34524 65932 34632
rect 66990 34620 66996 34672
rect 67048 34660 67054 34672
rect 75638 34660 75644 34672
rect 67048 34632 75644 34660
rect 67048 34620 67054 34632
rect 75638 34620 75644 34632
rect 75696 34620 75702 34672
rect 77754 34660 77760 34672
rect 77667 34632 77760 34660
rect 77754 34620 77760 34632
rect 77812 34660 77818 34672
rect 78766 34660 78772 34672
rect 77812 34632 78772 34660
rect 77812 34620 77818 34632
rect 78766 34620 78772 34632
rect 78824 34620 78830 34672
rect 79778 34620 79784 34672
rect 79836 34660 79842 34672
rect 79873 34663 79931 34669
rect 79873 34660 79885 34663
rect 79836 34632 79885 34660
rect 79836 34620 79842 34632
rect 79873 34629 79885 34632
rect 79919 34629 79931 34663
rect 79873 34623 79931 34629
rect 81526 34620 81532 34672
rect 81584 34660 81590 34672
rect 82173 34663 82231 34669
rect 82173 34660 82185 34663
rect 81584 34632 82185 34660
rect 81584 34620 81590 34632
rect 82173 34629 82185 34632
rect 82219 34629 82231 34663
rect 82538 34660 82544 34672
rect 82499 34632 82544 34660
rect 82173 34623 82231 34629
rect 82538 34620 82544 34632
rect 82596 34620 82602 34672
rect 85482 34620 85488 34672
rect 85540 34660 85546 34672
rect 85761 34663 85819 34669
rect 85761 34660 85773 34663
rect 85540 34632 85773 34660
rect 85540 34620 85546 34632
rect 85761 34629 85773 34632
rect 85807 34660 85819 34663
rect 86589 34663 86647 34669
rect 86589 34660 86601 34663
rect 85807 34632 86601 34660
rect 85807 34629 85819 34632
rect 85761 34623 85819 34629
rect 86589 34629 86601 34632
rect 86635 34629 86647 34663
rect 86589 34623 86647 34629
rect 87984 34660 88012 34700
rect 88150 34688 88156 34740
rect 88208 34728 88214 34740
rect 89257 34731 89315 34737
rect 89257 34728 89269 34731
rect 88208 34700 89269 34728
rect 88208 34688 88214 34700
rect 89257 34697 89269 34700
rect 89303 34697 89315 34731
rect 91278 34728 91284 34740
rect 91239 34700 91284 34728
rect 89257 34691 89315 34697
rect 91278 34688 91284 34700
rect 91336 34688 91342 34740
rect 88245 34663 88303 34669
rect 88245 34660 88257 34663
rect 87984 34632 88257 34660
rect 66254 34592 66260 34604
rect 66215 34564 66260 34592
rect 66254 34552 66260 34564
rect 66312 34552 66318 34604
rect 66346 34552 66352 34604
rect 66404 34592 66410 34604
rect 75086 34592 75092 34604
rect 66404 34564 75092 34592
rect 66404 34552 66410 34564
rect 75086 34552 75092 34564
rect 75144 34552 75150 34604
rect 76466 34592 76472 34604
rect 75196 34564 76328 34592
rect 76427 34564 76472 34592
rect 65981 34527 66039 34533
rect 65981 34524 65993 34527
rect 65904 34496 65993 34524
rect 65981 34493 65993 34496
rect 66027 34493 66039 34527
rect 75196 34524 75224 34564
rect 76190 34524 76196 34536
rect 65981 34487 66039 34493
rect 66088 34496 75224 34524
rect 76103 34496 76196 34524
rect 66088 34456 66116 34496
rect 76190 34484 76196 34496
rect 76248 34484 76254 34536
rect 76300 34524 76328 34564
rect 76466 34552 76472 34564
rect 76524 34552 76530 34604
rect 78490 34592 78496 34604
rect 76576 34564 78496 34592
rect 76576 34524 76604 34564
rect 78490 34552 78496 34564
rect 78548 34552 78554 34604
rect 78950 34592 78956 34604
rect 78911 34564 78956 34592
rect 78950 34552 78956 34564
rect 79008 34552 79014 34604
rect 81253 34595 81311 34601
rect 81253 34561 81265 34595
rect 81299 34592 81311 34595
rect 81342 34592 81348 34604
rect 81299 34564 81348 34592
rect 81299 34561 81311 34564
rect 81253 34555 81311 34561
rect 81342 34552 81348 34564
rect 81400 34552 81406 34604
rect 81618 34592 81624 34604
rect 81579 34564 81624 34592
rect 81618 34552 81624 34564
rect 81676 34552 81682 34604
rect 81805 34595 81863 34601
rect 81805 34561 81817 34595
rect 81851 34592 81863 34595
rect 83001 34595 83059 34601
rect 83001 34592 83013 34595
rect 81851 34564 83013 34592
rect 81851 34561 81863 34564
rect 81805 34555 81863 34561
rect 83001 34561 83013 34564
rect 83047 34561 83059 34595
rect 83001 34555 83059 34561
rect 84381 34595 84439 34601
rect 84381 34561 84393 34595
rect 84427 34592 84439 34595
rect 84427 34564 86540 34592
rect 84427 34561 84439 34564
rect 84381 34555 84439 34561
rect 76300 34496 76604 34524
rect 77110 34484 77116 34536
rect 77168 34524 77174 34536
rect 77754 34524 77760 34536
rect 77168 34496 77760 34524
rect 77168 34484 77174 34496
rect 77754 34484 77760 34496
rect 77812 34484 77818 34536
rect 78582 34484 78588 34536
rect 78640 34524 78646 34536
rect 78677 34527 78735 34533
rect 78677 34524 78689 34527
rect 78640 34496 78689 34524
rect 78640 34484 78646 34496
rect 78677 34493 78689 34496
rect 78723 34493 78735 34527
rect 78677 34487 78735 34493
rect 78858 34484 78864 34536
rect 78916 34524 78922 34536
rect 79781 34527 79839 34533
rect 79781 34524 79793 34527
rect 78916 34496 79793 34524
rect 78916 34484 78922 34496
rect 79781 34493 79793 34496
rect 79827 34493 79839 34527
rect 79781 34487 79839 34493
rect 80882 34484 80888 34536
rect 80940 34524 80946 34536
rect 80977 34527 81035 34533
rect 80977 34524 80989 34527
rect 80940 34496 80989 34524
rect 80940 34484 80946 34496
rect 80977 34493 80989 34496
rect 81023 34493 81035 34527
rect 81434 34524 81440 34536
rect 81395 34496 81440 34524
rect 80977 34487 81035 34493
rect 81434 34484 81440 34496
rect 81492 34484 81498 34536
rect 81721 34527 81779 34533
rect 81721 34493 81733 34527
rect 81767 34524 81779 34527
rect 82354 34524 82360 34536
rect 81767 34496 82216 34524
rect 82315 34496 82360 34524
rect 81767 34493 81779 34496
rect 81721 34487 81779 34493
rect 64064 34428 66116 34456
rect 62669 34419 62727 34425
rect 74626 34416 74632 34468
rect 74684 34456 74690 34468
rect 76009 34459 76067 34465
rect 76009 34456 76021 34459
rect 74684 34428 76021 34456
rect 74684 34416 74690 34428
rect 76009 34425 76021 34428
rect 76055 34456 76067 34459
rect 76208 34456 76236 34484
rect 78490 34456 78496 34468
rect 76055 34428 76236 34456
rect 77128 34428 78496 34456
rect 76055 34425 76067 34428
rect 76009 34419 76067 34425
rect 64141 34391 64199 34397
rect 64141 34388 64153 34391
rect 62408 34360 64153 34388
rect 64141 34357 64153 34360
rect 64187 34357 64199 34391
rect 64506 34388 64512 34400
rect 64419 34360 64512 34388
rect 64141 34351 64199 34357
rect 64506 34348 64512 34360
rect 64564 34388 64570 34400
rect 64693 34391 64751 34397
rect 64693 34388 64705 34391
rect 64564 34360 64705 34388
rect 64564 34348 64570 34360
rect 64693 34357 64705 34360
rect 64739 34388 64751 34391
rect 65978 34388 65984 34400
rect 64739 34360 65984 34388
rect 64739 34357 64751 34360
rect 64693 34351 64751 34357
rect 65978 34348 65984 34360
rect 66036 34348 66042 34400
rect 67358 34388 67364 34400
rect 67319 34360 67364 34388
rect 67358 34348 67364 34360
rect 67416 34388 67422 34400
rect 77128 34388 77156 34428
rect 78490 34416 78496 34428
rect 78548 34416 78554 34468
rect 78766 34416 78772 34468
rect 78824 34456 78830 34468
rect 81986 34456 81992 34468
rect 78824 34428 78869 34456
rect 81947 34428 81992 34456
rect 78824 34416 78830 34428
rect 81986 34416 81992 34428
rect 82044 34416 82050 34468
rect 82188 34456 82216 34496
rect 82354 34484 82360 34496
rect 82412 34484 82418 34536
rect 82538 34484 82544 34536
rect 82596 34524 82602 34536
rect 82725 34527 82783 34533
rect 82725 34524 82737 34527
rect 82596 34496 82737 34524
rect 82596 34484 82602 34496
rect 82725 34493 82737 34496
rect 82771 34493 82783 34527
rect 83458 34524 83464 34536
rect 82725 34487 82783 34493
rect 82832 34496 83464 34524
rect 82832 34456 82860 34496
rect 83458 34484 83464 34496
rect 83516 34484 83522 34536
rect 85393 34527 85451 34533
rect 85393 34493 85405 34527
rect 85439 34524 85451 34527
rect 85482 34524 85488 34536
rect 85439 34496 85488 34524
rect 85439 34493 85451 34496
rect 85393 34487 85451 34493
rect 85482 34484 85488 34496
rect 85540 34484 85546 34536
rect 86512 34533 86540 34564
rect 87984 34533 88012 34632
rect 88245 34629 88257 34632
rect 88291 34660 88303 34663
rect 88426 34660 88432 34672
rect 88291 34632 88432 34660
rect 88291 34629 88303 34632
rect 88245 34623 88303 34629
rect 88426 34620 88432 34632
rect 88484 34620 88490 34672
rect 88061 34595 88119 34601
rect 88061 34561 88073 34595
rect 88107 34592 88119 34595
rect 88334 34592 88340 34604
rect 88107 34564 88340 34592
rect 88107 34561 88119 34564
rect 88061 34555 88119 34561
rect 88334 34552 88340 34564
rect 88392 34592 88398 34604
rect 88797 34595 88855 34601
rect 88797 34592 88809 34595
rect 88392 34564 88809 34592
rect 88392 34552 88398 34564
rect 88797 34561 88809 34564
rect 88843 34561 88855 34595
rect 88797 34555 88855 34561
rect 86497 34527 86555 34533
rect 86497 34493 86509 34527
rect 86543 34493 86555 34527
rect 86497 34487 86555 34493
rect 87969 34527 88027 34533
rect 87969 34493 87981 34527
rect 88015 34493 88027 34527
rect 87969 34487 88027 34493
rect 88242 34484 88248 34536
rect 88300 34484 88306 34536
rect 88812 34524 88840 34555
rect 88978 34524 88984 34536
rect 88812 34496 88984 34524
rect 88978 34484 88984 34496
rect 89036 34484 89042 34536
rect 89165 34527 89223 34533
rect 89165 34493 89177 34527
rect 89211 34524 89223 34527
rect 90634 34524 90640 34536
rect 89211 34496 90640 34524
rect 89211 34493 89223 34496
rect 89165 34487 89223 34493
rect 90634 34484 90640 34496
rect 90692 34524 90698 34536
rect 91189 34527 91247 34533
rect 91189 34524 91201 34527
rect 90692 34496 91201 34524
rect 90692 34484 90698 34496
rect 91189 34493 91201 34496
rect 91235 34493 91247 34527
rect 91189 34487 91247 34493
rect 82188 34428 82860 34456
rect 88260 34456 88288 34484
rect 91005 34459 91063 34465
rect 91005 34456 91017 34459
rect 88260 34428 88932 34456
rect 85574 34388 85580 34400
rect 67416 34360 77156 34388
rect 85535 34360 85580 34388
rect 67416 34348 67422 34360
rect 85574 34348 85580 34360
rect 85632 34348 85638 34400
rect 88904 34388 88932 34428
rect 89088 34428 91017 34456
rect 89088 34388 89116 34428
rect 91005 34425 91017 34428
rect 91051 34425 91063 34459
rect 91005 34419 91063 34425
rect 88904 34360 89116 34388
rect 1104 34298 105616 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 50326 34298
rect 50378 34246 50390 34298
rect 50442 34246 50454 34298
rect 50506 34246 50518 34298
rect 50570 34246 81046 34298
rect 81098 34246 81110 34298
rect 81162 34246 81174 34298
rect 81226 34246 81238 34298
rect 81290 34246 105616 34298
rect 1104 34224 105616 34246
rect 5077 34187 5135 34193
rect 5077 34153 5089 34187
rect 5123 34184 5135 34187
rect 5534 34184 5540 34196
rect 5123 34156 5540 34184
rect 5123 34153 5135 34156
rect 5077 34147 5135 34153
rect 5534 34144 5540 34156
rect 5592 34144 5598 34196
rect 6086 34184 6092 34196
rect 6047 34156 6092 34184
rect 6086 34144 6092 34156
rect 6144 34144 6150 34196
rect 9766 34144 9772 34196
rect 9824 34184 9830 34196
rect 9861 34187 9919 34193
rect 9861 34184 9873 34187
rect 9824 34156 9873 34184
rect 9824 34144 9830 34156
rect 9861 34153 9873 34156
rect 9907 34153 9919 34187
rect 9861 34147 9919 34153
rect 10137 34187 10195 34193
rect 10137 34153 10149 34187
rect 10183 34184 10195 34187
rect 10226 34184 10232 34196
rect 10183 34156 10232 34184
rect 10183 34153 10195 34156
rect 10137 34147 10195 34153
rect 10226 34144 10232 34156
rect 10284 34144 10290 34196
rect 11514 34184 11520 34196
rect 11475 34156 11520 34184
rect 11514 34144 11520 34156
rect 11572 34144 11578 34196
rect 18046 34184 18052 34196
rect 13556 34156 18052 34184
rect 3786 34076 3792 34128
rect 3844 34116 3850 34128
rect 13556 34116 13584 34156
rect 18046 34144 18052 34156
rect 18104 34144 18110 34196
rect 27522 34144 27528 34196
rect 27580 34184 27586 34196
rect 37277 34187 37335 34193
rect 37277 34184 37289 34187
rect 27580 34156 37289 34184
rect 27580 34144 27586 34156
rect 37277 34153 37289 34156
rect 37323 34153 37335 34187
rect 37277 34147 37335 34153
rect 46845 34187 46903 34193
rect 46845 34153 46857 34187
rect 46891 34184 46903 34187
rect 56042 34184 56048 34196
rect 46891 34156 56048 34184
rect 46891 34153 46903 34156
rect 46845 34147 46903 34153
rect 56042 34144 56048 34156
rect 56100 34144 56106 34196
rect 13722 34116 13728 34128
rect 3844 34088 13584 34116
rect 13683 34088 13728 34116
rect 3844 34076 3850 34088
rect 13722 34076 13728 34088
rect 13780 34076 13786 34128
rect 15654 34076 15660 34128
rect 15712 34116 15718 34128
rect 21174 34116 21180 34128
rect 15712 34088 21180 34116
rect 15712 34076 15718 34088
rect 21174 34076 21180 34088
rect 21232 34076 21238 34128
rect 22741 34119 22799 34125
rect 22741 34085 22753 34119
rect 22787 34116 22799 34119
rect 24302 34116 24308 34128
rect 22787 34088 24308 34116
rect 22787 34085 22799 34088
rect 22741 34079 22799 34085
rect 24302 34076 24308 34088
rect 24360 34076 24366 34128
rect 24394 34076 24400 34128
rect 24452 34116 24458 34128
rect 48774 34116 48780 34128
rect 24452 34088 48780 34116
rect 24452 34076 24458 34088
rect 48774 34076 48780 34088
rect 48832 34076 48838 34128
rect 52362 34076 52368 34128
rect 52420 34116 52426 34128
rect 67358 34116 67364 34128
rect 52420 34088 67364 34116
rect 52420 34076 52426 34088
rect 67358 34076 67364 34088
rect 67416 34076 67422 34128
rect 4798 34008 4804 34060
rect 4856 34048 4862 34060
rect 4893 34051 4951 34057
rect 4893 34048 4905 34051
rect 4856 34020 4905 34048
rect 4856 34008 4862 34020
rect 4893 34017 4905 34020
rect 4939 34048 4951 34051
rect 5442 34048 5448 34060
rect 4939 34020 5448 34048
rect 4939 34017 4951 34020
rect 4893 34011 4951 34017
rect 5442 34008 5448 34020
rect 5500 34008 5506 34060
rect 6270 34048 6276 34060
rect 6231 34020 6276 34048
rect 6270 34008 6276 34020
rect 6328 34008 6334 34060
rect 6546 34048 6552 34060
rect 6507 34020 6552 34048
rect 6546 34008 6552 34020
rect 6604 34008 6610 34060
rect 9766 34008 9772 34060
rect 9824 34048 9830 34060
rect 10045 34051 10103 34057
rect 10045 34048 10057 34051
rect 9824 34020 10057 34048
rect 9824 34008 9830 34020
rect 10045 34017 10057 34020
rect 10091 34048 10103 34051
rect 10134 34048 10140 34060
rect 10091 34020 10140 34048
rect 10091 34017 10103 34020
rect 10045 34011 10103 34017
rect 10134 34008 10140 34020
rect 10192 34008 10198 34060
rect 11333 34051 11391 34057
rect 11333 34017 11345 34051
rect 11379 34048 11391 34051
rect 11974 34048 11980 34060
rect 11379 34020 11980 34048
rect 11379 34017 11391 34020
rect 11333 34011 11391 34017
rect 11974 34008 11980 34020
rect 12032 34008 12038 34060
rect 12621 34051 12679 34057
rect 12621 34017 12633 34051
rect 12667 34048 12679 34051
rect 13170 34048 13176 34060
rect 12667 34020 13176 34048
rect 12667 34017 12679 34020
rect 12621 34011 12679 34017
rect 13170 34008 13176 34020
rect 13228 34008 13234 34060
rect 13357 34051 13415 34057
rect 13357 34017 13369 34051
rect 13403 34048 13415 34051
rect 13906 34048 13912 34060
rect 13403 34020 13912 34048
rect 13403 34017 13415 34020
rect 13357 34011 13415 34017
rect 13906 34008 13912 34020
rect 13964 34008 13970 34060
rect 15286 34048 15292 34060
rect 15247 34020 15292 34048
rect 15286 34008 15292 34020
rect 15344 34008 15350 34060
rect 19613 34051 19671 34057
rect 19613 34017 19625 34051
rect 19659 34048 19671 34051
rect 19705 34051 19763 34057
rect 19705 34048 19717 34051
rect 19659 34020 19717 34048
rect 19659 34017 19671 34020
rect 19613 34011 19671 34017
rect 19705 34017 19717 34020
rect 19751 34048 19763 34051
rect 20162 34048 20168 34060
rect 19751 34020 20168 34048
rect 19751 34017 19763 34020
rect 19705 34011 19763 34017
rect 20162 34008 20168 34020
rect 20220 34008 20226 34060
rect 21450 34008 21456 34060
rect 21508 34048 21514 34060
rect 21508 34020 22048 34048
rect 21508 34008 21514 34020
rect 22020 33992 22048 34020
rect 23106 34008 23112 34060
rect 23164 34048 23170 34060
rect 24765 34051 24823 34057
rect 24765 34048 24777 34051
rect 23164 34020 24777 34048
rect 23164 34008 23170 34020
rect 24765 34017 24777 34020
rect 24811 34017 24823 34051
rect 24765 34011 24823 34017
rect 24857 34051 24915 34057
rect 24857 34017 24869 34051
rect 24903 34048 24915 34051
rect 56410 34048 56416 34060
rect 24903 34020 56416 34048
rect 24903 34017 24915 34020
rect 24857 34011 24915 34017
rect 56410 34008 56416 34020
rect 56468 34008 56474 34060
rect 12342 33980 12348 33992
rect 12255 33952 12348 33980
rect 12342 33940 12348 33952
rect 12400 33980 12406 33992
rect 12437 33983 12495 33989
rect 12437 33980 12449 33983
rect 12400 33952 12449 33980
rect 12400 33940 12406 33952
rect 12437 33949 12449 33952
rect 12483 33949 12495 33983
rect 12437 33943 12495 33949
rect 15838 33940 15844 33992
rect 15896 33980 15902 33992
rect 21085 33983 21143 33989
rect 15896 33952 20576 33980
rect 15896 33940 15902 33952
rect 11882 33872 11888 33924
rect 11940 33912 11946 33924
rect 20438 33912 20444 33924
rect 11940 33884 20444 33912
rect 11940 33872 11946 33884
rect 20438 33872 20444 33884
rect 20496 33872 20502 33924
rect 11238 33804 11244 33856
rect 11296 33844 11302 33856
rect 12710 33844 12716 33856
rect 11296 33816 12716 33844
rect 11296 33804 11302 33816
rect 12710 33804 12716 33816
rect 12768 33804 12774 33856
rect 13906 33844 13912 33856
rect 13867 33816 13912 33844
rect 13906 33804 13912 33816
rect 13964 33844 13970 33856
rect 15381 33847 15439 33853
rect 15381 33844 15393 33847
rect 13964 33816 15393 33844
rect 13964 33804 13970 33816
rect 15381 33813 15393 33816
rect 15427 33813 15439 33847
rect 15381 33807 15439 33813
rect 19889 33847 19947 33853
rect 19889 33813 19901 33847
rect 19935 33844 19947 33847
rect 19978 33844 19984 33856
rect 19935 33816 19984 33844
rect 19935 33813 19947 33816
rect 19889 33807 19947 33813
rect 19978 33804 19984 33816
rect 20036 33804 20042 33856
rect 20548 33844 20576 33952
rect 21085 33949 21097 33983
rect 21131 33980 21143 33983
rect 21266 33980 21272 33992
rect 21131 33952 21272 33980
rect 21131 33949 21143 33952
rect 21085 33943 21143 33949
rect 21266 33940 21272 33952
rect 21324 33940 21330 33992
rect 21358 33940 21364 33992
rect 21416 33980 21422 33992
rect 21416 33952 21461 33980
rect 21416 33940 21422 33952
rect 22002 33940 22008 33992
rect 22060 33980 22066 33992
rect 22925 33983 22983 33989
rect 22925 33980 22937 33983
rect 22060 33952 22937 33980
rect 22060 33940 22066 33952
rect 22925 33949 22937 33952
rect 22971 33980 22983 33983
rect 23658 33980 23664 33992
rect 22971 33952 23664 33980
rect 22971 33949 22983 33952
rect 22925 33943 22983 33949
rect 23658 33940 23664 33952
rect 23716 33940 23722 33992
rect 61746 33980 61752 33992
rect 24780 33952 61752 33980
rect 22462 33872 22468 33924
rect 22520 33912 22526 33924
rect 24394 33912 24400 33924
rect 22520 33884 24400 33912
rect 22520 33872 22526 33884
rect 24394 33872 24400 33884
rect 24452 33872 24458 33924
rect 24780 33912 24808 33952
rect 61746 33940 61752 33952
rect 61804 33940 61810 33992
rect 24504 33884 24808 33912
rect 25041 33915 25099 33921
rect 21726 33844 21732 33856
rect 20548 33816 21732 33844
rect 21726 33804 21732 33816
rect 21784 33804 21790 33856
rect 23198 33804 23204 33856
rect 23256 33844 23262 33856
rect 24504 33844 24532 33884
rect 25041 33881 25053 33915
rect 25087 33912 25099 33915
rect 62482 33912 62488 33924
rect 25087 33884 62488 33912
rect 25087 33881 25099 33884
rect 25041 33875 25099 33881
rect 62482 33872 62488 33884
rect 62540 33872 62546 33924
rect 23256 33816 24532 33844
rect 23256 33804 23262 33816
rect 24578 33804 24584 33856
rect 24636 33844 24642 33856
rect 49970 33844 49976 33856
rect 24636 33816 49976 33844
rect 24636 33804 24642 33816
rect 49970 33804 49976 33816
rect 50028 33804 50034 33856
rect 1104 33754 24656 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 24656 33754
rect 24762 33736 24768 33788
rect 24820 33776 24826 33788
rect 46566 33776 46572 33788
rect 24820 33748 46572 33776
rect 24820 33736 24826 33748
rect 46566 33736 46572 33748
rect 46624 33736 46630 33788
rect 1104 33680 24656 33702
rect 37277 33711 37335 33717
rect 37277 33677 37289 33711
rect 37323 33708 37335 33711
rect 46845 33711 46903 33717
rect 46845 33708 46857 33711
rect 37323 33680 46857 33708
rect 37323 33677 37335 33680
rect 37277 33671 37335 33677
rect 46845 33677 46857 33680
rect 46891 33677 46903 33711
rect 46845 33671 46903 33677
rect 4798 33640 4804 33652
rect 4759 33612 4804 33640
rect 4798 33600 4804 33612
rect 4856 33600 4862 33652
rect 9306 33600 9312 33652
rect 9364 33640 9370 33652
rect 21634 33640 21640 33652
rect 9364 33612 21640 33640
rect 9364 33600 9370 33612
rect 21634 33600 21640 33612
rect 21692 33600 21698 33652
rect 22186 33640 22192 33652
rect 22099 33612 22192 33640
rect 22186 33600 22192 33612
rect 22244 33640 22250 33652
rect 23842 33640 23848 33652
rect 22244 33612 23848 33640
rect 22244 33600 22250 33612
rect 23842 33600 23848 33612
rect 23900 33600 23906 33652
rect 24394 33600 24400 33652
rect 24452 33640 24458 33652
rect 24578 33640 24584 33652
rect 24452 33612 24584 33640
rect 24452 33600 24458 33612
rect 24578 33600 24584 33612
rect 24636 33600 24642 33652
rect 24854 33600 24860 33652
rect 24912 33640 24918 33652
rect 55950 33640 55956 33652
rect 24912 33612 55956 33640
rect 24912 33600 24918 33612
rect 55950 33600 55956 33612
rect 56008 33600 56014 33652
rect 11238 33572 11244 33584
rect 11199 33544 11244 33572
rect 11238 33532 11244 33544
rect 11296 33532 11302 33584
rect 54478 33572 54484 33584
rect 20548 33544 54484 33572
rect 11532 33476 15148 33504
rect 4062 33396 4068 33448
rect 4120 33436 4126 33448
rect 4617 33439 4675 33445
rect 4617 33436 4629 33439
rect 4120 33408 4629 33436
rect 4120 33396 4126 33408
rect 4617 33405 4629 33408
rect 4663 33436 4675 33439
rect 5626 33436 5632 33448
rect 4663 33408 5632 33436
rect 4663 33405 4675 33408
rect 4617 33399 4675 33405
rect 5626 33396 5632 33408
rect 5684 33396 5690 33448
rect 11057 33439 11115 33445
rect 11057 33405 11069 33439
rect 11103 33436 11115 33439
rect 11532 33436 11560 33476
rect 11103 33408 11560 33436
rect 11103 33405 11115 33408
rect 11057 33399 11115 33405
rect 11532 33309 11560 33408
rect 12253 33439 12311 33445
rect 12253 33405 12265 33439
rect 12299 33436 12311 33439
rect 12434 33436 12440 33448
rect 12299 33408 12440 33436
rect 12299 33405 12311 33408
rect 12253 33399 12311 33405
rect 12434 33396 12440 33408
rect 12492 33436 12498 33448
rect 12710 33436 12716 33448
rect 12492 33408 12585 33436
rect 12671 33408 12716 33436
rect 12492 33396 12498 33408
rect 12710 33396 12716 33408
rect 12768 33396 12774 33448
rect 11517 33303 11575 33309
rect 11517 33269 11529 33303
rect 11563 33300 11575 33303
rect 11698 33300 11704 33312
rect 11563 33272 11704 33300
rect 11563 33269 11575 33272
rect 11517 33263 11575 33269
rect 11698 33260 11704 33272
rect 11756 33260 11762 33312
rect 13722 33260 13728 33312
rect 13780 33300 13786 33312
rect 13817 33303 13875 33309
rect 13817 33300 13829 33303
rect 13780 33272 13829 33300
rect 13780 33260 13786 33272
rect 13817 33269 13829 33272
rect 13863 33269 13875 33303
rect 15120 33300 15148 33476
rect 20346 33464 20352 33516
rect 20404 33504 20410 33516
rect 20441 33507 20499 33513
rect 20441 33504 20453 33507
rect 20404 33476 20453 33504
rect 20404 33464 20410 33476
rect 20441 33473 20453 33476
rect 20487 33473 20499 33507
rect 20441 33467 20499 33473
rect 15194 33396 15200 33448
rect 15252 33436 15258 33448
rect 20548 33436 20576 33544
rect 54478 33532 54484 33544
rect 54536 33532 54542 33584
rect 21634 33464 21640 33516
rect 21692 33504 21698 33516
rect 30742 33504 30748 33516
rect 21692 33476 30748 33504
rect 21692 33464 21698 33476
rect 30742 33464 30748 33476
rect 30800 33464 30806 33516
rect 15252 33408 20576 33436
rect 20625 33439 20683 33445
rect 15252 33396 15258 33408
rect 20625 33405 20637 33439
rect 20671 33405 20683 33439
rect 20625 33399 20683 33405
rect 20346 33368 20352 33380
rect 20307 33340 20352 33368
rect 20346 33328 20352 33340
rect 20404 33328 20410 33380
rect 20640 33368 20668 33399
rect 20990 33396 20996 33448
rect 21048 33436 21054 33448
rect 21266 33445 21272 33448
rect 21085 33439 21143 33445
rect 21085 33436 21097 33439
rect 21048 33408 21097 33436
rect 21048 33396 21054 33408
rect 21085 33405 21097 33408
rect 21131 33405 21143 33439
rect 21265 33436 21272 33445
rect 21227 33408 21272 33436
rect 21085 33399 21143 33405
rect 21265 33399 21272 33408
rect 21266 33396 21272 33399
rect 21324 33396 21330 33448
rect 21542 33396 21548 33448
rect 21600 33436 21606 33448
rect 52086 33436 52092 33448
rect 21600 33408 52092 33436
rect 21600 33396 21606 33408
rect 52086 33396 52092 33408
rect 52144 33396 52150 33448
rect 20806 33368 20812 33380
rect 20640 33340 20812 33368
rect 20806 33328 20812 33340
rect 20864 33328 20870 33380
rect 21726 33328 21732 33380
rect 21784 33368 21790 33380
rect 54570 33368 54576 33380
rect 21784 33340 54576 33368
rect 21784 33328 21790 33340
rect 54570 33328 54576 33340
rect 54628 33328 54634 33380
rect 21266 33300 21272 33312
rect 15120 33272 21272 33300
rect 13817 33263 13875 33269
rect 21266 33260 21272 33272
rect 21324 33260 21330 33312
rect 21358 33260 21364 33312
rect 21416 33300 21422 33312
rect 21637 33303 21695 33309
rect 21637 33300 21649 33303
rect 21416 33272 21649 33300
rect 21416 33260 21422 33272
rect 21637 33269 21649 33272
rect 21683 33269 21695 33303
rect 21637 33263 21695 33269
rect 22005 33303 22063 33309
rect 22005 33269 22017 33303
rect 22051 33300 22063 33303
rect 22370 33300 22376 33312
rect 22051 33272 22376 33300
rect 22051 33269 22063 33272
rect 22005 33263 22063 33269
rect 22370 33260 22376 33272
rect 22428 33260 22434 33312
rect 22646 33260 22652 33312
rect 22704 33300 22710 33312
rect 24857 33303 24915 33309
rect 24857 33300 24869 33303
rect 22704 33272 24869 33300
rect 22704 33260 22710 33272
rect 24857 33269 24869 33272
rect 24903 33269 24915 33303
rect 24857 33263 24915 33269
rect 1104 33210 24656 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 24656 33210
rect 1104 33136 24656 33158
rect 3418 33056 3424 33108
rect 3476 33096 3482 33108
rect 6549 33099 6607 33105
rect 6549 33096 6561 33099
rect 3476 33068 6561 33096
rect 3476 33056 3482 33068
rect 6549 33065 6561 33068
rect 6595 33065 6607 33099
rect 6549 33059 6607 33065
rect 7006 33056 7012 33108
rect 7064 33096 7070 33108
rect 40034 33096 40040 33108
rect 7064 33068 40040 33096
rect 7064 33056 7070 33068
rect 40034 33056 40040 33068
rect 40092 33056 40098 33108
rect 52086 33056 52092 33108
rect 52144 33096 52150 33108
rect 54386 33096 54392 33108
rect 52144 33068 54392 33096
rect 52144 33056 52150 33068
rect 54386 33056 54392 33068
rect 54444 33056 54450 33108
rect 11422 32988 11428 33040
rect 11480 33028 11486 33040
rect 11480 33000 12296 33028
rect 11480 32988 11486 33000
rect 3510 32920 3516 32972
rect 3568 32960 3574 32972
rect 4065 32963 4123 32969
rect 4065 32960 4077 32963
rect 3568 32932 4077 32960
rect 3568 32920 3574 32932
rect 4065 32929 4077 32932
rect 4111 32960 4123 32963
rect 4341 32963 4399 32969
rect 4341 32960 4353 32963
rect 4111 32932 4353 32960
rect 4111 32929 4123 32932
rect 4065 32923 4123 32929
rect 4341 32929 4353 32932
rect 4387 32960 4399 32963
rect 4614 32960 4620 32972
rect 4387 32932 4620 32960
rect 4387 32929 4399 32932
rect 4341 32923 4399 32929
rect 4614 32920 4620 32932
rect 4672 32920 4678 32972
rect 5077 32963 5135 32969
rect 5077 32929 5089 32963
rect 5123 32960 5135 32963
rect 5169 32963 5227 32969
rect 5169 32960 5181 32963
rect 5123 32932 5181 32960
rect 5123 32929 5135 32932
rect 5077 32923 5135 32929
rect 5169 32929 5181 32932
rect 5215 32929 5227 32963
rect 5169 32923 5227 32929
rect 5445 32963 5503 32969
rect 5445 32929 5457 32963
rect 5491 32960 5503 32963
rect 6086 32960 6092 32972
rect 5491 32932 6092 32960
rect 5491 32929 5503 32932
rect 5445 32923 5503 32929
rect 6086 32920 6092 32932
rect 6144 32920 6150 32972
rect 11790 32960 11796 32972
rect 11751 32932 11796 32960
rect 11790 32920 11796 32932
rect 11848 32920 11854 32972
rect 12268 32969 12296 33000
rect 12710 32988 12716 33040
rect 12768 33028 12774 33040
rect 12897 33031 12955 33037
rect 12897 33028 12909 33031
rect 12768 33000 12909 33028
rect 12768 32988 12774 33000
rect 12897 32997 12909 33000
rect 12943 32997 12955 33031
rect 12897 32991 12955 32997
rect 13170 32988 13176 33040
rect 13228 33028 13234 33040
rect 13228 33000 17448 33028
rect 13228 32988 13234 33000
rect 12253 32963 12311 32969
rect 12253 32929 12265 32963
rect 12299 32929 12311 32963
rect 12253 32923 12311 32929
rect 12345 32963 12403 32969
rect 12345 32929 12357 32963
rect 12391 32960 12403 32963
rect 12526 32960 12532 32972
rect 12391 32932 12532 32960
rect 12391 32929 12403 32932
rect 12345 32923 12403 32929
rect 12526 32920 12532 32932
rect 12584 32920 12590 32972
rect 13817 32963 13875 32969
rect 13817 32929 13829 32963
rect 13863 32929 13875 32963
rect 15286 32960 15292 32972
rect 15247 32932 15292 32960
rect 13817 32923 13875 32929
rect 11517 32895 11575 32901
rect 11517 32861 11529 32895
rect 11563 32892 11575 32895
rect 11701 32895 11759 32901
rect 11701 32892 11713 32895
rect 11563 32864 11713 32892
rect 11563 32861 11575 32864
rect 11517 32855 11575 32861
rect 11701 32861 11713 32864
rect 11747 32861 11759 32895
rect 11701 32855 11759 32861
rect 3510 32784 3516 32836
rect 3568 32824 3574 32836
rect 3694 32824 3700 32836
rect 3568 32796 3700 32824
rect 3568 32784 3574 32796
rect 3694 32784 3700 32796
rect 3752 32784 3758 32836
rect 2406 32716 2412 32768
rect 2464 32756 2470 32768
rect 4062 32756 4068 32768
rect 2464 32728 4068 32756
rect 2464 32716 2470 32728
rect 4062 32716 4068 32728
rect 4120 32756 4126 32768
rect 4157 32759 4215 32765
rect 4157 32756 4169 32759
rect 4120 32728 4169 32756
rect 4120 32716 4126 32728
rect 4157 32725 4169 32728
rect 4203 32725 4215 32759
rect 4157 32719 4215 32725
rect 4798 32716 4804 32768
rect 4856 32756 4862 32768
rect 5077 32759 5135 32765
rect 5077 32756 5089 32759
rect 4856 32728 5089 32756
rect 4856 32716 4862 32728
rect 5077 32725 5089 32728
rect 5123 32756 5135 32759
rect 7009 32759 7067 32765
rect 7009 32756 7021 32759
rect 5123 32728 7021 32756
rect 5123 32725 5135 32728
rect 5077 32719 5135 32725
rect 7009 32725 7021 32728
rect 7055 32756 7067 32759
rect 8478 32756 8484 32768
rect 7055 32728 8484 32756
rect 7055 32725 7067 32728
rect 7009 32719 7067 32725
rect 8478 32716 8484 32728
rect 8536 32716 8542 32768
rect 11716 32756 11744 32855
rect 11974 32784 11980 32836
rect 12032 32824 12038 32836
rect 13832 32824 13860 32923
rect 15286 32920 15292 32932
rect 15344 32920 15350 32972
rect 17420 32969 17448 33000
rect 17494 32988 17500 33040
rect 17552 33028 17558 33040
rect 17552 33000 18184 33028
rect 17552 32988 17558 33000
rect 17405 32963 17463 32969
rect 17405 32929 17417 32963
rect 17451 32960 17463 32963
rect 17954 32960 17960 32972
rect 17451 32932 17960 32960
rect 17451 32929 17463 32932
rect 17405 32923 17463 32929
rect 17954 32920 17960 32932
rect 18012 32920 18018 32972
rect 18156 32969 18184 33000
rect 18322 32988 18328 33040
rect 18380 33028 18386 33040
rect 23569 33031 23627 33037
rect 18380 33000 19748 33028
rect 18380 32988 18386 33000
rect 18141 32963 18199 32969
rect 18141 32929 18153 32963
rect 18187 32960 18199 32963
rect 18693 32963 18751 32969
rect 18693 32960 18705 32963
rect 18187 32932 18705 32960
rect 18187 32929 18199 32932
rect 18141 32923 18199 32929
rect 18693 32929 18705 32932
rect 18739 32929 18751 32963
rect 19610 32960 19616 32972
rect 19571 32932 19616 32960
rect 18693 32923 18751 32929
rect 17221 32895 17279 32901
rect 17221 32861 17233 32895
rect 17267 32861 17279 32895
rect 18708 32892 18736 32923
rect 19610 32920 19616 32932
rect 19668 32920 19674 32972
rect 19720 32960 19748 33000
rect 23569 32997 23581 33031
rect 23615 33028 23627 33031
rect 24765 33031 24823 33037
rect 24765 33028 24777 33031
rect 23615 33000 24777 33028
rect 23615 32997 23627 33000
rect 23569 32991 23627 32997
rect 24765 32997 24777 33000
rect 24811 33028 24823 33031
rect 30926 33028 30932 33040
rect 24811 33000 30932 33028
rect 24811 32997 24823 33000
rect 24765 32991 24823 32997
rect 30926 32988 30932 33000
rect 30984 32988 30990 33040
rect 37274 32960 37280 32972
rect 19720 32932 37280 32960
rect 37274 32920 37280 32932
rect 37332 32920 37338 32972
rect 19705 32895 19763 32901
rect 19705 32892 19717 32895
rect 18708 32864 19717 32892
rect 17221 32855 17279 32861
rect 19705 32861 19717 32864
rect 19751 32861 19763 32895
rect 19705 32855 19763 32861
rect 12032 32796 13860 32824
rect 14001 32827 14059 32833
rect 12032 32784 12038 32796
rect 14001 32793 14013 32827
rect 14047 32824 14059 32827
rect 14274 32824 14280 32836
rect 14047 32796 14280 32824
rect 14047 32793 14059 32796
rect 14001 32787 14059 32793
rect 14274 32784 14280 32796
rect 14332 32784 14338 32836
rect 14458 32784 14464 32836
rect 14516 32824 14522 32836
rect 17236 32824 17264 32855
rect 14516 32796 17264 32824
rect 19720 32824 19748 32855
rect 21726 32852 21732 32904
rect 21784 32892 21790 32904
rect 21913 32895 21971 32901
rect 21913 32892 21925 32895
rect 21784 32864 21925 32892
rect 21784 32852 21790 32864
rect 21913 32861 21925 32864
rect 21959 32861 21971 32895
rect 22186 32892 22192 32904
rect 22147 32864 22192 32892
rect 21913 32855 21971 32861
rect 22186 32852 22192 32864
rect 22244 32852 22250 32904
rect 25133 32895 25191 32901
rect 25133 32861 25145 32895
rect 25179 32892 25191 32895
rect 31754 32892 31760 32904
rect 25179 32864 31760 32892
rect 25179 32861 25191 32864
rect 25133 32855 25191 32861
rect 31754 32852 31760 32864
rect 31812 32852 31818 32904
rect 25041 32827 25099 32833
rect 19720 32796 21864 32824
rect 14516 32784 14522 32796
rect 12342 32756 12348 32768
rect 11716 32728 12348 32756
rect 12342 32716 12348 32728
rect 12400 32756 12406 32768
rect 13814 32756 13820 32768
rect 12400 32728 13820 32756
rect 12400 32716 12406 32728
rect 13814 32716 13820 32728
rect 13872 32716 13878 32768
rect 15470 32756 15476 32768
rect 15431 32728 15476 32756
rect 15470 32716 15476 32728
rect 15528 32716 15534 32768
rect 17126 32756 17132 32768
rect 17087 32728 17132 32756
rect 17126 32716 17132 32728
rect 17184 32756 17190 32768
rect 17236 32756 17264 32796
rect 17184 32728 17264 32756
rect 17184 32716 17190 32728
rect 18046 32716 18052 32768
rect 18104 32756 18110 32768
rect 18417 32759 18475 32765
rect 18417 32756 18429 32759
rect 18104 32728 18429 32756
rect 18104 32716 18110 32728
rect 18417 32725 18429 32728
rect 18463 32725 18475 32759
rect 18417 32719 18475 32725
rect 19242 32716 19248 32768
rect 19300 32756 19306 32768
rect 19886 32756 19892 32768
rect 19300 32728 19892 32756
rect 19300 32716 19306 32728
rect 19886 32716 19892 32728
rect 19944 32716 19950 32768
rect 21726 32756 21732 32768
rect 21687 32728 21732 32756
rect 21726 32716 21732 32728
rect 21784 32716 21790 32768
rect 21836 32756 21864 32796
rect 23216 32796 23704 32824
rect 23216 32756 23244 32796
rect 21836 32728 23244 32756
rect 23676 32756 23704 32796
rect 25041 32793 25053 32827
rect 25087 32824 25099 32827
rect 34606 32824 34612 32836
rect 25087 32796 34612 32824
rect 25087 32793 25099 32796
rect 25041 32787 25099 32793
rect 34606 32784 34612 32796
rect 34664 32784 34670 32836
rect 37458 32756 37464 32768
rect 23676 32728 37464 32756
rect 37458 32716 37464 32728
rect 37516 32716 37522 32768
rect 37277 32691 37335 32697
rect 1104 32666 24656 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 24656 32666
rect 37277 32657 37289 32691
rect 37323 32688 37335 32691
rect 46845 32691 46903 32697
rect 46845 32688 46857 32691
rect 37323 32660 46857 32688
rect 37323 32657 37335 32660
rect 37277 32651 37335 32657
rect 46845 32657 46857 32660
rect 46891 32657 46903 32691
rect 46845 32651 46903 32657
rect 1104 32592 24656 32614
rect 28350 32580 28356 32632
rect 28408 32620 28414 32632
rect 48958 32620 48964 32632
rect 28408 32592 48964 32620
rect 28408 32580 28414 32592
rect 48958 32580 48964 32592
rect 49016 32580 49022 32632
rect 66162 32552 66168 32564
rect 4540 32524 66168 32552
rect 3694 32444 3700 32496
rect 3752 32484 3758 32496
rect 4540 32484 4568 32524
rect 66162 32512 66168 32524
rect 66220 32512 66226 32564
rect 3752 32456 4568 32484
rect 3752 32444 3758 32456
rect 4614 32444 4620 32496
rect 4672 32484 4678 32496
rect 5350 32484 5356 32496
rect 4672 32456 5356 32484
rect 4672 32444 4678 32456
rect 5350 32444 5356 32456
rect 5408 32444 5414 32496
rect 9769 32487 9827 32493
rect 9769 32453 9781 32487
rect 9815 32484 9827 32487
rect 10597 32487 10655 32493
rect 10597 32484 10609 32487
rect 9815 32456 10609 32484
rect 9815 32453 9827 32456
rect 9769 32447 9827 32453
rect 10597 32453 10609 32456
rect 10643 32484 10655 32487
rect 10643 32456 17264 32484
rect 10643 32453 10655 32456
rect 10597 32447 10655 32453
rect 2866 32376 2872 32428
rect 2924 32376 2930 32428
rect 2961 32419 3019 32425
rect 2961 32385 2973 32419
rect 3007 32416 3019 32419
rect 5810 32416 5816 32428
rect 3007 32388 5816 32416
rect 3007 32385 3019 32388
rect 2961 32379 3019 32385
rect 5810 32376 5816 32388
rect 5868 32376 5874 32428
rect 5902 32376 5908 32428
rect 5960 32416 5966 32428
rect 10318 32416 10324 32428
rect 5960 32388 10324 32416
rect 5960 32376 5966 32388
rect 10318 32376 10324 32388
rect 10376 32376 10382 32428
rect 11790 32376 11796 32428
rect 11848 32416 11854 32428
rect 12526 32416 12532 32428
rect 11848 32388 12532 32416
rect 11848 32376 11854 32388
rect 12526 32376 12532 32388
rect 12584 32376 12590 32428
rect 14093 32419 14151 32425
rect 14093 32385 14105 32419
rect 14139 32416 14151 32419
rect 17236 32416 17264 32456
rect 19886 32444 19892 32496
rect 19944 32484 19950 32496
rect 20441 32487 20499 32493
rect 20441 32484 20453 32487
rect 19944 32456 20453 32484
rect 19944 32444 19950 32456
rect 20441 32453 20453 32456
rect 20487 32484 20499 32487
rect 20806 32484 20812 32496
rect 20487 32456 20668 32484
rect 20767 32456 20812 32484
rect 20487 32453 20499 32456
rect 20441 32447 20499 32453
rect 19610 32416 19616 32428
rect 14139 32388 14504 32416
rect 17236 32388 18552 32416
rect 19571 32388 19616 32416
rect 14139 32385 14151 32388
rect 14093 32379 14151 32385
rect 2685 32351 2743 32357
rect 2685 32317 2697 32351
rect 2731 32317 2743 32351
rect 2884 32348 2912 32376
rect 3694 32348 3700 32360
rect 2884 32320 3700 32348
rect 2685 32311 2743 32317
rect 2700 32212 2728 32311
rect 3694 32308 3700 32320
rect 3752 32308 3758 32360
rect 4062 32308 4068 32360
rect 4120 32348 4126 32360
rect 5169 32351 5227 32357
rect 5169 32348 5181 32351
rect 4120 32320 5181 32348
rect 4120 32308 4126 32320
rect 5169 32317 5181 32320
rect 5215 32348 5227 32351
rect 5442 32348 5448 32360
rect 5215 32320 5448 32348
rect 5215 32317 5227 32320
rect 5169 32311 5227 32317
rect 5442 32308 5448 32320
rect 5500 32308 5506 32360
rect 5629 32351 5687 32357
rect 5629 32317 5641 32351
rect 5675 32317 5687 32351
rect 5629 32311 5687 32317
rect 4525 32283 4583 32289
rect 4525 32280 4537 32283
rect 3620 32252 4537 32280
rect 3620 32212 3648 32252
rect 4525 32249 4537 32252
rect 4571 32280 4583 32283
rect 4798 32280 4804 32292
rect 4571 32252 4804 32280
rect 4571 32249 4583 32252
rect 4525 32243 4583 32249
rect 4798 32240 4804 32252
rect 4856 32240 4862 32292
rect 5644 32280 5672 32311
rect 9674 32308 9680 32360
rect 9732 32348 9738 32360
rect 9953 32351 10011 32357
rect 9732 32320 9777 32348
rect 9732 32308 9738 32320
rect 9953 32317 9965 32351
rect 9999 32348 10011 32351
rect 11238 32348 11244 32360
rect 9999 32320 11244 32348
rect 9999 32317 10011 32320
rect 9953 32311 10011 32317
rect 11238 32308 11244 32320
rect 11296 32308 11302 32360
rect 11974 32308 11980 32360
rect 12032 32348 12038 32360
rect 12437 32351 12495 32357
rect 12437 32348 12449 32351
rect 12032 32320 12449 32348
rect 12032 32308 12038 32320
rect 12437 32317 12449 32320
rect 12483 32317 12495 32351
rect 12544 32348 12572 32376
rect 14476 32360 14504 32388
rect 14369 32351 14427 32357
rect 14369 32348 14381 32351
rect 12544 32320 14381 32348
rect 12437 32311 12495 32317
rect 14369 32317 14381 32320
rect 14415 32317 14427 32351
rect 14369 32311 14427 32317
rect 14458 32308 14464 32360
rect 14516 32348 14522 32360
rect 14921 32351 14979 32357
rect 14516 32320 14561 32348
rect 14516 32308 14522 32320
rect 14921 32317 14933 32351
rect 14967 32317 14979 32351
rect 14921 32311 14979 32317
rect 15105 32351 15163 32357
rect 15105 32317 15117 32351
rect 15151 32348 15163 32351
rect 15749 32351 15807 32357
rect 15749 32348 15761 32351
rect 15151 32320 15761 32348
rect 15151 32317 15163 32320
rect 15105 32311 15163 32317
rect 15749 32317 15761 32320
rect 15795 32348 15807 32351
rect 16942 32348 16948 32360
rect 15795 32320 16948 32348
rect 15795 32317 15807 32320
rect 15749 32311 15807 32317
rect 6089 32283 6147 32289
rect 6089 32280 6101 32283
rect 5644 32252 6101 32280
rect 6089 32249 6101 32252
rect 6135 32280 6147 32283
rect 14734 32280 14740 32292
rect 6135 32252 14740 32280
rect 6135 32249 6147 32252
rect 6089 32243 6147 32249
rect 14734 32240 14740 32252
rect 14792 32240 14798 32292
rect 14936 32280 14964 32311
rect 16942 32308 16948 32320
rect 17000 32308 17006 32360
rect 18138 32348 18144 32360
rect 18099 32320 18144 32348
rect 18138 32308 18144 32320
rect 18196 32308 18202 32360
rect 18411 32351 18469 32357
rect 18411 32348 18423 32351
rect 18248 32320 18423 32348
rect 16390 32280 16396 32292
rect 14936 32252 16396 32280
rect 16390 32240 16396 32252
rect 16448 32240 16454 32292
rect 18046 32240 18052 32292
rect 18104 32280 18110 32292
rect 18248 32280 18276 32320
rect 18411 32317 18423 32320
rect 18457 32317 18469 32351
rect 18524 32348 18552 32388
rect 19610 32376 19616 32388
rect 19668 32376 19674 32428
rect 20640 32357 20668 32456
rect 20806 32444 20812 32456
rect 20864 32444 20870 32496
rect 20898 32444 20904 32496
rect 20956 32484 20962 32496
rect 26881 32487 26939 32493
rect 26881 32484 26893 32487
rect 20956 32456 26893 32484
rect 20956 32444 20962 32456
rect 26881 32453 26893 32456
rect 26927 32453 26939 32487
rect 49602 32484 49608 32496
rect 26881 32447 26939 32453
rect 26988 32456 49608 32484
rect 21542 32376 21548 32428
rect 21600 32416 21606 32428
rect 22649 32419 22707 32425
rect 22649 32416 22661 32419
rect 21600 32388 22661 32416
rect 21600 32376 21606 32388
rect 22649 32385 22661 32388
rect 22695 32416 22707 32419
rect 24673 32419 24731 32425
rect 24673 32416 24685 32419
rect 22695 32388 24685 32416
rect 22695 32385 22707 32388
rect 22649 32379 22707 32385
rect 24673 32385 24685 32388
rect 24719 32385 24731 32419
rect 24673 32379 24731 32385
rect 24854 32376 24860 32428
rect 24912 32416 24918 32428
rect 26988 32416 27016 32456
rect 49602 32444 49608 32456
rect 49660 32444 49666 32496
rect 37277 32419 37335 32425
rect 37277 32416 37289 32419
rect 24912 32388 27016 32416
rect 31864 32388 37289 32416
rect 24912 32376 24918 32388
rect 20625 32351 20683 32357
rect 18524 32320 20484 32348
rect 18411 32311 18469 32317
rect 20456 32280 20484 32320
rect 20625 32317 20637 32351
rect 20671 32317 20683 32351
rect 20625 32311 20683 32317
rect 22557 32351 22615 32357
rect 22557 32317 22569 32351
rect 22603 32348 22615 32351
rect 24765 32351 24823 32357
rect 24765 32348 24777 32351
rect 22603 32320 24777 32348
rect 22603 32317 22615 32320
rect 22557 32311 22615 32317
rect 24765 32317 24777 32320
rect 24811 32317 24823 32351
rect 24765 32311 24823 32317
rect 25961 32351 26019 32357
rect 25961 32317 25973 32351
rect 26007 32348 26019 32351
rect 31864 32348 31892 32388
rect 37277 32385 37289 32388
rect 37323 32385 37335 32419
rect 37277 32379 37335 32385
rect 46845 32419 46903 32425
rect 46845 32385 46857 32419
rect 46891 32416 46903 32419
rect 62574 32416 62580 32428
rect 46891 32388 62580 32416
rect 46891 32385 46903 32388
rect 46845 32379 46903 32385
rect 62574 32376 62580 32388
rect 62632 32376 62638 32428
rect 26007 32320 31892 32348
rect 26007 32317 26019 32320
rect 25961 32311 26019 32317
rect 21818 32280 21824 32292
rect 18104 32252 18276 32280
rect 19076 32252 20392 32280
rect 20456 32252 21824 32280
rect 18104 32240 18110 32252
rect 2700 32184 3648 32212
rect 3878 32172 3884 32224
rect 3936 32212 3942 32224
rect 4065 32215 4123 32221
rect 4065 32212 4077 32215
rect 3936 32184 4077 32212
rect 3936 32172 3942 32184
rect 4065 32181 4077 32184
rect 4111 32181 4123 32215
rect 4065 32175 4123 32181
rect 5445 32215 5503 32221
rect 5445 32181 5457 32215
rect 5491 32212 5503 32215
rect 5534 32212 5540 32224
rect 5491 32184 5540 32212
rect 5491 32181 5503 32184
rect 5445 32175 5503 32181
rect 5534 32172 5540 32184
rect 5592 32172 5598 32224
rect 8570 32172 8576 32224
rect 8628 32212 8634 32224
rect 10137 32215 10195 32221
rect 10137 32212 10149 32215
rect 8628 32184 10149 32212
rect 8628 32172 8634 32184
rect 10137 32181 10149 32184
rect 10183 32181 10195 32215
rect 10137 32175 10195 32181
rect 12621 32215 12679 32221
rect 12621 32181 12633 32215
rect 12667 32212 12679 32215
rect 13170 32212 13176 32224
rect 12667 32184 13176 32212
rect 12667 32181 12679 32184
rect 12621 32175 12679 32181
rect 13170 32172 13176 32184
rect 13228 32172 13234 32224
rect 15381 32215 15439 32221
rect 15381 32181 15393 32215
rect 15427 32212 15439 32215
rect 15470 32212 15476 32224
rect 15427 32184 15476 32212
rect 15427 32181 15439 32184
rect 15381 32175 15439 32181
rect 15470 32172 15476 32184
rect 15528 32172 15534 32224
rect 15562 32172 15568 32224
rect 15620 32212 15626 32224
rect 19076 32212 19104 32252
rect 15620 32184 19104 32212
rect 19981 32215 20039 32221
rect 15620 32172 15626 32184
rect 19981 32181 19993 32215
rect 20027 32212 20039 32215
rect 20254 32212 20260 32224
rect 20027 32184 20260 32212
rect 20027 32181 20039 32184
rect 19981 32175 20039 32181
rect 20254 32172 20260 32184
rect 20312 32172 20318 32224
rect 20364 32212 20392 32252
rect 21818 32240 21824 32252
rect 21876 32240 21882 32292
rect 24949 32283 25007 32289
rect 24949 32249 24961 32283
rect 24995 32280 25007 32283
rect 46750 32280 46756 32292
rect 24995 32252 46756 32280
rect 24995 32249 25007 32252
rect 24949 32243 25007 32249
rect 46750 32240 46756 32252
rect 46808 32240 46814 32292
rect 63678 32212 63684 32224
rect 20364 32184 63684 32212
rect 63678 32172 63684 32184
rect 63736 32172 63742 32224
rect 1104 32122 24656 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 24656 32122
rect 1104 32048 24656 32070
rect 5442 31968 5448 32020
rect 5500 32008 5506 32020
rect 5813 32011 5871 32017
rect 5813 32008 5825 32011
rect 5500 31980 5825 32008
rect 5500 31968 5506 31980
rect 5813 31977 5825 31980
rect 5859 31977 5871 32011
rect 10870 32008 10876 32020
rect 10831 31980 10876 32008
rect 5813 31971 5871 31977
rect 10870 31968 10876 31980
rect 10928 31968 10934 32020
rect 13170 31968 13176 32020
rect 13228 32008 13234 32020
rect 13725 32011 13783 32017
rect 13725 32008 13737 32011
rect 13228 31980 13737 32008
rect 13228 31968 13234 31980
rect 13725 31977 13737 31980
rect 13771 31977 13783 32011
rect 13725 31971 13783 31977
rect 14001 32011 14059 32017
rect 14001 31977 14013 32011
rect 14047 32008 14059 32011
rect 14274 32008 14280 32020
rect 14047 31980 14280 32008
rect 14047 31977 14059 31980
rect 14001 31971 14059 31977
rect 14274 31968 14280 31980
rect 14332 31968 14338 32020
rect 14734 31968 14740 32020
rect 14792 32008 14798 32020
rect 15562 32008 15568 32020
rect 14792 31980 15568 32008
rect 14792 31968 14798 31980
rect 15562 31968 15568 31980
rect 15620 31968 15626 32020
rect 15657 32011 15715 32017
rect 15657 31977 15669 32011
rect 15703 32008 15715 32011
rect 16485 32011 16543 32017
rect 16485 32008 16497 32011
rect 15703 31980 16497 32008
rect 15703 31977 15715 31980
rect 15657 31971 15715 31977
rect 16485 31977 16497 31980
rect 16531 32008 16543 32011
rect 16574 32008 16580 32020
rect 16531 31980 16580 32008
rect 16531 31977 16543 31980
rect 16485 31971 16543 31977
rect 16574 31968 16580 31980
rect 16632 31968 16638 32020
rect 16850 31968 16856 32020
rect 16908 32008 16914 32020
rect 17770 32008 17776 32020
rect 16908 31980 17776 32008
rect 16908 31968 16914 31980
rect 17770 31968 17776 31980
rect 17828 31968 17834 32020
rect 18138 31968 18144 32020
rect 18196 32008 18202 32020
rect 20254 32008 20260 32020
rect 18196 31980 20260 32008
rect 18196 31968 18202 31980
rect 20254 31968 20260 31980
rect 20312 32008 20318 32020
rect 21726 32008 21732 32020
rect 20312 31980 21732 32008
rect 20312 31968 20318 31980
rect 21726 31968 21732 31980
rect 21784 31968 21790 32020
rect 21818 31968 21824 32020
rect 21876 32008 21882 32020
rect 52086 32008 52092 32020
rect 21876 31980 52092 32008
rect 21876 31968 21882 31980
rect 52086 31968 52092 31980
rect 52144 31968 52150 32020
rect 3329 31943 3387 31949
rect 3329 31909 3341 31943
rect 3375 31940 3387 31943
rect 3375 31912 9628 31940
rect 3375 31909 3387 31912
rect 3329 31903 3387 31909
rect 2685 31875 2743 31881
rect 2685 31841 2697 31875
rect 2731 31841 2743 31875
rect 2685 31835 2743 31841
rect 2961 31875 3019 31881
rect 2961 31841 2973 31875
rect 3007 31872 3019 31875
rect 3344 31872 3372 31903
rect 4062 31872 4068 31884
rect 3007 31844 3372 31872
rect 3975 31844 4068 31872
rect 3007 31841 3019 31844
rect 2961 31835 3019 31841
rect 2700 31736 2728 31835
rect 3142 31804 3148 31816
rect 3103 31776 3148 31804
rect 3142 31764 3148 31776
rect 3200 31764 3206 31816
rect 3786 31736 3792 31748
rect 2700 31708 3792 31736
rect 3786 31696 3792 31708
rect 3844 31736 3850 31748
rect 3988 31736 4016 31844
rect 4062 31832 4068 31844
rect 4120 31832 4126 31884
rect 4617 31875 4675 31881
rect 4617 31841 4629 31875
rect 4663 31841 4675 31875
rect 4617 31835 4675 31841
rect 4801 31875 4859 31881
rect 4801 31841 4813 31875
rect 4847 31872 4859 31875
rect 4982 31872 4988 31884
rect 4847 31844 4988 31872
rect 4847 31841 4859 31844
rect 4801 31835 4859 31841
rect 4632 31804 4660 31835
rect 4982 31832 4988 31844
rect 5040 31832 5046 31884
rect 5626 31872 5632 31884
rect 5587 31844 5632 31872
rect 5626 31832 5632 31844
rect 5684 31832 5690 31884
rect 8570 31872 8576 31884
rect 8531 31844 8576 31872
rect 8570 31832 8576 31844
rect 8628 31832 8634 31884
rect 9600 31872 9628 31912
rect 9674 31900 9680 31952
rect 9732 31940 9738 31952
rect 9732 31912 9777 31940
rect 9732 31900 9738 31912
rect 9950 31900 9956 31952
rect 10008 31940 10014 31952
rect 21634 31940 21640 31952
rect 10008 31912 21640 31940
rect 10008 31900 10014 31912
rect 21634 31900 21640 31912
rect 21692 31900 21698 31952
rect 10226 31872 10232 31884
rect 9600 31844 9904 31872
rect 10187 31844 10232 31872
rect 4893 31807 4951 31813
rect 4893 31804 4905 31807
rect 4632 31776 4905 31804
rect 4893 31773 4905 31776
rect 4939 31804 4951 31807
rect 8386 31804 8392 31816
rect 4939 31776 8392 31804
rect 4939 31773 4951 31776
rect 4893 31767 4951 31773
rect 8386 31764 8392 31776
rect 8444 31764 8450 31816
rect 3844 31708 4016 31736
rect 3844 31696 3850 31708
rect 4614 31696 4620 31748
rect 4672 31736 4678 31748
rect 9876 31736 9904 31844
rect 10226 31832 10232 31844
rect 10284 31832 10290 31884
rect 10505 31875 10563 31881
rect 10505 31841 10517 31875
rect 10551 31872 10563 31875
rect 10870 31872 10876 31884
rect 10551 31844 10876 31872
rect 10551 31841 10563 31844
rect 10505 31835 10563 31841
rect 10870 31832 10876 31844
rect 10928 31832 10934 31884
rect 13541 31875 13599 31881
rect 13541 31841 13553 31875
rect 13587 31872 13599 31875
rect 14274 31872 14280 31884
rect 13587 31844 14280 31872
rect 13587 31841 13599 31844
rect 13541 31835 13599 31841
rect 14274 31832 14280 31844
rect 14332 31832 14338 31884
rect 15286 31832 15292 31884
rect 15344 31872 15350 31884
rect 15470 31872 15476 31884
rect 15344 31844 15476 31872
rect 15344 31832 15350 31844
rect 15470 31832 15476 31844
rect 15528 31832 15534 31884
rect 16574 31832 16580 31884
rect 16632 31872 16638 31884
rect 17678 31872 17684 31884
rect 16632 31844 16677 31872
rect 17639 31844 17684 31872
rect 16632 31832 16638 31844
rect 17678 31832 17684 31844
rect 17736 31832 17742 31884
rect 21744 31872 21772 31968
rect 35618 31940 35624 31952
rect 22848 31912 35624 31940
rect 21913 31875 21971 31881
rect 21913 31872 21925 31875
rect 17788 31844 21036 31872
rect 21744 31844 21925 31872
rect 10318 31764 10324 31816
rect 10376 31804 10382 31816
rect 10689 31807 10747 31813
rect 10689 31804 10701 31807
rect 10376 31776 10701 31804
rect 10376 31764 10382 31776
rect 10689 31773 10701 31776
rect 10735 31773 10747 31807
rect 10689 31767 10747 31773
rect 15381 31807 15439 31813
rect 15381 31773 15393 31807
rect 15427 31804 15439 31807
rect 17034 31804 17040 31816
rect 15427 31776 17040 31804
rect 15427 31773 15439 31776
rect 15381 31767 15439 31773
rect 17034 31764 17040 31776
rect 17092 31764 17098 31816
rect 17788 31736 17816 31844
rect 17862 31764 17868 31816
rect 17920 31804 17926 31816
rect 18049 31807 18107 31813
rect 18049 31804 18061 31807
rect 17920 31776 18061 31804
rect 17920 31764 17926 31776
rect 18049 31773 18061 31776
rect 18095 31804 18107 31807
rect 20898 31804 20904 31816
rect 18095 31776 20904 31804
rect 18095 31773 18107 31776
rect 18049 31767 18107 31773
rect 20898 31764 20904 31776
rect 20956 31764 20962 31816
rect 21008 31804 21036 31844
rect 21913 31841 21925 31844
rect 21959 31841 21971 31875
rect 21913 31835 21971 31841
rect 22002 31832 22008 31884
rect 22060 31872 22066 31884
rect 22189 31875 22247 31881
rect 22189 31872 22201 31875
rect 22060 31844 22201 31872
rect 22060 31832 22066 31844
rect 22189 31841 22201 31844
rect 22235 31841 22247 31875
rect 22189 31835 22247 31841
rect 22278 31832 22284 31884
rect 22336 31872 22342 31884
rect 22848 31872 22876 31912
rect 35618 31900 35624 31912
rect 35676 31900 35682 31952
rect 22336 31844 22876 31872
rect 22336 31832 22342 31844
rect 23014 31832 23020 31884
rect 23072 31872 23078 31884
rect 25041 31875 25099 31881
rect 25041 31872 25053 31875
rect 23072 31844 25053 31872
rect 23072 31832 23078 31844
rect 25041 31841 25053 31844
rect 25087 31841 25099 31875
rect 25041 31835 25099 31841
rect 26881 31875 26939 31881
rect 26881 31841 26893 31875
rect 26927 31872 26939 31875
rect 51534 31872 51540 31884
rect 26927 31844 51540 31872
rect 26927 31841 26939 31844
rect 26881 31835 26939 31841
rect 51534 31832 51540 31844
rect 51592 31832 51598 31884
rect 55306 31804 55312 31816
rect 21008 31776 55312 31804
rect 55306 31764 55312 31776
rect 55364 31764 55370 31816
rect 62666 31736 62672 31748
rect 4672 31708 9812 31736
rect 9876 31708 17816 31736
rect 23216 31708 62672 31736
rect 4672 31696 4678 31708
rect 8662 31668 8668 31680
rect 8623 31640 8668 31668
rect 8662 31628 8668 31640
rect 8720 31628 8726 31680
rect 9784 31668 9812 31708
rect 15381 31671 15439 31677
rect 15381 31668 15393 31671
rect 9784 31640 15393 31668
rect 15381 31637 15393 31640
rect 15427 31637 15439 31671
rect 15381 31631 15439 31637
rect 16390 31628 16396 31680
rect 16448 31668 16454 31680
rect 16761 31671 16819 31677
rect 16761 31668 16773 31671
rect 16448 31640 16773 31668
rect 16448 31628 16454 31640
rect 16761 31637 16773 31640
rect 16807 31637 16819 31671
rect 16761 31631 16819 31637
rect 17034 31628 17040 31680
rect 17092 31668 17098 31680
rect 23216 31668 23244 31708
rect 62666 31696 62672 31708
rect 62724 31696 62730 31748
rect 81434 31696 81440 31748
rect 81492 31736 81498 31748
rect 81710 31736 81716 31748
rect 81492 31708 81716 31736
rect 81492 31696 81498 31708
rect 81710 31696 81716 31708
rect 81768 31696 81774 31748
rect 17092 31640 23244 31668
rect 17092 31628 17098 31640
rect 23290 31628 23296 31680
rect 23348 31668 23354 31680
rect 23477 31671 23535 31677
rect 23477 31668 23489 31671
rect 23348 31640 23489 31668
rect 23348 31628 23354 31640
rect 23477 31637 23489 31640
rect 23523 31668 23535 31671
rect 25133 31671 25191 31677
rect 25133 31668 25145 31671
rect 23523 31640 25145 31668
rect 23523 31637 23535 31640
rect 23477 31631 23535 31637
rect 25133 31637 25145 31640
rect 25179 31637 25191 31671
rect 51074 31668 51080 31680
rect 25133 31631 25191 31637
rect 43364 31640 51080 31668
rect 43364 31600 43392 31640
rect 51074 31628 51080 31640
rect 51132 31628 51138 31680
rect 54846 31668 54852 31680
rect 51184 31640 54852 31668
rect 51184 31600 51212 31640
rect 54846 31628 54852 31640
rect 54904 31628 54910 31680
rect 1104 31578 24656 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 24656 31578
rect 1104 31504 24656 31526
rect 26896 31572 43392 31600
rect 43456 31572 51212 31600
rect 4433 31467 4491 31473
rect 4433 31433 4445 31467
rect 4479 31464 4491 31467
rect 4614 31464 4620 31476
rect 4479 31436 4620 31464
rect 4479 31433 4491 31436
rect 4433 31427 4491 31433
rect 4614 31424 4620 31436
rect 4672 31424 4678 31476
rect 5997 31467 6055 31473
rect 5997 31433 6009 31467
rect 6043 31464 6055 31467
rect 11698 31464 11704 31476
rect 6043 31436 11560 31464
rect 11659 31436 11704 31464
rect 6043 31433 6055 31436
rect 5997 31427 6055 31433
rect 3804 31300 5120 31328
rect 3804 31272 3832 31300
rect 2406 31260 2412 31272
rect 2367 31232 2412 31260
rect 2406 31220 2412 31232
rect 2464 31220 2470 31272
rect 3786 31260 3792 31272
rect 3747 31232 3792 31260
rect 3786 31220 3792 31232
rect 3844 31220 3850 31272
rect 4065 31263 4123 31269
rect 4065 31229 4077 31263
rect 4111 31260 4123 31263
rect 4614 31260 4620 31272
rect 4111 31232 4620 31260
rect 4111 31229 4123 31232
rect 4065 31223 4123 31229
rect 4614 31220 4620 31232
rect 4672 31220 4678 31272
rect 5092 31269 5120 31300
rect 5077 31263 5135 31269
rect 5077 31229 5089 31263
rect 5123 31229 5135 31263
rect 5077 31223 5135 31229
rect 5629 31263 5687 31269
rect 5629 31229 5641 31263
rect 5675 31260 5687 31263
rect 6012 31260 6040 31427
rect 8662 31288 8668 31340
rect 8720 31328 8726 31340
rect 8757 31331 8815 31337
rect 8757 31328 8769 31331
rect 8720 31300 8769 31328
rect 8720 31288 8726 31300
rect 8757 31297 8769 31300
rect 8803 31297 8815 31331
rect 11532 31328 11560 31436
rect 11698 31424 11704 31436
rect 11756 31424 11762 31476
rect 11790 31424 11796 31476
rect 11848 31464 11854 31476
rect 26896 31464 26924 31572
rect 26970 31492 26976 31544
rect 27028 31532 27034 31544
rect 43456 31532 43484 31572
rect 51994 31560 52000 31612
rect 52052 31600 52058 31612
rect 55214 31600 55220 31612
rect 52052 31572 55220 31600
rect 52052 31560 52058 31572
rect 55214 31560 55220 31572
rect 55272 31560 55278 31612
rect 54294 31532 54300 31544
rect 27028 31504 43484 31532
rect 52288 31504 54300 31532
rect 27028 31492 27034 31504
rect 11848 31436 26924 31464
rect 11848 31424 11854 31436
rect 16942 31396 16948 31408
rect 16855 31368 16948 31396
rect 16942 31356 16948 31368
rect 17000 31396 17006 31408
rect 18322 31396 18328 31408
rect 17000 31368 18328 31396
rect 17000 31356 17006 31368
rect 18322 31356 18328 31368
rect 18380 31356 18386 31408
rect 21542 31396 21548 31408
rect 20364 31368 21548 31396
rect 14645 31331 14703 31337
rect 11532 31300 14504 31328
rect 8757 31291 8815 31297
rect 8478 31260 8484 31272
rect 5675 31232 6040 31260
rect 8391 31232 8484 31260
rect 5675 31229 5687 31232
rect 5629 31223 5687 31229
rect 8478 31220 8484 31232
rect 8536 31220 8542 31272
rect 9858 31220 9864 31272
rect 9916 31260 9922 31272
rect 10229 31263 10287 31269
rect 10229 31260 10241 31263
rect 9916 31232 10241 31260
rect 9916 31220 9922 31232
rect 10229 31229 10241 31232
rect 10275 31229 10287 31263
rect 10229 31223 10287 31229
rect 11149 31263 11207 31269
rect 11149 31229 11161 31263
rect 11195 31260 11207 31263
rect 11698 31260 11704 31272
rect 11195 31232 11704 31260
rect 11195 31229 11207 31232
rect 11149 31223 11207 31229
rect 11698 31220 11704 31232
rect 11756 31220 11762 31272
rect 14366 31260 14372 31272
rect 14327 31232 14372 31260
rect 14366 31220 14372 31232
rect 14424 31220 14430 31272
rect 14476 31260 14504 31300
rect 14645 31297 14657 31331
rect 14691 31328 14703 31331
rect 15378 31328 15384 31340
rect 14691 31300 15384 31328
rect 14691 31297 14703 31300
rect 14645 31291 14703 31297
rect 15378 31288 15384 31300
rect 15436 31288 15442 31340
rect 20070 31288 20076 31340
rect 20128 31328 20134 31340
rect 20364 31328 20392 31368
rect 21542 31356 21548 31368
rect 21600 31356 21606 31408
rect 22649 31399 22707 31405
rect 22649 31365 22661 31399
rect 22695 31396 22707 31399
rect 22738 31396 22744 31408
rect 22695 31368 22744 31396
rect 22695 31365 22707 31368
rect 22649 31359 22707 31365
rect 22738 31356 22744 31368
rect 22796 31356 22802 31408
rect 22925 31399 22983 31405
rect 22925 31365 22937 31399
rect 22971 31396 22983 31399
rect 23290 31396 23296 31408
rect 22971 31368 23296 31396
rect 22971 31365 22983 31368
rect 22925 31359 22983 31365
rect 22940 31328 22968 31359
rect 23290 31356 23296 31368
rect 23348 31356 23354 31408
rect 23382 31356 23388 31408
rect 23440 31396 23446 31408
rect 52288 31396 52316 31504
rect 54294 31492 54300 31504
rect 54352 31492 54358 31544
rect 53834 31424 53840 31476
rect 53892 31464 53898 31476
rect 54110 31464 54116 31476
rect 53892 31436 54116 31464
rect 53892 31424 53898 31436
rect 54110 31424 54116 31436
rect 54168 31424 54174 31476
rect 23440 31368 52316 31396
rect 23440 31356 23446 31368
rect 52362 31356 52368 31408
rect 52420 31396 52426 31408
rect 55398 31396 55404 31408
rect 52420 31368 55404 31396
rect 52420 31356 52426 31368
rect 55398 31356 55404 31368
rect 55456 31356 55462 31408
rect 20128 31300 20392 31328
rect 20128 31288 20134 31300
rect 14476 31232 15332 31260
rect 2593 31127 2651 31133
rect 2593 31093 2605 31127
rect 2639 31124 2651 31127
rect 2682 31124 2688 31136
rect 2639 31096 2688 31124
rect 2639 31093 2651 31096
rect 2593 31087 2651 31093
rect 2682 31084 2688 31096
rect 2740 31084 2746 31136
rect 3786 31124 3792 31136
rect 3747 31096 3792 31124
rect 3786 31084 3792 31096
rect 3844 31084 3850 31136
rect 4798 31084 4804 31136
rect 4856 31124 4862 31136
rect 5169 31127 5227 31133
rect 5169 31124 5181 31127
rect 4856 31096 5181 31124
rect 4856 31084 4862 31096
rect 5169 31093 5181 31096
rect 5215 31093 5227 31127
rect 8496 31124 8524 31220
rect 10134 31192 10140 31204
rect 10095 31164 10140 31192
rect 10134 31152 10140 31164
rect 10192 31152 10198 31204
rect 10962 31192 10968 31204
rect 10923 31164 10968 31192
rect 10962 31152 10968 31164
rect 11020 31152 11026 31204
rect 11517 31195 11575 31201
rect 11517 31161 11529 31195
rect 11563 31192 11575 31195
rect 11790 31192 11796 31204
rect 11563 31164 11796 31192
rect 11563 31161 11575 31164
rect 11517 31155 11575 31161
rect 11790 31152 11796 31164
rect 11848 31152 11854 31204
rect 15304 31192 15332 31232
rect 16022 31220 16028 31272
rect 16080 31260 16086 31272
rect 16853 31263 16911 31269
rect 16853 31260 16865 31263
rect 16080 31232 16865 31260
rect 16080 31220 16086 31232
rect 16853 31229 16865 31232
rect 16899 31229 16911 31263
rect 16853 31223 16911 31229
rect 19705 31263 19763 31269
rect 19705 31229 19717 31263
rect 19751 31260 19763 31263
rect 19981 31263 20039 31269
rect 19981 31260 19993 31263
rect 19751 31232 19993 31260
rect 19751 31229 19763 31232
rect 19705 31223 19763 31229
rect 19981 31229 19993 31232
rect 20027 31229 20039 31263
rect 20162 31260 20168 31272
rect 20123 31232 20168 31260
rect 19981 31223 20039 31229
rect 20162 31220 20168 31232
rect 20220 31220 20226 31272
rect 20364 31260 20392 31300
rect 22572 31300 22968 31328
rect 24765 31331 24823 31337
rect 22572 31272 22600 31300
rect 24765 31297 24777 31331
rect 24811 31328 24823 31331
rect 53834 31328 53840 31340
rect 24811 31300 53840 31328
rect 24811 31297 24823 31300
rect 24765 31291 24823 31297
rect 53834 31288 53840 31300
rect 53892 31328 53898 31340
rect 54018 31328 54024 31340
rect 53892 31300 54024 31328
rect 53892 31288 53898 31300
rect 54018 31288 54024 31300
rect 54076 31288 54082 31340
rect 20625 31263 20683 31269
rect 20625 31260 20637 31263
rect 20364 31232 20637 31260
rect 20625 31229 20637 31232
rect 20671 31229 20683 31263
rect 20625 31223 20683 31229
rect 20714 31220 20720 31272
rect 20772 31260 20778 31272
rect 22554 31260 22560 31272
rect 20772 31232 20817 31260
rect 21192 31232 21864 31260
rect 22467 31232 22560 31260
rect 20772 31220 20778 31232
rect 21192 31192 21220 31232
rect 15304 31164 21220 31192
rect 21269 31195 21327 31201
rect 21269 31161 21281 31195
rect 21315 31192 21327 31195
rect 21836 31192 21864 31232
rect 22554 31220 22560 31232
rect 22612 31220 22618 31272
rect 43438 31260 43444 31272
rect 22756 31232 43444 31260
rect 22756 31192 22784 31232
rect 43438 31220 43444 31232
rect 43496 31220 43502 31272
rect 56778 31220 56784 31272
rect 56836 31220 56842 31272
rect 21315 31164 21680 31192
rect 21836 31164 22784 31192
rect 41417 31195 41475 31201
rect 21315 31161 21327 31164
rect 21269 31155 21327 31161
rect 9858 31124 9864 31136
rect 8496 31096 9864 31124
rect 5169 31087 5227 31093
rect 9858 31084 9864 31096
rect 9916 31084 9922 31136
rect 15286 31084 15292 31136
rect 15344 31124 15350 31136
rect 15749 31127 15807 31133
rect 15749 31124 15761 31127
rect 15344 31096 15761 31124
rect 15344 31084 15350 31096
rect 15749 31093 15761 31096
rect 15795 31124 15807 31127
rect 16022 31124 16028 31136
rect 15795 31096 16028 31124
rect 15795 31093 15807 31096
rect 15749 31087 15807 31093
rect 16022 31084 16028 31096
rect 16080 31084 16086 31136
rect 16206 31124 16212 31136
rect 16167 31096 16212 31124
rect 16206 31084 16212 31096
rect 16264 31084 16270 31136
rect 19705 31127 19763 31133
rect 19705 31093 19717 31127
rect 19751 31124 19763 31127
rect 19889 31127 19947 31133
rect 19889 31124 19901 31127
rect 19751 31096 19901 31124
rect 19751 31093 19763 31096
rect 19705 31087 19763 31093
rect 19889 31093 19901 31096
rect 19935 31124 19947 31127
rect 20990 31124 20996 31136
rect 19935 31096 20996 31124
rect 19935 31093 19947 31096
rect 19889 31087 19947 31093
rect 20990 31084 20996 31096
rect 21048 31084 21054 31136
rect 21652 31124 21680 31164
rect 41417 31161 41429 31195
rect 41463 31192 41475 31195
rect 56796 31192 56824 31220
rect 41463 31164 56824 31192
rect 41463 31161 41475 31164
rect 41417 31155 41475 31161
rect 22186 31124 22192 31136
rect 21652 31096 22192 31124
rect 22186 31084 22192 31096
rect 22244 31084 22250 31136
rect 41325 31127 41383 31133
rect 41325 31124 41337 31127
rect 24688 31096 41337 31124
rect 1104 31034 24656 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 24656 31034
rect 1104 30960 24656 30982
rect 3418 30880 3424 30932
rect 3476 30920 3482 30932
rect 4157 30923 4215 30929
rect 4157 30920 4169 30923
rect 3476 30892 4169 30920
rect 3476 30880 3482 30892
rect 4157 30889 4169 30892
rect 4203 30889 4215 30923
rect 4157 30883 4215 30889
rect 4985 30923 5043 30929
rect 4985 30889 4997 30923
rect 5031 30920 5043 30923
rect 5074 30920 5080 30932
rect 5031 30892 5080 30920
rect 5031 30889 5043 30892
rect 4985 30883 5043 30889
rect 4062 30784 4068 30796
rect 4023 30756 4068 30784
rect 4062 30744 4068 30756
rect 4120 30744 4126 30796
rect 4617 30787 4675 30793
rect 4617 30753 4629 30787
rect 4663 30784 4675 30787
rect 5000 30784 5028 30883
rect 5074 30880 5080 30892
rect 5132 30880 5138 30932
rect 14277 30923 14335 30929
rect 14277 30889 14289 30923
rect 14323 30920 14335 30923
rect 15470 30920 15476 30932
rect 14323 30892 15476 30920
rect 14323 30889 14335 30892
rect 14277 30883 14335 30889
rect 15470 30880 15476 30892
rect 15528 30880 15534 30932
rect 20162 30880 20168 30932
rect 20220 30920 20226 30932
rect 20714 30920 20720 30932
rect 20220 30892 20720 30920
rect 20220 30880 20226 30892
rect 20714 30880 20720 30892
rect 20772 30880 20778 30932
rect 22094 30880 22100 30932
rect 22152 30920 22158 30932
rect 22373 30923 22431 30929
rect 22373 30920 22385 30923
rect 22152 30892 22385 30920
rect 22152 30880 22158 30892
rect 22373 30889 22385 30892
rect 22419 30889 22431 30923
rect 22373 30883 22431 30889
rect 22649 30923 22707 30929
rect 22649 30889 22661 30923
rect 22695 30920 22707 30923
rect 22738 30920 22744 30932
rect 22695 30892 22744 30920
rect 22695 30889 22707 30892
rect 22649 30883 22707 30889
rect 12069 30855 12127 30861
rect 12069 30852 12081 30855
rect 11716 30824 12081 30852
rect 4663 30756 5028 30784
rect 4663 30753 4675 30756
rect 4617 30747 4675 30753
rect 7558 30744 7564 30796
rect 7616 30784 7622 30796
rect 9677 30787 9735 30793
rect 9677 30784 9689 30787
rect 7616 30756 9689 30784
rect 7616 30744 7622 30756
rect 9677 30753 9689 30756
rect 9723 30753 9735 30787
rect 9677 30747 9735 30753
rect 9769 30787 9827 30793
rect 9769 30753 9781 30787
rect 9815 30784 9827 30787
rect 10318 30784 10324 30796
rect 9815 30756 10324 30784
rect 9815 30753 9827 30756
rect 9769 30747 9827 30753
rect 3050 30676 3056 30728
rect 3108 30716 3114 30728
rect 7006 30716 7012 30728
rect 3108 30688 7012 30716
rect 3108 30676 3114 30688
rect 7006 30676 7012 30688
rect 7064 30676 7070 30728
rect 9692 30716 9720 30747
rect 10318 30744 10324 30756
rect 10376 30784 10382 30796
rect 10962 30784 10968 30796
rect 10376 30756 10968 30784
rect 10376 30744 10382 30756
rect 10962 30744 10968 30756
rect 11020 30784 11026 30796
rect 11716 30793 11744 30824
rect 12069 30821 12081 30824
rect 12115 30852 12127 30855
rect 13998 30852 14004 30864
rect 12115 30824 14004 30852
rect 12115 30821 12127 30824
rect 12069 30815 12127 30821
rect 13998 30812 14004 30824
rect 14056 30812 14062 30864
rect 17954 30812 17960 30864
rect 18012 30852 18018 30864
rect 22554 30852 22560 30864
rect 18012 30824 22560 30852
rect 18012 30812 18018 30824
rect 22554 30812 22560 30824
rect 22612 30812 22618 30864
rect 11701 30787 11759 30793
rect 11020 30756 11560 30784
rect 11020 30744 11026 30756
rect 9953 30719 10011 30725
rect 9953 30716 9965 30719
rect 9692 30688 9965 30716
rect 9953 30685 9965 30688
rect 9999 30685 10011 30719
rect 9953 30679 10011 30685
rect 10873 30719 10931 30725
rect 10873 30685 10885 30719
rect 10919 30716 10931 30719
rect 11054 30716 11060 30728
rect 10919 30688 11060 30716
rect 10919 30685 10931 30688
rect 10873 30679 10931 30685
rect 11054 30676 11060 30688
rect 11112 30676 11118 30728
rect 11422 30716 11428 30728
rect 11383 30688 11428 30716
rect 11422 30676 11428 30688
rect 11480 30676 11486 30728
rect 11532 30716 11560 30756
rect 11701 30753 11713 30787
rect 11747 30753 11759 30787
rect 14182 30784 14188 30796
rect 14143 30756 14188 30784
rect 11701 30747 11759 30753
rect 14182 30744 14188 30756
rect 14240 30744 14246 30796
rect 20806 30744 20812 30796
rect 20864 30784 20870 30796
rect 21361 30787 21419 30793
rect 21361 30784 21373 30787
rect 20864 30756 21373 30784
rect 20864 30744 20870 30756
rect 21361 30753 21373 30756
rect 21407 30784 21419 30787
rect 21913 30787 21971 30793
rect 21913 30784 21925 30787
rect 21407 30756 21925 30784
rect 21407 30753 21419 30756
rect 21361 30747 21419 30753
rect 21913 30753 21925 30756
rect 21959 30753 21971 30787
rect 21913 30747 21971 30753
rect 22097 30787 22155 30793
rect 22097 30753 22109 30787
rect 22143 30784 22155 30787
rect 22664 30784 22692 30883
rect 22738 30880 22744 30892
rect 22796 30920 22802 30932
rect 24688 30920 24716 31096
rect 41325 31093 41337 31096
rect 41371 31093 41383 31127
rect 41325 31087 41383 31093
rect 26786 31016 26792 31068
rect 26844 31056 26850 31068
rect 53926 31056 53932 31068
rect 26844 31028 53932 31056
rect 26844 31016 26850 31028
rect 53926 31016 53932 31028
rect 53984 31016 53990 31068
rect 27062 30948 27068 31000
rect 27120 30988 27126 31000
rect 81802 30988 81808 31000
rect 27120 30960 81808 30988
rect 27120 30948 27126 30960
rect 81802 30948 81808 30960
rect 81860 30948 81866 31000
rect 22796 30892 24716 30920
rect 22796 30880 22802 30892
rect 26878 30880 26884 30932
rect 26936 30920 26942 30932
rect 81526 30920 81532 30932
rect 26936 30892 81532 30920
rect 26936 30880 26942 30892
rect 81526 30880 81532 30892
rect 81584 30880 81590 30932
rect 22143 30756 22692 30784
rect 22143 30753 22155 30756
rect 22097 30747 22155 30753
rect 11885 30719 11943 30725
rect 11885 30716 11897 30719
rect 11532 30688 11897 30716
rect 11885 30685 11897 30688
rect 11931 30685 11943 30719
rect 16206 30716 16212 30728
rect 16119 30688 16212 30716
rect 11885 30679 11943 30685
rect 16206 30676 16212 30688
rect 16264 30676 16270 30728
rect 16482 30716 16488 30728
rect 16443 30688 16488 30716
rect 16482 30676 16488 30688
rect 16540 30676 16546 30728
rect 21177 30719 21235 30725
rect 21177 30716 21189 30719
rect 21008 30688 21189 30716
rect 14366 30540 14372 30592
rect 14424 30580 14430 30592
rect 16025 30583 16083 30589
rect 16025 30580 16037 30583
rect 14424 30552 16037 30580
rect 14424 30540 14430 30552
rect 16025 30549 16037 30552
rect 16071 30580 16083 30583
rect 16224 30580 16252 30676
rect 21008 30592 21036 30688
rect 21177 30685 21189 30688
rect 21223 30685 21235 30719
rect 21177 30679 21235 30685
rect 22830 30676 22836 30728
rect 22888 30716 22894 30728
rect 25961 30719 26019 30725
rect 25961 30716 25973 30719
rect 22888 30688 25973 30716
rect 22888 30676 22894 30688
rect 25961 30685 25973 30688
rect 26007 30685 26019 30719
rect 25961 30679 26019 30685
rect 17586 30580 17592 30592
rect 16071 30552 16252 30580
rect 17547 30552 17592 30580
rect 16071 30549 16083 30552
rect 16025 30543 16083 30549
rect 17586 30540 17592 30552
rect 17644 30580 17650 30592
rect 17770 30580 17776 30592
rect 17644 30552 17776 30580
rect 17644 30540 17650 30552
rect 17770 30540 17776 30552
rect 17828 30540 17834 30592
rect 20990 30580 20996 30592
rect 20951 30552 20996 30580
rect 20990 30540 20996 30552
rect 21048 30540 21054 30592
rect 1104 30490 24656 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 24656 30490
rect 54018 30472 54024 30524
rect 54076 30512 54082 30524
rect 54846 30512 54852 30524
rect 54076 30484 54852 30512
rect 54076 30472 54082 30484
rect 54846 30472 54852 30484
rect 54904 30472 54910 30524
rect 1104 30416 24656 30438
rect 10980 30348 11192 30376
rect 4062 30268 4068 30320
rect 4120 30268 4126 30320
rect 5994 30308 6000 30320
rect 5955 30280 6000 30308
rect 5994 30268 6000 30280
rect 6052 30268 6058 30320
rect 9306 30308 9312 30320
rect 9267 30280 9312 30308
rect 9306 30268 9312 30280
rect 9364 30268 9370 30320
rect 10873 30311 10931 30317
rect 10873 30277 10885 30311
rect 10919 30308 10931 30311
rect 10980 30308 11008 30348
rect 10919 30280 11008 30308
rect 10919 30277 10931 30280
rect 10873 30271 10931 30277
rect 11054 30268 11060 30320
rect 11112 30268 11118 30320
rect 11164 30308 11192 30348
rect 11422 30336 11428 30388
rect 11480 30376 11486 30388
rect 12529 30379 12587 30385
rect 12529 30376 12541 30379
rect 11480 30348 12541 30376
rect 11480 30336 11486 30348
rect 12529 30345 12541 30348
rect 12575 30376 12587 30379
rect 12986 30376 12992 30388
rect 12575 30348 12992 30376
rect 12575 30345 12587 30348
rect 12529 30339 12587 30345
rect 12986 30336 12992 30348
rect 13044 30336 13050 30388
rect 16482 30376 16488 30388
rect 16443 30348 16488 30376
rect 16482 30336 16488 30348
rect 16540 30336 16546 30388
rect 16592 30348 22508 30376
rect 11701 30311 11759 30317
rect 11701 30308 11713 30311
rect 11164 30280 11713 30308
rect 11701 30277 11713 30280
rect 11747 30308 11759 30311
rect 11882 30308 11888 30320
rect 11747 30280 11888 30308
rect 11747 30277 11759 30280
rect 11701 30271 11759 30277
rect 11882 30268 11888 30280
rect 11940 30268 11946 30320
rect 4080 30240 4108 30268
rect 3804 30212 4752 30240
rect 2682 30132 2688 30184
rect 2740 30172 2746 30184
rect 3804 30181 3832 30212
rect 4724 30184 4752 30212
rect 3789 30175 3847 30181
rect 3789 30172 3801 30175
rect 2740 30144 3801 30172
rect 2740 30132 2746 30144
rect 3789 30141 3801 30144
rect 3835 30141 3847 30175
rect 3789 30135 3847 30141
rect 4065 30175 4123 30181
rect 4065 30141 4077 30175
rect 4111 30141 4123 30175
rect 4065 30135 4123 30141
rect 4080 30104 4108 30135
rect 4706 30132 4712 30184
rect 4764 30172 4770 30184
rect 5077 30175 5135 30181
rect 5077 30172 5089 30175
rect 4764 30144 5089 30172
rect 4764 30132 4770 30144
rect 5077 30141 5089 30144
rect 5123 30141 5135 30175
rect 5077 30135 5135 30141
rect 5629 30175 5687 30181
rect 5629 30141 5641 30175
rect 5675 30172 5687 30175
rect 6012 30172 6040 30268
rect 11072 30240 11100 30268
rect 10796 30212 11100 30240
rect 5675 30144 6040 30172
rect 9217 30175 9275 30181
rect 5675 30141 5687 30144
rect 5629 30135 5687 30141
rect 9217 30141 9229 30175
rect 9263 30172 9275 30175
rect 9398 30172 9404 30184
rect 9263 30144 9404 30172
rect 9263 30141 9275 30144
rect 9217 30135 9275 30141
rect 9398 30132 9404 30144
rect 9456 30172 9462 30184
rect 10594 30172 10600 30184
rect 9456 30144 10600 30172
rect 9456 30132 9462 30144
rect 10594 30132 10600 30144
rect 10652 30132 10658 30184
rect 10796 30181 10824 30212
rect 16482 30200 16488 30252
rect 16540 30240 16546 30252
rect 16592 30240 16620 30348
rect 16850 30308 16856 30320
rect 16811 30280 16856 30308
rect 16850 30268 16856 30280
rect 16908 30268 16914 30320
rect 16540 30212 16620 30240
rect 16540 30200 16546 30212
rect 10781 30175 10839 30181
rect 10781 30141 10793 30175
rect 10827 30141 10839 30175
rect 11054 30172 11060 30184
rect 10967 30144 11060 30172
rect 10781 30135 10839 30141
rect 11054 30132 11060 30144
rect 11112 30172 11118 30184
rect 11238 30172 11244 30184
rect 11112 30144 11244 30172
rect 11112 30132 11118 30144
rect 11238 30132 11244 30144
rect 11296 30132 11302 30184
rect 11422 30132 11428 30184
rect 11480 30172 11486 30184
rect 12437 30175 12495 30181
rect 12437 30172 12449 30175
rect 11480 30144 12449 30172
rect 11480 30132 11486 30144
rect 12437 30141 12449 30144
rect 12483 30172 12495 30175
rect 12713 30175 12771 30181
rect 12713 30172 12725 30175
rect 12483 30144 12725 30172
rect 12483 30141 12495 30144
rect 12437 30135 12495 30141
rect 12713 30141 12725 30144
rect 12759 30141 12771 30175
rect 15289 30175 15347 30181
rect 15289 30172 15301 30175
rect 12713 30135 12771 30141
rect 15212 30144 15301 30172
rect 4433 30107 4491 30113
rect 4433 30104 4445 30107
rect 4080 30076 4445 30104
rect 4433 30073 4445 30076
rect 4479 30104 4491 30107
rect 10870 30104 10876 30116
rect 4479 30076 10876 30104
rect 4479 30073 4491 30076
rect 4433 30067 4491 30073
rect 10870 30064 10876 30076
rect 10928 30064 10934 30116
rect 3602 30036 3608 30048
rect 3563 30008 3608 30036
rect 3602 29996 3608 30008
rect 3660 29996 3666 30048
rect 4706 29996 4712 30048
rect 4764 30036 4770 30048
rect 5169 30039 5227 30045
rect 5169 30036 5181 30039
rect 4764 30008 5181 30036
rect 4764 29996 4770 30008
rect 5169 30005 5181 30008
rect 5215 30005 5227 30039
rect 5169 29999 5227 30005
rect 9398 29996 9404 30048
rect 9456 30036 9462 30048
rect 9493 30039 9551 30045
rect 9493 30036 9505 30039
rect 9456 30008 9505 30036
rect 9456 29996 9462 30008
rect 9493 30005 9505 30008
rect 9539 30005 9551 30039
rect 9493 29999 9551 30005
rect 10686 29996 10692 30048
rect 10744 30036 10750 30048
rect 11241 30039 11299 30045
rect 11241 30036 11253 30039
rect 10744 30008 11253 30036
rect 10744 29996 10750 30008
rect 11241 30005 11253 30008
rect 11287 30005 11299 30039
rect 11241 29999 11299 30005
rect 14642 29996 14648 30048
rect 14700 30036 14706 30048
rect 15212 30045 15240 30144
rect 15289 30141 15301 30144
rect 15335 30141 15347 30175
rect 15470 30172 15476 30184
rect 15431 30144 15476 30172
rect 15289 30135 15347 30141
rect 15470 30132 15476 30144
rect 15528 30132 15534 30184
rect 16025 30175 16083 30181
rect 16025 30141 16037 30175
rect 16071 30141 16083 30175
rect 16025 30135 16083 30141
rect 16209 30175 16267 30181
rect 16209 30141 16221 30175
rect 16255 30172 16267 30175
rect 16868 30172 16896 30268
rect 18138 30200 18144 30252
rect 18196 30240 18202 30252
rect 21361 30243 21419 30249
rect 21361 30240 21373 30243
rect 18196 30212 21373 30240
rect 18196 30200 18202 30212
rect 21361 30209 21373 30212
rect 21407 30240 21419 30243
rect 22281 30243 22339 30249
rect 22281 30240 22293 30243
rect 21407 30212 22293 30240
rect 21407 30209 21419 30212
rect 21361 30203 21419 30209
rect 22281 30209 22293 30212
rect 22327 30209 22339 30243
rect 22480 30240 22508 30348
rect 22738 30336 22744 30388
rect 22796 30376 22802 30388
rect 23382 30376 23388 30388
rect 22796 30348 23388 30376
rect 22796 30336 22802 30348
rect 23382 30336 23388 30348
rect 23440 30336 23446 30388
rect 22557 30311 22615 30317
rect 22557 30277 22569 30311
rect 22603 30308 22615 30311
rect 22646 30308 22652 30320
rect 22603 30280 22652 30308
rect 22603 30277 22615 30280
rect 22557 30271 22615 30277
rect 22646 30268 22652 30280
rect 22704 30268 22710 30320
rect 24765 30311 24823 30317
rect 24765 30308 24777 30311
rect 22756 30280 24777 30308
rect 22756 30240 22784 30280
rect 24765 30277 24777 30280
rect 24811 30277 24823 30311
rect 24765 30271 24823 30277
rect 22480 30212 22784 30240
rect 22281 30203 22339 30209
rect 16255 30144 16896 30172
rect 19981 30175 20039 30181
rect 16255 30141 16267 30144
rect 16209 30135 16267 30141
rect 19981 30141 19993 30175
rect 20027 30141 20039 30175
rect 19981 30135 20039 30141
rect 20257 30175 20315 30181
rect 20257 30141 20269 30175
rect 20303 30172 20315 30175
rect 22094 30172 22100 30184
rect 20303 30144 22100 30172
rect 20303 30141 20315 30144
rect 20257 30135 20315 30141
rect 15488 30104 15516 30132
rect 16040 30104 16068 30135
rect 16390 30104 16396 30116
rect 15488 30076 16396 30104
rect 16390 30064 16396 30076
rect 16448 30064 16454 30116
rect 15197 30039 15255 30045
rect 15197 30036 15209 30039
rect 14700 30008 15209 30036
rect 14700 29996 14706 30008
rect 15197 30005 15209 30008
rect 15243 30036 15255 30039
rect 16298 30036 16304 30048
rect 15243 30008 16304 30036
rect 15243 30005 15255 30008
rect 15197 29999 15255 30005
rect 16298 29996 16304 30008
rect 16356 29996 16362 30048
rect 19889 30039 19947 30045
rect 19889 30005 19901 30039
rect 19935 30036 19947 30039
rect 19996 30036 20024 30135
rect 22094 30132 22100 30144
rect 22152 30132 22158 30184
rect 22296 30172 22324 30203
rect 24486 30200 24492 30252
rect 24544 30240 24550 30252
rect 26694 30240 26700 30252
rect 24544 30212 26700 30240
rect 24544 30200 24550 30212
rect 26694 30200 26700 30212
rect 26752 30200 26758 30252
rect 22465 30175 22523 30181
rect 22465 30172 22477 30175
rect 22296 30144 22477 30172
rect 22465 30141 22477 30144
rect 22511 30141 22523 30175
rect 22465 30135 22523 30141
rect 20254 30036 20260 30048
rect 19935 30008 20260 30036
rect 19935 30005 19947 30008
rect 19889 29999 19947 30005
rect 20254 29996 20260 30008
rect 20312 29996 20318 30048
rect 1104 29946 24656 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 24656 29946
rect 1104 29872 24656 29894
rect 3326 29832 3332 29844
rect 3287 29804 3332 29832
rect 3326 29792 3332 29804
rect 3384 29792 3390 29844
rect 8941 29835 8999 29841
rect 8941 29801 8953 29835
rect 8987 29832 8999 29835
rect 9306 29832 9312 29844
rect 8987 29804 9312 29832
rect 8987 29801 8999 29804
rect 8941 29795 8999 29801
rect 2682 29696 2688 29708
rect 2643 29668 2688 29696
rect 2682 29656 2688 29668
rect 2740 29656 2746 29708
rect 2869 29699 2927 29705
rect 2869 29665 2881 29699
rect 2915 29696 2927 29699
rect 3344 29696 3372 29792
rect 2915 29668 3372 29696
rect 4065 29699 4123 29705
rect 2915 29665 2927 29668
rect 2869 29659 2927 29665
rect 4065 29665 4077 29699
rect 4111 29696 4123 29699
rect 5813 29699 5871 29705
rect 5813 29696 5825 29699
rect 4111 29668 5825 29696
rect 4111 29665 4123 29668
rect 4065 29659 4123 29665
rect 5813 29665 5825 29668
rect 5859 29665 5871 29699
rect 5813 29659 5871 29665
rect 7561 29699 7619 29705
rect 7561 29665 7573 29699
rect 7607 29696 7619 29699
rect 7650 29696 7656 29708
rect 7607 29668 7656 29696
rect 7607 29665 7619 29668
rect 7561 29659 7619 29665
rect 2958 29628 2964 29640
rect 2919 29600 2964 29628
rect 2958 29588 2964 29600
rect 3016 29588 3022 29640
rect 2498 29520 2504 29572
rect 2556 29560 2562 29572
rect 4080 29560 4108 29659
rect 7650 29656 7656 29668
rect 7708 29696 7714 29708
rect 8113 29699 8171 29705
rect 8113 29696 8125 29699
rect 7708 29668 8125 29696
rect 7708 29656 7714 29668
rect 8113 29665 8125 29668
rect 8159 29665 8171 29699
rect 8113 29659 8171 29665
rect 8297 29699 8355 29705
rect 8297 29665 8309 29699
rect 8343 29696 8355 29699
rect 8956 29696 8984 29795
rect 9306 29792 9312 29804
rect 9364 29792 9370 29844
rect 14550 29792 14556 29844
rect 14608 29832 14614 29844
rect 16485 29835 16543 29841
rect 16485 29832 16497 29835
rect 14608 29804 16497 29832
rect 14608 29792 14614 29804
rect 16485 29801 16497 29804
rect 16531 29801 16543 29835
rect 16485 29795 16543 29801
rect 22094 29792 22100 29844
rect 22152 29832 22158 29844
rect 22465 29835 22523 29841
rect 22152 29804 22197 29832
rect 22152 29792 22158 29804
rect 22465 29801 22477 29835
rect 22511 29832 22523 29835
rect 22646 29832 22652 29844
rect 22511 29804 22652 29832
rect 22511 29801 22523 29804
rect 22465 29795 22523 29801
rect 22646 29792 22652 29804
rect 22704 29792 22710 29844
rect 10870 29724 10876 29776
rect 10928 29764 10934 29776
rect 26418 29764 26424 29776
rect 10928 29736 26424 29764
rect 10928 29724 10934 29736
rect 26418 29724 26424 29736
rect 26476 29724 26482 29776
rect 11609 29699 11667 29705
rect 11609 29696 11621 29699
rect 8343 29668 8984 29696
rect 9876 29668 11621 29696
rect 8343 29665 8355 29668
rect 8297 29659 8355 29665
rect 9876 29640 9904 29668
rect 11609 29665 11621 29668
rect 11655 29696 11667 29699
rect 14366 29696 14372 29708
rect 11655 29668 14372 29696
rect 11655 29665 11667 29668
rect 11609 29659 11667 29665
rect 14366 29656 14372 29668
rect 14424 29696 14430 29708
rect 14921 29699 14979 29705
rect 14424 29668 14780 29696
rect 14424 29656 14430 29668
rect 4341 29631 4399 29637
rect 4341 29597 4353 29631
rect 4387 29628 4399 29631
rect 5258 29628 5264 29640
rect 4387 29600 5264 29628
rect 4387 29597 4399 29600
rect 4341 29591 4399 29597
rect 5258 29588 5264 29600
rect 5316 29588 5322 29640
rect 7469 29631 7527 29637
rect 7469 29597 7481 29631
rect 7515 29597 7527 29631
rect 9858 29628 9864 29640
rect 9819 29600 9864 29628
rect 7469 29591 7527 29597
rect 2556 29532 4108 29560
rect 2556 29520 2562 29532
rect 4062 29452 4068 29504
rect 4120 29492 4126 29504
rect 5445 29495 5503 29501
rect 5445 29492 5457 29495
rect 4120 29464 5457 29492
rect 4120 29452 4126 29464
rect 5445 29461 5457 29464
rect 5491 29461 5503 29495
rect 7282 29492 7288 29504
rect 7195 29464 7288 29492
rect 5445 29455 5503 29461
rect 7282 29452 7288 29464
rect 7340 29492 7346 29504
rect 7484 29492 7512 29591
rect 9858 29588 9864 29600
rect 9916 29588 9922 29640
rect 10137 29631 10195 29637
rect 10137 29597 10149 29631
rect 10183 29628 10195 29631
rect 10778 29628 10784 29640
rect 10183 29600 10784 29628
rect 10183 29597 10195 29600
rect 10137 29591 10195 29597
rect 10778 29588 10784 29600
rect 10836 29588 10842 29640
rect 8478 29560 8484 29572
rect 8439 29532 8484 29560
rect 8478 29520 8484 29532
rect 8536 29520 8542 29572
rect 14642 29560 14648 29572
rect 10796 29532 14648 29560
rect 10796 29492 10824 29532
rect 14642 29520 14648 29532
rect 14700 29520 14706 29572
rect 7340 29464 10824 29492
rect 7340 29452 7346 29464
rect 11330 29452 11336 29504
rect 11388 29492 11394 29504
rect 14752 29501 14780 29668
rect 14921 29665 14933 29699
rect 14967 29665 14979 29699
rect 15286 29696 15292 29708
rect 15247 29668 15292 29696
rect 14921 29659 14979 29665
rect 14936 29560 14964 29659
rect 15286 29656 15292 29668
rect 15344 29656 15350 29708
rect 15378 29656 15384 29708
rect 15436 29696 15442 29708
rect 15473 29699 15531 29705
rect 15473 29696 15485 29699
rect 15436 29668 15485 29696
rect 15436 29656 15442 29668
rect 15473 29665 15485 29668
rect 15519 29665 15531 29699
rect 16025 29699 16083 29705
rect 16025 29696 16037 29699
rect 15473 29659 15531 29665
rect 15672 29668 16037 29696
rect 15010 29588 15016 29640
rect 15068 29628 15074 29640
rect 15672 29628 15700 29668
rect 16025 29665 16037 29668
rect 16071 29665 16083 29699
rect 16025 29659 16083 29665
rect 16209 29699 16267 29705
rect 16209 29665 16221 29699
rect 16255 29696 16267 29699
rect 16761 29699 16819 29705
rect 16761 29696 16773 29699
rect 16255 29668 16773 29696
rect 16255 29665 16267 29668
rect 16209 29659 16267 29665
rect 16761 29665 16773 29668
rect 16807 29696 16819 29699
rect 17494 29696 17500 29708
rect 16807 29668 17500 29696
rect 16807 29665 16819 29668
rect 16761 29659 16819 29665
rect 17494 29656 17500 29668
rect 17552 29656 17558 29708
rect 20806 29656 20812 29708
rect 20864 29696 20870 29708
rect 21085 29699 21143 29705
rect 21085 29696 21097 29699
rect 20864 29668 21097 29696
rect 20864 29656 20870 29668
rect 21085 29665 21097 29668
rect 21131 29696 21143 29699
rect 21637 29699 21695 29705
rect 21637 29696 21649 29699
rect 21131 29668 21649 29696
rect 21131 29665 21143 29668
rect 21085 29659 21143 29665
rect 21637 29665 21649 29668
rect 21683 29665 21695 29699
rect 21637 29659 21695 29665
rect 21821 29699 21879 29705
rect 21821 29665 21833 29699
rect 21867 29696 21879 29699
rect 22646 29696 22652 29708
rect 21867 29668 22652 29696
rect 21867 29665 21879 29668
rect 21821 29659 21879 29665
rect 22646 29656 22652 29668
rect 22704 29656 22710 29708
rect 20901 29631 20959 29637
rect 20901 29628 20913 29631
rect 15068 29600 15700 29628
rect 20824 29600 20913 29628
rect 15068 29588 15074 29600
rect 16390 29560 16396 29572
rect 14936 29532 16396 29560
rect 16390 29520 16396 29532
rect 16448 29520 16454 29572
rect 20824 29504 20852 29600
rect 20901 29597 20913 29600
rect 20947 29597 20959 29631
rect 20901 29591 20959 29597
rect 11425 29495 11483 29501
rect 11425 29492 11437 29495
rect 11388 29464 11437 29492
rect 11388 29452 11394 29464
rect 11425 29461 11437 29464
rect 11471 29461 11483 29495
rect 11425 29455 11483 29461
rect 14737 29495 14795 29501
rect 14737 29461 14749 29495
rect 14783 29492 14795 29495
rect 14918 29492 14924 29504
rect 14783 29464 14924 29492
rect 14783 29461 14795 29464
rect 14737 29455 14795 29461
rect 14918 29452 14924 29464
rect 14976 29452 14982 29504
rect 15010 29452 15016 29504
rect 15068 29492 15074 29504
rect 20717 29495 20775 29501
rect 15068 29464 15113 29492
rect 15068 29452 15074 29464
rect 20717 29461 20729 29495
rect 20763 29492 20775 29495
rect 20806 29492 20812 29504
rect 20763 29464 20812 29492
rect 20763 29461 20775 29464
rect 20717 29455 20775 29461
rect 20806 29452 20812 29464
rect 20864 29452 20870 29504
rect 53834 29452 53840 29504
rect 53892 29492 53898 29504
rect 54202 29492 54208 29504
rect 53892 29464 54208 29492
rect 53892 29452 53898 29464
rect 54202 29452 54208 29464
rect 54260 29452 54266 29504
rect 1104 29402 24656 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 24656 29402
rect 1104 29328 24656 29350
rect 10778 29288 10784 29300
rect 10739 29260 10784 29288
rect 10778 29248 10784 29260
rect 10836 29248 10842 29300
rect 13998 29248 14004 29300
rect 14056 29288 14062 29300
rect 15010 29288 15016 29300
rect 14056 29260 15016 29288
rect 14056 29248 14062 29260
rect 15010 29248 15016 29260
rect 15068 29248 15074 29300
rect 15105 29291 15163 29297
rect 15105 29257 15117 29291
rect 15151 29288 15163 29291
rect 15194 29288 15200 29300
rect 15151 29260 15200 29288
rect 15151 29257 15163 29260
rect 15105 29251 15163 29257
rect 15194 29248 15200 29260
rect 15252 29248 15258 29300
rect 15470 29220 15476 29232
rect 13924 29192 15476 29220
rect 2501 29155 2559 29161
rect 2501 29121 2513 29155
rect 2547 29152 2559 29155
rect 4249 29155 4307 29161
rect 4249 29152 4261 29155
rect 2547 29124 4261 29152
rect 2547 29121 2559 29124
rect 2501 29115 2559 29121
rect 4249 29121 4261 29124
rect 4295 29152 4307 29155
rect 8205 29155 8263 29161
rect 8205 29152 8217 29155
rect 4295 29124 8217 29152
rect 4295 29121 4307 29124
rect 4249 29115 4307 29121
rect 8205 29121 8217 29124
rect 8251 29121 8263 29155
rect 8478 29152 8484 29164
rect 8439 29124 8484 29152
rect 8205 29115 8263 29121
rect 2777 29087 2835 29093
rect 2777 29053 2789 29087
rect 2823 29084 2835 29087
rect 6914 29084 6920 29096
rect 2823 29056 6920 29084
rect 2823 29053 2835 29056
rect 2777 29047 2835 29053
rect 6914 29044 6920 29056
rect 6972 29044 6978 29096
rect 8220 29084 8248 29115
rect 8478 29112 8484 29124
rect 8536 29112 8542 29164
rect 9398 29112 9404 29164
rect 9456 29152 9462 29164
rect 9585 29155 9643 29161
rect 9585 29152 9597 29155
rect 9456 29124 9597 29152
rect 9456 29112 9462 29124
rect 9585 29121 9597 29124
rect 9631 29121 9643 29155
rect 9585 29115 9643 29121
rect 9858 29084 9864 29096
rect 8220 29056 9864 29084
rect 9858 29044 9864 29056
rect 9916 29084 9922 29096
rect 9953 29087 10011 29093
rect 9953 29084 9965 29087
rect 9916 29056 9965 29084
rect 9916 29044 9922 29056
rect 9953 29053 9965 29056
rect 9999 29053 10011 29087
rect 10686 29084 10692 29096
rect 10647 29056 10692 29084
rect 9953 29047 10011 29053
rect 10686 29044 10692 29056
rect 10744 29044 10750 29096
rect 12434 29044 12440 29096
rect 12492 29084 12498 29096
rect 13449 29087 13507 29093
rect 13449 29084 13461 29087
rect 12492 29056 13461 29084
rect 12492 29044 12498 29056
rect 13449 29053 13461 29056
rect 13495 29084 13507 29087
rect 13541 29087 13599 29093
rect 13541 29084 13553 29087
rect 13495 29056 13553 29084
rect 13495 29053 13507 29056
rect 13449 29047 13507 29053
rect 13541 29053 13553 29056
rect 13587 29053 13599 29087
rect 13541 29047 13599 29053
rect 13725 29087 13783 29093
rect 13725 29053 13737 29087
rect 13771 29084 13783 29087
rect 13924 29084 13952 29192
rect 15470 29180 15476 29192
rect 15528 29180 15534 29232
rect 19429 29155 19487 29161
rect 19429 29152 19441 29155
rect 19168 29124 19441 29152
rect 14277 29087 14335 29093
rect 14277 29084 14289 29087
rect 13771 29056 14289 29084
rect 13771 29053 13783 29056
rect 13725 29047 13783 29053
rect 14277 29053 14289 29056
rect 14323 29053 14335 29087
rect 14277 29047 14335 29053
rect 14461 29087 14519 29093
rect 14461 29053 14473 29087
rect 14507 29084 14519 29087
rect 15194 29084 15200 29096
rect 14507 29056 15200 29084
rect 14507 29053 14519 29056
rect 14461 29047 14519 29053
rect 15194 29044 15200 29056
rect 15252 29044 15258 29096
rect 17126 29044 17132 29096
rect 17184 29084 17190 29096
rect 19168 29093 19196 29124
rect 19429 29121 19441 29124
rect 19475 29121 19487 29155
rect 21637 29155 21695 29161
rect 21637 29152 21649 29155
rect 19429 29115 19487 29121
rect 20824 29124 21649 29152
rect 19153 29087 19211 29093
rect 19153 29084 19165 29087
rect 17184 29056 19165 29084
rect 17184 29044 17190 29056
rect 19153 29053 19165 29056
rect 19199 29053 19211 29087
rect 19153 29047 19211 29053
rect 19334 29044 19340 29096
rect 19392 29084 19398 29096
rect 19521 29087 19579 29093
rect 19521 29084 19533 29087
rect 19392 29056 19533 29084
rect 19392 29044 19398 29056
rect 19521 29053 19533 29056
rect 19567 29053 19579 29087
rect 19521 29047 19579 29053
rect 20073 29087 20131 29093
rect 20073 29053 20085 29087
rect 20119 29053 20131 29087
rect 20073 29047 20131 29053
rect 20257 29087 20315 29093
rect 20257 29053 20269 29087
rect 20303 29084 20315 29087
rect 20824 29084 20852 29124
rect 21637 29121 21649 29124
rect 21683 29121 21695 29155
rect 24762 29152 24768 29164
rect 21637 29115 21695 29121
rect 22388 29124 24768 29152
rect 20303 29056 20852 29084
rect 21545 29087 21603 29093
rect 20303 29053 20315 29056
rect 20257 29047 20315 29053
rect 21545 29053 21557 29087
rect 21591 29084 21603 29087
rect 21818 29084 21824 29096
rect 21591 29056 21824 29084
rect 21591 29053 21603 29056
rect 21545 29047 21603 29053
rect 3970 29016 3976 29028
rect 3712 28988 3976 29016
rect 2590 28908 2596 28960
rect 2648 28948 2654 28960
rect 3712 28948 3740 28988
rect 3970 28976 3976 28988
rect 4028 28976 4034 29028
rect 19536 29016 19564 29047
rect 20088 29016 20116 29047
rect 21818 29044 21824 29056
rect 21876 29084 21882 29096
rect 22388 29084 22416 29124
rect 24762 29112 24768 29124
rect 24820 29112 24826 29164
rect 22554 29084 22560 29096
rect 21876 29056 22416 29084
rect 22467 29056 22560 29084
rect 21876 29044 21882 29056
rect 22554 29044 22560 29056
rect 22612 29084 22618 29096
rect 23474 29084 23480 29096
rect 22612 29056 23480 29084
rect 22612 29044 22618 29056
rect 23474 29044 23480 29056
rect 23532 29044 23538 29096
rect 4172 28988 4384 29016
rect 3878 28948 3884 28960
rect 2648 28920 3740 28948
rect 3839 28920 3884 28948
rect 2648 28908 2654 28920
rect 3878 28908 3884 28920
rect 3936 28908 3942 28960
rect 4062 28908 4068 28960
rect 4120 28948 4126 28960
rect 4172 28948 4200 28988
rect 4120 28920 4200 28948
rect 4356 28948 4384 28988
rect 9508 28988 10088 29016
rect 9508 28948 9536 28988
rect 4356 28920 9536 28948
rect 10060 28948 10088 28988
rect 13280 28988 13492 29016
rect 13280 28948 13308 28988
rect 10060 28920 13308 28948
rect 13464 28948 13492 28988
rect 14568 28988 15148 29016
rect 14568 28948 14596 28988
rect 14734 28948 14740 28960
rect 13464 28920 14596 28948
rect 14695 28920 14740 28948
rect 4120 28908 4126 28920
rect 14734 28908 14740 28920
rect 14792 28908 14798 28960
rect 15120 28948 15148 28988
rect 19076 28988 19288 29016
rect 19536 28988 20116 29016
rect 20625 29019 20683 29025
rect 19076 28948 19104 28988
rect 15120 28920 19104 28948
rect 19260 28948 19288 28988
rect 20625 28985 20637 29019
rect 20671 29016 20683 29019
rect 20714 29016 20720 29028
rect 20671 28988 20720 29016
rect 20671 28985 20683 28988
rect 20625 28979 20683 28985
rect 20714 28976 20720 28988
rect 20772 28976 20778 29028
rect 22480 28988 22784 29016
rect 22480 28948 22508 28988
rect 22646 28948 22652 28960
rect 19260 28920 22508 28948
rect 22607 28920 22652 28948
rect 22646 28908 22652 28920
rect 22704 28908 22710 28960
rect 22756 28948 22784 28988
rect 27338 28948 27344 28960
rect 22756 28920 27344 28948
rect 27338 28908 27344 28920
rect 27396 28908 27402 28960
rect 1104 28858 24656 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 24656 28858
rect 1104 28784 24656 28806
rect 3970 28704 3976 28756
rect 4028 28744 4034 28756
rect 4157 28747 4215 28753
rect 4157 28744 4169 28747
rect 4028 28716 4169 28744
rect 4028 28704 4034 28716
rect 4157 28713 4169 28716
rect 4203 28713 4215 28747
rect 4157 28707 4215 28713
rect 4985 28747 5043 28753
rect 4985 28713 4997 28747
rect 5031 28744 5043 28747
rect 5031 28716 14964 28744
rect 5031 28713 5043 28716
rect 4985 28707 5043 28713
rect 4341 28611 4399 28617
rect 4341 28577 4353 28611
rect 4387 28608 4399 28611
rect 4522 28608 4528 28620
rect 4387 28580 4528 28608
rect 4387 28577 4399 28580
rect 4341 28571 4399 28577
rect 4522 28568 4528 28580
rect 4580 28568 4586 28620
rect 4617 28611 4675 28617
rect 4617 28577 4629 28611
rect 4663 28608 4675 28611
rect 5000 28608 5028 28707
rect 12912 28648 14320 28676
rect 12912 28617 12940 28648
rect 4663 28580 5028 28608
rect 12897 28611 12955 28617
rect 4663 28577 4675 28580
rect 4617 28571 4675 28577
rect 12897 28577 12909 28611
rect 12943 28577 12955 28611
rect 14185 28611 14243 28617
rect 14185 28608 14197 28611
rect 12897 28571 12955 28577
rect 14016 28580 14197 28608
rect 12805 28543 12863 28549
rect 12805 28509 12817 28543
rect 12851 28540 12863 28543
rect 13722 28540 13728 28552
rect 12851 28512 13728 28540
rect 12851 28509 12863 28512
rect 12805 28503 12863 28509
rect 13722 28500 13728 28512
rect 13780 28500 13786 28552
rect 10962 28432 10968 28484
rect 11020 28472 11026 28484
rect 14016 28481 14044 28580
rect 14185 28577 14197 28580
rect 14231 28577 14243 28611
rect 14185 28571 14243 28577
rect 14001 28475 14059 28481
rect 14001 28472 14013 28475
rect 11020 28444 14013 28472
rect 11020 28432 11026 28444
rect 14001 28441 14013 28444
rect 14047 28441 14059 28475
rect 14001 28435 14059 28441
rect 11790 28364 11796 28416
rect 11848 28404 11854 28416
rect 14292 28413 14320 28648
rect 14936 28472 14964 28716
rect 15194 28704 15200 28756
rect 15252 28744 15258 28756
rect 15381 28747 15439 28753
rect 15381 28744 15393 28747
rect 15252 28716 15393 28744
rect 15252 28704 15258 28716
rect 15381 28713 15393 28716
rect 15427 28713 15439 28747
rect 15381 28707 15439 28713
rect 19797 28747 19855 28753
rect 19797 28713 19809 28747
rect 19843 28744 19855 28747
rect 19843 28716 21128 28744
rect 19843 28713 19855 28716
rect 19797 28707 19855 28713
rect 19886 28636 19892 28688
rect 19944 28676 19950 28688
rect 20162 28676 20168 28688
rect 19944 28648 20168 28676
rect 19944 28636 19950 28648
rect 20162 28636 20168 28648
rect 20220 28636 20226 28688
rect 20346 28636 20352 28688
rect 20404 28676 20410 28688
rect 20530 28676 20536 28688
rect 20404 28648 20536 28676
rect 20404 28636 20410 28648
rect 20530 28636 20536 28648
rect 20588 28636 20594 28688
rect 15286 28608 15292 28620
rect 15247 28580 15292 28608
rect 15286 28568 15292 28580
rect 15344 28568 15350 28620
rect 16574 28608 16580 28620
rect 16535 28580 16580 28608
rect 16574 28568 16580 28580
rect 16632 28568 16638 28620
rect 18785 28611 18843 28617
rect 18785 28577 18797 28611
rect 18831 28608 18843 28611
rect 19334 28608 19340 28620
rect 18831 28580 19340 28608
rect 18831 28577 18843 28580
rect 18785 28571 18843 28577
rect 19334 28568 19340 28580
rect 19392 28568 19398 28620
rect 19518 28608 19524 28620
rect 19479 28580 19524 28608
rect 19518 28568 19524 28580
rect 19576 28568 19582 28620
rect 21100 28608 21128 28716
rect 21269 28611 21327 28617
rect 21269 28608 21281 28611
rect 21100 28580 21281 28608
rect 21269 28577 21281 28580
rect 21315 28577 21327 28611
rect 21269 28571 21327 28577
rect 18414 28500 18420 28552
rect 18472 28540 18478 28552
rect 18601 28543 18659 28549
rect 18601 28540 18613 28543
rect 18472 28512 18613 28540
rect 18472 28500 18478 28512
rect 18601 28509 18613 28512
rect 18647 28509 18659 28543
rect 18601 28503 18659 28509
rect 20346 28500 20352 28552
rect 20404 28540 20410 28552
rect 20993 28543 21051 28549
rect 20993 28540 21005 28543
rect 20404 28512 21005 28540
rect 20404 28500 20410 28512
rect 20993 28509 21005 28512
rect 21039 28509 21051 28543
rect 22554 28540 22560 28552
rect 22515 28512 22560 28540
rect 20993 28503 21051 28509
rect 22554 28500 22560 28512
rect 22612 28500 22618 28552
rect 14936 28444 20760 28472
rect 13081 28407 13139 28413
rect 13081 28404 13093 28407
rect 11848 28376 13093 28404
rect 11848 28364 11854 28376
rect 13081 28373 13093 28376
rect 13127 28373 13139 28407
rect 13081 28367 13139 28373
rect 14277 28407 14335 28413
rect 14277 28373 14289 28407
rect 14323 28404 14335 28407
rect 15378 28404 15384 28416
rect 14323 28376 15384 28404
rect 14323 28373 14335 28376
rect 14277 28367 14335 28373
rect 15378 28364 15384 28376
rect 15436 28404 15442 28416
rect 15654 28404 15660 28416
rect 15436 28376 15660 28404
rect 15436 28364 15442 28376
rect 15654 28364 15660 28376
rect 15712 28364 15718 28416
rect 16390 28404 16396 28416
rect 16351 28376 16396 28404
rect 16390 28364 16396 28376
rect 16448 28364 16454 28416
rect 18414 28404 18420 28416
rect 18375 28376 18420 28404
rect 18414 28364 18420 28376
rect 18472 28364 18478 28416
rect 20346 28364 20352 28416
rect 20404 28404 20410 28416
rect 20625 28407 20683 28413
rect 20625 28404 20637 28407
rect 20404 28376 20637 28404
rect 20404 28364 20410 28376
rect 20625 28373 20637 28376
rect 20671 28373 20683 28407
rect 20732 28404 20760 28444
rect 26510 28404 26516 28416
rect 20732 28376 26516 28404
rect 20625 28367 20683 28373
rect 26510 28364 26516 28376
rect 26568 28364 26574 28416
rect 54113 28407 54171 28413
rect 54113 28373 54125 28407
rect 54159 28404 54171 28407
rect 54294 28404 54300 28416
rect 54159 28376 54300 28404
rect 54159 28373 54171 28376
rect 54113 28367 54171 28373
rect 54294 28364 54300 28376
rect 54352 28364 54358 28416
rect 1104 28314 24656 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 24656 28314
rect 1104 28240 24656 28262
rect 13814 28160 13820 28212
rect 13872 28200 13878 28212
rect 18414 28200 18420 28212
rect 13872 28172 18420 28200
rect 13872 28160 13878 28172
rect 18414 28160 18420 28172
rect 18472 28160 18478 28212
rect 21818 28200 21824 28212
rect 21779 28172 21824 28200
rect 21818 28160 21824 28172
rect 21876 28160 21882 28212
rect 18785 28135 18843 28141
rect 18785 28101 18797 28135
rect 18831 28132 18843 28135
rect 20165 28135 20223 28141
rect 20165 28132 20177 28135
rect 18831 28104 20177 28132
rect 18831 28101 18843 28104
rect 18785 28095 18843 28101
rect 20165 28101 20177 28104
rect 20211 28101 20223 28135
rect 20165 28095 20223 28101
rect 2498 28064 2504 28076
rect 2459 28036 2504 28064
rect 2498 28024 2504 28036
rect 2556 28024 2562 28076
rect 7834 28024 7840 28076
rect 7892 28064 7898 28076
rect 8389 28067 8447 28073
rect 8389 28064 8401 28067
rect 7892 28036 8401 28064
rect 7892 28024 7898 28036
rect 8389 28033 8401 28036
rect 8435 28033 8447 28067
rect 8389 28027 8447 28033
rect 13817 28067 13875 28073
rect 13817 28033 13829 28067
rect 13863 28064 13875 28067
rect 14734 28064 14740 28076
rect 13863 28036 14740 28064
rect 13863 28033 13875 28036
rect 13817 28027 13875 28033
rect 14734 28024 14740 28036
rect 14792 28024 14798 28076
rect 20714 28064 20720 28076
rect 20675 28036 20720 28064
rect 20714 28024 20720 28036
rect 20772 28024 20778 28076
rect 2590 27956 2596 28008
rect 2648 27996 2654 28008
rect 2777 27999 2835 28005
rect 2777 27996 2789 27999
rect 2648 27968 2789 27996
rect 2648 27956 2654 27968
rect 2777 27965 2789 27968
rect 2823 27965 2835 27999
rect 7926 27996 7932 28008
rect 7887 27968 7932 27996
rect 2777 27959 2835 27965
rect 7926 27956 7932 27968
rect 7984 27956 7990 28008
rect 8021 27999 8079 28005
rect 8021 27965 8033 27999
rect 8067 27965 8079 27999
rect 8294 27996 8300 28008
rect 8255 27968 8300 27996
rect 8021 27959 8079 27965
rect 6914 27888 6920 27940
rect 6972 27928 6978 27940
rect 7285 27931 7343 27937
rect 7285 27928 7297 27931
rect 6972 27900 7297 27928
rect 6972 27888 6978 27900
rect 7285 27897 7297 27900
rect 7331 27897 7343 27931
rect 8036 27928 8064 27959
rect 8294 27956 8300 27968
rect 8352 27956 8358 28008
rect 11241 27999 11299 28005
rect 11241 27965 11253 27999
rect 11287 27996 11299 27999
rect 11974 27996 11980 28008
rect 11287 27968 11980 27996
rect 11287 27965 11299 27968
rect 11241 27959 11299 27965
rect 11974 27956 11980 27968
rect 12032 27956 12038 28008
rect 13541 27999 13599 28005
rect 13541 27965 13553 27999
rect 13587 27996 13599 27999
rect 14918 27996 14924 28008
rect 13587 27968 14924 27996
rect 13587 27965 13599 27968
rect 13541 27959 13599 27965
rect 14918 27956 14924 27968
rect 14976 27996 14982 28008
rect 15289 27999 15347 28005
rect 15289 27996 15301 27999
rect 14976 27968 15301 27996
rect 14976 27956 14982 27968
rect 15289 27965 15301 27968
rect 15335 27965 15347 27999
rect 15289 27959 15347 27965
rect 16390 27956 16396 28008
rect 16448 27996 16454 28008
rect 18969 27999 19027 28005
rect 18969 27996 18981 27999
rect 16448 27968 18981 27996
rect 16448 27956 16454 27968
rect 18969 27965 18981 27968
rect 19015 27965 19027 27999
rect 18969 27959 19027 27965
rect 20165 27999 20223 28005
rect 20165 27965 20177 27999
rect 20211 27996 20223 27999
rect 20346 27996 20352 28008
rect 20211 27968 20352 27996
rect 20211 27965 20223 27968
rect 20165 27959 20223 27965
rect 20346 27956 20352 27968
rect 20404 27996 20410 28008
rect 20441 27999 20499 28005
rect 20441 27996 20453 27999
rect 20404 27968 20453 27996
rect 20404 27956 20410 27968
rect 20441 27965 20453 27968
rect 20487 27965 20499 27999
rect 20441 27959 20499 27965
rect 11054 27928 11060 27940
rect 8036 27900 11060 27928
rect 7285 27891 7343 27897
rect 11054 27888 11060 27900
rect 11112 27888 11118 27940
rect 3878 27860 3884 27872
rect 3839 27832 3884 27860
rect 3878 27820 3884 27832
rect 3936 27820 3942 27872
rect 4341 27863 4399 27869
rect 4341 27829 4353 27863
rect 4387 27860 4399 27863
rect 4614 27860 4620 27872
rect 4387 27832 4620 27860
rect 4387 27829 4399 27832
rect 4341 27823 4399 27829
rect 4614 27820 4620 27832
rect 4672 27820 4678 27872
rect 11422 27860 11428 27872
rect 11383 27832 11428 27860
rect 11422 27820 11428 27832
rect 11480 27820 11486 27872
rect 14274 27820 14280 27872
rect 14332 27860 14338 27872
rect 14921 27863 14979 27869
rect 14921 27860 14933 27863
rect 14332 27832 14933 27860
rect 14332 27820 14338 27832
rect 14921 27829 14933 27832
rect 14967 27860 14979 27863
rect 15286 27860 15292 27872
rect 14967 27832 15292 27860
rect 14967 27829 14979 27832
rect 14921 27823 14979 27829
rect 15286 27820 15292 27832
rect 15344 27820 15350 27872
rect 20349 27863 20407 27869
rect 20349 27829 20361 27863
rect 20395 27860 20407 27863
rect 20456 27860 20484 27959
rect 20806 27860 20812 27872
rect 20395 27832 20812 27860
rect 20395 27829 20407 27832
rect 20349 27823 20407 27829
rect 20806 27820 20812 27832
rect 20864 27820 20870 27872
rect 21358 27820 21364 27872
rect 21416 27860 21422 27872
rect 24394 27860 24400 27872
rect 21416 27832 24400 27860
rect 21416 27820 21422 27832
rect 24394 27820 24400 27832
rect 24452 27820 24458 27872
rect 1104 27770 24656 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 24656 27770
rect 1104 27696 24656 27718
rect 9582 27656 9588 27668
rect 6932 27628 9588 27656
rect 6932 27461 6960 27628
rect 9582 27616 9588 27628
rect 9640 27616 9646 27668
rect 7760 27560 8524 27588
rect 7101 27523 7159 27529
rect 7101 27489 7113 27523
rect 7147 27520 7159 27523
rect 7650 27520 7656 27532
rect 7147 27492 7656 27520
rect 7147 27489 7159 27492
rect 7101 27483 7159 27489
rect 7650 27480 7656 27492
rect 7708 27480 7714 27532
rect 7760 27520 7788 27560
rect 8496 27532 8524 27560
rect 9490 27548 9496 27600
rect 9548 27588 9554 27600
rect 12526 27588 12532 27600
rect 9548 27560 9720 27588
rect 12487 27560 12532 27588
rect 9548 27548 9554 27560
rect 7828 27523 7886 27529
rect 7828 27520 7840 27523
rect 7760 27492 7840 27520
rect 7828 27489 7840 27492
rect 7874 27489 7886 27523
rect 8478 27520 8484 27532
rect 8439 27492 8484 27520
rect 7828 27483 7886 27489
rect 8478 27480 8484 27492
rect 8536 27480 8542 27532
rect 9692 27529 9720 27560
rect 12526 27548 12532 27560
rect 12584 27548 12590 27600
rect 15657 27591 15715 27597
rect 15657 27588 15669 27591
rect 15304 27560 15669 27588
rect 9677 27523 9735 27529
rect 9677 27489 9689 27523
rect 9723 27489 9735 27523
rect 9677 27483 9735 27489
rect 9766 27480 9772 27532
rect 9824 27520 9830 27532
rect 15304 27529 15332 27560
rect 15657 27557 15669 27560
rect 15703 27588 15715 27591
rect 15703 27560 18460 27588
rect 15703 27557 15715 27560
rect 15657 27551 15715 27557
rect 14369 27523 14427 27529
rect 9824 27492 13676 27520
rect 9824 27480 9830 27492
rect 6917 27455 6975 27461
rect 6917 27421 6929 27455
rect 6963 27421 6975 27455
rect 6917 27415 6975 27421
rect 6638 27276 6644 27328
rect 6696 27316 6702 27328
rect 6733 27319 6791 27325
rect 6733 27316 6745 27319
rect 6696 27288 6745 27316
rect 6696 27276 6702 27288
rect 6733 27285 6745 27288
rect 6779 27316 6791 27319
rect 6932 27316 6960 27415
rect 8386 27412 8392 27464
rect 8444 27452 8450 27464
rect 9490 27452 9496 27464
rect 8444 27424 9496 27452
rect 8444 27412 8450 27424
rect 9490 27412 9496 27424
rect 9548 27412 9554 27464
rect 12526 27412 12532 27464
rect 12584 27452 12590 27464
rect 12713 27455 12771 27461
rect 12713 27452 12725 27455
rect 12584 27424 12725 27452
rect 12584 27412 12590 27424
rect 12713 27421 12725 27424
rect 12759 27421 12771 27455
rect 12986 27452 12992 27464
rect 12947 27424 12992 27452
rect 12713 27415 12771 27421
rect 12986 27412 12992 27424
rect 13044 27412 13050 27464
rect 7098 27344 7104 27396
rect 7156 27384 7162 27396
rect 8021 27387 8079 27393
rect 8021 27384 8033 27387
rect 7156 27356 8033 27384
rect 7156 27344 7162 27356
rect 8021 27353 8033 27356
rect 8067 27353 8079 27387
rect 13648 27384 13676 27492
rect 14369 27489 14381 27523
rect 14415 27520 14427 27523
rect 15289 27523 15347 27529
rect 15289 27520 15301 27523
rect 14415 27492 15301 27520
rect 14415 27489 14427 27492
rect 14369 27483 14427 27489
rect 15289 27489 15301 27492
rect 15335 27489 15347 27523
rect 16298 27520 16304 27532
rect 16259 27492 16304 27520
rect 15289 27483 15347 27489
rect 16298 27480 16304 27492
rect 16356 27520 16362 27532
rect 16485 27523 16543 27529
rect 16485 27520 16497 27523
rect 16356 27492 16497 27520
rect 16356 27480 16362 27492
rect 16485 27489 16497 27492
rect 16531 27489 16543 27523
rect 16485 27483 16543 27489
rect 16669 27523 16727 27529
rect 16669 27489 16681 27523
rect 16715 27520 16727 27523
rect 17218 27520 17224 27532
rect 16715 27492 17224 27520
rect 16715 27489 16727 27492
rect 16669 27483 16727 27489
rect 17218 27480 17224 27492
rect 17276 27480 17282 27532
rect 17405 27523 17463 27529
rect 17405 27489 17417 27523
rect 17451 27520 17463 27523
rect 18322 27520 18328 27532
rect 17451 27492 18328 27520
rect 17451 27489 17463 27492
rect 17405 27483 17463 27489
rect 18322 27480 18328 27492
rect 18380 27480 18386 27532
rect 18432 27520 18460 27560
rect 53834 27548 53840 27600
rect 53892 27588 53898 27600
rect 54110 27588 54116 27600
rect 53892 27560 54116 27588
rect 53892 27548 53898 27560
rect 54110 27548 54116 27560
rect 54168 27548 54174 27600
rect 21358 27520 21364 27532
rect 18432 27492 21364 27520
rect 21358 27480 21364 27492
rect 21416 27480 21422 27532
rect 21450 27412 21456 27464
rect 21508 27452 21514 27464
rect 21637 27455 21695 27461
rect 21637 27452 21649 27455
rect 21508 27424 21649 27452
rect 21508 27412 21514 27424
rect 21637 27421 21649 27424
rect 21683 27421 21695 27455
rect 21910 27452 21916 27464
rect 21871 27424 21916 27452
rect 21637 27415 21695 27421
rect 21910 27412 21916 27424
rect 21968 27412 21974 27464
rect 22922 27412 22928 27464
rect 22980 27452 22986 27464
rect 23198 27452 23204 27464
rect 22980 27424 23204 27452
rect 22980 27412 22986 27424
rect 23198 27412 23204 27424
rect 23256 27412 23262 27464
rect 28350 27384 28356 27396
rect 13648 27356 21588 27384
rect 8021 27347 8079 27353
rect 6779 27288 6960 27316
rect 6779 27285 6791 27288
rect 6733 27279 6791 27285
rect 7650 27276 7656 27328
rect 7708 27316 7714 27328
rect 11422 27316 11428 27328
rect 7708 27288 11428 27316
rect 7708 27276 7714 27288
rect 11422 27276 11428 27288
rect 11480 27276 11486 27328
rect 13078 27276 13084 27328
rect 13136 27316 13142 27328
rect 15381 27319 15439 27325
rect 15381 27316 15393 27319
rect 13136 27288 15393 27316
rect 13136 27276 13142 27288
rect 15381 27285 15393 27288
rect 15427 27285 15439 27319
rect 15381 27279 15439 27285
rect 17681 27319 17739 27325
rect 17681 27285 17693 27319
rect 17727 27316 17739 27319
rect 17862 27316 17868 27328
rect 17727 27288 17868 27316
rect 17727 27285 17739 27288
rect 17681 27279 17739 27285
rect 17862 27276 17868 27288
rect 17920 27276 17926 27328
rect 20806 27276 20812 27328
rect 20864 27316 20870 27328
rect 21450 27316 21456 27328
rect 20864 27288 21456 27316
rect 20864 27276 20870 27288
rect 21450 27276 21456 27288
rect 21508 27276 21514 27328
rect 21560 27316 21588 27356
rect 23032 27356 28356 27384
rect 23032 27316 23060 27356
rect 28350 27344 28356 27356
rect 28408 27344 28414 27396
rect 23198 27316 23204 27328
rect 21560 27288 23060 27316
rect 23159 27288 23204 27316
rect 23198 27276 23204 27288
rect 23256 27276 23262 27328
rect 1104 27226 24656 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 24656 27226
rect 1104 27152 24656 27174
rect 2774 27072 2780 27124
rect 2832 27112 2838 27124
rect 3418 27112 3424 27124
rect 2832 27084 3424 27112
rect 2832 27072 2838 27084
rect 3418 27072 3424 27084
rect 3476 27072 3482 27124
rect 4062 27072 4068 27124
rect 4120 27112 4126 27124
rect 25682 27112 25688 27124
rect 4120 27084 25688 27112
rect 4120 27072 4126 27084
rect 25682 27072 25688 27084
rect 25740 27072 25746 27124
rect 4341 27047 4399 27053
rect 4341 27013 4353 27047
rect 4387 27044 4399 27047
rect 4614 27044 4620 27056
rect 4387 27016 4620 27044
rect 4387 27013 4399 27016
rect 4341 27007 4399 27013
rect 4614 27004 4620 27016
rect 4672 27044 4678 27056
rect 6822 27044 6828 27056
rect 4672 27016 6828 27044
rect 4672 27004 4678 27016
rect 6822 27004 6828 27016
rect 6880 27004 6886 27056
rect 7760 27016 12848 27044
rect 2498 26976 2504 26988
rect 2459 26948 2504 26976
rect 2498 26936 2504 26948
rect 2556 26936 2562 26988
rect 2777 26979 2835 26985
rect 2777 26945 2789 26979
rect 2823 26976 2835 26979
rect 3602 26976 3608 26988
rect 2823 26948 3608 26976
rect 2823 26945 2835 26948
rect 2777 26939 2835 26945
rect 3602 26936 3608 26948
rect 3660 26936 3666 26988
rect 4062 26936 4068 26988
rect 4120 26976 4126 26988
rect 7098 26976 7104 26988
rect 4120 26948 6960 26976
rect 7059 26948 7104 26976
rect 4120 26936 4126 26948
rect 5721 26911 5779 26917
rect 5721 26877 5733 26911
rect 5767 26877 5779 26911
rect 6822 26908 6828 26920
rect 6783 26880 6828 26908
rect 5721 26871 5779 26877
rect 5736 26840 5764 26871
rect 6822 26868 6828 26880
rect 6880 26868 6886 26920
rect 6932 26908 6960 26948
rect 7098 26936 7104 26948
rect 7156 26936 7162 26988
rect 7760 26908 7788 27016
rect 12253 26979 12311 26985
rect 12253 26945 12265 26979
rect 12299 26976 12311 26979
rect 12437 26979 12495 26985
rect 12437 26976 12449 26979
rect 12299 26948 12449 26976
rect 12299 26945 12311 26948
rect 12253 26939 12311 26945
rect 12437 26945 12449 26948
rect 12483 26976 12495 26979
rect 12483 26948 12756 26976
rect 12483 26945 12495 26948
rect 12437 26939 12495 26945
rect 6932 26880 7788 26908
rect 11422 26868 11428 26920
rect 11480 26908 11486 26920
rect 12575 26911 12633 26917
rect 12575 26908 12587 26911
rect 11480 26880 12587 26908
rect 11480 26868 11486 26880
rect 12575 26877 12587 26880
rect 12621 26877 12633 26911
rect 12575 26871 12633 26877
rect 12728 26852 12756 26948
rect 6914 26840 6920 26852
rect 5736 26812 6920 26840
rect 6914 26800 6920 26812
rect 6972 26800 6978 26852
rect 12710 26800 12716 26852
rect 12768 26800 12774 26852
rect 12820 26840 12848 27016
rect 12986 27004 12992 27056
rect 13044 27044 13050 27056
rect 13541 27047 13599 27053
rect 13541 27044 13553 27047
rect 13044 27016 13553 27044
rect 13044 27004 13050 27016
rect 13541 27013 13553 27016
rect 13587 27013 13599 27047
rect 18322 27044 18328 27056
rect 18283 27016 18328 27044
rect 13541 27007 13599 27013
rect 18322 27004 18328 27016
rect 18380 27004 18386 27056
rect 19886 27004 19892 27056
rect 19944 27044 19950 27056
rect 20622 27044 20628 27056
rect 19944 27016 20628 27044
rect 19944 27004 19950 27016
rect 20622 27004 20628 27016
rect 20680 27004 20686 27056
rect 19904 26976 19932 27004
rect 21177 26979 21235 26985
rect 18156 26948 20116 26976
rect 12986 26868 12992 26920
rect 13044 26908 13050 26920
rect 13081 26911 13139 26917
rect 13081 26908 13093 26911
rect 13044 26880 13093 26908
rect 13044 26868 13050 26880
rect 13081 26877 13093 26880
rect 13127 26877 13139 26911
rect 13081 26871 13139 26877
rect 13170 26868 13176 26920
rect 13228 26908 13234 26920
rect 18156 26908 18184 26948
rect 13228 26880 18184 26908
rect 18233 26911 18291 26917
rect 13228 26868 13234 26880
rect 18233 26877 18245 26911
rect 18279 26908 18291 26911
rect 19242 26908 19248 26920
rect 18279 26880 19248 26908
rect 18279 26877 18291 26880
rect 18233 26871 18291 26877
rect 19242 26868 19248 26880
rect 19300 26868 19306 26920
rect 20088 26917 20116 26948
rect 21177 26945 21189 26979
rect 21223 26976 21235 26979
rect 21910 26976 21916 26988
rect 21223 26948 21916 26976
rect 21223 26945 21235 26948
rect 21177 26939 21235 26945
rect 21910 26936 21916 26948
rect 21968 26936 21974 26988
rect 19889 26911 19947 26917
rect 19889 26877 19901 26911
rect 19935 26877 19947 26911
rect 19889 26871 19947 26877
rect 20073 26911 20131 26917
rect 20073 26877 20085 26911
rect 20119 26877 20131 26911
rect 20073 26871 20131 26877
rect 18690 26840 18696 26852
rect 12820 26812 18696 26840
rect 18690 26800 18696 26812
rect 18748 26800 18754 26852
rect 3418 26732 3424 26784
rect 3476 26772 3482 26784
rect 3602 26772 3608 26784
rect 3476 26744 3608 26772
rect 3476 26732 3482 26744
rect 3602 26732 3608 26744
rect 3660 26732 3666 26784
rect 3878 26772 3884 26784
rect 3839 26744 3884 26772
rect 3878 26732 3884 26744
rect 3936 26732 3942 26784
rect 5813 26775 5871 26781
rect 5813 26741 5825 26775
rect 5859 26772 5871 26775
rect 6730 26772 6736 26784
rect 5859 26744 6736 26772
rect 5859 26741 5871 26744
rect 5813 26735 5871 26741
rect 6730 26732 6736 26744
rect 6788 26732 6794 26784
rect 8386 26772 8392 26784
rect 8347 26744 8392 26772
rect 8386 26732 8392 26744
rect 8444 26732 8450 26784
rect 8570 26772 8576 26784
rect 8531 26744 8576 26772
rect 8570 26732 8576 26744
rect 8628 26732 8634 26784
rect 13722 26732 13728 26784
rect 13780 26772 13786 26784
rect 17218 26772 17224 26784
rect 13780 26744 17224 26772
rect 13780 26732 13786 26744
rect 17218 26732 17224 26744
rect 17276 26732 17282 26784
rect 19797 26775 19855 26781
rect 19797 26741 19809 26775
rect 19843 26772 19855 26775
rect 19904 26772 19932 26871
rect 20622 26868 20628 26920
rect 20680 26908 20686 26920
rect 20809 26911 20867 26917
rect 20680 26880 20725 26908
rect 20680 26868 20686 26880
rect 20809 26877 20821 26911
rect 20855 26908 20867 26911
rect 20855 26880 21496 26908
rect 20855 26877 20867 26880
rect 20809 26871 20867 26877
rect 20162 26800 20168 26852
rect 20220 26840 20226 26852
rect 20824 26840 20852 26871
rect 20220 26812 20852 26840
rect 20220 26800 20226 26812
rect 20714 26772 20720 26784
rect 19843 26744 20720 26772
rect 19843 26741 19855 26744
rect 19797 26735 19855 26741
rect 20714 26732 20720 26744
rect 20772 26732 20778 26784
rect 21468 26781 21496 26880
rect 21453 26775 21511 26781
rect 21453 26741 21465 26775
rect 21499 26772 21511 26775
rect 23290 26772 23296 26784
rect 21499 26744 23296 26772
rect 21499 26741 21511 26744
rect 21453 26735 21511 26741
rect 23290 26732 23296 26744
rect 23348 26732 23354 26784
rect 1104 26682 24656 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 24656 26682
rect 1104 26608 24656 26630
rect 3326 26528 3332 26580
rect 3384 26568 3390 26580
rect 3510 26568 3516 26580
rect 3384 26540 3516 26568
rect 3384 26528 3390 26540
rect 3510 26528 3516 26540
rect 3568 26528 3574 26580
rect 10781 26571 10839 26577
rect 10781 26537 10793 26571
rect 10827 26568 10839 26571
rect 10962 26568 10968 26580
rect 10827 26540 10968 26568
rect 10827 26537 10839 26540
rect 10781 26531 10839 26537
rect 10962 26528 10968 26540
rect 11020 26528 11026 26580
rect 11701 26571 11759 26577
rect 11701 26537 11713 26571
rect 11747 26568 11759 26571
rect 12526 26568 12532 26580
rect 11747 26540 12532 26568
rect 11747 26537 11759 26540
rect 11701 26531 11759 26537
rect 8297 26503 8355 26509
rect 8297 26469 8309 26503
rect 8343 26500 8355 26503
rect 8570 26500 8576 26512
rect 8343 26472 8576 26500
rect 8343 26469 8355 26472
rect 8297 26463 8355 26469
rect 6730 26432 6736 26444
rect 6691 26404 6736 26432
rect 6730 26392 6736 26404
rect 6788 26392 6794 26444
rect 6457 26367 6515 26373
rect 6457 26333 6469 26367
rect 6503 26364 6515 26367
rect 6822 26364 6828 26376
rect 6503 26336 6828 26364
rect 6503 26333 6515 26336
rect 6457 26327 6515 26333
rect 6822 26324 6828 26336
rect 6880 26364 6886 26376
rect 8312 26364 8340 26463
rect 8570 26460 8576 26472
rect 8628 26500 8634 26512
rect 11716 26500 11744 26531
rect 12526 26528 12532 26540
rect 12584 26528 12590 26580
rect 24302 26568 24308 26580
rect 15488 26540 24308 26568
rect 8628 26472 11744 26500
rect 8628 26460 8634 26472
rect 12434 26460 12440 26512
rect 12492 26500 12498 26512
rect 12805 26503 12863 26509
rect 12805 26500 12817 26503
rect 12492 26472 12817 26500
rect 12492 26460 12498 26472
rect 12805 26469 12817 26472
rect 12851 26500 12863 26503
rect 15381 26503 15439 26509
rect 15381 26500 15393 26503
rect 12851 26472 13032 26500
rect 12851 26469 12863 26472
rect 12805 26463 12863 26469
rect 10597 26435 10655 26441
rect 10597 26432 10609 26435
rect 6880 26336 8340 26364
rect 10428 26404 10609 26432
rect 6880 26324 6886 26336
rect 10226 26256 10232 26308
rect 10284 26296 10290 26308
rect 10428 26305 10456 26404
rect 10597 26401 10609 26404
rect 10643 26401 10655 26435
rect 10597 26395 10655 26401
rect 11885 26435 11943 26441
rect 11885 26401 11897 26435
rect 11931 26432 11943 26435
rect 12342 26432 12348 26444
rect 11931 26404 12348 26432
rect 11931 26401 11943 26404
rect 11885 26395 11943 26401
rect 12342 26392 12348 26404
rect 12400 26392 12406 26444
rect 13004 26441 13032 26472
rect 13924 26472 15393 26500
rect 12989 26435 13047 26441
rect 12989 26401 13001 26435
rect 13035 26401 13047 26435
rect 12989 26395 13047 26401
rect 13173 26435 13231 26441
rect 13173 26401 13185 26435
rect 13219 26432 13231 26435
rect 13722 26432 13728 26444
rect 13219 26404 13728 26432
rect 13219 26401 13231 26404
rect 13173 26395 13231 26401
rect 13722 26392 13728 26404
rect 13780 26392 13786 26444
rect 13924 26441 13952 26472
rect 15381 26469 15393 26472
rect 15427 26469 15439 26503
rect 15381 26463 15439 26469
rect 13909 26435 13967 26441
rect 13909 26401 13921 26435
rect 13955 26401 13967 26435
rect 15286 26432 15292 26444
rect 15199 26404 15292 26432
rect 13909 26395 13967 26401
rect 15286 26392 15292 26404
rect 15344 26432 15350 26444
rect 15488 26432 15516 26540
rect 24302 26528 24308 26540
rect 24360 26528 24366 26580
rect 19242 26500 19248 26512
rect 19155 26472 19248 26500
rect 19242 26460 19248 26472
rect 19300 26500 19306 26512
rect 23382 26500 23388 26512
rect 19300 26472 23388 26500
rect 19300 26460 19306 26472
rect 23382 26460 23388 26472
rect 23440 26460 23446 26512
rect 17862 26432 17868 26444
rect 15344 26404 15516 26432
rect 17823 26404 17868 26432
rect 15344 26392 15350 26404
rect 17862 26392 17868 26404
rect 17920 26392 17926 26444
rect 19334 26392 19340 26444
rect 19392 26432 19398 26444
rect 20530 26432 20536 26444
rect 19392 26404 20536 26432
rect 19392 26392 19398 26404
rect 20530 26392 20536 26404
rect 20588 26432 20594 26444
rect 20901 26435 20959 26441
rect 20901 26432 20913 26435
rect 20588 26404 20913 26432
rect 20588 26392 20594 26404
rect 20901 26401 20913 26404
rect 20947 26401 20959 26435
rect 23198 26432 23204 26444
rect 23159 26404 23204 26432
rect 20901 26395 20959 26401
rect 23198 26392 23204 26404
rect 23256 26392 23262 26444
rect 23290 26392 23296 26444
rect 23348 26432 23354 26444
rect 24854 26432 24860 26444
rect 23348 26404 24860 26432
rect 23348 26392 23354 26404
rect 24854 26392 24860 26404
rect 24912 26392 24918 26444
rect 17589 26367 17647 26373
rect 17589 26333 17601 26367
rect 17635 26364 17647 26367
rect 19426 26364 19432 26376
rect 17635 26336 19432 26364
rect 17635 26333 17647 26336
rect 17589 26327 17647 26333
rect 19426 26324 19432 26336
rect 19484 26324 19490 26376
rect 10413 26299 10471 26305
rect 10413 26296 10425 26299
rect 10284 26268 10425 26296
rect 10284 26256 10290 26268
rect 10413 26265 10425 26268
rect 10459 26265 10471 26299
rect 10413 26259 10471 26265
rect 13814 26256 13820 26308
rect 13872 26296 13878 26308
rect 14093 26299 14151 26305
rect 14093 26296 14105 26299
rect 13872 26268 14105 26296
rect 13872 26256 13878 26268
rect 14093 26265 14105 26268
rect 14139 26265 14151 26299
rect 14093 26259 14151 26265
rect 8018 26228 8024 26240
rect 7979 26200 8024 26228
rect 8018 26188 8024 26200
rect 8076 26188 8082 26240
rect 12434 26188 12440 26240
rect 12492 26228 12498 26240
rect 18230 26228 18236 26240
rect 12492 26200 18236 26228
rect 12492 26188 12498 26200
rect 18230 26188 18236 26200
rect 18288 26188 18294 26240
rect 21082 26228 21088 26240
rect 21043 26200 21088 26228
rect 21082 26188 21088 26200
rect 21140 26188 21146 26240
rect 1104 26138 24656 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 24656 26138
rect 1104 26064 24656 26086
rect 4062 25984 4068 26036
rect 4120 26024 4126 26036
rect 12434 26024 12440 26036
rect 4120 25996 12440 26024
rect 4120 25984 4126 25996
rect 12434 25984 12440 25996
rect 12492 25984 12498 26036
rect 12526 25984 12532 26036
rect 12584 26024 12590 26036
rect 13357 26027 13415 26033
rect 13357 26024 13369 26027
rect 12584 25996 13369 26024
rect 12584 25984 12590 25996
rect 13357 25993 13369 25996
rect 13403 25993 13415 26027
rect 13357 25987 13415 25993
rect 15105 26027 15163 26033
rect 15105 25993 15117 26027
rect 15151 26024 15163 26027
rect 15286 26024 15292 26036
rect 15151 25996 15292 26024
rect 15151 25993 15163 25996
rect 15105 25987 15163 25993
rect 4341 25959 4399 25965
rect 4341 25925 4353 25959
rect 4387 25956 4399 25959
rect 4614 25956 4620 25968
rect 4387 25928 4620 25956
rect 4387 25925 4399 25928
rect 4341 25919 4399 25925
rect 2777 25891 2835 25897
rect 2777 25857 2789 25891
rect 2823 25888 2835 25891
rect 2958 25888 2964 25900
rect 2823 25860 2964 25888
rect 2823 25857 2835 25860
rect 2777 25851 2835 25857
rect 2958 25848 2964 25860
rect 3016 25848 3022 25900
rect 2498 25820 2504 25832
rect 2411 25792 2504 25820
rect 2498 25780 2504 25792
rect 2556 25820 2562 25832
rect 4356 25820 4384 25919
rect 4614 25916 4620 25928
rect 4672 25916 4678 25968
rect 12621 25959 12679 25965
rect 12621 25925 12633 25959
rect 12667 25925 12679 25959
rect 12621 25919 12679 25925
rect 7834 25848 7840 25900
rect 7892 25888 7898 25900
rect 7892 25860 8156 25888
rect 7892 25848 7898 25860
rect 8128 25829 8156 25860
rect 2556 25792 4384 25820
rect 7929 25823 7987 25829
rect 2556 25780 2562 25792
rect 7929 25789 7941 25823
rect 7975 25789 7987 25823
rect 7929 25783 7987 25789
rect 8113 25823 8171 25829
rect 8113 25789 8125 25823
rect 8159 25789 8171 25823
rect 8113 25783 8171 25789
rect 7944 25752 7972 25783
rect 12434 25780 12440 25832
rect 12492 25820 12498 25832
rect 12636 25820 12664 25919
rect 13372 25888 13400 25987
rect 15286 25984 15292 25996
rect 15344 25984 15350 26036
rect 13541 25891 13599 25897
rect 13541 25888 13553 25891
rect 13372 25860 13553 25888
rect 13541 25857 13553 25860
rect 13587 25857 13599 25891
rect 13814 25888 13820 25900
rect 13775 25860 13820 25888
rect 13541 25851 13599 25857
rect 13814 25848 13820 25860
rect 13872 25848 13878 25900
rect 13998 25888 14004 25900
rect 13924 25860 14004 25888
rect 13924 25820 13952 25860
rect 13998 25848 14004 25860
rect 14056 25848 14062 25900
rect 12492 25792 12537 25820
rect 12636 25792 13952 25820
rect 12492 25780 12498 25792
rect 19426 25780 19432 25832
rect 19484 25820 19490 25832
rect 19613 25823 19671 25829
rect 19613 25820 19625 25823
rect 19484 25792 19625 25820
rect 19484 25780 19490 25792
rect 19613 25789 19625 25792
rect 19659 25789 19671 25823
rect 19886 25820 19892 25832
rect 19847 25792 19892 25820
rect 19613 25783 19671 25789
rect 8018 25752 8024 25764
rect 7931 25724 8024 25752
rect 8018 25712 8024 25724
rect 8076 25752 8082 25764
rect 8076 25724 8616 25752
rect 8076 25712 8082 25724
rect 8588 25696 8616 25724
rect 3878 25684 3884 25696
rect 3839 25656 3884 25684
rect 3878 25644 3884 25656
rect 3936 25644 3942 25696
rect 7926 25684 7932 25696
rect 7887 25656 7932 25684
rect 7926 25644 7932 25656
rect 7984 25644 7990 25696
rect 8570 25684 8576 25696
rect 8531 25656 8576 25684
rect 8570 25644 8576 25656
rect 8628 25644 8634 25696
rect 19521 25687 19579 25693
rect 19521 25653 19533 25687
rect 19567 25684 19579 25687
rect 19628 25684 19656 25783
rect 19886 25780 19892 25792
rect 19944 25780 19950 25832
rect 20806 25684 20812 25696
rect 19567 25656 20812 25684
rect 19567 25653 19579 25656
rect 19521 25647 19579 25653
rect 20806 25644 20812 25656
rect 20864 25644 20870 25696
rect 20898 25644 20904 25696
rect 20956 25684 20962 25696
rect 20993 25687 21051 25693
rect 20993 25684 21005 25687
rect 20956 25656 21005 25684
rect 20956 25644 20962 25656
rect 20993 25653 21005 25656
rect 21039 25684 21051 25687
rect 24762 25684 24768 25696
rect 21039 25656 24768 25684
rect 21039 25653 21051 25656
rect 20993 25647 21051 25653
rect 24762 25644 24768 25656
rect 24820 25644 24826 25696
rect 1104 25594 24656 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 24656 25594
rect 1104 25520 24656 25542
rect 8570 25440 8576 25492
rect 8628 25480 8634 25492
rect 21082 25480 21088 25492
rect 8628 25452 18644 25480
rect 8628 25440 8634 25452
rect 7377 25415 7435 25421
rect 7377 25381 7389 25415
rect 7423 25412 7435 25415
rect 7466 25412 7472 25424
rect 7423 25384 7472 25412
rect 7423 25381 7435 25384
rect 7377 25375 7435 25381
rect 7466 25372 7472 25384
rect 7524 25372 7530 25424
rect 10226 25372 10232 25424
rect 10284 25412 10290 25424
rect 12805 25415 12863 25421
rect 12805 25412 12817 25415
rect 10284 25384 12817 25412
rect 10284 25372 10290 25384
rect 12805 25381 12817 25384
rect 12851 25412 12863 25415
rect 13541 25415 13599 25421
rect 12851 25384 13216 25412
rect 12851 25381 12863 25384
rect 12805 25375 12863 25381
rect 3510 25304 3516 25356
rect 3568 25344 3574 25356
rect 3970 25344 3976 25356
rect 3568 25316 3976 25344
rect 3568 25304 3574 25316
rect 3970 25304 3976 25316
rect 4028 25304 4034 25356
rect 11701 25347 11759 25353
rect 11701 25313 11713 25347
rect 11747 25313 11759 25347
rect 11882 25344 11888 25356
rect 11843 25316 11888 25344
rect 11701 25307 11759 25313
rect 5721 25279 5779 25285
rect 5721 25245 5733 25279
rect 5767 25245 5779 25279
rect 5994 25276 6000 25288
rect 5955 25248 6000 25276
rect 5721 25239 5779 25245
rect 5736 25140 5764 25239
rect 5994 25236 6000 25248
rect 6052 25236 6058 25288
rect 11716 25208 11744 25307
rect 11882 25304 11888 25316
rect 11940 25344 11946 25356
rect 13188 25353 13216 25384
rect 13541 25381 13553 25415
rect 13587 25412 13599 25415
rect 14182 25412 14188 25424
rect 13587 25384 14188 25412
rect 13587 25381 13599 25384
rect 13541 25375 13599 25381
rect 14182 25372 14188 25384
rect 14240 25372 14246 25424
rect 12989 25347 13047 25353
rect 12989 25344 13001 25347
rect 11940 25316 13001 25344
rect 11940 25304 11946 25316
rect 12989 25313 13001 25316
rect 13035 25313 13047 25347
rect 12989 25307 13047 25313
rect 13173 25347 13231 25353
rect 13173 25313 13185 25347
rect 13219 25313 13231 25347
rect 13173 25307 13231 25313
rect 14553 25347 14611 25353
rect 14553 25313 14565 25347
rect 14599 25344 14611 25347
rect 16574 25344 16580 25356
rect 14599 25316 16580 25344
rect 14599 25313 14611 25316
rect 14553 25307 14611 25313
rect 16574 25304 16580 25316
rect 16632 25304 16638 25356
rect 17218 25304 17224 25356
rect 17276 25344 17282 25356
rect 18509 25347 18567 25353
rect 18509 25344 18521 25347
rect 17276 25316 18521 25344
rect 17276 25304 17282 25316
rect 18509 25313 18521 25316
rect 18555 25313 18567 25347
rect 18509 25307 18567 25313
rect 11974 25276 11980 25288
rect 11935 25248 11980 25276
rect 11974 25236 11980 25248
rect 12032 25236 12038 25288
rect 12710 25236 12716 25288
rect 12768 25276 12774 25288
rect 18233 25279 18291 25285
rect 18233 25276 18245 25279
rect 12768 25248 18245 25276
rect 12768 25236 12774 25248
rect 18233 25245 18245 25248
rect 18279 25276 18291 25279
rect 18325 25279 18383 25285
rect 18325 25276 18337 25279
rect 18279 25248 18337 25276
rect 18279 25245 18291 25248
rect 18233 25239 18291 25245
rect 18325 25245 18337 25248
rect 18371 25245 18383 25279
rect 18325 25239 18383 25245
rect 12253 25211 12311 25217
rect 12253 25208 12265 25211
rect 11716 25180 12265 25208
rect 12253 25177 12265 25180
rect 12299 25177 12311 25211
rect 12253 25171 12311 25177
rect 7561 25143 7619 25149
rect 7561 25140 7573 25143
rect 5736 25112 7573 25140
rect 7561 25109 7573 25112
rect 7607 25140 7619 25143
rect 7926 25140 7932 25152
rect 7607 25112 7932 25140
rect 7607 25109 7619 25112
rect 7561 25103 7619 25109
rect 7926 25100 7932 25112
rect 7984 25100 7990 25152
rect 12268 25140 12296 25171
rect 12342 25168 12348 25220
rect 12400 25208 12406 25220
rect 14369 25211 14427 25217
rect 14369 25208 14381 25211
rect 12400 25180 14381 25208
rect 12400 25168 12406 25180
rect 14369 25177 14381 25180
rect 14415 25177 14427 25211
rect 18616 25208 18644 25452
rect 19076 25452 21088 25480
rect 19076 25353 19104 25452
rect 21082 25440 21088 25452
rect 21140 25440 21146 25492
rect 19613 25415 19671 25421
rect 19613 25381 19625 25415
rect 19659 25412 19671 25415
rect 19886 25412 19892 25424
rect 19659 25384 19892 25412
rect 19659 25381 19671 25384
rect 19613 25375 19671 25381
rect 19886 25372 19892 25384
rect 19944 25372 19950 25424
rect 19061 25347 19119 25353
rect 19061 25313 19073 25347
rect 19107 25313 19119 25347
rect 19061 25307 19119 25313
rect 19245 25347 19303 25353
rect 19245 25313 19257 25347
rect 19291 25344 19303 25347
rect 20622 25344 20628 25356
rect 19291 25316 20628 25344
rect 19291 25313 19303 25316
rect 19245 25307 19303 25313
rect 20622 25304 20628 25316
rect 20680 25304 20686 25356
rect 21082 25344 21088 25356
rect 20995 25316 21088 25344
rect 21082 25304 21088 25316
rect 21140 25344 21146 25356
rect 21542 25344 21548 25356
rect 21140 25316 21548 25344
rect 21140 25304 21146 25316
rect 21542 25304 21548 25316
rect 21600 25344 21606 25356
rect 21637 25347 21695 25353
rect 21637 25344 21649 25347
rect 21600 25316 21649 25344
rect 21600 25304 21606 25316
rect 21637 25313 21649 25316
rect 21683 25313 21695 25347
rect 21818 25344 21824 25356
rect 21779 25316 21824 25344
rect 21637 25307 21695 25313
rect 21818 25304 21824 25316
rect 21876 25304 21882 25356
rect 20714 25236 20720 25288
rect 20772 25276 20778 25288
rect 20901 25279 20959 25285
rect 20901 25276 20913 25279
rect 20772 25248 20913 25276
rect 20772 25236 20778 25248
rect 20901 25245 20913 25248
rect 20947 25245 20959 25279
rect 20901 25239 20959 25245
rect 22002 25208 22008 25220
rect 18616 25180 22008 25208
rect 14369 25171 14427 25177
rect 22002 25168 22008 25180
rect 22060 25168 22066 25220
rect 12710 25140 12716 25152
rect 12268 25112 12716 25140
rect 12710 25100 12716 25112
rect 12768 25100 12774 25152
rect 20714 25140 20720 25152
rect 20675 25112 20720 25140
rect 20714 25100 20720 25112
rect 20772 25100 20778 25152
rect 22094 25100 22100 25152
rect 22152 25140 22158 25152
rect 22152 25112 22197 25140
rect 22152 25100 22158 25112
rect 1104 25050 24656 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 24656 25050
rect 1104 24976 24656 24998
rect 2777 24803 2835 24809
rect 2777 24769 2789 24803
rect 2823 24800 2835 24803
rect 4341 24803 4399 24809
rect 4341 24800 4353 24803
rect 2823 24772 4353 24800
rect 2823 24769 2835 24772
rect 2777 24763 2835 24769
rect 4341 24769 4353 24772
rect 4387 24800 4399 24803
rect 4890 24800 4896 24812
rect 4387 24772 4896 24800
rect 4387 24769 4399 24772
rect 4341 24763 4399 24769
rect 4890 24760 4896 24772
rect 4948 24760 4954 24812
rect 6825 24803 6883 24809
rect 6825 24769 6837 24803
rect 6871 24800 6883 24803
rect 7926 24800 7932 24812
rect 6871 24772 7932 24800
rect 6871 24769 6883 24772
rect 6825 24763 6883 24769
rect 2498 24732 2504 24744
rect 2459 24704 2504 24732
rect 2498 24692 2504 24704
rect 2556 24692 2562 24744
rect 4525 24735 4583 24741
rect 4525 24701 4537 24735
rect 4571 24732 4583 24735
rect 6840 24732 6868 24763
rect 7926 24760 7932 24772
rect 7984 24760 7990 24812
rect 8478 24800 8484 24812
rect 8391 24772 8484 24800
rect 8478 24760 8484 24772
rect 8536 24800 8542 24812
rect 21361 24803 21419 24809
rect 8536 24772 21220 24800
rect 8536 24760 8542 24772
rect 7098 24732 7104 24744
rect 4571 24704 6868 24732
rect 7059 24704 7104 24732
rect 4571 24701 4583 24704
rect 4525 24695 4583 24701
rect 7098 24692 7104 24704
rect 7156 24692 7162 24744
rect 11425 24735 11483 24741
rect 11425 24701 11437 24735
rect 11471 24732 11483 24735
rect 12342 24732 12348 24744
rect 11471 24704 12348 24732
rect 11471 24701 11483 24704
rect 11425 24695 11483 24701
rect 12342 24692 12348 24704
rect 12400 24692 12406 24744
rect 12437 24735 12495 24741
rect 12437 24701 12449 24735
rect 12483 24732 12495 24735
rect 12618 24732 12624 24744
rect 12483 24704 12624 24732
rect 12483 24701 12495 24704
rect 12437 24695 12495 24701
rect 12618 24692 12624 24704
rect 12676 24692 12682 24744
rect 13541 24735 13599 24741
rect 13541 24701 13553 24735
rect 13587 24701 13599 24735
rect 13541 24695 13599 24701
rect 15289 24735 15347 24741
rect 15289 24701 15301 24735
rect 15335 24732 15347 24735
rect 15657 24735 15715 24741
rect 15657 24732 15669 24735
rect 15335 24704 15669 24732
rect 15335 24701 15347 24704
rect 15289 24695 15347 24701
rect 15657 24701 15669 24704
rect 15703 24732 15715 24735
rect 16482 24732 16488 24744
rect 15703 24704 16488 24732
rect 15703 24701 15715 24704
rect 15657 24695 15715 24701
rect 4062 24624 4068 24676
rect 4120 24664 4126 24676
rect 13446 24664 13452 24676
rect 4120 24636 4568 24664
rect 4120 24624 4126 24636
rect 3234 24556 3240 24608
rect 3292 24596 3298 24608
rect 3881 24599 3939 24605
rect 3881 24596 3893 24599
rect 3292 24568 3893 24596
rect 3292 24556 3298 24568
rect 3881 24565 3893 24568
rect 3927 24565 3939 24599
rect 4540 24596 4568 24636
rect 7760 24636 13308 24664
rect 13359 24636 13452 24664
rect 7760 24596 7788 24636
rect 4540 24568 7788 24596
rect 3881 24559 3939 24565
rect 7926 24556 7932 24608
rect 7984 24596 7990 24608
rect 8665 24599 8723 24605
rect 8665 24596 8677 24599
rect 7984 24568 8677 24596
rect 7984 24556 7990 24568
rect 8665 24565 8677 24568
rect 8711 24596 8723 24599
rect 9030 24596 9036 24608
rect 8711 24568 9036 24596
rect 8711 24565 8723 24568
rect 8665 24559 8723 24565
rect 9030 24556 9036 24568
rect 9088 24596 9094 24608
rect 11241 24599 11299 24605
rect 11241 24596 11253 24599
rect 9088 24568 11253 24596
rect 9088 24556 9094 24568
rect 11241 24565 11253 24568
rect 11287 24596 11299 24599
rect 11422 24596 11428 24608
rect 11287 24568 11428 24596
rect 11287 24565 11299 24568
rect 11241 24559 11299 24565
rect 11422 24556 11428 24568
rect 11480 24556 11486 24608
rect 12526 24596 12532 24608
rect 12487 24568 12532 24596
rect 12526 24556 12532 24568
rect 12584 24556 12590 24608
rect 12618 24556 12624 24608
rect 12676 24596 12682 24608
rect 12713 24599 12771 24605
rect 12713 24596 12725 24599
rect 12676 24568 12725 24596
rect 12676 24556 12682 24568
rect 12713 24565 12725 24568
rect 12759 24565 12771 24599
rect 13280 24596 13308 24636
rect 13446 24624 13452 24636
rect 13504 24664 13510 24676
rect 13556 24664 13584 24695
rect 16482 24692 16488 24704
rect 16540 24692 16546 24744
rect 19337 24735 19395 24741
rect 19337 24701 19349 24735
rect 19383 24701 19395 24735
rect 21085 24735 21143 24741
rect 21085 24732 21097 24735
rect 19337 24695 19395 24701
rect 20916 24704 21097 24732
rect 19352 24664 19380 24695
rect 13504 24636 19380 24664
rect 13504 24624 13510 24636
rect 19352 24608 19380 24636
rect 13538 24596 13544 24608
rect 13280 24568 13544 24596
rect 12713 24559 12771 24565
rect 13538 24556 13544 24568
rect 13596 24556 13602 24608
rect 13722 24596 13728 24608
rect 13683 24568 13728 24596
rect 13722 24556 13728 24568
rect 13780 24556 13786 24608
rect 14642 24556 14648 24608
rect 14700 24596 14706 24608
rect 15381 24599 15439 24605
rect 15381 24596 15393 24599
rect 14700 24568 15393 24596
rect 14700 24556 14706 24568
rect 15381 24565 15393 24568
rect 15427 24565 15439 24599
rect 15381 24559 15439 24565
rect 19245 24599 19303 24605
rect 19245 24565 19257 24599
rect 19291 24596 19303 24599
rect 19334 24596 19340 24608
rect 19291 24568 19340 24596
rect 19291 24565 19303 24568
rect 19245 24559 19303 24565
rect 19334 24556 19340 24568
rect 19392 24556 19398 24608
rect 19521 24599 19579 24605
rect 19521 24565 19533 24599
rect 19567 24596 19579 24599
rect 20530 24596 20536 24608
rect 19567 24568 20536 24596
rect 19567 24565 19579 24568
rect 19521 24559 19579 24565
rect 20530 24556 20536 24568
rect 20588 24556 20594 24608
rect 20806 24556 20812 24608
rect 20864 24596 20870 24608
rect 20916 24605 20944 24704
rect 21085 24701 21097 24704
rect 21131 24701 21143 24735
rect 21192 24732 21220 24772
rect 21361 24769 21373 24803
rect 21407 24800 21419 24803
rect 22094 24800 22100 24812
rect 21407 24772 22100 24800
rect 21407 24769 21419 24772
rect 21361 24763 21419 24769
rect 22094 24760 22100 24772
rect 22152 24760 22158 24812
rect 26786 24732 26792 24744
rect 21192 24704 26792 24732
rect 21085 24695 21143 24701
rect 26786 24692 26792 24704
rect 26844 24692 26850 24744
rect 22741 24667 22799 24673
rect 22741 24633 22753 24667
rect 22787 24664 22799 24667
rect 23566 24664 23572 24676
rect 22787 24636 23572 24664
rect 22787 24633 22799 24636
rect 22741 24627 22799 24633
rect 23566 24624 23572 24636
rect 23624 24624 23630 24676
rect 20901 24599 20959 24605
rect 20901 24596 20913 24599
rect 20864 24568 20913 24596
rect 20864 24556 20870 24568
rect 20901 24565 20913 24568
rect 20947 24565 20959 24599
rect 20901 24559 20959 24565
rect 1104 24506 24656 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 24656 24506
rect 1104 24432 24656 24454
rect 5994 24352 6000 24404
rect 6052 24392 6058 24404
rect 6457 24395 6515 24401
rect 6457 24392 6469 24395
rect 6052 24364 6469 24392
rect 6052 24352 6058 24364
rect 6457 24361 6469 24364
rect 6503 24361 6515 24395
rect 6457 24355 6515 24361
rect 7377 24395 7435 24401
rect 7377 24361 7389 24395
rect 7423 24392 7435 24395
rect 7466 24392 7472 24404
rect 7423 24364 7472 24392
rect 7423 24361 7435 24364
rect 7377 24355 7435 24361
rect 7466 24352 7472 24364
rect 7524 24352 7530 24404
rect 12342 24352 12348 24404
rect 12400 24392 12406 24404
rect 13446 24392 13452 24404
rect 12400 24364 13452 24392
rect 12400 24352 12406 24364
rect 13446 24352 13452 24364
rect 13504 24352 13510 24404
rect 13538 24352 13544 24404
rect 13596 24392 13602 24404
rect 17310 24392 17316 24404
rect 13596 24364 17316 24392
rect 13596 24352 13602 24364
rect 17310 24352 17316 24364
rect 17368 24352 17374 24404
rect 19521 24395 19579 24401
rect 19521 24361 19533 24395
rect 19567 24392 19579 24395
rect 20162 24392 20168 24404
rect 19567 24364 20168 24392
rect 19567 24361 19579 24364
rect 19521 24355 19579 24361
rect 7006 24324 7012 24336
rect 6196 24296 7012 24324
rect 5445 24259 5503 24265
rect 5445 24225 5457 24259
rect 5491 24256 5503 24259
rect 5997 24259 6055 24265
rect 5997 24256 6009 24259
rect 5491 24228 6009 24256
rect 5491 24225 5503 24228
rect 5445 24219 5503 24225
rect 5997 24225 6009 24228
rect 6043 24256 6055 24259
rect 6086 24256 6092 24268
rect 6043 24228 6092 24256
rect 6043 24225 6055 24228
rect 5997 24219 6055 24225
rect 6086 24216 6092 24228
rect 6144 24216 6150 24268
rect 6196 24265 6224 24296
rect 7006 24284 7012 24296
rect 7064 24324 7070 24336
rect 7561 24327 7619 24333
rect 7561 24324 7573 24327
rect 7064 24296 7573 24324
rect 7064 24284 7070 24296
rect 7561 24293 7573 24296
rect 7607 24293 7619 24327
rect 7561 24287 7619 24293
rect 12710 24284 12716 24336
rect 12768 24324 12774 24336
rect 18322 24324 18328 24336
rect 12768 24296 15424 24324
rect 12768 24284 12774 24296
rect 6181 24259 6239 24265
rect 6181 24225 6193 24259
rect 6227 24225 6239 24259
rect 7466 24256 7472 24268
rect 7427 24228 7472 24256
rect 6181 24219 6239 24225
rect 7466 24216 7472 24228
rect 7524 24216 7530 24268
rect 10873 24259 10931 24265
rect 10873 24225 10885 24259
rect 10919 24256 10931 24259
rect 11422 24256 11428 24268
rect 10919 24228 11428 24256
rect 10919 24225 10931 24228
rect 10873 24219 10931 24225
rect 11422 24216 11428 24228
rect 11480 24256 11486 24268
rect 15396 24256 15424 24296
rect 17788 24296 18328 24324
rect 17788 24265 17816 24296
rect 18322 24284 18328 24296
rect 18380 24324 18386 24336
rect 18380 24296 19196 24324
rect 18380 24284 18386 24296
rect 17773 24259 17831 24265
rect 17773 24256 17785 24259
rect 11480 24228 12756 24256
rect 15396 24228 17785 24256
rect 11480 24216 11486 24228
rect 5169 24191 5227 24197
rect 5169 24157 5181 24191
rect 5215 24188 5227 24191
rect 5353 24191 5411 24197
rect 5353 24188 5365 24191
rect 5215 24160 5365 24188
rect 5215 24157 5227 24160
rect 5169 24151 5227 24157
rect 5353 24157 5365 24160
rect 5399 24157 5411 24191
rect 5353 24151 5411 24157
rect 11149 24191 11207 24197
rect 11149 24157 11161 24191
rect 11195 24188 11207 24191
rect 11238 24188 11244 24200
rect 11195 24160 11244 24188
rect 11195 24157 11207 24160
rect 11149 24151 11207 24157
rect 5368 24120 5396 24151
rect 11238 24148 11244 24160
rect 11296 24148 11302 24200
rect 6638 24120 6644 24132
rect 5368 24092 6644 24120
rect 6638 24080 6644 24092
rect 6696 24120 6702 24132
rect 6822 24120 6828 24132
rect 6696 24092 6828 24120
rect 6696 24080 6702 24092
rect 6822 24080 6828 24092
rect 6880 24080 6886 24132
rect 12437 24055 12495 24061
rect 12437 24021 12449 24055
rect 12483 24052 12495 24055
rect 12618 24052 12624 24064
rect 12483 24024 12624 24052
rect 12483 24021 12495 24024
rect 12437 24015 12495 24021
rect 12618 24012 12624 24024
rect 12676 24012 12682 24064
rect 12728 24061 12756 24228
rect 17773 24225 17785 24228
rect 17819 24225 17831 24259
rect 17773 24219 17831 24225
rect 18049 24259 18107 24265
rect 18049 24225 18061 24259
rect 18095 24256 18107 24259
rect 18414 24256 18420 24268
rect 18095 24228 18420 24256
rect 18095 24225 18107 24228
rect 18049 24219 18107 24225
rect 18414 24216 18420 24228
rect 18472 24256 18478 24268
rect 19168 24265 19196 24296
rect 18785 24259 18843 24265
rect 18785 24256 18797 24259
rect 18472 24228 18797 24256
rect 18472 24216 18478 24228
rect 18785 24225 18797 24228
rect 18831 24225 18843 24259
rect 18785 24219 18843 24225
rect 19153 24259 19211 24265
rect 19153 24225 19165 24259
rect 19199 24225 19211 24259
rect 19153 24219 19211 24225
rect 19337 24259 19395 24265
rect 19337 24225 19349 24259
rect 19383 24256 19395 24259
rect 19536 24256 19564 24355
rect 20162 24352 20168 24364
rect 20220 24352 20226 24404
rect 20622 24352 20628 24404
rect 20680 24392 20686 24404
rect 20993 24395 21051 24401
rect 20993 24392 21005 24395
rect 20680 24364 21005 24392
rect 20680 24352 20686 24364
rect 20993 24361 21005 24364
rect 21039 24361 21051 24395
rect 20993 24355 21051 24361
rect 21818 24352 21824 24404
rect 21876 24392 21882 24404
rect 22005 24395 22063 24401
rect 22005 24392 22017 24395
rect 21876 24364 22017 24392
rect 21876 24352 21882 24364
rect 22005 24361 22017 24364
rect 22051 24361 22063 24395
rect 22005 24355 22063 24361
rect 23566 24324 23572 24336
rect 23032 24296 23572 24324
rect 20898 24256 20904 24268
rect 19383 24228 19564 24256
rect 20859 24228 20904 24256
rect 19383 24225 19395 24228
rect 19337 24219 19395 24225
rect 20898 24216 20904 24228
rect 20956 24216 20962 24268
rect 21913 24259 21971 24265
rect 21913 24225 21925 24259
rect 21959 24256 21971 24259
rect 23032 24256 23060 24296
rect 23566 24284 23572 24296
rect 23624 24284 23630 24336
rect 21959 24228 23060 24256
rect 23109 24259 23167 24265
rect 21959 24225 21971 24228
rect 21913 24219 21971 24225
rect 23109 24225 23121 24259
rect 23155 24225 23167 24259
rect 23109 24219 23167 24225
rect 23385 24259 23443 24265
rect 23385 24225 23397 24259
rect 23431 24256 23443 24259
rect 23474 24256 23480 24268
rect 23431 24228 23480 24256
rect 23431 24225 23443 24228
rect 23385 24219 23443 24225
rect 15289 24191 15347 24197
rect 15289 24188 15301 24191
rect 15028 24160 15301 24188
rect 12713 24055 12771 24061
rect 12713 24021 12725 24055
rect 12759 24052 12771 24055
rect 12894 24052 12900 24064
rect 12759 24024 12900 24052
rect 12759 24021 12771 24024
rect 12713 24015 12771 24021
rect 12894 24012 12900 24024
rect 12952 24052 12958 24064
rect 15028 24061 15056 24160
rect 15289 24157 15301 24160
rect 15335 24157 15347 24191
rect 15562 24188 15568 24200
rect 15523 24160 15568 24188
rect 15289 24151 15347 24157
rect 15562 24148 15568 24160
rect 15620 24148 15626 24200
rect 16482 24148 16488 24200
rect 16540 24188 16546 24200
rect 16669 24191 16727 24197
rect 16669 24188 16681 24191
rect 16540 24160 16681 24188
rect 16540 24148 16546 24160
rect 16669 24157 16681 24160
rect 16715 24157 16727 24191
rect 16669 24151 16727 24157
rect 17034 24148 17040 24200
rect 17092 24188 17098 24200
rect 18141 24191 18199 24197
rect 18141 24188 18153 24191
rect 17092 24160 18153 24188
rect 17092 24148 17098 24160
rect 18141 24157 18153 24160
rect 18187 24157 18199 24191
rect 18874 24188 18880 24200
rect 18835 24160 18880 24188
rect 18141 24151 18199 24157
rect 18874 24148 18880 24160
rect 18932 24148 18938 24200
rect 23124 24188 23152 24219
rect 23474 24216 23480 24228
rect 23532 24216 23538 24268
rect 53834 24216 53840 24268
rect 53892 24256 53898 24268
rect 54754 24256 54760 24268
rect 53892 24228 54760 24256
rect 53892 24216 53898 24228
rect 54754 24216 54760 24228
rect 54812 24216 54818 24268
rect 24118 24188 24124 24200
rect 23124 24160 24124 24188
rect 24118 24148 24124 24160
rect 24176 24148 24182 24200
rect 16574 24080 16580 24132
rect 16632 24120 16638 24132
rect 22925 24123 22983 24129
rect 22925 24120 22937 24123
rect 16632 24092 22937 24120
rect 16632 24080 16638 24092
rect 22925 24089 22937 24092
rect 22971 24089 22983 24123
rect 22925 24083 22983 24089
rect 15013 24055 15071 24061
rect 15013 24052 15025 24055
rect 12952 24024 15025 24052
rect 12952 24012 12958 24024
rect 15013 24021 15025 24024
rect 15059 24021 15071 24055
rect 15013 24015 15071 24021
rect 22278 24012 22284 24064
rect 22336 24052 22342 24064
rect 23477 24055 23535 24061
rect 23477 24052 23489 24055
rect 22336 24024 23489 24052
rect 22336 24012 22342 24024
rect 23477 24021 23489 24024
rect 23523 24021 23535 24055
rect 23477 24015 23535 24021
rect 1104 23962 24656 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 24656 23962
rect 1104 23888 24656 23910
rect 7653 23851 7711 23857
rect 7653 23817 7665 23851
rect 7699 23848 7711 23851
rect 8478 23848 8484 23860
rect 7699 23820 8484 23848
rect 7699 23817 7711 23820
rect 7653 23811 7711 23817
rect 2774 23672 2780 23724
rect 2832 23712 2838 23724
rect 2832 23684 2877 23712
rect 2832 23672 2838 23684
rect 2498 23644 2504 23656
rect 2459 23616 2504 23644
rect 2498 23604 2504 23616
rect 2556 23604 2562 23656
rect 7285 23647 7343 23653
rect 7285 23613 7297 23647
rect 7331 23644 7343 23647
rect 7668 23644 7696 23811
rect 8478 23808 8484 23820
rect 8536 23808 8542 23860
rect 12250 23848 12256 23860
rect 8588 23820 12256 23848
rect 8018 23740 8024 23792
rect 8076 23780 8082 23792
rect 8588 23780 8616 23820
rect 12250 23808 12256 23820
rect 12308 23808 12314 23860
rect 12621 23851 12679 23857
rect 12621 23817 12633 23851
rect 12667 23848 12679 23851
rect 12710 23848 12716 23860
rect 12667 23820 12716 23848
rect 12667 23817 12679 23820
rect 12621 23811 12679 23817
rect 12710 23808 12716 23820
rect 12768 23808 12774 23860
rect 14921 23851 14979 23857
rect 14921 23817 14933 23851
rect 14967 23848 14979 23851
rect 15562 23848 15568 23860
rect 14967 23820 15568 23848
rect 14967 23817 14979 23820
rect 14921 23811 14979 23817
rect 15562 23808 15568 23820
rect 15620 23808 15626 23860
rect 18782 23808 18788 23860
rect 18840 23848 18846 23860
rect 20990 23848 20996 23860
rect 18840 23820 20996 23848
rect 18840 23808 18846 23820
rect 20990 23808 20996 23820
rect 21048 23848 21054 23860
rect 21177 23851 21235 23857
rect 21177 23848 21189 23851
rect 21048 23820 21189 23848
rect 21048 23808 21054 23820
rect 21177 23817 21189 23820
rect 21223 23817 21235 23851
rect 21177 23811 21235 23817
rect 8076 23752 8616 23780
rect 10045 23783 10103 23789
rect 8076 23740 8082 23752
rect 10045 23749 10057 23783
rect 10091 23780 10103 23783
rect 12802 23780 12808 23792
rect 10091 23752 12808 23780
rect 10091 23749 10103 23752
rect 10045 23743 10103 23749
rect 10244 23721 10272 23752
rect 12802 23740 12808 23752
rect 12860 23740 12866 23792
rect 20714 23780 20720 23792
rect 18064 23752 20720 23780
rect 10229 23715 10287 23721
rect 10229 23681 10241 23715
rect 10275 23681 10287 23715
rect 11333 23715 11391 23721
rect 11333 23712 11345 23715
rect 10229 23675 10287 23681
rect 11256 23684 11345 23712
rect 11256 23656 11284 23684
rect 11333 23681 11345 23684
rect 11379 23681 11391 23715
rect 11333 23675 11391 23681
rect 12250 23672 12256 23724
rect 12308 23712 12314 23724
rect 13541 23715 13599 23721
rect 13541 23712 13553 23715
rect 12308 23684 13553 23712
rect 12308 23672 12314 23684
rect 13541 23681 13553 23684
rect 13587 23712 13599 23715
rect 13630 23712 13636 23724
rect 13587 23684 13636 23712
rect 13587 23681 13599 23684
rect 13541 23675 13599 23681
rect 13630 23672 13636 23684
rect 13688 23712 13694 23724
rect 13725 23715 13783 23721
rect 13725 23712 13737 23715
rect 13688 23684 13737 23712
rect 13688 23672 13694 23684
rect 13725 23681 13737 23684
rect 13771 23681 13783 23715
rect 13725 23675 13783 23681
rect 17770 23672 17776 23724
rect 17828 23712 17834 23724
rect 18064 23721 18092 23752
rect 20714 23740 20720 23752
rect 20772 23740 20778 23792
rect 18049 23715 18107 23721
rect 18049 23712 18061 23715
rect 17828 23684 18061 23712
rect 17828 23672 17834 23684
rect 18049 23681 18061 23684
rect 18095 23681 18107 23715
rect 21192 23712 21220 23811
rect 21361 23715 21419 23721
rect 21361 23712 21373 23715
rect 21192 23684 21373 23712
rect 18049 23675 18107 23681
rect 21361 23681 21373 23684
rect 21407 23681 21419 23715
rect 21361 23675 21419 23681
rect 7331 23616 7696 23644
rect 7331 23613 7343 23616
rect 7285 23607 7343 23613
rect 9858 23604 9864 23656
rect 9916 23644 9922 23656
rect 10321 23647 10379 23653
rect 10321 23644 10333 23647
rect 9916 23616 10333 23644
rect 9916 23604 9922 23616
rect 10321 23613 10333 23616
rect 10367 23644 10379 23647
rect 10870 23644 10876 23656
rect 10367 23616 10876 23644
rect 10367 23613 10379 23616
rect 10321 23607 10379 23613
rect 10870 23604 10876 23616
rect 10928 23604 10934 23656
rect 11057 23647 11115 23653
rect 11057 23613 11069 23647
rect 11103 23613 11115 23647
rect 11057 23607 11115 23613
rect 11072 23576 11100 23607
rect 11238 23604 11244 23656
rect 11296 23604 11302 23656
rect 12434 23604 12440 23656
rect 12492 23644 12498 23656
rect 12802 23644 12808 23656
rect 12492 23616 12808 23644
rect 12492 23604 12498 23616
rect 12802 23604 12808 23616
rect 12860 23604 12866 23656
rect 13909 23647 13967 23653
rect 13909 23613 13921 23647
rect 13955 23613 13967 23647
rect 13909 23607 13967 23613
rect 12526 23576 12532 23588
rect 11072 23548 12532 23576
rect 12526 23536 12532 23548
rect 12584 23536 12590 23588
rect 13924 23576 13952 23607
rect 14458 23604 14464 23656
rect 14516 23644 14522 23656
rect 14642 23644 14648 23656
rect 14516 23616 14561 23644
rect 14603 23616 14648 23644
rect 14516 23604 14522 23616
rect 14642 23604 14648 23616
rect 14700 23604 14706 23656
rect 18233 23647 18291 23653
rect 18233 23644 18245 23647
rect 17052 23616 18245 23644
rect 14476 23576 14504 23604
rect 13464 23548 13860 23576
rect 13924 23548 14504 23576
rect 3878 23508 3884 23520
rect 3839 23480 3884 23508
rect 3878 23468 3884 23480
rect 3936 23468 3942 23520
rect 4341 23511 4399 23517
rect 4341 23477 4353 23511
rect 4387 23508 4399 23511
rect 4614 23508 4620 23520
rect 4387 23480 4620 23508
rect 4387 23477 4399 23480
rect 4341 23471 4399 23477
rect 4614 23468 4620 23480
rect 4672 23468 4678 23520
rect 6914 23468 6920 23520
rect 6972 23508 6978 23520
rect 7377 23511 7435 23517
rect 7377 23508 7389 23511
rect 6972 23480 7389 23508
rect 6972 23468 6978 23480
rect 7377 23477 7389 23480
rect 7423 23477 7435 23511
rect 7377 23471 7435 23477
rect 10870 23468 10876 23520
rect 10928 23508 10934 23520
rect 13464 23508 13492 23548
rect 10928 23480 13492 23508
rect 13832 23508 13860 23548
rect 17052 23508 17080 23616
rect 18233 23613 18245 23616
rect 18279 23613 18291 23647
rect 18233 23607 18291 23613
rect 18785 23647 18843 23653
rect 18785 23613 18797 23647
rect 18831 23613 18843 23647
rect 18785 23607 18843 23613
rect 18248 23576 18276 23607
rect 18598 23576 18604 23588
rect 18248 23548 18604 23576
rect 18598 23536 18604 23548
rect 18656 23576 18662 23588
rect 18800 23576 18828 23607
rect 18874 23604 18880 23656
rect 18932 23644 18938 23656
rect 18969 23647 19027 23653
rect 18969 23644 18981 23647
rect 18932 23616 18981 23644
rect 18932 23604 18938 23616
rect 18969 23613 18981 23616
rect 19015 23613 19027 23647
rect 18969 23607 19027 23613
rect 18656 23548 18828 23576
rect 18984 23576 19012 23607
rect 20162 23604 20168 23656
rect 20220 23644 20226 23656
rect 20257 23647 20315 23653
rect 20257 23644 20269 23647
rect 20220 23616 20269 23644
rect 20220 23604 20226 23616
rect 20257 23613 20269 23616
rect 20303 23613 20315 23647
rect 21542 23644 21548 23656
rect 21455 23616 21548 23644
rect 20257 23607 20315 23613
rect 21542 23604 21548 23616
rect 21600 23604 21606 23656
rect 22097 23647 22155 23653
rect 22097 23613 22109 23647
rect 22143 23613 22155 23647
rect 22278 23644 22284 23656
rect 22239 23616 22284 23644
rect 22097 23607 22155 23613
rect 20349 23579 20407 23585
rect 20349 23576 20361 23579
rect 18984 23548 20361 23576
rect 18656 23536 18662 23548
rect 20349 23545 20361 23548
rect 20395 23545 20407 23579
rect 21560 23576 21588 23604
rect 22112 23576 22140 23607
rect 22278 23604 22284 23616
rect 22336 23604 22342 23656
rect 21560 23548 22140 23576
rect 20349 23539 20407 23545
rect 17770 23508 17776 23520
rect 13832 23480 17080 23508
rect 17731 23480 17776 23508
rect 10928 23468 10934 23480
rect 17770 23468 17776 23480
rect 17828 23468 17834 23520
rect 19242 23508 19248 23520
rect 19203 23480 19248 23508
rect 19242 23468 19248 23480
rect 19300 23468 19306 23520
rect 20162 23508 20168 23520
rect 20123 23480 20168 23508
rect 20162 23468 20168 23480
rect 20220 23468 20226 23520
rect 22554 23508 22560 23520
rect 22515 23480 22560 23508
rect 22554 23468 22560 23480
rect 22612 23468 22618 23520
rect 1104 23418 24656 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 24656 23418
rect 1104 23344 24656 23366
rect 4062 23264 4068 23316
rect 4120 23304 4126 23316
rect 23014 23304 23020 23316
rect 4120 23276 23020 23304
rect 4120 23264 4126 23276
rect 23014 23264 23020 23276
rect 23072 23264 23078 23316
rect 6733 23239 6791 23245
rect 6733 23205 6745 23239
rect 6779 23236 6791 23239
rect 7098 23236 7104 23248
rect 6779 23208 7104 23236
rect 6779 23205 6791 23208
rect 6733 23199 6791 23205
rect 7098 23196 7104 23208
rect 7156 23196 7162 23248
rect 11701 23239 11759 23245
rect 11701 23205 11713 23239
rect 11747 23236 11759 23239
rect 12618 23236 12624 23248
rect 11747 23208 12624 23236
rect 11747 23205 11759 23208
rect 11701 23199 11759 23205
rect 5629 23171 5687 23177
rect 5629 23137 5641 23171
rect 5675 23168 5687 23171
rect 6178 23168 6184 23180
rect 5675 23140 6184 23168
rect 5675 23137 5687 23140
rect 5629 23131 5687 23137
rect 6178 23128 6184 23140
rect 6236 23128 6242 23180
rect 6365 23171 6423 23177
rect 6365 23137 6377 23171
rect 6411 23168 6423 23171
rect 6914 23168 6920 23180
rect 6411 23140 6920 23168
rect 6411 23137 6423 23140
rect 6365 23131 6423 23137
rect 6914 23128 6920 23140
rect 6972 23128 6978 23180
rect 7653 23171 7711 23177
rect 7653 23137 7665 23171
rect 7699 23168 7711 23171
rect 7742 23168 7748 23180
rect 7699 23140 7748 23168
rect 7699 23137 7711 23140
rect 7653 23131 7711 23137
rect 7742 23128 7748 23140
rect 7800 23128 7806 23180
rect 9677 23171 9735 23177
rect 9677 23137 9689 23171
rect 9723 23168 9735 23171
rect 11882 23168 11888 23180
rect 9723 23140 11888 23168
rect 9723 23137 9735 23140
rect 9677 23131 9735 23137
rect 11882 23128 11888 23140
rect 11940 23128 11946 23180
rect 12452 23177 12480 23208
rect 12618 23196 12624 23208
rect 12676 23196 12682 23248
rect 19705 23239 19763 23245
rect 19705 23205 19717 23239
rect 19751 23236 19763 23239
rect 20162 23236 20168 23248
rect 19751 23208 20168 23236
rect 19751 23205 19763 23208
rect 19705 23199 19763 23205
rect 20162 23196 20168 23208
rect 20220 23196 20226 23248
rect 12437 23171 12495 23177
rect 12437 23137 12449 23171
rect 12483 23168 12495 23171
rect 12802 23168 12808 23180
rect 12483 23140 12517 23168
rect 12763 23140 12808 23168
rect 12483 23137 12495 23140
rect 12437 23131 12495 23137
rect 12802 23128 12808 23140
rect 12860 23128 12866 23180
rect 12986 23168 12992 23180
rect 12947 23140 12992 23168
rect 12986 23128 12992 23140
rect 13044 23128 13050 23180
rect 18325 23171 18383 23177
rect 18325 23137 18337 23171
rect 18371 23168 18383 23171
rect 19242 23168 19248 23180
rect 18371 23140 19248 23168
rect 18371 23137 18383 23140
rect 18325 23131 18383 23137
rect 19242 23128 19248 23140
rect 19300 23128 19306 23180
rect 22189 23171 22247 23177
rect 22189 23137 22201 23171
rect 22235 23168 22247 23171
rect 22554 23168 22560 23180
rect 22235 23140 22560 23168
rect 22235 23137 22247 23140
rect 22189 23131 22247 23137
rect 22554 23128 22560 23140
rect 22612 23128 22618 23180
rect 5258 23060 5264 23112
rect 5316 23100 5322 23112
rect 5353 23103 5411 23109
rect 5353 23100 5365 23103
rect 5316 23072 5365 23100
rect 5316 23060 5322 23072
rect 5353 23069 5365 23072
rect 5399 23100 5411 23103
rect 5537 23103 5595 23109
rect 5537 23100 5549 23103
rect 5399 23072 5549 23100
rect 5399 23069 5411 23072
rect 5353 23063 5411 23069
rect 5537 23069 5549 23072
rect 5583 23069 5595 23103
rect 12526 23100 12532 23112
rect 12487 23072 12532 23100
rect 5537 23063 5595 23069
rect 5552 23032 5580 23063
rect 12526 23060 12532 23072
rect 12584 23060 12590 23112
rect 18049 23103 18107 23109
rect 18049 23069 18061 23103
rect 18095 23100 18107 23103
rect 19610 23100 19616 23112
rect 18095 23072 19616 23100
rect 18095 23069 18107 23072
rect 18049 23063 18107 23069
rect 19610 23060 19616 23072
rect 19668 23100 19674 23112
rect 19889 23103 19947 23109
rect 19889 23100 19901 23103
rect 19668 23072 19901 23100
rect 19668 23060 19674 23072
rect 19889 23069 19901 23072
rect 19935 23100 19947 23103
rect 20806 23100 20812 23112
rect 19935 23072 20812 23100
rect 19935 23069 19947 23072
rect 19889 23063 19947 23069
rect 20806 23060 20812 23072
rect 20864 23100 20870 23112
rect 21634 23100 21640 23112
rect 20864 23072 21640 23100
rect 20864 23060 20870 23072
rect 21634 23060 21640 23072
rect 21692 23100 21698 23112
rect 21729 23103 21787 23109
rect 21729 23100 21741 23103
rect 21692 23072 21741 23100
rect 21692 23060 21698 23072
rect 21729 23069 21741 23072
rect 21775 23100 21787 23103
rect 21913 23103 21971 23109
rect 21913 23100 21925 23103
rect 21775 23072 21925 23100
rect 21775 23069 21787 23072
rect 21729 23063 21787 23069
rect 21913 23069 21925 23072
rect 21959 23069 21971 23103
rect 21913 23063 21971 23069
rect 7282 23032 7288 23044
rect 5552 23004 7288 23032
rect 7282 22992 7288 23004
rect 7340 22992 7346 23044
rect 6178 22924 6184 22976
rect 6236 22964 6242 22976
rect 7466 22964 7472 22976
rect 6236 22936 7472 22964
rect 6236 22924 6242 22936
rect 7466 22924 7472 22936
rect 7524 22964 7530 22976
rect 7837 22967 7895 22973
rect 7837 22964 7849 22967
rect 7524 22936 7849 22964
rect 7524 22924 7530 22936
rect 7837 22933 7849 22936
rect 7883 22933 7895 22967
rect 9766 22964 9772 22976
rect 9727 22936 9772 22964
rect 7837 22927 7895 22933
rect 9766 22924 9772 22936
rect 9824 22924 9830 22976
rect 12066 22964 12072 22976
rect 12027 22936 12072 22964
rect 12066 22924 12072 22936
rect 12124 22924 12130 22976
rect 23474 22964 23480 22976
rect 23435 22936 23480 22964
rect 23474 22924 23480 22936
rect 23532 22924 23538 22976
rect 1104 22874 24656 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 24656 22874
rect 81618 22856 81624 22908
rect 81676 22896 81682 22908
rect 82262 22896 82268 22908
rect 81676 22868 82268 22896
rect 81676 22856 81682 22868
rect 82262 22856 82268 22868
rect 82320 22856 82326 22908
rect 1104 22800 24656 22822
rect 3142 22720 3148 22772
rect 3200 22760 3206 22772
rect 3881 22763 3939 22769
rect 3881 22760 3893 22763
rect 3200 22732 3893 22760
rect 3200 22720 3206 22732
rect 3881 22729 3893 22732
rect 3927 22729 3939 22763
rect 3881 22723 3939 22729
rect 4525 22763 4583 22769
rect 4525 22729 4537 22763
rect 4571 22760 4583 22763
rect 4614 22760 4620 22772
rect 4571 22732 4620 22760
rect 4571 22729 4583 22732
rect 4525 22723 4583 22729
rect 4614 22720 4620 22732
rect 4672 22760 4678 22772
rect 9030 22760 9036 22772
rect 4672 22732 9036 22760
rect 4672 22720 4678 22732
rect 7300 22633 7328 22732
rect 9030 22720 9036 22732
rect 9088 22720 9094 22772
rect 9674 22760 9680 22772
rect 9635 22732 9680 22760
rect 9674 22720 9680 22732
rect 9732 22720 9738 22772
rect 13817 22763 13875 22769
rect 13817 22729 13829 22763
rect 13863 22760 13875 22763
rect 13906 22760 13912 22772
rect 13863 22732 13912 22760
rect 13863 22729 13875 22732
rect 13817 22723 13875 22729
rect 7285 22627 7343 22633
rect 7285 22593 7297 22627
rect 7331 22593 7343 22627
rect 7285 22587 7343 22593
rect 12526 22584 12532 22636
rect 12584 22624 12590 22636
rect 12802 22624 12808 22636
rect 12584 22596 12808 22624
rect 12584 22584 12590 22596
rect 12802 22584 12808 22596
rect 12860 22624 12866 22636
rect 13173 22627 13231 22633
rect 12860 22596 13124 22624
rect 12860 22584 12866 22596
rect 2498 22556 2504 22568
rect 2459 22528 2504 22556
rect 2498 22516 2504 22528
rect 2556 22516 2562 22568
rect 2777 22559 2835 22565
rect 2777 22525 2789 22559
rect 2823 22556 2835 22559
rect 7561 22559 7619 22565
rect 2823 22528 4384 22556
rect 2823 22525 2835 22528
rect 2777 22519 2835 22525
rect 4356 22497 4384 22528
rect 7561 22525 7573 22559
rect 7607 22556 7619 22559
rect 7926 22556 7932 22568
rect 7607 22528 7932 22556
rect 7607 22525 7619 22528
rect 7561 22519 7619 22525
rect 7926 22516 7932 22528
rect 7984 22516 7990 22568
rect 8941 22559 8999 22565
rect 8941 22525 8953 22559
rect 8987 22556 8999 22559
rect 9674 22556 9680 22568
rect 8987 22528 9680 22556
rect 8987 22525 8999 22528
rect 8941 22519 8999 22525
rect 9674 22516 9680 22528
rect 9732 22556 9738 22568
rect 13096 22565 13124 22596
rect 13173 22593 13185 22627
rect 13219 22624 13231 22627
rect 13832 22624 13860 22723
rect 13906 22720 13912 22732
rect 13964 22720 13970 22772
rect 13219 22596 13860 22624
rect 19521 22627 19579 22633
rect 13219 22593 13231 22596
rect 13173 22587 13231 22593
rect 19521 22593 19533 22627
rect 19567 22624 19579 22627
rect 19610 22624 19616 22636
rect 19567 22596 19616 22624
rect 19567 22593 19579 22596
rect 19521 22587 19579 22593
rect 19610 22584 19616 22596
rect 19668 22584 19674 22636
rect 9769 22559 9827 22565
rect 9769 22556 9781 22559
rect 9732 22528 9781 22556
rect 9732 22516 9738 22528
rect 9769 22525 9781 22528
rect 9815 22525 9827 22559
rect 9769 22519 9827 22525
rect 13081 22559 13139 22565
rect 13081 22525 13093 22559
rect 13127 22525 13139 22559
rect 13081 22519 13139 22525
rect 13449 22559 13507 22565
rect 13449 22525 13461 22559
rect 13495 22525 13507 22559
rect 13449 22519 13507 22525
rect 13633 22559 13691 22565
rect 13633 22525 13645 22559
rect 13679 22556 13691 22559
rect 14642 22556 14648 22568
rect 13679 22528 14648 22556
rect 13679 22525 13691 22528
rect 13633 22519 13691 22525
rect 4341 22491 4399 22497
rect 4341 22457 4353 22491
rect 4387 22488 4399 22491
rect 5626 22488 5632 22500
rect 4387 22460 5632 22488
rect 4387 22457 4399 22460
rect 4341 22451 4399 22457
rect 5626 22448 5632 22460
rect 5684 22448 5690 22500
rect 12434 22448 12440 22500
rect 12492 22488 12498 22500
rect 12492 22460 12537 22488
rect 12492 22448 12498 22460
rect 12618 22448 12624 22500
rect 12676 22488 12682 22500
rect 13464 22488 13492 22519
rect 14642 22516 14648 22528
rect 14700 22516 14706 22568
rect 19886 22556 19892 22568
rect 19847 22528 19892 22556
rect 19886 22516 19892 22528
rect 19944 22516 19950 22568
rect 18414 22488 18420 22500
rect 12676 22460 18420 22488
rect 12676 22448 12682 22460
rect 18414 22448 18420 22460
rect 18472 22448 18478 22500
rect 21266 22488 21272 22500
rect 21227 22460 21272 22488
rect 21266 22448 21272 22460
rect 21324 22448 21330 22500
rect 9861 22423 9919 22429
rect 9861 22389 9873 22423
rect 9907 22420 9919 22423
rect 9950 22420 9956 22432
rect 9907 22392 9956 22420
rect 9907 22389 9919 22392
rect 9861 22383 9919 22389
rect 9950 22380 9956 22392
rect 10008 22380 10014 22432
rect 12253 22423 12311 22429
rect 12253 22389 12265 22423
rect 12299 22420 12311 22423
rect 12636 22420 12664 22448
rect 12299 22392 12664 22420
rect 12299 22389 12311 22392
rect 12253 22383 12311 22389
rect 1104 22330 24656 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 24656 22330
rect 1104 22256 24656 22278
rect 4614 22216 4620 22228
rect 4172 22188 4620 22216
rect 4065 22083 4123 22089
rect 4065 22049 4077 22083
rect 4111 22080 4123 22083
rect 4172 22080 4200 22188
rect 4614 22176 4620 22188
rect 4672 22216 4678 22228
rect 7926 22216 7932 22228
rect 4672 22188 5028 22216
rect 7887 22188 7932 22216
rect 4672 22176 4678 22188
rect 4111 22052 4200 22080
rect 4341 22083 4399 22089
rect 4111 22049 4123 22052
rect 4065 22043 4123 22049
rect 4341 22049 4353 22083
rect 4387 22080 4399 22083
rect 4706 22080 4712 22092
rect 4387 22052 4712 22080
rect 4387 22049 4399 22052
rect 4341 22043 4399 22049
rect 4706 22040 4712 22052
rect 4764 22040 4770 22092
rect 5000 22080 5028 22188
rect 7926 22176 7932 22188
rect 7984 22176 7990 22228
rect 12437 22219 12495 22225
rect 12437 22185 12449 22219
rect 12483 22216 12495 22219
rect 12710 22216 12716 22228
rect 12483 22188 12716 22216
rect 12483 22185 12495 22188
rect 12437 22179 12495 22185
rect 12710 22176 12716 22188
rect 12768 22176 12774 22228
rect 18322 22216 18328 22228
rect 18283 22188 18328 22216
rect 18322 22176 18328 22188
rect 18380 22176 18386 22228
rect 19981 22219 20039 22225
rect 19981 22185 19993 22219
rect 20027 22216 20039 22219
rect 20070 22216 20076 22228
rect 20027 22188 20076 22216
rect 20027 22185 20039 22188
rect 19981 22179 20039 22185
rect 7742 22148 7748 22160
rect 6932 22120 7748 22148
rect 6932 22089 6960 22120
rect 7742 22108 7748 22120
rect 7800 22108 7806 22160
rect 5813 22083 5871 22089
rect 5813 22080 5825 22083
rect 5000 22052 5825 22080
rect 5813 22049 5825 22052
rect 5859 22049 5871 22083
rect 5813 22043 5871 22049
rect 6917 22083 6975 22089
rect 6917 22049 6929 22083
rect 6963 22080 6975 22083
rect 7466 22080 7472 22092
rect 6963 22052 6997 22080
rect 7427 22052 7472 22080
rect 6963 22049 6975 22052
rect 6917 22043 6975 22049
rect 7466 22040 7472 22052
rect 7524 22040 7530 22092
rect 7653 22083 7711 22089
rect 7653 22049 7665 22083
rect 7699 22080 7711 22083
rect 7699 22052 7972 22080
rect 7699 22049 7711 22052
rect 7653 22043 7711 22049
rect 6733 22015 6791 22021
rect 6733 21981 6745 22015
rect 6779 21981 6791 22015
rect 6733 21975 6791 21981
rect 4062 21836 4068 21888
rect 4120 21876 4126 21888
rect 5445 21879 5503 21885
rect 5445 21876 5457 21879
rect 4120 21848 5457 21876
rect 4120 21836 4126 21848
rect 5445 21845 5457 21848
rect 5491 21845 5503 21879
rect 6638 21876 6644 21888
rect 6599 21848 6644 21876
rect 5445 21839 5503 21845
rect 6638 21836 6644 21848
rect 6696 21876 6702 21888
rect 6748 21876 6776 21975
rect 6696 21848 6776 21876
rect 7944 21876 7972 22052
rect 9122 22040 9128 22092
rect 9180 22080 9186 22092
rect 9677 22083 9735 22089
rect 9677 22080 9689 22083
rect 9180 22052 9689 22080
rect 9180 22040 9186 22052
rect 9677 22049 9689 22052
rect 9723 22049 9735 22083
rect 9677 22043 9735 22049
rect 11517 22083 11575 22089
rect 11517 22049 11529 22083
rect 11563 22080 11575 22083
rect 12434 22080 12440 22092
rect 11563 22052 12440 22080
rect 11563 22049 11575 22052
rect 11517 22043 11575 22049
rect 12434 22040 12440 22052
rect 12492 22040 12498 22092
rect 12728 22080 12756 22176
rect 13262 22148 13268 22160
rect 13004 22120 13268 22148
rect 13004 22089 13032 22120
rect 13262 22108 13268 22120
rect 13320 22108 13326 22160
rect 18340 22148 18368 22176
rect 18690 22148 18696 22160
rect 18340 22120 18696 22148
rect 18690 22108 18696 22120
rect 18748 22148 18754 22160
rect 18748 22120 19656 22148
rect 18748 22108 18754 22120
rect 12989 22083 13047 22089
rect 12989 22080 13001 22083
rect 12728 22052 13001 22080
rect 12989 22049 13001 22052
rect 13035 22049 13047 22083
rect 12989 22043 13047 22049
rect 13173 22083 13231 22089
rect 13173 22049 13185 22083
rect 13219 22049 13231 22083
rect 13173 22043 13231 22049
rect 13449 22083 13507 22089
rect 13449 22049 13461 22083
rect 13495 22080 13507 22083
rect 13814 22080 13820 22092
rect 13495 22052 13820 22080
rect 13495 22049 13507 22052
rect 13449 22043 13507 22049
rect 9490 21972 9496 22024
rect 9548 22012 9554 22024
rect 12529 22015 12587 22021
rect 9548 21984 12480 22012
rect 9548 21972 9554 21984
rect 9858 21944 9864 21956
rect 9819 21916 9864 21944
rect 9858 21904 9864 21916
rect 9916 21904 9922 21956
rect 12452 21944 12480 21984
rect 12529 21981 12541 22015
rect 12575 22012 12587 22015
rect 12710 22012 12716 22024
rect 12575 21984 12716 22012
rect 12575 21981 12587 21984
rect 12529 21975 12587 21981
rect 12710 21972 12716 21984
rect 12768 21972 12774 22024
rect 12802 21972 12808 22024
rect 12860 22012 12866 22024
rect 13188 22012 13216 22043
rect 13814 22040 13820 22052
rect 13872 22040 13878 22092
rect 14001 22083 14059 22089
rect 14001 22049 14013 22083
rect 14047 22080 14059 22083
rect 14182 22080 14188 22092
rect 14047 22052 14188 22080
rect 14047 22049 14059 22052
rect 14001 22043 14059 22049
rect 14182 22040 14188 22052
rect 14240 22040 14246 22092
rect 14458 22040 14464 22092
rect 14516 22080 14522 22092
rect 17313 22083 17371 22089
rect 17313 22080 17325 22083
rect 14516 22052 17325 22080
rect 14516 22040 14522 22052
rect 17313 22049 17325 22052
rect 17359 22049 17371 22083
rect 17313 22043 17371 22049
rect 18414 22040 18420 22092
rect 18472 22080 18478 22092
rect 19628 22089 19656 22120
rect 18509 22083 18567 22089
rect 18509 22080 18521 22083
rect 18472 22052 18521 22080
rect 18472 22040 18478 22052
rect 18509 22049 18521 22052
rect 18555 22080 18567 22083
rect 19245 22083 19303 22089
rect 19245 22080 19257 22083
rect 18555 22052 19257 22080
rect 18555 22049 18567 22052
rect 18509 22043 18567 22049
rect 19245 22049 19257 22052
rect 19291 22049 19303 22083
rect 19245 22043 19303 22049
rect 19613 22083 19671 22089
rect 19613 22049 19625 22083
rect 19659 22049 19671 22083
rect 19613 22043 19671 22049
rect 19797 22083 19855 22089
rect 19797 22049 19809 22083
rect 19843 22080 19855 22083
rect 19996 22080 20024 22179
rect 20070 22176 20076 22188
rect 20128 22176 20134 22228
rect 21266 22148 21272 22160
rect 20916 22120 21272 22148
rect 20916 22089 20944 22120
rect 21266 22108 21272 22120
rect 21324 22108 21330 22160
rect 19843 22052 20024 22080
rect 20901 22083 20959 22089
rect 19843 22049 19855 22052
rect 19797 22043 19855 22049
rect 20901 22049 20913 22083
rect 20947 22049 20959 22083
rect 20901 22043 20959 22049
rect 24029 22083 24087 22089
rect 24029 22049 24041 22083
rect 24075 22080 24087 22083
rect 24305 22083 24363 22089
rect 24305 22080 24317 22083
rect 24075 22052 24317 22080
rect 24075 22049 24087 22052
rect 24029 22043 24087 22049
rect 24305 22049 24317 22052
rect 24351 22080 24363 22083
rect 24486 22080 24492 22092
rect 24351 22052 24492 22080
rect 24351 22049 24363 22052
rect 24305 22043 24363 22049
rect 24486 22040 24492 22052
rect 24544 22040 24550 22092
rect 12860 21984 13216 22012
rect 13725 22015 13783 22021
rect 12860 21972 12866 21984
rect 13725 21981 13737 22015
rect 13771 22012 13783 22015
rect 14090 22012 14096 22024
rect 13771 21984 14096 22012
rect 13771 21981 13783 21984
rect 13725 21975 13783 21981
rect 14090 21972 14096 21984
rect 14148 21972 14154 22024
rect 18046 21972 18052 22024
rect 18104 22012 18110 22024
rect 18601 22015 18659 22021
rect 18601 22012 18613 22015
rect 18104 21984 18613 22012
rect 18104 21972 18110 21984
rect 18601 21981 18613 21984
rect 18647 21981 18659 22015
rect 18601 21975 18659 21981
rect 19058 21972 19064 22024
rect 19116 22012 19122 22024
rect 19153 22015 19211 22021
rect 19153 22012 19165 22015
rect 19116 21984 19165 22012
rect 19116 21972 19122 21984
rect 19153 21981 19165 21984
rect 19199 22012 19211 22015
rect 20993 22015 21051 22021
rect 20993 22012 21005 22015
rect 19199 21984 21005 22012
rect 19199 21981 19211 21984
rect 19153 21975 19211 21981
rect 20993 21981 21005 21984
rect 21039 21981 21051 22015
rect 20993 21975 21051 21981
rect 28442 21944 28448 21956
rect 12452 21916 28448 21944
rect 28442 21904 28448 21916
rect 28500 21904 28506 21956
rect 9950 21876 9956 21888
rect 7944 21848 9956 21876
rect 6696 21836 6702 21848
rect 9950 21836 9956 21848
rect 10008 21836 10014 21888
rect 11609 21879 11667 21885
rect 11609 21845 11621 21879
rect 11655 21876 11667 21879
rect 11698 21876 11704 21888
rect 11655 21848 11704 21876
rect 11655 21845 11667 21848
rect 11609 21839 11667 21845
rect 11698 21836 11704 21848
rect 11756 21836 11762 21888
rect 12250 21876 12256 21888
rect 12211 21848 12256 21876
rect 12250 21836 12256 21848
rect 12308 21836 12314 21888
rect 14090 21836 14096 21888
rect 14148 21876 14154 21888
rect 14185 21879 14243 21885
rect 14185 21876 14197 21879
rect 14148 21848 14197 21876
rect 14148 21836 14154 21848
rect 14185 21845 14197 21848
rect 14231 21876 14243 21879
rect 15838 21876 15844 21888
rect 14231 21848 15844 21876
rect 14231 21845 14243 21848
rect 14185 21839 14243 21845
rect 15838 21836 15844 21848
rect 15896 21836 15902 21888
rect 17497 21879 17555 21885
rect 17497 21845 17509 21879
rect 17543 21876 17555 21879
rect 19150 21876 19156 21888
rect 17543 21848 19156 21876
rect 17543 21845 17555 21848
rect 17497 21839 17555 21845
rect 19150 21836 19156 21848
rect 19208 21836 19214 21888
rect 24118 21876 24124 21888
rect 24079 21848 24124 21876
rect 24118 21836 24124 21848
rect 24176 21836 24182 21888
rect 1104 21786 24656 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 24656 21786
rect 1104 21712 24656 21734
rect 4341 21675 4399 21681
rect 4341 21641 4353 21675
rect 4387 21672 4399 21675
rect 5166 21672 5172 21684
rect 4387 21644 5172 21672
rect 4387 21641 4399 21644
rect 4341 21635 4399 21641
rect 2777 21539 2835 21545
rect 2777 21505 2789 21539
rect 2823 21536 2835 21539
rect 4356 21536 4384 21635
rect 5166 21632 5172 21644
rect 5224 21632 5230 21684
rect 7742 21632 7748 21684
rect 7800 21672 7806 21684
rect 9306 21672 9312 21684
rect 7800 21644 9312 21672
rect 7800 21632 7806 21644
rect 9306 21632 9312 21644
rect 9364 21632 9370 21684
rect 17126 21672 17132 21684
rect 9416 21644 17132 21672
rect 4525 21607 4583 21613
rect 4525 21573 4537 21607
rect 4571 21604 4583 21607
rect 4614 21604 4620 21616
rect 4571 21576 4620 21604
rect 4571 21573 4583 21576
rect 4525 21567 4583 21573
rect 2823 21508 4384 21536
rect 2823 21505 2835 21508
rect 2777 21499 2835 21505
rect 2498 21468 2504 21480
rect 2411 21440 2504 21468
rect 2498 21428 2504 21440
rect 2556 21468 2562 21480
rect 4540 21468 4568 21567
rect 4614 21564 4620 21576
rect 4672 21564 4678 21616
rect 6638 21564 6644 21616
rect 6696 21604 6702 21616
rect 9416 21604 9444 21644
rect 17126 21632 17132 21644
rect 17184 21632 17190 21684
rect 19613 21675 19671 21681
rect 19613 21641 19625 21675
rect 19659 21672 19671 21675
rect 19886 21672 19892 21684
rect 19659 21644 19892 21672
rect 19659 21641 19671 21644
rect 19613 21635 19671 21641
rect 19886 21632 19892 21644
rect 19944 21632 19950 21684
rect 6696 21576 9444 21604
rect 12253 21607 12311 21613
rect 6696 21564 6702 21576
rect 12253 21573 12265 21607
rect 12299 21604 12311 21607
rect 14001 21607 14059 21613
rect 12299 21576 12480 21604
rect 12299 21573 12311 21576
rect 12253 21567 12311 21573
rect 12452 21548 12480 21576
rect 14001 21573 14013 21607
rect 14047 21604 14059 21607
rect 14090 21604 14096 21616
rect 14047 21576 14096 21604
rect 14047 21573 14059 21576
rect 14001 21567 14059 21573
rect 14090 21564 14096 21576
rect 14148 21564 14154 21616
rect 5626 21496 5632 21548
rect 5684 21536 5690 21548
rect 6178 21536 6184 21548
rect 5684 21508 6184 21536
rect 5684 21496 5690 21508
rect 6178 21496 6184 21508
rect 6236 21536 6242 21548
rect 7929 21539 7987 21545
rect 7929 21536 7941 21539
rect 6236 21508 7941 21536
rect 6236 21496 6242 21508
rect 7929 21505 7941 21508
rect 7975 21505 7987 21539
rect 9766 21536 9772 21548
rect 7929 21499 7987 21505
rect 8036 21508 9772 21536
rect 2556 21440 4568 21468
rect 2556 21428 2562 21440
rect 5718 21428 5724 21480
rect 5776 21468 5782 21480
rect 8036 21477 8064 21508
rect 9766 21496 9772 21508
rect 9824 21496 9830 21548
rect 12434 21496 12440 21548
rect 12492 21536 12498 21548
rect 12710 21536 12716 21548
rect 12492 21508 12537 21536
rect 12671 21508 12716 21536
rect 12492 21496 12498 21508
rect 12710 21496 12716 21508
rect 12768 21496 12774 21548
rect 22370 21496 22376 21548
rect 22428 21536 22434 21548
rect 22922 21536 22928 21548
rect 22428 21508 22928 21536
rect 22428 21496 22434 21508
rect 22922 21496 22928 21508
rect 22980 21496 22986 21548
rect 6825 21471 6883 21477
rect 6825 21468 6837 21471
rect 5776 21440 6837 21468
rect 5776 21428 5782 21440
rect 6825 21437 6837 21440
rect 6871 21437 6883 21471
rect 8021 21471 8079 21477
rect 8021 21468 8033 21471
rect 6825 21431 6883 21437
rect 6932 21440 8033 21468
rect 6730 21360 6736 21412
rect 6788 21400 6794 21412
rect 6932 21400 6960 21440
rect 8021 21437 8033 21440
rect 8067 21437 8079 21471
rect 9122 21468 9128 21480
rect 9083 21440 9128 21468
rect 8021 21431 8079 21437
rect 9122 21428 9128 21440
rect 9180 21428 9186 21480
rect 9306 21428 9312 21480
rect 9364 21468 9370 21480
rect 14458 21468 14464 21480
rect 9364 21440 14464 21468
rect 9364 21428 9370 21440
rect 14458 21428 14464 21440
rect 14516 21428 14522 21480
rect 18417 21471 18475 21477
rect 18417 21437 18429 21471
rect 18463 21437 18475 21471
rect 18598 21468 18604 21480
rect 18559 21440 18604 21468
rect 18417 21431 18475 21437
rect 12526 21400 12532 21412
rect 6788 21372 6960 21400
rect 7024 21372 12532 21400
rect 6788 21360 6794 21372
rect 3142 21292 3148 21344
rect 3200 21332 3206 21344
rect 7024 21341 7052 21372
rect 12526 21360 12532 21372
rect 12584 21360 12590 21412
rect 3881 21335 3939 21341
rect 3881 21332 3893 21335
rect 3200 21304 3893 21332
rect 3200 21292 3206 21304
rect 3881 21301 3893 21304
rect 3927 21301 3939 21335
rect 3881 21295 3939 21301
rect 7009 21335 7067 21341
rect 7009 21301 7021 21335
rect 7055 21301 7067 21335
rect 7009 21295 7067 21301
rect 7929 21335 7987 21341
rect 7929 21301 7941 21335
rect 7975 21332 7987 21335
rect 8205 21335 8263 21341
rect 8205 21332 8217 21335
rect 7975 21304 8217 21332
rect 7975 21301 7987 21304
rect 7929 21295 7987 21301
rect 8205 21301 8217 21304
rect 8251 21332 8263 21335
rect 12250 21332 12256 21344
rect 8251 21304 12256 21332
rect 8251 21301 8263 21304
rect 8205 21295 8263 21301
rect 12250 21292 12256 21304
rect 12308 21332 12314 21344
rect 12710 21332 12716 21344
rect 12308 21304 12716 21332
rect 12308 21292 12314 21304
rect 12710 21292 12716 21304
rect 12768 21292 12774 21344
rect 18325 21335 18383 21341
rect 18325 21301 18337 21335
rect 18371 21332 18383 21335
rect 18432 21332 18460 21431
rect 18598 21428 18604 21440
rect 18656 21428 18662 21480
rect 19058 21468 19064 21480
rect 19019 21440 19064 21468
rect 19058 21428 19064 21440
rect 19116 21428 19122 21480
rect 19150 21428 19156 21480
rect 19208 21468 19214 21480
rect 21174 21468 21180 21480
rect 19208 21440 21180 21468
rect 19208 21428 19214 21440
rect 21174 21428 21180 21440
rect 21232 21428 21238 21480
rect 22189 21471 22247 21477
rect 22189 21437 22201 21471
rect 22235 21468 22247 21471
rect 22462 21468 22468 21480
rect 22235 21440 22468 21468
rect 22235 21437 22247 21440
rect 22189 21431 22247 21437
rect 22462 21428 22468 21440
rect 22520 21468 22526 21480
rect 22520 21440 22600 21468
rect 22520 21428 22526 21440
rect 22572 21344 22600 21440
rect 18782 21332 18788 21344
rect 18371 21304 18788 21332
rect 18371 21301 18383 21304
rect 18325 21295 18383 21301
rect 18782 21292 18788 21304
rect 18840 21292 18846 21344
rect 22278 21332 22284 21344
rect 22239 21304 22284 21332
rect 22278 21292 22284 21304
rect 22336 21292 22342 21344
rect 22554 21332 22560 21344
rect 22515 21304 22560 21332
rect 22554 21292 22560 21304
rect 22612 21292 22618 21344
rect 1104 21242 24656 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 24656 21242
rect 1104 21168 24656 21190
rect 7098 21088 7104 21140
rect 7156 21128 7162 21140
rect 7377 21131 7435 21137
rect 7377 21128 7389 21131
rect 7156 21100 7389 21128
rect 7156 21088 7162 21100
rect 7377 21097 7389 21100
rect 7423 21097 7435 21131
rect 22370 21128 22376 21140
rect 7377 21091 7435 21097
rect 21744 21100 22376 21128
rect 7009 21063 7067 21069
rect 7009 21029 7021 21063
rect 7055 21060 7067 21063
rect 7469 21063 7527 21069
rect 7469 21060 7481 21063
rect 7055 21032 7481 21060
rect 7055 21029 7067 21032
rect 7009 21023 7067 21029
rect 7469 21029 7481 21032
rect 7515 21060 7527 21063
rect 7558 21060 7564 21072
rect 7515 21032 7564 21060
rect 7515 21029 7527 21032
rect 7469 21023 7527 21029
rect 7558 21020 7564 21032
rect 7616 21020 7622 21072
rect 7834 21060 7840 21072
rect 7795 21032 7840 21060
rect 7834 21020 7840 21032
rect 7892 21020 7898 21072
rect 7282 20992 7288 21004
rect 7243 20964 7288 20992
rect 7282 20952 7288 20964
rect 7340 20952 7346 21004
rect 15286 20992 15292 21004
rect 15199 20964 15292 20992
rect 15286 20952 15292 20964
rect 15344 20992 15350 21004
rect 15654 20992 15660 21004
rect 15344 20964 15660 20992
rect 15344 20952 15350 20964
rect 15654 20952 15660 20964
rect 15712 20952 15718 21004
rect 21545 20995 21603 21001
rect 21545 20961 21557 20995
rect 21591 20992 21603 20995
rect 21634 20992 21640 21004
rect 21591 20964 21640 20992
rect 21591 20961 21603 20964
rect 21545 20955 21603 20961
rect 21634 20952 21640 20964
rect 21692 20952 21698 21004
rect 7101 20927 7159 20933
rect 7101 20893 7113 20927
rect 7147 20924 7159 20927
rect 7190 20924 7196 20936
rect 7147 20896 7196 20924
rect 7147 20893 7159 20896
rect 7101 20887 7159 20893
rect 7190 20884 7196 20896
rect 7248 20884 7254 20936
rect 12434 20884 12440 20936
rect 12492 20924 12498 20936
rect 12713 20927 12771 20933
rect 12713 20924 12725 20927
rect 12492 20896 12725 20924
rect 12492 20884 12498 20896
rect 12713 20893 12725 20896
rect 12759 20893 12771 20927
rect 12986 20924 12992 20936
rect 12947 20896 12992 20924
rect 12713 20887 12771 20893
rect 12621 20791 12679 20797
rect 12621 20757 12633 20791
rect 12667 20788 12679 20791
rect 12728 20788 12756 20887
rect 12986 20884 12992 20896
rect 13044 20884 13050 20936
rect 14369 20927 14427 20933
rect 14369 20893 14381 20927
rect 14415 20924 14427 20927
rect 14550 20924 14556 20936
rect 14415 20896 14556 20924
rect 14415 20893 14427 20896
rect 14369 20887 14427 20893
rect 14550 20884 14556 20896
rect 14608 20924 14614 20936
rect 21744 20924 21772 21100
rect 22370 21088 22376 21100
rect 22428 21088 22434 21140
rect 22554 21088 22560 21140
rect 22612 21128 22618 21140
rect 23017 21131 23075 21137
rect 23017 21128 23029 21131
rect 22612 21100 23029 21128
rect 22612 21088 22618 21100
rect 23017 21097 23029 21100
rect 23063 21097 23075 21131
rect 23017 21091 23075 21097
rect 21910 20924 21916 20936
rect 14608 20896 21772 20924
rect 21871 20896 21916 20924
rect 14608 20884 14614 20896
rect 21910 20884 21916 20896
rect 21968 20884 21974 20936
rect 13814 20816 13820 20868
rect 13872 20856 13878 20868
rect 15473 20859 15531 20865
rect 15473 20856 15485 20859
rect 13872 20828 15485 20856
rect 13872 20816 13878 20828
rect 15473 20825 15485 20828
rect 15519 20825 15531 20859
rect 15473 20819 15531 20825
rect 12894 20788 12900 20800
rect 12667 20760 12900 20788
rect 12667 20757 12679 20760
rect 12621 20751 12679 20757
rect 12894 20748 12900 20760
rect 12952 20788 12958 20800
rect 13722 20788 13728 20800
rect 12952 20760 13728 20788
rect 12952 20748 12958 20760
rect 13722 20748 13728 20760
rect 13780 20748 13786 20800
rect 1104 20698 24656 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 24656 20698
rect 1104 20624 24656 20646
rect 4341 20587 4399 20593
rect 4341 20553 4353 20587
rect 4387 20584 4399 20587
rect 4614 20584 4620 20596
rect 4387 20556 4620 20584
rect 4387 20553 4399 20556
rect 4341 20547 4399 20553
rect 4614 20544 4620 20556
rect 4672 20544 4678 20596
rect 8205 20587 8263 20593
rect 8205 20553 8217 20587
rect 8251 20584 8263 20587
rect 8754 20584 8760 20596
rect 8251 20556 8760 20584
rect 8251 20553 8263 20556
rect 8205 20547 8263 20553
rect 2498 20448 2504 20460
rect 2459 20420 2504 20448
rect 2498 20408 2504 20420
rect 2556 20408 2562 20460
rect 2777 20451 2835 20457
rect 2777 20417 2789 20451
rect 2823 20448 2835 20451
rect 3510 20448 3516 20460
rect 2823 20420 3516 20448
rect 2823 20417 2835 20420
rect 2777 20411 2835 20417
rect 3510 20408 3516 20420
rect 3568 20408 3574 20460
rect 6914 20380 6920 20392
rect 6875 20352 6920 20380
rect 6914 20340 6920 20352
rect 6972 20340 6978 20392
rect 7469 20383 7527 20389
rect 7469 20349 7481 20383
rect 7515 20349 7527 20383
rect 7469 20343 7527 20349
rect 7837 20383 7895 20389
rect 7837 20349 7849 20383
rect 7883 20380 7895 20383
rect 8110 20380 8116 20392
rect 7883 20352 8116 20380
rect 7883 20349 7895 20352
rect 7837 20343 7895 20349
rect 3878 20244 3884 20256
rect 3839 20216 3884 20244
rect 3878 20204 3884 20216
rect 3936 20204 3942 20256
rect 7484 20244 7512 20343
rect 8110 20340 8116 20352
rect 8168 20380 8174 20392
rect 8220 20380 8248 20547
rect 8754 20544 8760 20556
rect 8812 20544 8818 20596
rect 15378 20584 15384 20596
rect 15339 20556 15384 20584
rect 15378 20544 15384 20556
rect 15436 20544 15442 20596
rect 19705 20587 19763 20593
rect 19705 20553 19717 20587
rect 19751 20584 19763 20587
rect 19889 20587 19947 20593
rect 19889 20584 19901 20587
rect 19751 20556 19901 20584
rect 19751 20553 19763 20556
rect 19705 20547 19763 20553
rect 19889 20553 19901 20556
rect 19935 20584 19947 20587
rect 19978 20584 19984 20596
rect 19935 20556 19984 20584
rect 19935 20553 19947 20556
rect 19889 20547 19947 20553
rect 19978 20544 19984 20556
rect 20036 20544 20042 20596
rect 22741 20587 22799 20593
rect 22741 20553 22753 20587
rect 22787 20584 22799 20587
rect 23106 20584 23112 20596
rect 22787 20556 23112 20584
rect 22787 20553 22799 20556
rect 22741 20547 22799 20553
rect 13722 20448 13728 20460
rect 13635 20420 13728 20448
rect 13722 20408 13728 20420
rect 13780 20448 13786 20460
rect 13817 20451 13875 20457
rect 13817 20448 13829 20451
rect 13780 20420 13829 20448
rect 13780 20408 13786 20420
rect 13817 20417 13829 20420
rect 13863 20417 13875 20451
rect 20165 20451 20223 20457
rect 20165 20448 20177 20451
rect 13817 20411 13875 20417
rect 19904 20420 20177 20448
rect 8168 20352 8248 20380
rect 8168 20340 8174 20352
rect 13906 20340 13912 20392
rect 13964 20380 13970 20392
rect 14093 20383 14151 20389
rect 14093 20380 14105 20383
rect 13964 20352 14105 20380
rect 13964 20340 13970 20352
rect 14093 20349 14105 20352
rect 14139 20349 14151 20383
rect 14093 20343 14151 20349
rect 8018 20312 8024 20324
rect 7979 20284 8024 20312
rect 8018 20272 8024 20284
rect 8076 20272 8082 20324
rect 8389 20247 8447 20253
rect 8389 20244 8401 20247
rect 7484 20216 8401 20244
rect 8389 20213 8401 20216
rect 8435 20244 8447 20247
rect 8478 20244 8484 20256
rect 8435 20216 8484 20244
rect 8435 20213 8447 20216
rect 8389 20207 8447 20213
rect 8478 20204 8484 20216
rect 8536 20204 8542 20256
rect 19426 20204 19432 20256
rect 19484 20244 19490 20256
rect 19904 20244 19932 20420
rect 20165 20417 20177 20420
rect 20211 20417 20223 20451
rect 20165 20411 20223 20417
rect 19978 20340 19984 20392
rect 20036 20380 20042 20392
rect 20349 20383 20407 20389
rect 20349 20380 20361 20383
rect 20036 20352 20361 20380
rect 20036 20340 20042 20352
rect 20349 20349 20361 20352
rect 20395 20349 20407 20383
rect 20806 20380 20812 20392
rect 20767 20352 20812 20380
rect 20349 20343 20407 20349
rect 20364 20312 20392 20343
rect 20806 20340 20812 20352
rect 20864 20340 20870 20392
rect 20901 20383 20959 20389
rect 20901 20349 20913 20383
rect 20947 20349 20959 20383
rect 20901 20343 20959 20349
rect 22373 20383 22431 20389
rect 22373 20349 22385 20383
rect 22419 20380 22431 20383
rect 22554 20380 22560 20392
rect 22419 20352 22560 20380
rect 22419 20349 22431 20352
rect 22373 20343 22431 20349
rect 20916 20312 20944 20343
rect 22554 20340 22560 20352
rect 22612 20380 22618 20392
rect 22756 20380 22784 20547
rect 23106 20544 23112 20556
rect 23164 20544 23170 20596
rect 22612 20352 22784 20380
rect 22612 20340 22618 20352
rect 22465 20315 22523 20321
rect 22465 20312 22477 20315
rect 20364 20284 20944 20312
rect 21192 20284 22477 20312
rect 19981 20247 20039 20253
rect 19981 20244 19993 20247
rect 19484 20216 19993 20244
rect 19484 20204 19490 20216
rect 19981 20213 19993 20216
rect 20027 20244 20039 20247
rect 20622 20244 20628 20256
rect 20027 20216 20628 20244
rect 20027 20213 20039 20216
rect 19981 20207 20039 20213
rect 20622 20204 20628 20216
rect 20680 20204 20686 20256
rect 20806 20204 20812 20256
rect 20864 20244 20870 20256
rect 21192 20244 21220 20284
rect 22465 20281 22477 20284
rect 22511 20281 22523 20315
rect 22465 20275 22523 20281
rect 20864 20216 21220 20244
rect 20864 20204 20870 20216
rect 21266 20204 21272 20256
rect 21324 20244 21330 20256
rect 21361 20247 21419 20253
rect 21361 20244 21373 20247
rect 21324 20216 21373 20244
rect 21324 20204 21330 20216
rect 21361 20213 21373 20216
rect 21407 20213 21419 20247
rect 21361 20207 21419 20213
rect 1104 20154 24656 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 24656 20154
rect 1104 20080 24656 20102
rect 6178 20040 6184 20052
rect 5644 20012 6184 20040
rect 5644 19981 5672 20012
rect 6178 20000 6184 20012
rect 6236 20000 6242 20052
rect 8110 20040 8116 20052
rect 8071 20012 8116 20040
rect 8110 20000 8116 20012
rect 8168 20000 8174 20052
rect 14550 20040 14556 20052
rect 14511 20012 14556 20040
rect 14550 20000 14556 20012
rect 14608 20000 14614 20052
rect 22554 20040 22560 20052
rect 22515 20012 22560 20040
rect 22554 20000 22560 20012
rect 22612 20000 22618 20052
rect 5629 19975 5687 19981
rect 5629 19941 5641 19975
rect 5675 19941 5687 19975
rect 5629 19935 5687 19941
rect 5997 19975 6055 19981
rect 5997 19941 6009 19975
rect 6043 19972 6055 19975
rect 9122 19972 9128 19984
rect 6043 19944 9128 19972
rect 6043 19941 6055 19944
rect 5997 19935 6055 19941
rect 9122 19932 9128 19944
rect 9180 19932 9186 19984
rect 12897 19975 12955 19981
rect 12897 19941 12909 19975
rect 12943 19972 12955 19975
rect 12986 19972 12992 19984
rect 12943 19944 12992 19972
rect 12943 19941 12955 19944
rect 12897 19935 12955 19941
rect 12986 19932 12992 19944
rect 13044 19932 13050 19984
rect 14568 19972 14596 20000
rect 13372 19944 14044 19972
rect 5445 19907 5503 19913
rect 5445 19873 5457 19907
rect 5491 19873 5503 19907
rect 5445 19867 5503 19873
rect 5537 19907 5595 19913
rect 5537 19873 5549 19907
rect 5583 19904 5595 19907
rect 6546 19904 6552 19916
rect 5583 19876 6552 19904
rect 5583 19873 5595 19876
rect 5537 19867 5595 19873
rect 5261 19839 5319 19845
rect 5261 19805 5273 19839
rect 5307 19836 5319 19839
rect 5350 19836 5356 19848
rect 5307 19808 5356 19836
rect 5307 19805 5319 19808
rect 5261 19799 5319 19805
rect 5350 19796 5356 19808
rect 5408 19796 5414 19848
rect 5460 19836 5488 19867
rect 6546 19864 6552 19876
rect 6604 19864 6610 19916
rect 7006 19904 7012 19916
rect 6967 19876 7012 19904
rect 7006 19864 7012 19876
rect 7064 19864 7070 19916
rect 7377 19907 7435 19913
rect 7377 19873 7389 19907
rect 7423 19904 7435 19907
rect 7745 19907 7803 19913
rect 7423 19876 7696 19904
rect 7423 19873 7435 19876
rect 7377 19867 7435 19873
rect 7282 19836 7288 19848
rect 5460 19808 7288 19836
rect 7282 19796 7288 19808
rect 7340 19836 7346 19848
rect 7466 19836 7472 19848
rect 7340 19808 7472 19836
rect 7340 19796 7346 19808
rect 7466 19796 7472 19808
rect 7524 19796 7530 19848
rect 7668 19768 7696 19876
rect 7745 19873 7757 19907
rect 7791 19904 7803 19907
rect 8110 19904 8116 19916
rect 7791 19876 8116 19904
rect 7791 19873 7803 19876
rect 7745 19867 7803 19873
rect 8110 19864 8116 19876
rect 8168 19904 8174 19916
rect 9306 19904 9312 19916
rect 8168 19876 9312 19904
rect 8168 19864 8174 19876
rect 9306 19864 9312 19876
rect 9364 19864 9370 19916
rect 13372 19913 13400 19944
rect 13357 19907 13415 19913
rect 13357 19904 13369 19907
rect 12544 19876 13369 19904
rect 7834 19836 7840 19848
rect 7795 19808 7840 19836
rect 7834 19796 7840 19808
rect 7892 19796 7898 19848
rect 7668 19740 7880 19768
rect 7852 19700 7880 19740
rect 8205 19703 8263 19709
rect 8205 19700 8217 19703
rect 7852 19672 8217 19700
rect 8205 19669 8217 19672
rect 8251 19700 8263 19703
rect 8478 19700 8484 19712
rect 8251 19672 8484 19700
rect 8251 19669 8263 19672
rect 8205 19663 8263 19669
rect 8478 19660 8484 19672
rect 8536 19700 8542 19712
rect 10778 19700 10784 19712
rect 8536 19672 10784 19700
rect 8536 19660 8542 19672
rect 10778 19660 10784 19672
rect 10836 19660 10842 19712
rect 12544 19700 12572 19876
rect 13357 19873 13369 19876
rect 13403 19873 13415 19907
rect 13630 19904 13636 19916
rect 13591 19876 13636 19904
rect 13357 19867 13415 19873
rect 13630 19864 13636 19876
rect 13688 19864 13694 19916
rect 13814 19904 13820 19916
rect 13775 19876 13820 19904
rect 13814 19864 13820 19876
rect 13872 19864 13878 19916
rect 12621 19839 12679 19845
rect 12621 19805 12633 19839
rect 12667 19836 12679 19839
rect 12710 19836 12716 19848
rect 12667 19808 12716 19836
rect 12667 19805 12679 19808
rect 12621 19799 12679 19805
rect 12710 19796 12716 19808
rect 12768 19836 12774 19848
rect 13648 19836 13676 19864
rect 12768 19808 13676 19836
rect 14016 19836 14044 19944
rect 14108 19944 14596 19972
rect 14108 19913 14136 19944
rect 14093 19907 14151 19913
rect 14093 19873 14105 19907
rect 14139 19873 14151 19907
rect 14093 19867 14151 19873
rect 14182 19864 14188 19916
rect 14240 19904 14246 19916
rect 14369 19907 14427 19913
rect 14369 19904 14381 19907
rect 14240 19876 14381 19904
rect 14240 19864 14246 19876
rect 14369 19873 14381 19876
rect 14415 19904 14427 19907
rect 14918 19904 14924 19916
rect 14415 19876 14924 19904
rect 14415 19873 14427 19876
rect 14369 19867 14427 19873
rect 14918 19864 14924 19876
rect 14976 19864 14982 19916
rect 15286 19904 15292 19916
rect 15247 19876 15292 19904
rect 15286 19864 15292 19876
rect 15344 19864 15350 19916
rect 21266 19904 21272 19916
rect 21227 19876 21272 19904
rect 21266 19864 21272 19876
rect 21324 19864 21330 19916
rect 19426 19836 19432 19848
rect 14016 19808 19432 19836
rect 12768 19796 12774 19808
rect 19426 19796 19432 19808
rect 19484 19796 19490 19848
rect 20717 19839 20775 19845
rect 20717 19805 20729 19839
rect 20763 19836 20775 19839
rect 20990 19836 20996 19848
rect 20763 19808 20996 19836
rect 20763 19805 20775 19808
rect 20717 19799 20775 19805
rect 20990 19796 20996 19808
rect 21048 19796 21054 19848
rect 12710 19700 12716 19712
rect 12544 19672 12716 19700
rect 12710 19660 12716 19672
rect 12768 19660 12774 19712
rect 15378 19660 15384 19712
rect 15436 19700 15442 19712
rect 15473 19703 15531 19709
rect 15473 19700 15485 19703
rect 15436 19672 15485 19700
rect 15436 19660 15442 19672
rect 15473 19669 15485 19672
rect 15519 19669 15531 19703
rect 15473 19663 15531 19669
rect 1104 19610 24656 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 24656 19610
rect 1104 19536 24656 19558
rect 15197 19499 15255 19505
rect 15197 19465 15209 19499
rect 15243 19496 15255 19499
rect 15286 19496 15292 19508
rect 15243 19468 15292 19496
rect 15243 19465 15255 19468
rect 15197 19459 15255 19465
rect 15286 19456 15292 19468
rect 15344 19456 15350 19508
rect 19978 19496 19984 19508
rect 19939 19468 19984 19496
rect 19978 19456 19984 19468
rect 20036 19496 20042 19508
rect 20073 19499 20131 19505
rect 20073 19496 20085 19499
rect 20036 19468 20085 19496
rect 20036 19456 20042 19468
rect 20073 19465 20085 19468
rect 20119 19496 20131 19499
rect 21637 19499 21695 19505
rect 20119 19468 20668 19496
rect 20119 19465 20131 19468
rect 20073 19459 20131 19465
rect 14550 19388 14556 19440
rect 14608 19428 14614 19440
rect 15657 19431 15715 19437
rect 15657 19428 15669 19431
rect 14608 19400 15669 19428
rect 14608 19388 14614 19400
rect 15657 19397 15669 19400
rect 15703 19397 15715 19431
rect 15657 19391 15715 19397
rect 8294 19320 8300 19372
rect 8352 19360 8358 19372
rect 9309 19363 9367 19369
rect 9309 19360 9321 19363
rect 8352 19332 9321 19360
rect 8352 19320 8358 19332
rect 9309 19329 9321 19332
rect 9355 19329 9367 19363
rect 9309 19323 9367 19329
rect 10873 19363 10931 19369
rect 10873 19329 10885 19363
rect 10919 19360 10931 19363
rect 12342 19360 12348 19372
rect 10919 19332 12348 19360
rect 10919 19329 10931 19332
rect 10873 19323 10931 19329
rect 12342 19320 12348 19332
rect 12400 19320 12406 19372
rect 13814 19320 13820 19372
rect 13872 19360 13878 19372
rect 14918 19360 14924 19372
rect 13872 19332 14412 19360
rect 14879 19332 14924 19360
rect 13872 19320 13878 19332
rect 14384 19304 14412 19332
rect 14918 19320 14924 19332
rect 14976 19320 14982 19372
rect 7190 19292 7196 19304
rect 7024 19264 7196 19292
rect 7024 19236 7052 19264
rect 7190 19252 7196 19264
rect 7248 19252 7254 19304
rect 8386 19292 8392 19304
rect 7392 19264 8392 19292
rect 7006 19224 7012 19236
rect 6967 19196 7012 19224
rect 7006 19184 7012 19196
rect 7064 19184 7070 19236
rect 7098 19184 7104 19236
rect 7156 19224 7162 19236
rect 7392 19233 7420 19264
rect 8386 19252 8392 19264
rect 8444 19252 8450 19304
rect 8662 19252 8668 19304
rect 8720 19292 8726 19304
rect 8757 19295 8815 19301
rect 8757 19292 8769 19295
rect 8720 19264 8769 19292
rect 8720 19252 8726 19264
rect 8757 19261 8769 19264
rect 8803 19261 8815 19295
rect 8757 19255 8815 19261
rect 8925 19295 8983 19301
rect 8925 19261 8937 19295
rect 8971 19292 8983 19295
rect 9398 19292 9404 19304
rect 8971 19264 9404 19292
rect 8971 19261 8983 19264
rect 8925 19255 8983 19261
rect 9398 19252 9404 19264
rect 9456 19252 9462 19304
rect 9766 19252 9772 19304
rect 9824 19292 9830 19304
rect 12437 19295 12495 19301
rect 9824 19264 10548 19292
rect 9824 19252 9830 19264
rect 7285 19227 7343 19233
rect 7285 19224 7297 19227
rect 7156 19196 7297 19224
rect 7156 19184 7162 19196
rect 7285 19193 7297 19196
rect 7331 19193 7343 19227
rect 7285 19187 7343 19193
rect 7377 19227 7435 19233
rect 7377 19193 7389 19227
rect 7423 19193 7435 19227
rect 7377 19187 7435 19193
rect 7650 19184 7656 19236
rect 7708 19224 7714 19236
rect 7745 19227 7803 19233
rect 7745 19224 7757 19227
rect 7708 19196 7757 19224
rect 7708 19184 7714 19196
rect 7745 19193 7757 19196
rect 7791 19193 7803 19227
rect 7745 19187 7803 19193
rect 8478 19184 8484 19236
rect 8536 19224 8542 19236
rect 10520 19233 10548 19264
rect 12437 19261 12449 19295
rect 12483 19292 12495 19295
rect 12618 19292 12624 19304
rect 12483 19264 12624 19292
rect 12483 19261 12495 19264
rect 12437 19255 12495 19261
rect 12618 19252 12624 19264
rect 12676 19292 12682 19304
rect 12805 19295 12863 19301
rect 12805 19292 12817 19295
rect 12676 19264 12817 19292
rect 12676 19252 12682 19264
rect 12805 19261 12817 19264
rect 12851 19261 12863 19295
rect 12805 19255 12863 19261
rect 13541 19295 13599 19301
rect 13541 19261 13553 19295
rect 13587 19292 13599 19295
rect 13906 19292 13912 19304
rect 13587 19264 13912 19292
rect 13587 19261 13599 19264
rect 13541 19255 13599 19261
rect 13906 19252 13912 19264
rect 13964 19252 13970 19304
rect 14090 19292 14096 19304
rect 14051 19264 14096 19292
rect 14090 19252 14096 19264
rect 14148 19252 14154 19304
rect 14185 19295 14243 19301
rect 14185 19261 14197 19295
rect 14231 19261 14243 19295
rect 14366 19292 14372 19304
rect 14279 19264 14372 19292
rect 14185 19255 14243 19261
rect 8573 19227 8631 19233
rect 8573 19224 8585 19227
rect 8536 19196 8585 19224
rect 8536 19184 8542 19196
rect 8573 19193 8585 19196
rect 8619 19224 8631 19227
rect 10137 19227 10195 19233
rect 10137 19224 10149 19227
rect 8619 19196 10149 19224
rect 8619 19193 8631 19196
rect 8573 19187 8631 19193
rect 10137 19193 10149 19196
rect 10183 19193 10195 19227
rect 10413 19227 10471 19233
rect 10413 19224 10425 19227
rect 10137 19187 10195 19193
rect 10244 19196 10425 19224
rect 5902 19116 5908 19168
rect 5960 19156 5966 19168
rect 7193 19159 7251 19165
rect 7193 19156 7205 19159
rect 5960 19128 7205 19156
rect 5960 19116 5966 19128
rect 7193 19125 7205 19128
rect 7239 19156 7251 19159
rect 8662 19156 8668 19168
rect 7239 19128 8668 19156
rect 7239 19125 7251 19128
rect 7193 19119 7251 19125
rect 8662 19116 8668 19128
rect 8720 19116 8726 19168
rect 8846 19156 8852 19168
rect 8807 19128 8852 19156
rect 8846 19116 8852 19128
rect 8904 19156 8910 19168
rect 10244 19156 10272 19196
rect 10413 19193 10425 19196
rect 10459 19193 10471 19227
rect 10413 19187 10471 19193
rect 10505 19227 10563 19233
rect 10505 19193 10517 19227
rect 10551 19193 10563 19227
rect 10505 19187 10563 19193
rect 13265 19227 13323 19233
rect 13265 19193 13277 19227
rect 13311 19224 13323 19227
rect 13630 19224 13636 19236
rect 13311 19196 13636 19224
rect 13311 19193 13323 19196
rect 13265 19187 13323 19193
rect 13630 19184 13636 19196
rect 13688 19224 13694 19236
rect 14200 19224 14228 19255
rect 14366 19252 14372 19264
rect 14424 19252 14430 19304
rect 14829 19295 14887 19301
rect 14829 19261 14841 19295
rect 14875 19292 14887 19295
rect 15194 19292 15200 19304
rect 14875 19264 15200 19292
rect 14875 19261 14887 19264
rect 14829 19255 14887 19261
rect 15194 19252 15200 19264
rect 15252 19252 15258 19304
rect 15672 19292 15700 19391
rect 20441 19363 20499 19369
rect 20441 19329 20453 19363
rect 20487 19329 20499 19363
rect 20441 19323 20499 19329
rect 15841 19295 15899 19301
rect 15841 19292 15853 19295
rect 15672 19264 15853 19292
rect 15841 19261 15853 19264
rect 15887 19261 15899 19295
rect 15841 19255 15899 19261
rect 15933 19295 15991 19301
rect 15933 19261 15945 19295
rect 15979 19261 15991 19295
rect 18046 19292 18052 19304
rect 18007 19264 18052 19292
rect 15933 19255 15991 19261
rect 13688 19196 14228 19224
rect 14384 19224 14412 19252
rect 15948 19224 15976 19255
rect 18046 19252 18052 19264
rect 18104 19252 18110 19304
rect 14384 19196 15976 19224
rect 13688 19184 13694 19196
rect 16114 19184 16120 19236
rect 16172 19224 16178 19236
rect 16393 19227 16451 19233
rect 16393 19224 16405 19227
rect 16172 19196 16405 19224
rect 16172 19184 16178 19196
rect 16393 19193 16405 19196
rect 16439 19193 16451 19227
rect 20257 19227 20315 19233
rect 20257 19224 20269 19227
rect 16393 19187 16451 19193
rect 16500 19196 20269 19224
rect 8904 19128 10272 19156
rect 8904 19116 8910 19128
rect 10318 19116 10324 19168
rect 10376 19156 10382 19168
rect 10376 19128 10421 19156
rect 10376 19116 10382 19128
rect 12526 19116 12532 19168
rect 12584 19156 12590 19168
rect 12621 19159 12679 19165
rect 12621 19156 12633 19159
rect 12584 19128 12633 19156
rect 12584 19116 12590 19128
rect 12621 19125 12633 19128
rect 12667 19125 12679 19159
rect 13446 19156 13452 19168
rect 13407 19128 13452 19156
rect 12621 19119 12679 19125
rect 13446 19116 13452 19128
rect 13504 19156 13510 19168
rect 14090 19156 14096 19168
rect 13504 19128 14096 19156
rect 13504 19116 13510 19128
rect 14090 19116 14096 19128
rect 14148 19156 14154 19168
rect 16500 19156 16528 19196
rect 20257 19193 20269 19196
rect 20303 19224 20315 19227
rect 20456 19224 20484 19323
rect 20640 19301 20668 19468
rect 21637 19465 21649 19499
rect 21683 19496 21695 19499
rect 21910 19496 21916 19508
rect 21683 19468 21916 19496
rect 21683 19465 21695 19468
rect 21637 19459 21695 19465
rect 21910 19456 21916 19468
rect 21968 19456 21974 19508
rect 54110 19360 54116 19372
rect 54071 19332 54116 19360
rect 54110 19320 54116 19332
rect 54168 19320 54174 19372
rect 20625 19295 20683 19301
rect 20625 19261 20637 19295
rect 20671 19292 20683 19295
rect 21177 19295 21235 19301
rect 21177 19292 21189 19295
rect 20671 19264 21189 19292
rect 20671 19261 20683 19264
rect 20625 19255 20683 19261
rect 21177 19261 21189 19264
rect 21223 19261 21235 19295
rect 21177 19255 21235 19261
rect 21361 19295 21419 19301
rect 21361 19261 21373 19295
rect 21407 19292 21419 19295
rect 22278 19292 22284 19304
rect 21407 19264 22284 19292
rect 21407 19261 21419 19264
rect 21361 19255 21419 19261
rect 22278 19252 22284 19264
rect 22336 19252 22342 19304
rect 20303 19196 20484 19224
rect 20303 19193 20315 19196
rect 20257 19187 20315 19193
rect 18138 19156 18144 19168
rect 14148 19128 16528 19156
rect 18099 19128 18144 19156
rect 14148 19116 14154 19128
rect 18138 19116 18144 19128
rect 18196 19116 18202 19168
rect 20456 19156 20484 19196
rect 20714 19156 20720 19168
rect 20456 19128 20720 19156
rect 20714 19116 20720 19128
rect 20772 19116 20778 19168
rect 1104 19066 24656 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 24656 19066
rect 1104 18992 24656 19014
rect 3326 18912 3332 18964
rect 3384 18952 3390 18964
rect 22830 18952 22836 18964
rect 3384 18924 22836 18952
rect 3384 18912 3390 18924
rect 22830 18912 22836 18924
rect 22888 18912 22894 18964
rect 5350 18844 5356 18896
rect 5408 18884 5414 18896
rect 5721 18887 5779 18893
rect 5721 18884 5733 18887
rect 5408 18856 5733 18884
rect 5408 18844 5414 18856
rect 5721 18853 5733 18856
rect 5767 18853 5779 18887
rect 5721 18847 5779 18853
rect 6089 18887 6147 18893
rect 6089 18853 6101 18887
rect 6135 18884 6147 18887
rect 6730 18884 6736 18896
rect 6135 18856 6736 18884
rect 6135 18853 6147 18856
rect 6089 18847 6147 18853
rect 6730 18844 6736 18856
rect 6788 18844 6794 18896
rect 8941 18887 8999 18893
rect 8941 18884 8953 18887
rect 8312 18856 8953 18884
rect 5902 18816 5908 18828
rect 5863 18788 5908 18816
rect 5902 18776 5908 18788
rect 5960 18776 5966 18828
rect 5994 18776 6000 18828
rect 6052 18816 6058 18828
rect 7098 18816 7104 18828
rect 6052 18788 7104 18816
rect 6052 18776 6058 18788
rect 7098 18776 7104 18788
rect 7156 18776 7162 18828
rect 7650 18816 7656 18828
rect 7611 18788 7656 18816
rect 7650 18776 7656 18788
rect 7708 18776 7714 18828
rect 7834 18816 7840 18828
rect 7795 18788 7840 18816
rect 7834 18776 7840 18788
rect 7892 18776 7898 18828
rect 8110 18816 8116 18828
rect 8071 18788 8116 18816
rect 8110 18776 8116 18788
rect 8168 18776 8174 18828
rect 8312 18825 8340 18856
rect 8941 18853 8953 18856
rect 8987 18884 8999 18887
rect 9030 18884 9036 18896
rect 8987 18856 9036 18884
rect 8987 18853 8999 18856
rect 8941 18847 8999 18853
rect 9030 18844 9036 18856
rect 9088 18884 9094 18896
rect 16574 18884 16580 18896
rect 9088 18856 16580 18884
rect 9088 18844 9094 18856
rect 16574 18844 16580 18856
rect 16632 18844 16638 18896
rect 18601 18887 18659 18893
rect 18601 18884 18613 18887
rect 17972 18856 18613 18884
rect 17972 18828 18000 18856
rect 18601 18853 18613 18856
rect 18647 18853 18659 18887
rect 18601 18847 18659 18853
rect 8297 18819 8355 18825
rect 8297 18785 8309 18819
rect 8343 18785 8355 18819
rect 8297 18779 8355 18785
rect 13449 18819 13507 18825
rect 13449 18785 13461 18819
rect 13495 18785 13507 18819
rect 13630 18816 13636 18828
rect 13591 18788 13636 18816
rect 13449 18779 13507 18785
rect 6454 18748 6460 18760
rect 6415 18720 6460 18748
rect 6454 18708 6460 18720
rect 6512 18708 6518 18760
rect 7285 18751 7343 18757
rect 7285 18717 7297 18751
rect 7331 18748 7343 18751
rect 12897 18751 12955 18757
rect 12897 18748 12909 18751
rect 7331 18720 12909 18748
rect 7331 18717 7343 18720
rect 7285 18711 7343 18717
rect 12897 18717 12909 18720
rect 12943 18717 12955 18751
rect 13464 18748 13492 18779
rect 13630 18776 13636 18788
rect 13688 18776 13694 18828
rect 13817 18819 13875 18825
rect 13817 18785 13829 18819
rect 13863 18785 13875 18819
rect 13998 18816 14004 18828
rect 13959 18788 14004 18816
rect 13817 18779 13875 18785
rect 13832 18748 13860 18779
rect 13998 18776 14004 18788
rect 14056 18776 14062 18828
rect 14366 18816 14372 18828
rect 14327 18788 14372 18816
rect 14366 18776 14372 18788
rect 14424 18776 14430 18828
rect 15378 18816 15384 18828
rect 15339 18788 15384 18816
rect 15378 18776 15384 18788
rect 15436 18776 15442 18828
rect 17954 18816 17960 18828
rect 17915 18788 17960 18816
rect 17954 18776 17960 18788
rect 18012 18776 18018 18828
rect 18046 18776 18052 18828
rect 18104 18816 18110 18828
rect 18104 18788 18149 18816
rect 18104 18776 18110 18788
rect 15289 18751 15347 18757
rect 13464 18720 13584 18748
rect 13832 18720 14044 18748
rect 12897 18711 12955 18717
rect 7466 18640 7472 18692
rect 7524 18680 7530 18692
rect 10318 18680 10324 18692
rect 7524 18652 10324 18680
rect 7524 18640 7530 18652
rect 10318 18640 10324 18652
rect 10376 18640 10382 18692
rect 7742 18572 7748 18624
rect 7800 18612 7806 18624
rect 8665 18615 8723 18621
rect 8665 18612 8677 18615
rect 7800 18584 8677 18612
rect 7800 18572 7806 18584
rect 8665 18581 8677 18584
rect 8711 18581 8723 18615
rect 9122 18612 9128 18624
rect 9083 18584 9128 18612
rect 8665 18575 8723 18581
rect 9122 18572 9128 18584
rect 9180 18572 9186 18624
rect 13556 18612 13584 18720
rect 14016 18692 14044 18720
rect 15289 18717 15301 18751
rect 15335 18748 15347 18751
rect 15838 18748 15844 18760
rect 15335 18720 15844 18748
rect 15335 18717 15347 18720
rect 15289 18711 15347 18717
rect 15838 18708 15844 18720
rect 15896 18748 15902 18760
rect 15933 18751 15991 18757
rect 15933 18748 15945 18751
rect 15896 18720 15945 18748
rect 15896 18708 15902 18720
rect 15933 18717 15945 18720
rect 15979 18717 15991 18751
rect 15933 18711 15991 18717
rect 21726 18708 21732 18760
rect 21784 18748 21790 18760
rect 21821 18751 21879 18757
rect 21821 18748 21833 18751
rect 21784 18720 21833 18748
rect 21784 18708 21790 18720
rect 21821 18717 21833 18720
rect 21867 18748 21879 18751
rect 21913 18751 21971 18757
rect 21913 18748 21925 18751
rect 21867 18720 21925 18748
rect 21867 18717 21879 18720
rect 21821 18711 21879 18717
rect 21913 18717 21925 18720
rect 21959 18717 21971 18751
rect 22186 18748 22192 18760
rect 22147 18720 22192 18748
rect 21913 18711 21971 18717
rect 22186 18708 22192 18720
rect 22244 18708 22250 18760
rect 13998 18640 14004 18692
rect 14056 18640 14062 18692
rect 14366 18612 14372 18624
rect 13556 18584 14372 18612
rect 14366 18572 14372 18584
rect 14424 18612 14430 18624
rect 14461 18615 14519 18621
rect 14461 18612 14473 18615
rect 14424 18584 14473 18612
rect 14424 18572 14430 18584
rect 14461 18581 14473 18584
rect 14507 18581 14519 18615
rect 15562 18612 15568 18624
rect 15523 18584 15568 18612
rect 14461 18575 14519 18581
rect 15562 18572 15568 18584
rect 15620 18572 15626 18624
rect 18230 18612 18236 18624
rect 18191 18584 18236 18612
rect 18230 18572 18236 18584
rect 18288 18572 18294 18624
rect 23477 18615 23535 18621
rect 23477 18581 23489 18615
rect 23523 18612 23535 18615
rect 24765 18615 24823 18621
rect 24765 18612 24777 18615
rect 23523 18584 24777 18612
rect 23523 18581 23535 18584
rect 23477 18575 23535 18581
rect 24765 18581 24777 18584
rect 24811 18581 24823 18615
rect 24765 18575 24823 18581
rect 1104 18522 24656 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 24656 18522
rect 1104 18448 24656 18470
rect 4341 18411 4399 18417
rect 4341 18377 4353 18411
rect 4387 18408 4399 18411
rect 4982 18408 4988 18420
rect 4387 18380 4988 18408
rect 4387 18377 4399 18380
rect 4341 18371 4399 18377
rect 2501 18275 2559 18281
rect 2501 18241 2513 18275
rect 2547 18272 2559 18275
rect 4246 18272 4252 18284
rect 2547 18244 4252 18272
rect 2547 18241 2559 18244
rect 2501 18235 2559 18241
rect 4246 18232 4252 18244
rect 4304 18232 4310 18284
rect 2777 18207 2835 18213
rect 2777 18173 2789 18207
rect 2823 18204 2835 18207
rect 4356 18204 4384 18371
rect 4982 18368 4988 18380
rect 5040 18368 5046 18420
rect 5813 18411 5871 18417
rect 5813 18377 5825 18411
rect 5859 18408 5871 18411
rect 5994 18408 6000 18420
rect 5859 18380 6000 18408
rect 5859 18377 5871 18380
rect 5813 18371 5871 18377
rect 5994 18368 6000 18380
rect 6052 18368 6058 18420
rect 9030 18408 9036 18420
rect 8991 18380 9036 18408
rect 9030 18368 9036 18380
rect 9088 18368 9094 18420
rect 10965 18411 11023 18417
rect 10965 18377 10977 18411
rect 11011 18408 11023 18411
rect 12618 18408 12624 18420
rect 11011 18380 12624 18408
rect 11011 18377 11023 18380
rect 10965 18371 11023 18377
rect 12618 18368 12624 18380
rect 12676 18368 12682 18420
rect 15286 18368 15292 18420
rect 15344 18408 15350 18420
rect 16117 18411 16175 18417
rect 16117 18408 16129 18411
rect 15344 18380 16129 18408
rect 15344 18368 15350 18380
rect 16117 18377 16129 18380
rect 16163 18408 16175 18411
rect 16209 18411 16267 18417
rect 16209 18408 16221 18411
rect 16163 18380 16221 18408
rect 16163 18377 16175 18380
rect 16117 18371 16175 18377
rect 16209 18377 16221 18380
rect 16255 18377 16267 18411
rect 18690 18408 18696 18420
rect 18651 18380 18696 18408
rect 16209 18371 16267 18377
rect 18690 18368 18696 18380
rect 18748 18368 18754 18420
rect 22186 18408 22192 18420
rect 22147 18380 22192 18408
rect 22186 18368 22192 18380
rect 22244 18368 22250 18420
rect 6454 18300 6460 18352
rect 6512 18340 6518 18352
rect 9674 18340 9680 18352
rect 6512 18312 9680 18340
rect 6512 18300 6518 18312
rect 9674 18300 9680 18312
rect 9732 18300 9738 18352
rect 10778 18300 10784 18352
rect 10836 18340 10842 18352
rect 12526 18340 12532 18352
rect 10836 18312 12532 18340
rect 10836 18300 10842 18312
rect 12526 18300 12532 18312
rect 12584 18340 12590 18352
rect 18785 18343 18843 18349
rect 18785 18340 18797 18343
rect 12584 18312 18797 18340
rect 12584 18300 12590 18312
rect 18785 18309 18797 18312
rect 18831 18309 18843 18343
rect 20162 18340 20168 18352
rect 18785 18303 18843 18309
rect 19628 18312 20168 18340
rect 7469 18275 7527 18281
rect 7469 18241 7481 18275
rect 7515 18272 7527 18275
rect 13265 18275 13323 18281
rect 13265 18272 13277 18275
rect 7515 18244 13277 18272
rect 7515 18241 7527 18244
rect 7469 18235 7527 18241
rect 13265 18241 13277 18244
rect 13311 18241 13323 18275
rect 13265 18235 13323 18241
rect 13630 18232 13636 18284
rect 13688 18272 13694 18284
rect 16117 18275 16175 18281
rect 13688 18244 13952 18272
rect 13688 18232 13694 18244
rect 5626 18204 5632 18216
rect 2823 18176 4384 18204
rect 5587 18176 5632 18204
rect 2823 18173 2835 18176
rect 2777 18167 2835 18173
rect 5626 18164 5632 18176
rect 5684 18164 5690 18216
rect 7837 18207 7895 18213
rect 7837 18173 7849 18207
rect 7883 18173 7895 18207
rect 8018 18204 8024 18216
rect 7979 18176 8024 18204
rect 7837 18167 7895 18173
rect 7852 18136 7880 18167
rect 8018 18164 8024 18176
rect 8076 18164 8082 18216
rect 8205 18207 8263 18213
rect 8205 18173 8217 18207
rect 8251 18204 8263 18207
rect 8481 18207 8539 18213
rect 8251 18176 8432 18204
rect 8251 18173 8263 18176
rect 8205 18167 8263 18173
rect 8294 18136 8300 18148
rect 7852 18108 8300 18136
rect 8294 18096 8300 18108
rect 8352 18096 8358 18148
rect 3878 18068 3884 18080
rect 3839 18040 3884 18068
rect 3878 18028 3884 18040
rect 3936 18028 3942 18080
rect 4246 18028 4252 18080
rect 4304 18068 4310 18080
rect 4525 18071 4583 18077
rect 4525 18068 4537 18071
rect 4304 18040 4537 18068
rect 4304 18028 4310 18040
rect 4525 18037 4537 18040
rect 4571 18068 4583 18071
rect 4982 18068 4988 18080
rect 4571 18040 4988 18068
rect 4571 18037 4583 18040
rect 4525 18031 4583 18037
rect 4982 18028 4988 18040
rect 5040 18028 5046 18080
rect 8404 18068 8432 18176
rect 8481 18173 8493 18207
rect 8527 18204 8539 18207
rect 9030 18204 9036 18216
rect 8527 18176 9036 18204
rect 8527 18173 8539 18176
rect 8481 18167 8539 18173
rect 9030 18164 9036 18176
rect 9088 18164 9094 18216
rect 9214 18164 9220 18216
rect 9272 18204 9278 18216
rect 10781 18207 10839 18213
rect 10781 18204 10793 18207
rect 9272 18176 10793 18204
rect 9272 18164 9278 18176
rect 10781 18173 10793 18176
rect 10827 18173 10839 18207
rect 10781 18167 10839 18173
rect 13078 18164 13084 18216
rect 13136 18204 13142 18216
rect 13648 18204 13676 18232
rect 13924 18213 13952 18244
rect 16117 18241 16129 18275
rect 16163 18272 16175 18275
rect 16393 18275 16451 18281
rect 16393 18272 16405 18275
rect 16163 18244 16405 18272
rect 16163 18241 16175 18244
rect 16117 18235 16175 18241
rect 16393 18241 16405 18244
rect 16439 18241 16451 18275
rect 16393 18235 16451 18241
rect 13136 18176 13676 18204
rect 13817 18207 13875 18213
rect 13136 18164 13142 18176
rect 13817 18173 13829 18207
rect 13863 18173 13875 18207
rect 13817 18167 13875 18173
rect 13909 18207 13967 18213
rect 13909 18173 13921 18207
rect 13955 18173 13967 18207
rect 13909 18167 13967 18173
rect 8941 18139 8999 18145
rect 8941 18105 8953 18139
rect 8987 18136 8999 18139
rect 9398 18136 9404 18148
rect 8987 18108 9404 18136
rect 8987 18105 8999 18108
rect 8941 18099 8999 18105
rect 9398 18096 9404 18108
rect 9456 18096 9462 18148
rect 8570 18068 8576 18080
rect 8404 18040 8576 18068
rect 8570 18028 8576 18040
rect 8628 18068 8634 18080
rect 9309 18071 9367 18077
rect 9309 18068 9321 18071
rect 8628 18040 9321 18068
rect 8628 18028 8634 18040
rect 9309 18037 9321 18040
rect 9355 18068 9367 18071
rect 9490 18068 9496 18080
rect 9355 18040 9496 18068
rect 9355 18037 9367 18040
rect 9309 18031 9367 18037
rect 9490 18028 9496 18040
rect 9548 18028 9554 18080
rect 13832 18068 13860 18167
rect 13998 18164 14004 18216
rect 14056 18204 14062 18216
rect 14093 18207 14151 18213
rect 14093 18204 14105 18207
rect 14056 18176 14105 18204
rect 14056 18164 14062 18176
rect 14093 18173 14105 18176
rect 14139 18173 14151 18207
rect 14093 18167 14151 18173
rect 14553 18207 14611 18213
rect 14553 18173 14565 18207
rect 14599 18173 14611 18207
rect 14553 18167 14611 18173
rect 14737 18207 14795 18213
rect 14737 18173 14749 18207
rect 14783 18204 14795 18207
rect 15378 18204 15384 18216
rect 14783 18176 15384 18204
rect 14783 18173 14795 18176
rect 14737 18167 14795 18173
rect 14090 18068 14096 18080
rect 13832 18040 14096 18068
rect 14090 18028 14096 18040
rect 14148 18028 14154 18080
rect 14568 18068 14596 18167
rect 15378 18164 15384 18176
rect 15436 18204 15442 18216
rect 16485 18207 16543 18213
rect 16485 18204 16497 18207
rect 15436 18176 16497 18204
rect 15436 18164 15442 18176
rect 16485 18173 16497 18176
rect 16531 18204 16543 18207
rect 18046 18204 18052 18216
rect 16531 18176 18052 18204
rect 16531 18173 16543 18176
rect 16485 18167 16543 18173
rect 18046 18164 18052 18176
rect 18104 18164 18110 18216
rect 18800 18204 18828 18303
rect 19628 18213 19656 18312
rect 20162 18300 20168 18312
rect 20220 18300 20226 18352
rect 21174 18300 21180 18352
rect 21232 18340 21238 18352
rect 21818 18340 21824 18352
rect 21232 18312 21824 18340
rect 21232 18300 21238 18312
rect 21818 18300 21824 18312
rect 21876 18300 21882 18352
rect 19705 18275 19763 18281
rect 19705 18241 19717 18275
rect 19751 18272 19763 18275
rect 19751 18244 21404 18272
rect 19751 18241 19763 18244
rect 19705 18235 19763 18241
rect 19613 18207 19671 18213
rect 19613 18204 19625 18207
rect 18800 18176 19625 18204
rect 19613 18173 19625 18176
rect 19659 18173 19671 18207
rect 19935 18207 19993 18213
rect 19935 18204 19947 18207
rect 19613 18167 19671 18173
rect 19720 18176 19947 18204
rect 16942 18136 16948 18148
rect 16903 18108 16948 18136
rect 16942 18096 16948 18108
rect 17000 18096 17006 18148
rect 18690 18096 18696 18148
rect 18748 18136 18754 18148
rect 19720 18136 19748 18176
rect 19935 18173 19947 18176
rect 19981 18173 19993 18207
rect 19935 18167 19993 18173
rect 20165 18207 20223 18213
rect 20165 18173 20177 18207
rect 20211 18173 20223 18207
rect 20165 18167 20223 18173
rect 18748 18108 19748 18136
rect 20180 18136 20208 18167
rect 20714 18164 20720 18216
rect 20772 18204 20778 18216
rect 20993 18207 21051 18213
rect 20993 18204 21005 18207
rect 20772 18176 21005 18204
rect 20772 18164 20778 18176
rect 20993 18173 21005 18176
rect 21039 18173 21051 18207
rect 21174 18204 21180 18216
rect 21135 18176 21180 18204
rect 20993 18167 21051 18173
rect 21174 18164 21180 18176
rect 21232 18164 21238 18216
rect 21376 18204 21404 18244
rect 21634 18204 21640 18216
rect 21376 18176 21640 18204
rect 21634 18164 21640 18176
rect 21692 18164 21698 18216
rect 21729 18207 21787 18213
rect 21729 18173 21741 18207
rect 21775 18204 21787 18207
rect 21818 18204 21824 18216
rect 21775 18176 21824 18204
rect 21775 18173 21787 18176
rect 21729 18167 21787 18173
rect 21818 18164 21824 18176
rect 21876 18164 21882 18216
rect 22278 18136 22284 18148
rect 20180 18108 22284 18136
rect 18748 18096 18754 18108
rect 14921 18071 14979 18077
rect 14921 18068 14933 18071
rect 14568 18040 14933 18068
rect 14921 18037 14933 18040
rect 14967 18068 14979 18071
rect 17586 18068 17592 18080
rect 14967 18040 17592 18068
rect 14967 18037 14979 18040
rect 14921 18031 14979 18037
rect 17586 18028 17592 18040
rect 17644 18028 17650 18080
rect 19245 18071 19303 18077
rect 19245 18037 19257 18071
rect 19291 18068 19303 18071
rect 19426 18068 19432 18080
rect 19291 18040 19432 18068
rect 19291 18037 19303 18040
rect 19245 18031 19303 18037
rect 19426 18028 19432 18040
rect 19484 18028 19490 18080
rect 19720 18068 19748 18108
rect 22278 18096 22284 18108
rect 22336 18096 22342 18148
rect 19978 18068 19984 18080
rect 19720 18040 19984 18068
rect 19978 18028 19984 18040
rect 20036 18028 20042 18080
rect 20714 18028 20720 18080
rect 20772 18068 20778 18080
rect 20809 18071 20867 18077
rect 20809 18068 20821 18071
rect 20772 18040 20821 18068
rect 20772 18028 20778 18040
rect 20809 18037 20821 18040
rect 20855 18037 20867 18071
rect 20809 18031 20867 18037
rect 24765 18003 24823 18009
rect 1104 17978 24656 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 24656 17978
rect 24765 17969 24777 18003
rect 24811 17969 24823 18003
rect 24765 17963 24823 17969
rect 1104 17904 24656 17926
rect 24780 17932 24808 17963
rect 26970 17932 26976 17944
rect 24780 17904 26976 17932
rect 6546 17824 6552 17876
rect 6604 17864 6610 17876
rect 12986 17864 12992 17876
rect 6604 17836 12992 17864
rect 6604 17824 6610 17836
rect 12986 17824 12992 17836
rect 13044 17864 13050 17876
rect 13998 17864 14004 17876
rect 13044 17836 14004 17864
rect 13044 17824 13050 17836
rect 13998 17824 14004 17836
rect 14056 17824 14062 17876
rect 21634 17824 21640 17876
rect 21692 17864 21698 17876
rect 22833 17867 22891 17873
rect 22833 17864 22845 17867
rect 21692 17836 22845 17864
rect 21692 17824 21698 17836
rect 22833 17833 22845 17836
rect 22879 17833 22891 17867
rect 22833 17827 22891 17833
rect 23109 17867 23167 17873
rect 23109 17833 23121 17867
rect 23155 17864 23167 17867
rect 24780 17864 24808 17904
rect 26970 17892 26976 17904
rect 27028 17892 27034 17944
rect 23155 17836 24808 17864
rect 23155 17833 23167 17836
rect 23109 17827 23167 17833
rect 5460 17768 6776 17796
rect 4341 17731 4399 17737
rect 4341 17697 4353 17731
rect 4387 17728 4399 17731
rect 4614 17728 4620 17740
rect 4387 17700 4620 17728
rect 4387 17697 4399 17700
rect 4341 17691 4399 17697
rect 4614 17688 4620 17700
rect 4672 17688 4678 17740
rect 5460 17737 5488 17768
rect 6748 17740 6776 17768
rect 5445 17731 5503 17737
rect 5445 17697 5457 17731
rect 5491 17697 5503 17731
rect 6546 17728 6552 17740
rect 6507 17700 6552 17728
rect 5445 17691 5503 17697
rect 6546 17688 6552 17700
rect 6604 17688 6610 17740
rect 6730 17688 6736 17740
rect 6788 17728 6794 17740
rect 6825 17731 6883 17737
rect 6825 17728 6837 17731
rect 6788 17700 6837 17728
rect 6788 17688 6794 17700
rect 6825 17697 6837 17700
rect 6871 17697 6883 17731
rect 8205 17731 8263 17737
rect 8205 17728 8217 17731
rect 6825 17691 6883 17697
rect 7208 17700 8217 17728
rect 4525 17595 4583 17601
rect 4525 17561 4537 17595
rect 4571 17592 4583 17595
rect 5902 17592 5908 17604
rect 4571 17564 5908 17592
rect 4571 17561 4583 17564
rect 4525 17555 4583 17561
rect 5902 17552 5908 17564
rect 5960 17592 5966 17604
rect 6641 17595 6699 17601
rect 6641 17592 6653 17595
rect 5960 17564 6653 17592
rect 5960 17552 5966 17564
rect 6641 17561 6653 17564
rect 6687 17592 6699 17595
rect 7208 17592 7236 17700
rect 8205 17697 8217 17700
rect 8251 17697 8263 17731
rect 8205 17691 8263 17697
rect 12066 17688 12072 17740
rect 12124 17728 12130 17740
rect 13081 17731 13139 17737
rect 13081 17728 13093 17731
rect 12124 17700 13093 17728
rect 12124 17688 12130 17700
rect 13081 17697 13093 17700
rect 13127 17697 13139 17731
rect 13081 17691 13139 17697
rect 18046 17688 18052 17740
rect 18104 17728 18110 17740
rect 18233 17731 18291 17737
rect 18233 17728 18245 17731
rect 18104 17700 18245 17728
rect 18104 17688 18110 17700
rect 18233 17697 18245 17700
rect 18279 17697 18291 17731
rect 18233 17691 18291 17697
rect 19426 17688 19432 17740
rect 19484 17728 19490 17740
rect 19521 17731 19579 17737
rect 19521 17728 19533 17731
rect 19484 17700 19533 17728
rect 19484 17688 19490 17700
rect 19521 17697 19533 17700
rect 19567 17697 19579 17731
rect 19521 17691 19579 17697
rect 22741 17731 22799 17737
rect 22741 17697 22753 17731
rect 22787 17728 22799 17731
rect 23124 17728 23152 17827
rect 22787 17700 23152 17728
rect 22787 17697 22799 17700
rect 22741 17691 22799 17697
rect 7285 17663 7343 17669
rect 7285 17629 7297 17663
rect 7331 17629 7343 17663
rect 7285 17623 7343 17629
rect 6687 17564 7236 17592
rect 7300 17592 7328 17623
rect 8018 17620 8024 17672
rect 8076 17660 8082 17672
rect 8113 17663 8171 17669
rect 8113 17660 8125 17663
rect 8076 17632 8125 17660
rect 8076 17620 8082 17632
rect 8113 17629 8125 17632
rect 8159 17629 8171 17663
rect 8113 17623 8171 17629
rect 18141 17663 18199 17669
rect 18141 17629 18153 17663
rect 18187 17660 18199 17663
rect 18322 17660 18328 17672
rect 18187 17632 18328 17660
rect 18187 17629 18199 17632
rect 18141 17623 18199 17629
rect 18322 17620 18328 17632
rect 18380 17660 18386 17672
rect 18785 17663 18843 17669
rect 18785 17660 18797 17663
rect 18380 17632 18797 17660
rect 18380 17620 18386 17632
rect 18785 17629 18797 17632
rect 18831 17629 18843 17663
rect 18785 17623 18843 17629
rect 9122 17592 9128 17604
rect 7300 17564 9128 17592
rect 6687 17561 6699 17564
rect 6641 17555 6699 17561
rect 9122 17552 9128 17564
rect 9180 17552 9186 17604
rect 12066 17552 12072 17604
rect 12124 17592 12130 17604
rect 15930 17592 15936 17604
rect 12124 17564 15936 17592
rect 12124 17552 12130 17564
rect 15930 17552 15936 17564
rect 15988 17552 15994 17604
rect 16666 17552 16672 17604
rect 16724 17592 16730 17604
rect 19613 17595 19671 17601
rect 19613 17592 19625 17595
rect 16724 17564 19625 17592
rect 16724 17552 16730 17564
rect 19613 17561 19625 17564
rect 19659 17561 19671 17595
rect 19613 17555 19671 17561
rect 5629 17527 5687 17533
rect 5629 17493 5641 17527
rect 5675 17524 5687 17527
rect 7006 17524 7012 17536
rect 5675 17496 7012 17524
rect 5675 17493 5687 17496
rect 5629 17487 5687 17493
rect 7006 17484 7012 17496
rect 7064 17524 7070 17536
rect 7650 17524 7656 17536
rect 7064 17496 7656 17524
rect 7064 17484 7070 17496
rect 7650 17484 7656 17496
rect 7708 17484 7714 17536
rect 8294 17484 8300 17536
rect 8352 17524 8358 17536
rect 8389 17527 8447 17533
rect 8389 17524 8401 17527
rect 8352 17496 8401 17524
rect 8352 17484 8358 17496
rect 8389 17493 8401 17496
rect 8435 17524 8447 17527
rect 13078 17524 13084 17536
rect 8435 17496 13084 17524
rect 8435 17493 8447 17496
rect 8389 17487 8447 17493
rect 13078 17484 13084 17496
rect 13136 17484 13142 17536
rect 13173 17527 13231 17533
rect 13173 17493 13185 17527
rect 13219 17524 13231 17527
rect 14182 17524 14188 17536
rect 13219 17496 14188 17524
rect 13219 17493 13231 17496
rect 13173 17487 13231 17493
rect 14182 17484 14188 17496
rect 14240 17484 14246 17536
rect 18414 17524 18420 17536
rect 18375 17496 18420 17524
rect 18414 17484 18420 17496
rect 18472 17484 18478 17536
rect 1104 17434 24656 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 24656 17434
rect 1104 17360 24656 17382
rect 4065 17323 4123 17329
rect 4065 17289 4077 17323
rect 4111 17320 4123 17323
rect 6546 17320 6552 17332
rect 4111 17292 6552 17320
rect 4111 17289 4123 17292
rect 4065 17283 4123 17289
rect 6546 17280 6552 17292
rect 6604 17280 6610 17332
rect 15562 17320 15568 17332
rect 14660 17292 15568 17320
rect 5810 17212 5816 17264
rect 5868 17252 5874 17264
rect 10226 17252 10232 17264
rect 5868 17224 10232 17252
rect 5868 17212 5874 17224
rect 10226 17212 10232 17224
rect 10284 17212 10290 17264
rect 5718 17184 5724 17196
rect 5679 17156 5724 17184
rect 5718 17144 5724 17156
rect 5776 17144 5782 17196
rect 7929 17187 7987 17193
rect 7929 17184 7941 17187
rect 7300 17156 7941 17184
rect 2869 17119 2927 17125
rect 2869 17085 2881 17119
rect 2915 17085 2927 17119
rect 3878 17116 3884 17128
rect 3839 17088 3884 17116
rect 2869 17079 2927 17085
rect 2884 16992 2912 17079
rect 3878 17076 3884 17088
rect 3936 17116 3942 17128
rect 4985 17119 5043 17125
rect 4985 17116 4997 17119
rect 3936 17088 4997 17116
rect 3936 17076 3942 17088
rect 4985 17085 4997 17088
rect 5031 17085 5043 17119
rect 4985 17079 5043 17085
rect 5077 17119 5135 17125
rect 5077 17085 5089 17119
rect 5123 17085 5135 17119
rect 5077 17079 5135 17085
rect 5261 17119 5319 17125
rect 5261 17085 5273 17119
rect 5307 17116 5319 17119
rect 5350 17116 5356 17128
rect 5307 17088 5356 17116
rect 5307 17085 5319 17088
rect 5261 17079 5319 17085
rect 2961 17051 3019 17057
rect 2961 17017 2973 17051
rect 3007 17048 3019 17051
rect 4614 17048 4620 17060
rect 3007 17020 4620 17048
rect 3007 17017 3019 17020
rect 2961 17011 3019 17017
rect 4614 17008 4620 17020
rect 4672 17008 4678 17060
rect 2777 16983 2835 16989
rect 2777 16949 2789 16983
rect 2823 16980 2835 16983
rect 2866 16980 2872 16992
rect 2823 16952 2872 16980
rect 2823 16949 2835 16952
rect 2777 16943 2835 16949
rect 2866 16940 2872 16952
rect 2924 16980 2930 16992
rect 4801 16983 4859 16989
rect 4801 16980 4813 16983
rect 2924 16952 4813 16980
rect 2924 16940 2930 16952
rect 4801 16949 4813 16952
rect 4847 16980 4859 16983
rect 5092 16980 5120 17079
rect 5350 17076 5356 17088
rect 5408 17076 5414 17128
rect 7006 17076 7012 17128
rect 7064 17116 7070 17128
rect 7300 17125 7328 17156
rect 7929 17153 7941 17156
rect 7975 17153 7987 17187
rect 14182 17184 14188 17196
rect 14143 17156 14188 17184
rect 7929 17147 7987 17153
rect 14182 17144 14188 17156
rect 14240 17144 14246 17196
rect 14660 17184 14688 17292
rect 15562 17280 15568 17292
rect 15620 17280 15626 17332
rect 15930 17280 15936 17332
rect 15988 17320 15994 17332
rect 19429 17323 19487 17329
rect 19429 17320 19441 17323
rect 15988 17292 19441 17320
rect 15988 17280 15994 17292
rect 19429 17289 19441 17292
rect 19475 17289 19487 17323
rect 19978 17320 19984 17332
rect 19939 17292 19984 17320
rect 19429 17283 19487 17289
rect 19978 17280 19984 17292
rect 20036 17280 20042 17332
rect 20162 17320 20168 17332
rect 20123 17292 20168 17320
rect 20162 17280 20168 17292
rect 20220 17320 20226 17332
rect 27062 17320 27068 17332
rect 20220 17292 21404 17320
rect 20220 17280 20226 17292
rect 15841 17255 15899 17261
rect 15841 17221 15853 17255
rect 15887 17252 15899 17255
rect 16482 17252 16488 17264
rect 15887 17224 16488 17252
rect 15887 17221 15899 17224
rect 15841 17215 15899 17221
rect 15856 17184 15884 17215
rect 16482 17212 16488 17224
rect 16540 17252 16546 17264
rect 19886 17252 19892 17264
rect 16540 17224 19380 17252
rect 19847 17224 19892 17252
rect 16540 17212 16546 17224
rect 14568 17156 14688 17184
rect 15028 17156 15884 17184
rect 18049 17187 18107 17193
rect 7285 17119 7343 17125
rect 7285 17116 7297 17119
rect 7064 17088 7297 17116
rect 7064 17076 7070 17088
rect 7285 17085 7297 17088
rect 7331 17085 7343 17119
rect 7466 17116 7472 17128
rect 7427 17088 7472 17116
rect 7285 17079 7343 17085
rect 7466 17076 7472 17088
rect 7524 17076 7530 17128
rect 7650 17116 7656 17128
rect 7611 17088 7656 17116
rect 7650 17076 7656 17088
rect 7708 17076 7714 17128
rect 8294 17116 8300 17128
rect 8255 17088 8300 17116
rect 8294 17076 8300 17088
rect 8352 17076 8358 17128
rect 9122 17116 9128 17128
rect 9083 17088 9128 17116
rect 9122 17076 9128 17088
rect 9180 17076 9186 17128
rect 10962 17116 10968 17128
rect 10923 17088 10968 17116
rect 10962 17076 10968 17088
rect 11020 17076 11026 17128
rect 11146 17125 11152 17128
rect 11098 17119 11152 17125
rect 11098 17085 11110 17119
rect 11144 17085 11152 17119
rect 11098 17079 11152 17085
rect 11146 17076 11152 17079
rect 11204 17076 11210 17128
rect 14568 17125 14596 17156
rect 14553 17119 14611 17125
rect 14553 17085 14565 17119
rect 14599 17085 14611 17119
rect 14734 17116 14740 17128
rect 14695 17088 14740 17116
rect 14553 17079 14611 17085
rect 14734 17076 14740 17088
rect 14792 17076 14798 17128
rect 15028 17125 15056 17156
rect 18049 17153 18061 17187
rect 18095 17184 18107 17187
rect 18138 17184 18144 17196
rect 18095 17156 18144 17184
rect 18095 17153 18107 17156
rect 18049 17147 18107 17153
rect 18138 17144 18144 17156
rect 18196 17144 18202 17196
rect 19150 17184 19156 17196
rect 18892 17156 19156 17184
rect 15013 17119 15071 17125
rect 15013 17085 15025 17119
rect 15059 17085 15071 17119
rect 15194 17116 15200 17128
rect 15107 17088 15200 17116
rect 15013 17079 15071 17085
rect 15194 17076 15200 17088
rect 15252 17116 15258 17128
rect 16945 17119 17003 17125
rect 15252 17088 15332 17116
rect 15252 17076 15258 17088
rect 6825 17051 6883 17057
rect 6825 17017 6837 17051
rect 6871 17048 6883 17051
rect 11164 17048 11192 17076
rect 11514 17048 11520 17060
rect 6871 17020 11192 17048
rect 11475 17020 11520 17048
rect 6871 17017 6883 17020
rect 6825 17011 6883 17017
rect 11514 17008 11520 17020
rect 11572 17008 11578 17060
rect 15304 17048 15332 17088
rect 16945 17085 16957 17119
rect 16991 17116 17003 17119
rect 17034 17116 17040 17128
rect 16991 17088 17040 17116
rect 16991 17085 17003 17088
rect 16945 17079 17003 17085
rect 17034 17076 17040 17088
rect 17092 17076 17098 17128
rect 18230 17116 18236 17128
rect 18191 17088 18236 17116
rect 18230 17076 18236 17088
rect 18288 17076 18294 17128
rect 18598 17116 18604 17128
rect 18559 17088 18604 17116
rect 18598 17076 18604 17088
rect 18656 17076 18662 17128
rect 18892 17125 18920 17156
rect 19150 17144 19156 17156
rect 19208 17144 19214 17196
rect 18877 17119 18935 17125
rect 18877 17085 18889 17119
rect 18923 17085 18935 17119
rect 19058 17116 19064 17128
rect 19019 17088 19064 17116
rect 18877 17079 18935 17085
rect 19058 17076 19064 17088
rect 19116 17076 19122 17128
rect 18966 17048 18972 17060
rect 15304 17020 18972 17048
rect 18966 17008 18972 17020
rect 19024 17008 19030 17060
rect 19352 17048 19380 17224
rect 19886 17212 19892 17224
rect 19944 17212 19950 17264
rect 19996 17252 20024 17280
rect 19996 17224 21036 17252
rect 20806 17184 20812 17196
rect 20767 17156 20812 17184
rect 20806 17144 20812 17156
rect 20864 17144 20870 17196
rect 19426 17076 19432 17128
rect 19484 17116 19490 17128
rect 21008 17125 21036 17224
rect 21376 17125 21404 17292
rect 21652 17292 27068 17320
rect 20349 17119 20407 17125
rect 20349 17116 20361 17119
rect 19484 17088 20361 17116
rect 19484 17076 19490 17088
rect 20349 17085 20361 17088
rect 20395 17085 20407 17119
rect 20349 17079 20407 17085
rect 20993 17119 21051 17125
rect 20993 17085 21005 17119
rect 21039 17085 21051 17119
rect 20993 17079 21051 17085
rect 21361 17119 21419 17125
rect 21361 17085 21373 17119
rect 21407 17085 21419 17119
rect 21542 17116 21548 17128
rect 21503 17088 21548 17116
rect 21361 17079 21419 17085
rect 21542 17076 21548 17088
rect 21600 17076 21606 17128
rect 21652 17048 21680 17292
rect 27062 17280 27068 17292
rect 27120 17280 27126 17332
rect 21818 17212 21824 17264
rect 21876 17252 21882 17264
rect 23293 17255 23351 17261
rect 23293 17252 23305 17255
rect 21876 17224 23305 17252
rect 21876 17212 21882 17224
rect 23293 17221 23305 17224
rect 23339 17221 23351 17255
rect 23293 17215 23351 17221
rect 23477 17119 23535 17125
rect 23477 17085 23489 17119
rect 23523 17116 23535 17119
rect 24118 17116 24124 17128
rect 23523 17088 24124 17116
rect 23523 17085 23535 17088
rect 23477 17079 23535 17085
rect 24118 17076 24124 17088
rect 24176 17076 24182 17128
rect 19352 17020 21680 17048
rect 7834 16980 7840 16992
rect 4847 16952 7840 16980
rect 4847 16949 4859 16952
rect 4801 16943 4859 16949
rect 7834 16940 7840 16952
rect 7892 16940 7898 16992
rect 9306 16980 9312 16992
rect 9267 16952 9312 16980
rect 9306 16940 9312 16952
rect 9364 16940 9370 16992
rect 10873 16983 10931 16989
rect 10873 16949 10885 16983
rect 10919 16980 10931 16983
rect 10962 16980 10968 16992
rect 10919 16952 10968 16980
rect 10919 16949 10931 16952
rect 10873 16943 10931 16949
rect 10962 16940 10968 16952
rect 11020 16980 11026 16992
rect 12434 16980 12440 16992
rect 11020 16952 12440 16980
rect 11020 16940 11026 16952
rect 12434 16940 12440 16952
rect 12492 16940 12498 16992
rect 15562 16980 15568 16992
rect 15523 16952 15568 16980
rect 15562 16940 15568 16952
rect 15620 16940 15626 16992
rect 17037 16983 17095 16989
rect 17037 16949 17049 16983
rect 17083 16980 17095 16983
rect 18046 16980 18052 16992
rect 17083 16952 18052 16980
rect 17083 16949 17095 16952
rect 17037 16943 17095 16949
rect 18046 16940 18052 16952
rect 18104 16940 18110 16992
rect 19058 16940 19064 16992
rect 19116 16980 19122 16992
rect 19613 16983 19671 16989
rect 19613 16980 19625 16983
rect 19116 16952 19625 16980
rect 19116 16940 19122 16952
rect 19613 16949 19625 16952
rect 19659 16949 19671 16983
rect 19613 16943 19671 16949
rect 1104 16890 24656 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 24656 16890
rect 1104 16816 24656 16838
rect 3053 16779 3111 16785
rect 3053 16745 3065 16779
rect 3099 16776 3111 16779
rect 3878 16776 3884 16788
rect 3099 16748 3884 16776
rect 3099 16745 3111 16748
rect 3053 16739 3111 16745
rect 3878 16736 3884 16748
rect 3936 16736 3942 16788
rect 5350 16736 5356 16788
rect 5408 16776 5414 16788
rect 7282 16776 7288 16788
rect 5408 16748 7288 16776
rect 5408 16736 5414 16748
rect 7282 16736 7288 16748
rect 7340 16776 7346 16788
rect 8018 16776 8024 16788
rect 7340 16748 8024 16776
rect 7340 16736 7346 16748
rect 8018 16736 8024 16748
rect 8076 16736 8082 16788
rect 14734 16736 14740 16788
rect 14792 16776 14798 16788
rect 17218 16776 17224 16788
rect 14792 16748 17224 16776
rect 14792 16736 14798 16748
rect 17218 16736 17224 16748
rect 17276 16736 17282 16788
rect 21542 16736 21548 16788
rect 21600 16776 21606 16788
rect 22649 16779 22707 16785
rect 22649 16776 22661 16779
rect 21600 16748 22661 16776
rect 21600 16736 21606 16748
rect 22649 16745 22661 16748
rect 22695 16745 22707 16779
rect 22649 16739 22707 16745
rect 4614 16668 4620 16720
rect 4672 16708 4678 16720
rect 7193 16711 7251 16717
rect 4672 16680 6592 16708
rect 4672 16668 4678 16680
rect 2869 16643 2927 16649
rect 2869 16609 2881 16643
rect 2915 16640 2927 16643
rect 2961 16643 3019 16649
rect 2961 16640 2973 16643
rect 2915 16612 2973 16640
rect 2915 16609 2927 16612
rect 2869 16603 2927 16609
rect 2961 16609 2973 16612
rect 3007 16640 3019 16643
rect 4525 16643 4583 16649
rect 4525 16640 4537 16643
rect 3007 16612 4537 16640
rect 3007 16609 3019 16612
rect 2961 16603 3019 16609
rect 4525 16609 4537 16612
rect 4571 16640 4583 16643
rect 4890 16640 4896 16652
rect 4571 16612 4896 16640
rect 4571 16609 4583 16612
rect 4525 16603 4583 16609
rect 4890 16600 4896 16612
rect 4948 16600 4954 16652
rect 5000 16649 5028 16680
rect 4985 16643 5043 16649
rect 4985 16609 4997 16643
rect 5031 16609 5043 16643
rect 4985 16603 5043 16609
rect 5169 16643 5227 16649
rect 5169 16609 5181 16643
rect 5215 16609 5227 16643
rect 5169 16603 5227 16609
rect 5184 16572 5212 16603
rect 5626 16600 5632 16652
rect 5684 16640 5690 16652
rect 6564 16649 6592 16680
rect 7193 16677 7205 16711
rect 7239 16708 7251 16711
rect 9214 16708 9220 16720
rect 7239 16680 9220 16708
rect 7239 16677 7251 16680
rect 7193 16671 7251 16677
rect 9214 16668 9220 16680
rect 9272 16668 9278 16720
rect 10321 16711 10379 16717
rect 10321 16677 10333 16711
rect 10367 16708 10379 16711
rect 11330 16708 11336 16720
rect 10367 16680 11336 16708
rect 10367 16677 10379 16680
rect 10321 16671 10379 16677
rect 11330 16668 11336 16680
rect 11388 16668 11394 16720
rect 11790 16668 11796 16720
rect 11848 16668 11854 16720
rect 18322 16668 18328 16720
rect 18380 16708 18386 16720
rect 21818 16708 21824 16720
rect 18380 16680 21824 16708
rect 18380 16668 18386 16680
rect 21818 16668 21824 16680
rect 21876 16668 21882 16720
rect 6457 16643 6515 16649
rect 6457 16640 6469 16643
rect 5684 16612 6469 16640
rect 5684 16600 5690 16612
rect 6457 16609 6469 16612
rect 6503 16609 6515 16643
rect 6457 16603 6515 16609
rect 6549 16643 6607 16649
rect 6549 16609 6561 16643
rect 6595 16609 6607 16643
rect 6730 16640 6736 16652
rect 6691 16612 6736 16640
rect 6549 16603 6607 16609
rect 4816 16544 5212 16572
rect 5537 16575 5595 16581
rect 4816 16448 4844 16544
rect 5537 16541 5549 16575
rect 5583 16572 5595 16575
rect 5810 16572 5816 16584
rect 5583 16544 5816 16572
rect 5583 16541 5595 16544
rect 5537 16535 5595 16541
rect 5810 16532 5816 16544
rect 5868 16532 5874 16584
rect 6472 16572 6500 16603
rect 6730 16600 6736 16612
rect 6788 16600 6794 16652
rect 7834 16640 7840 16652
rect 7795 16612 7840 16640
rect 7834 16600 7840 16612
rect 7892 16640 7898 16652
rect 8021 16643 8079 16649
rect 8021 16640 8033 16643
rect 7892 16612 8033 16640
rect 7892 16600 7898 16612
rect 8021 16609 8033 16612
rect 8067 16609 8079 16643
rect 8021 16603 8079 16609
rect 9306 16600 9312 16652
rect 9364 16640 9370 16652
rect 10137 16643 10195 16649
rect 10137 16640 10149 16643
rect 9364 16612 10149 16640
rect 9364 16600 9370 16612
rect 10137 16609 10149 16612
rect 10183 16640 10195 16643
rect 10229 16643 10287 16649
rect 10229 16640 10241 16643
rect 10183 16612 10241 16640
rect 10183 16609 10195 16612
rect 10137 16603 10195 16609
rect 10229 16609 10241 16612
rect 10275 16609 10287 16643
rect 10229 16603 10287 16609
rect 11054 16600 11060 16652
rect 11112 16640 11118 16652
rect 11425 16643 11483 16649
rect 11425 16640 11437 16643
rect 11112 16612 11437 16640
rect 11112 16600 11118 16612
rect 11425 16609 11437 16612
rect 11471 16609 11483 16643
rect 11425 16603 11483 16609
rect 11514 16600 11520 16652
rect 11572 16649 11578 16652
rect 11572 16643 11630 16649
rect 11572 16609 11584 16643
rect 11618 16609 11630 16643
rect 11572 16603 11630 16609
rect 11572 16600 11578 16603
rect 7006 16572 7012 16584
rect 6472 16544 7012 16572
rect 7006 16532 7012 16544
rect 7064 16532 7070 16584
rect 11808 16581 11836 16668
rect 13078 16640 13084 16652
rect 13039 16612 13084 16640
rect 13078 16600 13084 16612
rect 13136 16600 13142 16652
rect 16666 16640 16672 16652
rect 16627 16612 16672 16640
rect 16666 16600 16672 16612
rect 16724 16600 16730 16652
rect 16942 16640 16948 16652
rect 16903 16612 16948 16640
rect 16942 16600 16948 16612
rect 17000 16600 17006 16652
rect 17218 16640 17224 16652
rect 17179 16612 17224 16640
rect 17218 16600 17224 16612
rect 17276 16600 17282 16652
rect 17310 16600 17316 16652
rect 17368 16640 17374 16652
rect 17405 16643 17463 16649
rect 17405 16640 17417 16643
rect 17368 16612 17417 16640
rect 17368 16600 17374 16612
rect 17405 16609 17417 16612
rect 17451 16609 17463 16643
rect 17586 16640 17592 16652
rect 17547 16612 17592 16640
rect 17405 16603 17463 16609
rect 11793 16575 11851 16581
rect 11793 16541 11805 16575
rect 11839 16541 11851 16575
rect 11793 16535 11851 16541
rect 11882 16532 11888 16584
rect 11940 16572 11946 16584
rect 12986 16572 12992 16584
rect 11940 16544 11985 16572
rect 12947 16544 12992 16572
rect 11940 16532 11946 16544
rect 12986 16532 12992 16544
rect 13044 16532 13050 16584
rect 13538 16572 13544 16584
rect 13499 16544 13544 16572
rect 13538 16532 13544 16544
rect 13596 16532 13602 16584
rect 17420 16572 17448 16603
rect 17586 16600 17592 16612
rect 17644 16600 17650 16652
rect 18506 16640 18512 16652
rect 17696 16612 18512 16640
rect 17696 16572 17724 16612
rect 18506 16600 18512 16612
rect 18564 16600 18570 16652
rect 18966 16640 18972 16652
rect 18927 16612 18972 16640
rect 18966 16600 18972 16612
rect 19024 16600 19030 16652
rect 22557 16643 22615 16649
rect 22557 16609 22569 16643
rect 22603 16640 22615 16643
rect 22646 16640 22652 16652
rect 22603 16612 22652 16640
rect 22603 16609 22615 16612
rect 22557 16603 22615 16609
rect 22646 16600 22652 16612
rect 22704 16640 22710 16652
rect 22833 16643 22891 16649
rect 22833 16640 22845 16643
rect 22704 16612 22845 16640
rect 22704 16600 22710 16612
rect 22833 16609 22845 16612
rect 22879 16640 22891 16643
rect 23566 16640 23572 16652
rect 22879 16612 23572 16640
rect 22879 16609 22891 16612
rect 22833 16603 22891 16609
rect 23566 16600 23572 16612
rect 23624 16600 23630 16652
rect 17954 16572 17960 16584
rect 17420 16544 17724 16572
rect 17915 16544 17960 16572
rect 17954 16532 17960 16544
rect 18012 16532 18018 16584
rect 7466 16464 7472 16516
rect 7524 16504 7530 16516
rect 8205 16507 8263 16513
rect 8205 16504 8217 16507
rect 7524 16476 8217 16504
rect 7524 16464 7530 16476
rect 8205 16473 8217 16476
rect 8251 16473 8263 16507
rect 11698 16504 11704 16516
rect 11659 16476 11704 16504
rect 8205 16467 8263 16473
rect 11698 16464 11704 16476
rect 11756 16464 11762 16516
rect 12434 16464 12440 16516
rect 12492 16504 12498 16516
rect 26878 16504 26884 16516
rect 12492 16476 26884 16504
rect 12492 16464 12498 16476
rect 26878 16464 26884 16476
rect 26936 16464 26942 16516
rect 4798 16436 4804 16448
rect 4759 16408 4804 16436
rect 4798 16396 4804 16408
rect 4856 16396 4862 16448
rect 16574 16396 16580 16448
rect 16632 16436 16638 16448
rect 17586 16436 17592 16448
rect 16632 16408 17592 16436
rect 16632 16396 16638 16408
rect 17586 16396 17592 16408
rect 17644 16436 17650 16448
rect 18233 16439 18291 16445
rect 18233 16436 18245 16439
rect 17644 16408 18245 16436
rect 17644 16396 17650 16408
rect 18233 16405 18245 16408
rect 18279 16436 18291 16439
rect 19058 16436 19064 16448
rect 18279 16408 19064 16436
rect 18279 16405 18291 16408
rect 18233 16399 18291 16405
rect 19058 16396 19064 16408
rect 19116 16436 19122 16448
rect 19153 16439 19211 16445
rect 19153 16436 19165 16439
rect 19116 16408 19165 16436
rect 19116 16396 19122 16408
rect 19153 16405 19165 16408
rect 19199 16405 19211 16439
rect 19153 16399 19211 16405
rect 1104 16346 24656 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 24656 16346
rect 1104 16272 24656 16294
rect 5169 16235 5227 16241
rect 5169 16201 5181 16235
rect 5215 16232 5227 16235
rect 5350 16232 5356 16244
rect 5215 16204 5356 16232
rect 5215 16201 5227 16204
rect 5169 16195 5227 16201
rect 5350 16192 5356 16204
rect 5408 16192 5414 16244
rect 20622 16192 20628 16244
rect 20680 16232 20686 16244
rect 20717 16235 20775 16241
rect 20717 16232 20729 16235
rect 20680 16204 20729 16232
rect 20680 16192 20686 16204
rect 20717 16201 20729 16204
rect 20763 16201 20775 16235
rect 20717 16195 20775 16201
rect 7101 16167 7159 16173
rect 7101 16133 7113 16167
rect 7147 16164 7159 16167
rect 7466 16164 7472 16176
rect 7147 16136 7472 16164
rect 7147 16133 7159 16136
rect 7101 16127 7159 16133
rect 7466 16124 7472 16136
rect 7524 16124 7530 16176
rect 9769 16099 9827 16105
rect 9769 16065 9781 16099
rect 9815 16096 9827 16099
rect 9950 16096 9956 16108
rect 9815 16068 9956 16096
rect 9815 16065 9827 16068
rect 9769 16059 9827 16065
rect 9950 16056 9956 16068
rect 10008 16056 10014 16108
rect 10778 16096 10784 16108
rect 10152 16068 10784 16096
rect 2498 16028 2504 16040
rect 2459 16000 2504 16028
rect 2498 15988 2504 16000
rect 2556 15988 2562 16040
rect 2777 16031 2835 16037
rect 2777 15997 2789 16031
rect 2823 16028 2835 16031
rect 3050 16028 3056 16040
rect 2823 16000 3056 16028
rect 2823 15997 2835 16000
rect 2777 15991 2835 15997
rect 3050 15988 3056 16000
rect 3108 16028 3114 16040
rect 4249 16031 4307 16037
rect 4249 16028 4261 16031
rect 3108 16000 4261 16028
rect 3108 15988 3114 16000
rect 4249 15997 4261 16000
rect 4295 15997 4307 16031
rect 4249 15991 4307 15997
rect 4985 16031 5043 16037
rect 4985 15997 4997 16031
rect 5031 16028 5043 16031
rect 7006 16028 7012 16040
rect 5031 16000 5065 16028
rect 6967 16000 7012 16028
rect 5031 15997 5043 16000
rect 4985 15991 5043 15997
rect 4798 15920 4804 15972
rect 4856 15960 4862 15972
rect 4893 15963 4951 15969
rect 4893 15960 4905 15963
rect 4856 15932 4905 15960
rect 4856 15920 4862 15932
rect 4893 15929 4905 15932
rect 4939 15960 4951 15963
rect 5000 15960 5028 15991
rect 7006 15988 7012 16000
rect 7064 15988 7070 16040
rect 7282 16028 7288 16040
rect 7243 16000 7288 16028
rect 7282 15988 7288 16000
rect 7340 15988 7346 16040
rect 10152 16037 10180 16068
rect 10778 16056 10784 16068
rect 10836 16056 10842 16108
rect 11146 16056 11152 16108
rect 11204 16096 11210 16108
rect 18046 16096 18052 16108
rect 11204 16068 12572 16096
rect 18007 16068 18052 16096
rect 11204 16056 11210 16068
rect 10137 16031 10195 16037
rect 10137 15997 10149 16031
rect 10183 15997 10195 16031
rect 10410 16028 10416 16040
rect 10371 16000 10416 16028
rect 10137 15991 10195 15997
rect 10410 15988 10416 16000
rect 10468 15988 10474 16040
rect 12544 16037 12572 16068
rect 18046 16056 18052 16068
rect 18104 16056 18110 16108
rect 20732 16096 20760 16195
rect 20901 16099 20959 16105
rect 20901 16096 20913 16099
rect 20732 16068 20913 16096
rect 20901 16065 20913 16068
rect 20947 16065 20959 16099
rect 20901 16059 20959 16065
rect 12437 16031 12495 16037
rect 12437 15997 12449 16031
rect 12483 15997 12495 16031
rect 12437 15991 12495 15997
rect 12529 16031 12587 16037
rect 12529 15997 12541 16031
rect 12575 16028 12587 16031
rect 15194 16028 15200 16040
rect 12575 16000 15200 16028
rect 12575 15997 12587 16000
rect 12529 15991 12587 15997
rect 5350 15960 5356 15972
rect 4939 15932 5356 15960
rect 4939 15929 4951 15932
rect 4893 15923 4951 15929
rect 5350 15920 5356 15932
rect 5408 15920 5414 15972
rect 7745 15963 7803 15969
rect 7745 15929 7757 15963
rect 7791 15960 7803 15963
rect 7926 15960 7932 15972
rect 7791 15932 7932 15960
rect 7791 15929 7803 15932
rect 7745 15923 7803 15929
rect 7926 15920 7932 15932
rect 7984 15920 7990 15972
rect 10686 15960 10692 15972
rect 10647 15932 10692 15960
rect 10686 15920 10692 15932
rect 10744 15920 10750 15972
rect 3878 15892 3884 15904
rect 3839 15864 3884 15892
rect 3878 15852 3884 15864
rect 3936 15852 3942 15904
rect 4525 15895 4583 15901
rect 4525 15861 4537 15895
rect 4571 15892 4583 15895
rect 4614 15892 4620 15904
rect 4571 15864 4620 15892
rect 4571 15861 4583 15864
rect 4525 15855 4583 15861
rect 4614 15852 4620 15864
rect 4672 15892 4678 15904
rect 4982 15892 4988 15904
rect 4672 15864 4988 15892
rect 4672 15852 4678 15864
rect 4982 15852 4988 15864
rect 5040 15852 5046 15904
rect 12452 15892 12480 15991
rect 15194 15988 15200 16000
rect 15252 15988 15258 16040
rect 18414 16028 18420 16040
rect 18375 16000 18420 16028
rect 18414 15988 18420 16000
rect 18472 15988 18478 16040
rect 18598 16028 18604 16040
rect 18511 16000 18604 16028
rect 18598 15988 18604 16000
rect 18656 15988 18662 16040
rect 18785 16031 18843 16037
rect 18785 15997 18797 16031
rect 18831 15997 18843 16031
rect 18966 16028 18972 16040
rect 18927 16000 18972 16028
rect 18785 15991 18843 15997
rect 12986 15960 12992 15972
rect 12947 15932 12992 15960
rect 12986 15920 12992 15932
rect 13044 15920 13050 15972
rect 17218 15920 17224 15972
rect 17276 15960 17282 15972
rect 18616 15960 18644 15988
rect 17276 15932 18644 15960
rect 18800 15960 18828 15991
rect 18966 15988 18972 16000
rect 19024 15988 19030 16040
rect 21082 16028 21088 16040
rect 21043 16000 21088 16028
rect 21082 15988 21088 16000
rect 21140 15988 21146 16040
rect 21542 16028 21548 16040
rect 21503 16000 21548 16028
rect 21542 15988 21548 16000
rect 21600 15988 21606 16040
rect 21637 16031 21695 16037
rect 21637 15997 21649 16031
rect 21683 15997 21695 16031
rect 21637 15991 21695 15997
rect 19705 15963 19763 15969
rect 19705 15960 19717 15963
rect 18800 15932 19717 15960
rect 17276 15920 17282 15932
rect 19705 15929 19717 15932
rect 19751 15960 19763 15963
rect 19886 15960 19892 15972
rect 19751 15932 19892 15960
rect 19751 15929 19763 15932
rect 19705 15923 19763 15929
rect 19886 15920 19892 15932
rect 19944 15920 19950 15972
rect 21100 15960 21128 15988
rect 21652 15960 21680 15991
rect 22186 15960 22192 15972
rect 21100 15932 21680 15960
rect 22147 15932 22192 15960
rect 22186 15920 22192 15932
rect 22244 15920 22250 15972
rect 13173 15895 13231 15901
rect 13173 15892 13185 15895
rect 12452 15864 13185 15892
rect 13173 15861 13185 15864
rect 13219 15892 13231 15895
rect 13262 15892 13268 15904
rect 13219 15864 13268 15892
rect 13219 15861 13231 15864
rect 13173 15855 13231 15861
rect 13262 15852 13268 15864
rect 13320 15852 13326 15904
rect 17862 15852 17868 15904
rect 17920 15892 17926 15904
rect 19429 15895 19487 15901
rect 19429 15892 19441 15895
rect 17920 15864 19441 15892
rect 17920 15852 17926 15864
rect 19429 15861 19441 15864
rect 19475 15861 19487 15895
rect 19429 15855 19487 15861
rect 1104 15802 24656 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 24656 15802
rect 1104 15728 24656 15750
rect 3694 15648 3700 15700
rect 3752 15688 3758 15700
rect 5445 15691 5503 15697
rect 5445 15688 5457 15691
rect 3752 15660 5457 15688
rect 3752 15648 3758 15660
rect 5445 15657 5457 15660
rect 5491 15657 5503 15691
rect 8665 15691 8723 15697
rect 8665 15688 8677 15691
rect 5445 15651 5503 15657
rect 7760 15660 8677 15688
rect 3786 15620 3792 15632
rect 3747 15592 3792 15620
rect 3786 15580 3792 15592
rect 3844 15580 3850 15632
rect 3804 15552 3832 15580
rect 4341 15555 4399 15561
rect 4341 15552 4353 15555
rect 3804 15524 4353 15552
rect 4341 15521 4353 15524
rect 4387 15521 4399 15555
rect 4341 15515 4399 15521
rect 5442 15512 5448 15564
rect 5500 15552 5506 15564
rect 6365 15555 6423 15561
rect 6365 15552 6377 15555
rect 5500 15524 6377 15552
rect 5500 15512 5506 15524
rect 6365 15521 6377 15524
rect 6411 15552 6423 15555
rect 6549 15555 6607 15561
rect 6549 15552 6561 15555
rect 6411 15524 6561 15552
rect 6411 15521 6423 15524
rect 6365 15515 6423 15521
rect 6549 15521 6561 15524
rect 6595 15521 6607 15555
rect 7760 15552 7788 15660
rect 8665 15657 8677 15660
rect 8711 15688 8723 15691
rect 10134 15688 10140 15700
rect 8711 15660 10140 15688
rect 8711 15657 8723 15660
rect 8665 15651 8723 15657
rect 10134 15648 10140 15660
rect 10192 15648 10198 15700
rect 13814 15648 13820 15700
rect 13872 15688 13878 15700
rect 13909 15691 13967 15697
rect 13909 15688 13921 15691
rect 13872 15660 13921 15688
rect 13872 15648 13878 15660
rect 13909 15657 13921 15660
rect 13955 15688 13967 15691
rect 14642 15688 14648 15700
rect 13955 15660 14648 15688
rect 13955 15657 13967 15660
rect 13909 15651 13967 15657
rect 14642 15648 14648 15660
rect 14700 15648 14706 15700
rect 15102 15688 15108 15700
rect 15015 15660 15108 15688
rect 15102 15648 15108 15660
rect 15160 15688 15166 15700
rect 16390 15688 16396 15700
rect 15160 15660 16396 15688
rect 15160 15648 15166 15660
rect 16390 15648 16396 15660
rect 16448 15648 16454 15700
rect 20990 15648 20996 15700
rect 21048 15688 21054 15700
rect 21729 15691 21787 15697
rect 21729 15688 21741 15691
rect 21048 15660 21741 15688
rect 21048 15648 21054 15660
rect 21729 15657 21741 15660
rect 21775 15657 21787 15691
rect 21729 15651 21787 15657
rect 7926 15620 7932 15632
rect 7887 15592 7932 15620
rect 7926 15580 7932 15592
rect 7984 15620 7990 15632
rect 10410 15620 10416 15632
rect 7984 15592 10416 15620
rect 7984 15580 7990 15592
rect 9968 15561 9996 15592
rect 10410 15580 10416 15592
rect 10468 15580 10474 15632
rect 10686 15580 10692 15632
rect 10744 15620 10750 15632
rect 12989 15623 13047 15629
rect 12989 15620 13001 15623
rect 10744 15592 13001 15620
rect 10744 15580 10750 15592
rect 12989 15589 13001 15592
rect 13035 15589 13047 15623
rect 18049 15623 18107 15629
rect 18049 15620 18061 15623
rect 12989 15583 13047 15589
rect 16040 15592 18061 15620
rect 8113 15555 8171 15561
rect 8113 15552 8125 15555
rect 7760 15524 8125 15552
rect 6549 15515 6607 15521
rect 8113 15521 8125 15524
rect 8159 15521 8171 15555
rect 8113 15515 8171 15521
rect 9953 15555 10011 15561
rect 9953 15521 9965 15555
rect 9999 15521 10011 15555
rect 9953 15515 10011 15521
rect 10045 15555 10103 15561
rect 10045 15521 10057 15555
rect 10091 15552 10103 15555
rect 11609 15555 11667 15561
rect 11609 15552 11621 15555
rect 10091 15524 11621 15552
rect 10091 15521 10103 15524
rect 10045 15515 10103 15521
rect 11609 15521 11621 15524
rect 11655 15521 11667 15555
rect 11609 15515 11667 15521
rect 11977 15555 12035 15561
rect 11977 15521 11989 15555
rect 12023 15552 12035 15555
rect 12802 15552 12808 15564
rect 12023 15524 12808 15552
rect 12023 15521 12035 15524
rect 11977 15515 12035 15521
rect 12802 15512 12808 15524
rect 12860 15512 12866 15564
rect 13538 15552 13544 15564
rect 12912 15524 13544 15552
rect 2498 15444 2504 15496
rect 2556 15484 2562 15496
rect 4065 15487 4123 15493
rect 4065 15484 4077 15487
rect 2556 15456 4077 15484
rect 2556 15444 2562 15456
rect 4065 15453 4077 15456
rect 4111 15484 4123 15487
rect 4522 15484 4528 15496
rect 4111 15456 4528 15484
rect 4111 15453 4123 15456
rect 4065 15447 4123 15453
rect 4522 15444 4528 15456
rect 4580 15444 4586 15496
rect 8386 15484 8392 15496
rect 8347 15456 8392 15484
rect 8386 15444 8392 15456
rect 8444 15444 8450 15496
rect 11330 15444 11336 15496
rect 11388 15484 11394 15496
rect 11517 15487 11575 15493
rect 11517 15484 11529 15487
rect 11388 15456 11529 15484
rect 11388 15444 11394 15456
rect 11517 15453 11529 15456
rect 11563 15453 11575 15487
rect 11517 15447 11575 15453
rect 12069 15487 12127 15493
rect 12069 15453 12081 15487
rect 12115 15484 12127 15487
rect 12526 15484 12532 15496
rect 12115 15456 12532 15484
rect 12115 15453 12127 15456
rect 12069 15447 12127 15453
rect 12526 15444 12532 15456
rect 12584 15484 12590 15496
rect 12912 15484 12940 15524
rect 13538 15512 13544 15524
rect 13596 15512 13602 15564
rect 16040 15561 16068 15592
rect 18049 15589 18061 15592
rect 18095 15589 18107 15623
rect 18049 15583 18107 15589
rect 16025 15555 16083 15561
rect 16025 15521 16037 15555
rect 16071 15521 16083 15555
rect 16025 15515 16083 15521
rect 16114 15512 16120 15564
rect 16172 15552 16178 15564
rect 16390 15552 16396 15564
rect 16172 15524 16217 15552
rect 16351 15524 16396 15552
rect 16172 15512 16178 15524
rect 16390 15512 16396 15524
rect 16448 15512 16454 15564
rect 16574 15552 16580 15564
rect 16535 15524 16580 15552
rect 16574 15512 16580 15524
rect 16632 15552 16638 15564
rect 16669 15555 16727 15561
rect 16669 15552 16681 15555
rect 16632 15524 16681 15552
rect 16632 15512 16638 15524
rect 16669 15521 16681 15524
rect 16715 15521 16727 15555
rect 16669 15515 16727 15521
rect 17957 15555 18015 15561
rect 17957 15521 17969 15555
rect 18003 15552 18015 15555
rect 19426 15552 19432 15564
rect 18003 15524 19432 15552
rect 18003 15521 18015 15524
rect 17957 15515 18015 15521
rect 19426 15512 19432 15524
rect 19484 15512 19490 15564
rect 19521 15555 19579 15561
rect 19521 15521 19533 15555
rect 19567 15552 19579 15555
rect 19886 15552 19892 15564
rect 19567 15524 19892 15552
rect 19567 15521 19579 15524
rect 19521 15515 19579 15521
rect 19886 15512 19892 15524
rect 19944 15512 19950 15564
rect 21744 15552 21772 15651
rect 23566 15620 23572 15632
rect 23527 15592 23572 15620
rect 23566 15580 23572 15592
rect 23624 15580 23630 15632
rect 21913 15555 21971 15561
rect 21913 15552 21925 15555
rect 21744 15524 21925 15552
rect 21913 15521 21925 15524
rect 21959 15521 21971 15555
rect 22186 15552 22192 15564
rect 22147 15524 22192 15552
rect 21913 15515 21971 15521
rect 22186 15512 22192 15524
rect 22244 15512 22250 15564
rect 12584 15456 12940 15484
rect 12584 15444 12590 15456
rect 12986 15444 12992 15496
rect 13044 15484 13050 15496
rect 13136 15487 13194 15493
rect 13136 15484 13148 15487
rect 13044 15456 13148 15484
rect 13044 15444 13050 15456
rect 13136 15453 13148 15456
rect 13182 15453 13194 15487
rect 13354 15484 13360 15496
rect 13315 15456 13360 15484
rect 13136 15447 13194 15453
rect 13354 15444 13360 15456
rect 13412 15444 13418 15496
rect 13630 15444 13636 15496
rect 13688 15484 13694 15496
rect 15381 15487 15439 15493
rect 15381 15484 15393 15487
rect 13688 15456 15393 15484
rect 13688 15444 13694 15456
rect 15381 15453 15393 15456
rect 15427 15453 15439 15487
rect 15381 15447 15439 15453
rect 11054 15416 11060 15428
rect 11015 15388 11060 15416
rect 11054 15376 11060 15388
rect 11112 15376 11118 15428
rect 11146 15376 11152 15428
rect 11204 15416 11210 15428
rect 13449 15419 13507 15425
rect 13449 15416 13461 15419
rect 11204 15388 13461 15416
rect 11204 15376 11210 15388
rect 13449 15385 13461 15388
rect 13495 15385 13507 15419
rect 13449 15379 13507 15385
rect 5442 15308 5448 15360
rect 5500 15348 5506 15360
rect 5813 15351 5871 15357
rect 5813 15348 5825 15351
rect 5500 15320 5825 15348
rect 5500 15308 5506 15320
rect 5813 15317 5825 15320
rect 5859 15317 5871 15351
rect 5813 15311 5871 15317
rect 6733 15351 6791 15357
rect 6733 15317 6745 15351
rect 6779 15348 6791 15351
rect 7098 15348 7104 15360
rect 6779 15320 7104 15348
rect 6779 15317 6791 15320
rect 6733 15311 6791 15317
rect 7098 15308 7104 15320
rect 7156 15308 7162 15360
rect 13265 15351 13323 15357
rect 13265 15317 13277 15351
rect 13311 15348 13323 15351
rect 13814 15348 13820 15360
rect 13311 15320 13820 15348
rect 13311 15317 13323 15320
rect 13265 15311 13323 15317
rect 13814 15308 13820 15320
rect 13872 15308 13878 15360
rect 19426 15308 19432 15360
rect 19484 15348 19490 15360
rect 19904 15357 19932 15512
rect 19613 15351 19671 15357
rect 19613 15348 19625 15351
rect 19484 15320 19625 15348
rect 19484 15308 19490 15320
rect 19613 15317 19625 15320
rect 19659 15317 19671 15351
rect 19613 15311 19671 15317
rect 19889 15351 19947 15357
rect 19889 15317 19901 15351
rect 19935 15348 19947 15351
rect 21910 15348 21916 15360
rect 19935 15320 21916 15348
rect 19935 15317 19947 15320
rect 19889 15311 19947 15317
rect 21910 15308 21916 15320
rect 21968 15308 21974 15360
rect 1104 15258 24656 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 24656 15258
rect 1104 15184 24656 15206
rect 5353 15147 5411 15153
rect 5353 15113 5365 15147
rect 5399 15144 5411 15147
rect 7006 15144 7012 15156
rect 5399 15116 7012 15144
rect 5399 15113 5411 15116
rect 5353 15107 5411 15113
rect 7006 15104 7012 15116
rect 7064 15104 7070 15156
rect 7558 15104 7564 15156
rect 7616 15144 7622 15156
rect 8389 15147 8447 15153
rect 8389 15144 8401 15147
rect 7616 15116 8401 15144
rect 7616 15104 7622 15116
rect 8389 15113 8401 15116
rect 8435 15113 8447 15147
rect 8389 15107 8447 15113
rect 8662 15104 8668 15156
rect 8720 15144 8726 15156
rect 11149 15147 11207 15153
rect 8720 15116 11100 15144
rect 8720 15104 8726 15116
rect 4341 15079 4399 15085
rect 4341 15045 4353 15079
rect 4387 15076 4399 15079
rect 5534 15076 5540 15088
rect 4387 15048 5540 15076
rect 4387 15045 4399 15048
rect 4341 15039 4399 15045
rect 2498 15008 2504 15020
rect 2459 14980 2504 15008
rect 2498 14968 2504 14980
rect 2556 14968 2562 15020
rect 2777 15011 2835 15017
rect 2777 14977 2789 15011
rect 2823 15008 2835 15011
rect 4356 15008 4384 15039
rect 5534 15036 5540 15048
rect 5592 15036 5598 15088
rect 11072 15076 11100 15116
rect 11149 15113 11161 15147
rect 11195 15144 11207 15147
rect 11238 15144 11244 15156
rect 11195 15116 11244 15144
rect 11195 15113 11207 15116
rect 11149 15107 11207 15113
rect 11238 15104 11244 15116
rect 11296 15104 11302 15156
rect 20346 15144 20352 15156
rect 11348 15116 20352 15144
rect 11348 15076 11376 15116
rect 20346 15104 20352 15116
rect 20404 15104 20410 15156
rect 21910 15144 21916 15156
rect 21871 15116 21916 15144
rect 21910 15104 21916 15116
rect 21968 15104 21974 15156
rect 11072 15048 11376 15076
rect 13078 15036 13084 15088
rect 13136 15076 13142 15088
rect 13265 15079 13323 15085
rect 13265 15076 13277 15079
rect 13136 15048 13277 15076
rect 13136 15036 13142 15048
rect 13265 15045 13277 15048
rect 13311 15076 13323 15079
rect 15746 15076 15752 15088
rect 13311 15048 15752 15076
rect 13311 15045 13323 15048
rect 13265 15039 13323 15045
rect 15746 15036 15752 15048
rect 15804 15036 15810 15088
rect 2823 14980 4384 15008
rect 4525 15011 4583 15017
rect 2823 14977 2835 14980
rect 2777 14971 2835 14977
rect 4525 14977 4537 15011
rect 4571 15008 4583 15011
rect 4614 15008 4620 15020
rect 4571 14980 4620 15008
rect 4571 14977 4583 14980
rect 4525 14971 4583 14977
rect 4614 14968 4620 14980
rect 4672 15008 4678 15020
rect 5442 15008 5448 15020
rect 4672 14980 5448 15008
rect 4672 14968 4678 14980
rect 5442 14968 5448 14980
rect 5500 14968 5506 15020
rect 11882 15008 11888 15020
rect 8220 14980 11888 15008
rect 4982 14900 4988 14952
rect 5040 14940 5046 14952
rect 5169 14943 5227 14949
rect 5169 14940 5181 14943
rect 5040 14912 5181 14940
rect 5040 14900 5046 14912
rect 5169 14909 5181 14912
rect 5215 14909 5227 14943
rect 5169 14903 5227 14909
rect 7653 14943 7711 14949
rect 7653 14909 7665 14943
rect 7699 14940 7711 14943
rect 7926 14940 7932 14952
rect 7699 14912 7932 14940
rect 7699 14909 7711 14912
rect 7653 14903 7711 14909
rect 7926 14900 7932 14912
rect 7984 14900 7990 14952
rect 8220 14949 8248 14980
rect 11882 14968 11888 14980
rect 11940 14968 11946 15020
rect 12618 14968 12624 15020
rect 12676 15008 12682 15020
rect 13170 15008 13176 15020
rect 12676 14980 13176 15008
rect 12676 14968 12682 14980
rect 13170 14968 13176 14980
rect 13228 15008 13234 15020
rect 14737 15011 14795 15017
rect 14737 15008 14749 15011
rect 13228 14980 14749 15008
rect 13228 14968 13234 14980
rect 14737 14977 14749 14980
rect 14783 15008 14795 15011
rect 14921 15011 14979 15017
rect 14921 15008 14933 15011
rect 14783 14980 14933 15008
rect 14783 14977 14795 14980
rect 14737 14971 14795 14977
rect 14921 14977 14933 14980
rect 14967 14977 14979 15011
rect 14921 14971 14979 14977
rect 20257 15011 20315 15017
rect 20257 14977 20269 15011
rect 20303 15008 20315 15011
rect 20349 15011 20407 15017
rect 20349 15008 20361 15011
rect 20303 14980 20361 15008
rect 20303 14977 20315 14980
rect 20257 14971 20315 14977
rect 20349 14977 20361 14980
rect 20395 15008 20407 15011
rect 20990 15008 20996 15020
rect 20395 14980 20996 15008
rect 20395 14977 20407 14980
rect 20349 14971 20407 14977
rect 8205 14943 8263 14949
rect 8205 14909 8217 14943
rect 8251 14909 8263 14943
rect 10410 14940 10416 14952
rect 10371 14912 10416 14940
rect 8205 14903 8263 14909
rect 10410 14900 10416 14912
rect 10468 14900 10474 14952
rect 10597 14943 10655 14949
rect 10597 14909 10609 14943
rect 10643 14940 10655 14943
rect 11238 14940 11244 14952
rect 10643 14912 11244 14940
rect 10643 14909 10655 14912
rect 10597 14903 10655 14909
rect 11238 14900 11244 14912
rect 11296 14900 11302 14952
rect 13449 14943 13507 14949
rect 13449 14909 13461 14943
rect 13495 14909 13507 14943
rect 13449 14903 13507 14909
rect 8113 14875 8171 14881
rect 8113 14841 8125 14875
rect 8159 14872 8171 14875
rect 8386 14872 8392 14884
rect 8159 14844 8392 14872
rect 8159 14841 8171 14844
rect 8113 14835 8171 14841
rect 8386 14832 8392 14844
rect 8444 14832 8450 14884
rect 13464 14872 13492 14903
rect 13538 14900 13544 14952
rect 13596 14940 13602 14952
rect 15105 14943 15163 14949
rect 13596 14912 13641 14940
rect 13596 14900 13602 14912
rect 15105 14909 15117 14943
rect 15151 14940 15163 14943
rect 15194 14940 15200 14952
rect 15151 14912 15200 14940
rect 15151 14909 15163 14912
rect 15105 14903 15163 14909
rect 15194 14900 15200 14912
rect 15252 14900 15258 14952
rect 15286 14900 15292 14952
rect 15344 14940 15350 14952
rect 15565 14943 15623 14949
rect 15565 14940 15577 14943
rect 15344 14912 15577 14940
rect 15344 14900 15350 14912
rect 15565 14909 15577 14912
rect 15611 14909 15623 14943
rect 15565 14903 15623 14909
rect 15657 14943 15715 14949
rect 15657 14909 15669 14943
rect 15703 14909 15715 14943
rect 15657 14903 15715 14909
rect 14918 14872 14924 14884
rect 13464 14844 14924 14872
rect 14918 14832 14924 14844
rect 14976 14832 14982 14884
rect 15212 14872 15240 14900
rect 15672 14872 15700 14903
rect 15746 14900 15752 14952
rect 15804 14940 15810 14952
rect 20272 14940 20300 14971
rect 20990 14968 20996 14980
rect 21048 14968 21054 15020
rect 20622 14940 20628 14952
rect 15804 14912 20300 14940
rect 20583 14912 20628 14940
rect 15804 14900 15810 14912
rect 20622 14900 20628 14912
rect 20680 14900 20686 14952
rect 15212 14844 15700 14872
rect 3878 14804 3884 14816
rect 3839 14776 3884 14804
rect 3878 14764 3884 14776
rect 3936 14764 3942 14816
rect 4982 14804 4988 14816
rect 4943 14776 4988 14804
rect 4982 14764 4988 14776
rect 5040 14764 5046 14816
rect 7098 14764 7104 14816
rect 7156 14804 7162 14816
rect 7653 14807 7711 14813
rect 7653 14804 7665 14807
rect 7156 14776 7665 14804
rect 7156 14764 7162 14776
rect 7653 14773 7665 14776
rect 7699 14804 7711 14807
rect 7745 14807 7803 14813
rect 7745 14804 7757 14807
rect 7699 14776 7757 14804
rect 7699 14773 7711 14776
rect 7653 14767 7711 14773
rect 7745 14773 7757 14776
rect 7791 14773 7803 14807
rect 7745 14767 7803 14773
rect 10594 14764 10600 14816
rect 10652 14804 10658 14816
rect 10689 14807 10747 14813
rect 10689 14804 10701 14807
rect 10652 14776 10701 14804
rect 10652 14764 10658 14776
rect 10689 14773 10701 14776
rect 10735 14773 10747 14807
rect 10689 14767 10747 14773
rect 13725 14807 13783 14813
rect 13725 14773 13737 14807
rect 13771 14804 13783 14807
rect 13906 14804 13912 14816
rect 13771 14776 13912 14804
rect 13771 14773 13783 14776
rect 13725 14767 13783 14773
rect 13906 14764 13912 14776
rect 13964 14804 13970 14816
rect 14734 14804 14740 14816
rect 13964 14776 14740 14804
rect 13964 14764 13970 14776
rect 14734 14764 14740 14776
rect 14792 14764 14798 14816
rect 16114 14804 16120 14816
rect 16075 14776 16120 14804
rect 16114 14764 16120 14776
rect 16172 14764 16178 14816
rect 1104 14714 24656 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 24656 14714
rect 1104 14640 24656 14662
rect 5537 14603 5595 14609
rect 5537 14569 5549 14603
rect 5583 14600 5595 14603
rect 6730 14600 6736 14612
rect 5583 14572 6736 14600
rect 5583 14569 5595 14572
rect 5537 14563 5595 14569
rect 6730 14560 6736 14572
rect 6788 14560 6794 14612
rect 7926 14560 7932 14612
rect 7984 14600 7990 14612
rect 10229 14603 10287 14609
rect 10229 14600 10241 14603
rect 7984 14572 10241 14600
rect 7984 14560 7990 14572
rect 10229 14569 10241 14572
rect 10275 14569 10287 14603
rect 10229 14563 10287 14569
rect 14277 14603 14335 14609
rect 14277 14569 14289 14603
rect 14323 14600 14335 14603
rect 15286 14600 15292 14612
rect 14323 14572 15292 14600
rect 14323 14569 14335 14572
rect 14277 14563 14335 14569
rect 5350 14424 5356 14476
rect 5408 14464 5414 14476
rect 5445 14467 5503 14473
rect 5445 14464 5457 14467
rect 5408 14436 5457 14464
rect 5408 14424 5414 14436
rect 5445 14433 5457 14436
rect 5491 14433 5503 14467
rect 5445 14427 5503 14433
rect 8573 14467 8631 14473
rect 8573 14433 8585 14467
rect 8619 14464 8631 14467
rect 10244 14464 10272 14563
rect 15286 14560 15292 14572
rect 15344 14560 15350 14612
rect 15746 14600 15752 14612
rect 15707 14572 15752 14600
rect 15746 14560 15752 14572
rect 15804 14560 15810 14612
rect 16482 14600 16488 14612
rect 15948 14572 16488 14600
rect 10594 14532 10600 14544
rect 10555 14504 10600 14532
rect 10594 14492 10600 14504
rect 10652 14492 10658 14544
rect 12989 14535 13047 14541
rect 12989 14501 13001 14535
rect 13035 14532 13047 14535
rect 13354 14532 13360 14544
rect 13035 14504 13360 14532
rect 13035 14501 13047 14504
rect 12989 14495 13047 14501
rect 13354 14492 13360 14504
rect 13412 14492 13418 14544
rect 14553 14535 14611 14541
rect 14553 14501 14565 14535
rect 14599 14532 14611 14535
rect 15948 14532 15976 14572
rect 16482 14560 16488 14572
rect 16540 14600 16546 14612
rect 17221 14603 17279 14609
rect 17221 14600 17233 14603
rect 16540 14572 17233 14600
rect 16540 14560 16546 14572
rect 17221 14569 17233 14572
rect 17267 14569 17279 14603
rect 17221 14563 17279 14569
rect 17770 14560 17776 14612
rect 17828 14600 17834 14612
rect 18325 14603 18383 14609
rect 18325 14600 18337 14603
rect 17828 14572 18337 14600
rect 17828 14560 17834 14572
rect 18325 14569 18337 14572
rect 18371 14600 18383 14603
rect 18417 14603 18475 14609
rect 18417 14600 18429 14603
rect 18371 14572 18429 14600
rect 18371 14569 18383 14572
rect 18325 14563 18383 14569
rect 18417 14569 18429 14572
rect 18463 14569 18475 14603
rect 18417 14563 18475 14569
rect 14599 14504 15976 14532
rect 19889 14535 19947 14541
rect 14599 14501 14611 14504
rect 14553 14495 14611 14501
rect 19889 14501 19901 14535
rect 19935 14532 19947 14535
rect 20622 14532 20628 14544
rect 19935 14504 20628 14532
rect 19935 14501 19947 14504
rect 19889 14495 19947 14501
rect 10413 14467 10471 14473
rect 10413 14464 10425 14467
rect 8619 14436 8984 14464
rect 10244 14436 10425 14464
rect 8619 14433 8631 14436
rect 8573 14427 8631 14433
rect 5350 14260 5356 14272
rect 5311 14232 5356 14260
rect 5350 14220 5356 14232
rect 5408 14220 5414 14272
rect 8662 14260 8668 14272
rect 8623 14232 8668 14260
rect 8662 14220 8668 14232
rect 8720 14220 8726 14272
rect 8956 14269 8984 14436
rect 10413 14433 10425 14436
rect 10459 14433 10471 14467
rect 10413 14427 10471 14433
rect 10689 14467 10747 14473
rect 10689 14433 10701 14467
rect 10735 14464 10747 14467
rect 11146 14464 11152 14476
rect 10735 14436 11152 14464
rect 10735 14433 10747 14436
rect 10689 14427 10747 14433
rect 11146 14424 11152 14436
rect 11204 14424 11210 14476
rect 12526 14464 12532 14476
rect 12487 14436 12532 14464
rect 12526 14424 12532 14436
rect 12584 14424 12590 14476
rect 14185 14467 14243 14473
rect 14185 14433 14197 14467
rect 14231 14464 14243 14467
rect 14568 14464 14596 14495
rect 20622 14492 20628 14504
rect 20680 14492 20686 14544
rect 14231 14436 14596 14464
rect 14231 14433 14243 14436
rect 14185 14427 14243 14433
rect 15194 14424 15200 14476
rect 15252 14464 15258 14476
rect 16114 14464 16120 14476
rect 15252 14436 15976 14464
rect 16075 14436 16120 14464
rect 15252 14424 15258 14436
rect 12437 14399 12495 14405
rect 12437 14365 12449 14399
rect 12483 14396 12495 14399
rect 13630 14396 13636 14408
rect 12483 14368 13636 14396
rect 12483 14365 12495 14368
rect 12437 14359 12495 14365
rect 13630 14356 13636 14368
rect 13688 14356 13694 14408
rect 15746 14356 15752 14408
rect 15804 14396 15810 14408
rect 15841 14399 15899 14405
rect 15841 14396 15853 14399
rect 15804 14368 15853 14396
rect 15804 14356 15810 14368
rect 15841 14365 15853 14368
rect 15887 14365 15899 14399
rect 15948 14396 15976 14436
rect 16114 14424 16120 14436
rect 16172 14424 16178 14476
rect 18785 14467 18843 14473
rect 18785 14464 18797 14467
rect 16224 14436 18797 14464
rect 16224 14396 16252 14436
rect 18785 14433 18797 14436
rect 18831 14464 18843 14467
rect 19337 14467 19395 14473
rect 19337 14464 19349 14467
rect 18831 14436 19349 14464
rect 18831 14433 18843 14436
rect 18785 14427 18843 14433
rect 19337 14433 19349 14436
rect 19383 14433 19395 14467
rect 19337 14427 19395 14433
rect 19426 14424 19432 14476
rect 19484 14464 19490 14476
rect 19521 14467 19579 14473
rect 19521 14464 19533 14467
rect 19484 14436 19533 14464
rect 19484 14424 19490 14436
rect 19521 14433 19533 14436
rect 19567 14433 19579 14467
rect 19521 14427 19579 14433
rect 22741 14467 22799 14473
rect 22741 14433 22753 14467
rect 22787 14464 22799 14467
rect 23474 14464 23480 14476
rect 22787 14436 23480 14464
rect 22787 14433 22799 14436
rect 22741 14427 22799 14433
rect 23474 14424 23480 14436
rect 23532 14424 23538 14476
rect 15948 14368 16252 14396
rect 18325 14399 18383 14405
rect 15841 14359 15899 14365
rect 18325 14365 18337 14399
rect 18371 14396 18383 14399
rect 18601 14399 18659 14405
rect 18601 14396 18613 14399
rect 18371 14368 18613 14396
rect 18371 14365 18383 14368
rect 18325 14359 18383 14365
rect 18601 14365 18613 14368
rect 18647 14365 18659 14399
rect 18601 14359 18659 14365
rect 10318 14288 10324 14340
rect 10376 14328 10382 14340
rect 10376 14300 10916 14328
rect 10376 14288 10382 14300
rect 8941 14263 8999 14269
rect 8941 14229 8953 14263
rect 8987 14260 8999 14263
rect 9582 14260 9588 14272
rect 8987 14232 9588 14260
rect 8987 14229 8999 14232
rect 8941 14223 8999 14229
rect 9582 14220 9588 14232
rect 9640 14220 9646 14272
rect 10888 14269 10916 14300
rect 10873 14263 10931 14269
rect 10873 14229 10885 14263
rect 10919 14229 10931 14263
rect 10873 14223 10931 14229
rect 15470 14220 15476 14272
rect 15528 14260 15534 14272
rect 18782 14260 18788 14272
rect 15528 14232 18788 14260
rect 15528 14220 15534 14232
rect 18782 14220 18788 14232
rect 18840 14220 18846 14272
rect 21818 14220 21824 14272
rect 21876 14260 21882 14272
rect 22833 14263 22891 14269
rect 22833 14260 22845 14263
rect 21876 14232 22845 14260
rect 21876 14220 21882 14232
rect 22833 14229 22845 14232
rect 22879 14229 22891 14263
rect 22833 14223 22891 14229
rect 1104 14170 24656 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 24656 14170
rect 1104 14096 24656 14118
rect 4341 14059 4399 14065
rect 4341 14025 4353 14059
rect 4387 14056 4399 14059
rect 4706 14056 4712 14068
rect 4387 14028 4712 14056
rect 4387 14025 4399 14028
rect 4341 14019 4399 14025
rect 2777 13923 2835 13929
rect 2777 13889 2789 13923
rect 2823 13920 2835 13923
rect 4356 13920 4384 14019
rect 4706 14016 4712 14028
rect 4764 14016 4770 14068
rect 5442 14016 5448 14068
rect 5500 14056 5506 14068
rect 7929 14059 7987 14065
rect 7929 14056 7941 14059
rect 5500 14028 7941 14056
rect 5500 14016 5506 14028
rect 7929 14025 7941 14028
rect 7975 14056 7987 14059
rect 9582 14056 9588 14068
rect 7975 14028 8984 14056
rect 9495 14028 9588 14056
rect 7975 14025 7987 14028
rect 7929 14019 7987 14025
rect 8956 13988 8984 14028
rect 9582 14016 9588 14028
rect 9640 14056 9646 14068
rect 10870 14056 10876 14068
rect 9640 14028 10876 14056
rect 9640 14016 9646 14028
rect 10870 14016 10876 14028
rect 10928 14016 10934 14068
rect 10962 14016 10968 14068
rect 11020 14056 11026 14068
rect 13078 14056 13084 14068
rect 11020 14028 13084 14056
rect 11020 14016 11026 14028
rect 13078 14016 13084 14028
rect 13136 14016 13142 14068
rect 14918 14016 14924 14068
rect 14976 14056 14982 14068
rect 15105 14059 15163 14065
rect 15105 14056 15117 14059
rect 14976 14028 15117 14056
rect 14976 14016 14982 14028
rect 15105 14025 15117 14028
rect 15151 14025 15163 14059
rect 15105 14019 15163 14025
rect 18417 14059 18475 14065
rect 18417 14025 18429 14059
rect 18463 14056 18475 14059
rect 19150 14056 19156 14068
rect 18463 14028 19156 14056
rect 18463 14025 18475 14028
rect 18417 14019 18475 14025
rect 9861 13991 9919 13997
rect 9861 13988 9873 13991
rect 8956 13960 9873 13988
rect 9861 13957 9873 13960
rect 9907 13988 9919 13991
rect 10594 13988 10600 14000
rect 9907 13960 10600 13988
rect 9907 13957 9919 13960
rect 9861 13951 9919 13957
rect 10594 13948 10600 13960
rect 10652 13948 10658 14000
rect 10689 13991 10747 13997
rect 10689 13957 10701 13991
rect 10735 13988 10747 13991
rect 15194 13988 15200 14000
rect 10735 13960 15200 13988
rect 10735 13957 10747 13960
rect 10689 13951 10747 13957
rect 15194 13948 15200 13960
rect 15252 13988 15258 14000
rect 18322 13988 18328 14000
rect 15252 13960 15608 13988
rect 15252 13948 15258 13960
rect 6086 13920 6092 13932
rect 2823 13892 4384 13920
rect 5736 13892 6092 13920
rect 2823 13889 2835 13892
rect 2777 13883 2835 13889
rect 2501 13855 2559 13861
rect 2501 13821 2513 13855
rect 2547 13852 2559 13855
rect 4433 13855 4491 13861
rect 4433 13852 4445 13855
rect 2547 13824 4445 13852
rect 2547 13821 2559 13824
rect 2501 13815 2559 13821
rect 4433 13821 4445 13824
rect 4479 13852 4491 13855
rect 4522 13852 4528 13864
rect 4479 13824 4528 13852
rect 4479 13821 4491 13824
rect 4433 13815 4491 13821
rect 4522 13812 4528 13824
rect 4580 13812 4586 13864
rect 5736 13861 5764 13892
rect 6086 13880 6092 13892
rect 6144 13920 6150 13932
rect 13262 13920 13268 13932
rect 6144 13892 13268 13920
rect 6144 13880 6150 13892
rect 13262 13880 13268 13892
rect 13320 13880 13326 13932
rect 15013 13923 15071 13929
rect 15013 13889 15025 13923
rect 15059 13920 15071 13923
rect 15470 13920 15476 13932
rect 15059 13892 15476 13920
rect 15059 13889 15071 13892
rect 15013 13883 15071 13889
rect 5721 13855 5779 13861
rect 5721 13821 5733 13855
rect 5767 13821 5779 13855
rect 5721 13815 5779 13821
rect 7929 13855 7987 13861
rect 7929 13821 7941 13855
rect 7975 13852 7987 13855
rect 8021 13855 8079 13861
rect 8021 13852 8033 13855
rect 7975 13824 8033 13852
rect 7975 13821 7987 13824
rect 7929 13815 7987 13821
rect 8021 13821 8033 13824
rect 8067 13821 8079 13855
rect 8294 13852 8300 13864
rect 8255 13824 8300 13852
rect 8021 13815 8079 13821
rect 8294 13812 8300 13824
rect 8352 13812 8358 13864
rect 9674 13812 9680 13864
rect 9732 13852 9738 13864
rect 10505 13855 10563 13861
rect 10505 13852 10517 13855
rect 9732 13824 10517 13852
rect 9732 13812 9738 13824
rect 10505 13821 10517 13824
rect 10551 13821 10563 13855
rect 10505 13815 10563 13821
rect 12158 13812 12164 13864
rect 12216 13852 12222 13864
rect 15028 13852 15056 13883
rect 15470 13880 15476 13892
rect 15528 13880 15534 13932
rect 15580 13861 15608 13960
rect 15672 13960 18328 13988
rect 12216 13824 15056 13852
rect 15289 13855 15347 13861
rect 12216 13812 12222 13824
rect 15289 13821 15301 13855
rect 15335 13852 15347 13855
rect 15565 13855 15623 13861
rect 15335 13824 15516 13852
rect 15335 13821 15347 13824
rect 15289 13815 15347 13821
rect 5534 13744 5540 13796
rect 5592 13784 5598 13796
rect 6638 13784 6644 13796
rect 5592 13756 6644 13784
rect 5592 13744 5598 13756
rect 6638 13744 6644 13756
rect 6696 13744 6702 13796
rect 15488 13784 15516 13824
rect 15565 13821 15577 13855
rect 15611 13821 15623 13855
rect 15565 13815 15623 13821
rect 15672 13784 15700 13960
rect 18322 13948 18328 13960
rect 18380 13948 18386 14000
rect 18141 13923 18199 13929
rect 18141 13920 18153 13923
rect 16868 13892 18153 13920
rect 15746 13812 15752 13864
rect 15804 13852 15810 13864
rect 16117 13855 16175 13861
rect 16117 13852 16129 13855
rect 15804 13824 16129 13852
rect 15804 13812 15810 13824
rect 16117 13821 16129 13824
rect 16163 13821 16175 13855
rect 16117 13815 16175 13821
rect 16301 13855 16359 13861
rect 16301 13821 16313 13855
rect 16347 13852 16359 13855
rect 16868 13852 16896 13892
rect 18141 13889 18153 13892
rect 18187 13889 18199 13923
rect 18141 13883 18199 13889
rect 16347 13824 16896 13852
rect 18049 13855 18107 13861
rect 16347 13821 16359 13824
rect 16301 13815 16359 13821
rect 18049 13821 18061 13855
rect 18095 13852 18107 13855
rect 18230 13852 18236 13864
rect 18095 13824 18236 13852
rect 18095 13821 18107 13824
rect 18049 13815 18107 13821
rect 18230 13812 18236 13824
rect 18288 13852 18294 13864
rect 18432 13852 18460 14019
rect 19150 14016 19156 14028
rect 19208 14016 19214 14068
rect 19334 14016 19340 14068
rect 19392 14056 19398 14068
rect 19429 14059 19487 14065
rect 19429 14056 19441 14059
rect 19392 14028 19441 14056
rect 19392 14016 19398 14028
rect 19429 14025 19441 14028
rect 19475 14025 19487 14059
rect 20714 14056 20720 14068
rect 20675 14028 20720 14056
rect 19429 14019 19487 14025
rect 18288 13824 18460 13852
rect 19444 13852 19472 14019
rect 20714 14016 20720 14028
rect 20772 14016 20778 14068
rect 19797 13991 19855 13997
rect 19797 13957 19809 13991
rect 19843 13957 19855 13991
rect 19797 13951 19855 13957
rect 19613 13855 19671 13861
rect 19613 13852 19625 13855
rect 19444 13824 19625 13852
rect 18288 13812 18294 13824
rect 19613 13821 19625 13824
rect 19659 13821 19671 13855
rect 19812 13852 19840 13951
rect 20732 13920 20760 14016
rect 20901 13923 20959 13929
rect 20901 13920 20913 13923
rect 20732 13892 20913 13920
rect 20901 13889 20913 13892
rect 20947 13889 20959 13923
rect 20901 13883 20959 13889
rect 20806 13852 20812 13864
rect 19812 13824 20812 13852
rect 19613 13815 19671 13821
rect 20806 13812 20812 13824
rect 20864 13852 20870 13864
rect 21085 13855 21143 13861
rect 21085 13852 21097 13855
rect 20864 13824 21097 13852
rect 20864 13812 20870 13824
rect 21085 13821 21097 13824
rect 21131 13821 21143 13855
rect 21085 13815 21143 13821
rect 21637 13855 21695 13861
rect 21637 13821 21649 13855
rect 21683 13821 21695 13855
rect 21818 13852 21824 13864
rect 21779 13824 21824 13852
rect 21637 13815 21695 13821
rect 16666 13784 16672 13796
rect 15488 13756 15700 13784
rect 16627 13756 16672 13784
rect 16666 13744 16672 13756
rect 16724 13744 16730 13796
rect 21100 13784 21128 13815
rect 21652 13784 21680 13815
rect 21818 13812 21824 13824
rect 21876 13812 21882 13864
rect 22186 13784 22192 13796
rect 21100 13756 21680 13784
rect 22147 13756 22192 13784
rect 22186 13744 22192 13756
rect 22244 13744 22250 13796
rect 3878 13716 3884 13728
rect 3839 13688 3884 13716
rect 3878 13676 3884 13688
rect 3936 13676 3942 13728
rect 5810 13716 5816 13728
rect 5771 13688 5816 13716
rect 5810 13676 5816 13688
rect 5868 13676 5874 13728
rect 1104 13626 24656 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 24656 13626
rect 1104 13552 24656 13574
rect 6086 13512 6092 13524
rect 6047 13484 6092 13512
rect 6086 13472 6092 13484
rect 6144 13472 6150 13524
rect 7282 13512 7288 13524
rect 7195 13484 7288 13512
rect 7282 13472 7288 13484
rect 7340 13512 7346 13524
rect 7834 13512 7840 13524
rect 7340 13484 7840 13512
rect 7340 13472 7346 13484
rect 7834 13472 7840 13484
rect 7892 13472 7898 13524
rect 8294 13472 8300 13524
rect 8352 13512 8358 13524
rect 8573 13515 8631 13521
rect 8573 13512 8585 13515
rect 8352 13484 8585 13512
rect 8352 13472 8358 13484
rect 8573 13481 8585 13484
rect 8619 13481 8631 13515
rect 12710 13512 12716 13524
rect 8573 13475 8631 13481
rect 11532 13484 12716 13512
rect 11333 13447 11391 13453
rect 11333 13444 11345 13447
rect 7484 13416 11345 13444
rect 4062 13336 4068 13388
rect 4120 13376 4126 13388
rect 7484 13376 7512 13416
rect 11333 13413 11345 13416
rect 11379 13444 11391 13447
rect 11532 13444 11560 13484
rect 12710 13472 12716 13484
rect 12768 13472 12774 13524
rect 14093 13515 14151 13521
rect 14093 13481 14105 13515
rect 14139 13512 14151 13515
rect 15102 13512 15108 13524
rect 14139 13484 15108 13512
rect 14139 13481 14151 13484
rect 14093 13475 14151 13481
rect 13817 13447 13875 13453
rect 13817 13444 13829 13447
rect 11379 13416 11560 13444
rect 11379 13413 11391 13416
rect 11333 13407 11391 13413
rect 4120 13348 7512 13376
rect 7561 13379 7619 13385
rect 4120 13336 4126 13348
rect 7561 13345 7573 13379
rect 7607 13376 7619 13379
rect 8113 13379 8171 13385
rect 8113 13376 8125 13379
rect 7607 13348 8125 13376
rect 7607 13345 7619 13348
rect 7561 13339 7619 13345
rect 8113 13345 8125 13348
rect 8159 13345 8171 13379
rect 8113 13339 8171 13345
rect 8297 13379 8355 13385
rect 8297 13345 8309 13379
rect 8343 13376 8355 13379
rect 8662 13376 8668 13388
rect 8343 13348 8668 13376
rect 8343 13345 8355 13348
rect 8297 13339 8355 13345
rect 4522 13308 4528 13320
rect 4483 13280 4528 13308
rect 4522 13268 4528 13280
rect 4580 13268 4586 13320
rect 4801 13311 4859 13317
rect 4801 13277 4813 13311
rect 4847 13308 4859 13311
rect 5718 13308 5724 13320
rect 4847 13280 5724 13308
rect 4847 13277 4859 13280
rect 4801 13271 4859 13277
rect 5718 13268 5724 13280
rect 5776 13268 5782 13320
rect 7282 13268 7288 13320
rect 7340 13308 7346 13320
rect 7377 13311 7435 13317
rect 7377 13308 7389 13311
rect 7340 13280 7389 13308
rect 7340 13268 7346 13280
rect 7377 13277 7389 13280
rect 7423 13277 7435 13311
rect 7377 13271 7435 13277
rect 7466 13268 7472 13320
rect 7524 13308 7530 13320
rect 7576 13308 7604 13339
rect 8662 13336 8668 13348
rect 8720 13336 8726 13388
rect 9674 13376 9680 13388
rect 9635 13348 9680 13376
rect 9674 13336 9680 13348
rect 9732 13336 9738 13388
rect 11532 13385 11560 13416
rect 12452 13416 13829 13444
rect 11517 13379 11575 13385
rect 11517 13345 11529 13379
rect 11563 13345 11575 13379
rect 11698 13376 11704 13388
rect 11659 13348 11704 13376
rect 11517 13339 11575 13345
rect 11698 13336 11704 13348
rect 11756 13376 11762 13388
rect 12452 13385 12480 13416
rect 13817 13413 13829 13416
rect 13863 13413 13875 13447
rect 13817 13407 13875 13413
rect 12253 13379 12311 13385
rect 12253 13376 12265 13379
rect 11756 13348 12265 13376
rect 11756 13336 11762 13348
rect 12253 13345 12265 13348
rect 12299 13345 12311 13379
rect 12253 13339 12311 13345
rect 12437 13379 12495 13385
rect 12437 13345 12449 13379
rect 12483 13345 12495 13379
rect 12437 13339 12495 13345
rect 13725 13379 13783 13385
rect 13725 13345 13737 13379
rect 13771 13376 13783 13379
rect 13998 13376 14004 13388
rect 13771 13348 14004 13376
rect 13771 13345 13783 13348
rect 13725 13339 13783 13345
rect 13998 13336 14004 13348
rect 14056 13376 14062 13388
rect 14108 13376 14136 13475
rect 15102 13472 15108 13484
rect 15160 13472 15166 13524
rect 21726 13512 21732 13524
rect 21687 13484 21732 13512
rect 21726 13472 21732 13484
rect 21784 13472 21790 13524
rect 23474 13512 23480 13524
rect 23435 13484 23480 13512
rect 23474 13472 23480 13484
rect 23532 13472 23538 13524
rect 18230 13444 18236 13456
rect 18191 13416 18236 13444
rect 18230 13404 18236 13416
rect 18288 13404 18294 13456
rect 14918 13376 14924 13388
rect 14056 13348 14136 13376
rect 14879 13348 14924 13376
rect 14056 13336 14062 13348
rect 14918 13336 14924 13348
rect 14976 13336 14982 13388
rect 16666 13336 16672 13388
rect 16724 13376 16730 13388
rect 16853 13379 16911 13385
rect 16853 13376 16865 13379
rect 16724 13348 16865 13376
rect 16724 13336 16730 13348
rect 16853 13345 16865 13348
rect 16899 13345 16911 13379
rect 21744 13376 21772 13472
rect 21913 13379 21971 13385
rect 21913 13376 21925 13379
rect 21744 13348 21925 13376
rect 16853 13339 16911 13345
rect 21913 13345 21925 13348
rect 21959 13376 21971 13379
rect 22002 13376 22008 13388
rect 21959 13348 22008 13376
rect 21959 13345 21971 13348
rect 21913 13339 21971 13345
rect 22002 13336 22008 13348
rect 22060 13336 22066 13388
rect 22186 13376 22192 13388
rect 22147 13348 22192 13376
rect 22186 13336 22192 13348
rect 22244 13336 22250 13388
rect 16577 13311 16635 13317
rect 16577 13308 16589 13311
rect 7524 13280 7604 13308
rect 7524 13268 7530 13280
rect 4540 13172 4568 13268
rect 7576 13240 7604 13280
rect 16408 13280 16589 13308
rect 9858 13240 9864 13252
rect 7576 13212 9864 13240
rect 9858 13200 9864 13212
rect 9916 13200 9922 13252
rect 6273 13175 6331 13181
rect 6273 13172 6285 13175
rect 4540 13144 6285 13172
rect 6273 13141 6285 13144
rect 6319 13141 6331 13175
rect 12710 13172 12716 13184
rect 12671 13144 12716 13172
rect 6273 13135 6331 13141
rect 12710 13132 12716 13144
rect 12768 13132 12774 13184
rect 14737 13175 14795 13181
rect 14737 13141 14749 13175
rect 14783 13172 14795 13175
rect 15378 13172 15384 13184
rect 14783 13144 15384 13172
rect 14783 13141 14795 13144
rect 14737 13135 14795 13141
rect 15378 13132 15384 13144
rect 15436 13172 15442 13184
rect 16408 13181 16436 13280
rect 16577 13277 16589 13280
rect 16623 13277 16635 13311
rect 16577 13271 16635 13277
rect 16393 13175 16451 13181
rect 16393 13172 16405 13175
rect 15436 13144 16405 13172
rect 15436 13132 15442 13144
rect 16393 13141 16405 13144
rect 16439 13141 16451 13175
rect 16393 13135 16451 13141
rect 1104 13082 24656 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 24656 13082
rect 1104 13008 24656 13030
rect 4433 12971 4491 12977
rect 4433 12937 4445 12971
rect 4479 12968 4491 12971
rect 5534 12968 5540 12980
rect 4479 12940 5540 12968
rect 4479 12937 4491 12940
rect 4433 12931 4491 12937
rect 4632 12841 4660 12940
rect 5534 12928 5540 12940
rect 5592 12928 5598 12980
rect 5718 12968 5724 12980
rect 5679 12940 5724 12968
rect 5718 12928 5724 12940
rect 5776 12928 5782 12980
rect 7929 12971 7987 12977
rect 7929 12937 7941 12971
rect 7975 12968 7987 12971
rect 8386 12968 8392 12980
rect 7975 12940 8392 12968
rect 7975 12937 7987 12940
rect 7929 12931 7987 12937
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12801 4675 12835
rect 4617 12795 4675 12801
rect 4709 12767 4767 12773
rect 4709 12733 4721 12767
rect 4755 12733 4767 12767
rect 4709 12727 4767 12733
rect 4724 12696 4752 12727
rect 5258 12724 5264 12776
rect 5316 12764 5322 12776
rect 5445 12767 5503 12773
rect 5316 12736 5361 12764
rect 5316 12724 5322 12736
rect 5445 12733 5457 12767
rect 5491 12764 5503 12767
rect 5810 12764 5816 12776
rect 5491 12736 5816 12764
rect 5491 12733 5503 12736
rect 5445 12727 5503 12733
rect 5810 12724 5816 12736
rect 5868 12724 5874 12776
rect 7561 12767 7619 12773
rect 7561 12733 7573 12767
rect 7607 12764 7619 12767
rect 7944 12764 7972 12931
rect 8386 12928 8392 12940
rect 8444 12968 8450 12980
rect 8570 12968 8576 12980
rect 8444 12940 8576 12968
rect 8444 12928 8450 12940
rect 8570 12928 8576 12940
rect 8628 12928 8634 12980
rect 10505 12971 10563 12977
rect 10505 12937 10517 12971
rect 10551 12968 10563 12971
rect 11698 12968 11704 12980
rect 10551 12940 11704 12968
rect 10551 12937 10563 12940
rect 10505 12931 10563 12937
rect 11698 12928 11704 12940
rect 11756 12968 11762 12980
rect 20530 12968 20536 12980
rect 11756 12940 15056 12968
rect 20491 12940 20536 12968
rect 11756 12928 11762 12940
rect 13998 12900 14004 12912
rect 13959 12872 14004 12900
rect 13998 12860 14004 12872
rect 14056 12860 14062 12912
rect 12710 12832 12716 12844
rect 12671 12804 12716 12832
rect 12710 12792 12716 12804
rect 12768 12792 12774 12844
rect 13078 12792 13084 12844
rect 13136 12832 13142 12844
rect 14185 12835 14243 12841
rect 14185 12832 14197 12835
rect 13136 12804 14197 12832
rect 13136 12792 13142 12804
rect 14185 12801 14197 12804
rect 14231 12801 14243 12835
rect 15028 12832 15056 12940
rect 20530 12928 20536 12940
rect 20588 12928 20594 12980
rect 20548 12832 20576 12928
rect 20625 12835 20683 12841
rect 20625 12832 20637 12835
rect 15028 12804 15240 12832
rect 20548 12804 20637 12832
rect 14185 12795 14243 12801
rect 7607 12736 7972 12764
rect 7607 12733 7619 12736
rect 7561 12727 7619 12733
rect 9858 12724 9864 12776
rect 9916 12764 9922 12776
rect 10321 12767 10379 12773
rect 10321 12764 10333 12767
rect 9916 12736 10333 12764
rect 9916 12724 9922 12736
rect 10321 12733 10333 12736
rect 10367 12733 10379 12767
rect 10321 12727 10379 12733
rect 12437 12767 12495 12773
rect 12437 12733 12449 12767
rect 12483 12764 12495 12767
rect 13096 12764 13124 12792
rect 15212 12773 15240 12804
rect 20625 12801 20637 12804
rect 20671 12801 20683 12835
rect 20625 12795 20683 12801
rect 15013 12767 15071 12773
rect 15013 12764 15025 12767
rect 12483 12736 13124 12764
rect 14844 12736 15025 12764
rect 12483 12733 12495 12736
rect 12437 12727 12495 12733
rect 4890 12696 4896 12708
rect 4724 12668 4896 12696
rect 4890 12656 4896 12668
rect 4948 12696 4954 12708
rect 7466 12696 7472 12708
rect 4948 12668 7472 12696
rect 4948 12656 4954 12668
rect 7466 12656 7472 12668
rect 7524 12656 7530 12708
rect 6914 12588 6920 12640
rect 6972 12628 6978 12640
rect 7653 12631 7711 12637
rect 7653 12628 7665 12631
rect 6972 12600 7665 12628
rect 6972 12588 6978 12600
rect 7653 12597 7665 12600
rect 7699 12597 7711 12631
rect 7653 12591 7711 12597
rect 12342 12588 12348 12640
rect 12400 12628 12406 12640
rect 13446 12628 13452 12640
rect 12400 12600 13452 12628
rect 12400 12588 12406 12600
rect 13446 12588 13452 12600
rect 13504 12628 13510 12640
rect 14844 12637 14872 12736
rect 15013 12733 15025 12736
rect 15059 12733 15071 12767
rect 15013 12727 15071 12733
rect 15197 12767 15255 12773
rect 15197 12733 15209 12767
rect 15243 12764 15255 12767
rect 15746 12764 15752 12776
rect 15243 12736 15752 12764
rect 15243 12733 15255 12736
rect 15197 12727 15255 12733
rect 15746 12724 15752 12736
rect 15804 12724 15810 12776
rect 15933 12767 15991 12773
rect 15933 12733 15945 12767
rect 15979 12764 15991 12767
rect 16574 12764 16580 12776
rect 15979 12736 16580 12764
rect 15979 12733 15991 12736
rect 15933 12727 15991 12733
rect 16574 12724 16580 12736
rect 16632 12724 16638 12776
rect 20806 12764 20812 12776
rect 20767 12736 20812 12764
rect 20806 12724 20812 12736
rect 20864 12724 20870 12776
rect 21361 12767 21419 12773
rect 21361 12733 21373 12767
rect 21407 12733 21419 12767
rect 21361 12727 21419 12733
rect 21545 12767 21603 12773
rect 21545 12733 21557 12767
rect 21591 12764 21603 12767
rect 22278 12764 22284 12776
rect 21591 12736 22284 12764
rect 21591 12733 21603 12736
rect 21545 12727 21603 12733
rect 20824 12696 20852 12724
rect 21376 12696 21404 12727
rect 22278 12724 22284 12736
rect 22336 12724 22342 12776
rect 20824 12668 21404 12696
rect 14829 12631 14887 12637
rect 14829 12628 14841 12631
rect 13504 12600 14841 12628
rect 13504 12588 13510 12600
rect 14829 12597 14841 12600
rect 14875 12597 14887 12631
rect 16206 12628 16212 12640
rect 16167 12600 16212 12628
rect 14829 12591 14887 12597
rect 16206 12588 16212 12600
rect 16264 12588 16270 12640
rect 21818 12628 21824 12640
rect 21779 12600 21824 12628
rect 21818 12588 21824 12600
rect 21876 12588 21882 12640
rect 1104 12538 24656 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 24656 12538
rect 1104 12464 24656 12486
rect 5077 12427 5135 12433
rect 5077 12393 5089 12427
rect 5123 12424 5135 12427
rect 5258 12424 5264 12436
rect 5123 12396 5264 12424
rect 5123 12393 5135 12396
rect 5077 12387 5135 12393
rect 5258 12384 5264 12396
rect 5316 12384 5322 12436
rect 8478 12424 8484 12436
rect 8439 12396 8484 12424
rect 8478 12384 8484 12396
rect 8536 12384 8542 12436
rect 11974 12384 11980 12436
rect 12032 12424 12038 12436
rect 17954 12424 17960 12436
rect 12032 12396 17960 12424
rect 12032 12384 12038 12396
rect 17954 12384 17960 12396
rect 18012 12384 18018 12436
rect 21361 12427 21419 12433
rect 21361 12393 21373 12427
rect 21407 12424 21419 12427
rect 22002 12424 22008 12436
rect 21407 12396 22008 12424
rect 21407 12393 21419 12396
rect 21361 12387 21419 12393
rect 4890 12288 4896 12300
rect 4851 12260 4896 12288
rect 4890 12248 4896 12260
rect 4948 12248 4954 12300
rect 5258 12248 5264 12300
rect 5316 12288 5322 12300
rect 6181 12291 6239 12297
rect 6181 12288 6193 12291
rect 5316 12260 6193 12288
rect 5316 12248 5322 12260
rect 6181 12257 6193 12260
rect 6227 12288 6239 12291
rect 6730 12288 6736 12300
rect 6227 12260 6736 12288
rect 6227 12257 6239 12260
rect 6181 12251 6239 12257
rect 6730 12248 6736 12260
rect 6788 12248 6794 12300
rect 6914 12288 6920 12300
rect 6875 12260 6920 12288
rect 6914 12248 6920 12260
rect 6972 12248 6978 12300
rect 8205 12291 8263 12297
rect 8205 12257 8217 12291
rect 8251 12288 8263 12291
rect 8496 12288 8524 12384
rect 17310 12356 17316 12368
rect 17271 12328 17316 12356
rect 17310 12316 17316 12328
rect 17368 12316 17374 12368
rect 8251 12260 8524 12288
rect 15933 12291 15991 12297
rect 8251 12257 8263 12260
rect 8205 12251 8263 12257
rect 15933 12257 15945 12291
rect 15979 12288 15991 12291
rect 16206 12288 16212 12300
rect 15979 12260 16212 12288
rect 15979 12257 15991 12260
rect 15933 12251 15991 12257
rect 16206 12248 16212 12260
rect 16264 12248 16270 12300
rect 18322 12288 18328 12300
rect 18283 12260 18328 12288
rect 18322 12248 18328 12260
rect 18380 12248 18386 12300
rect 21358 12248 21364 12300
rect 21416 12288 21422 12300
rect 21468 12297 21496 12396
rect 22002 12384 22008 12396
rect 22060 12384 22066 12436
rect 23109 12359 23167 12365
rect 23109 12325 23121 12359
rect 23155 12356 23167 12359
rect 23382 12356 23388 12368
rect 23155 12328 23388 12356
rect 23155 12325 23167 12328
rect 23109 12319 23167 12325
rect 23382 12316 23388 12328
rect 23440 12316 23446 12368
rect 21453 12291 21511 12297
rect 21453 12288 21465 12291
rect 21416 12260 21465 12288
rect 21416 12248 21422 12260
rect 21453 12257 21465 12260
rect 21499 12257 21511 12291
rect 21453 12251 21511 12257
rect 21729 12291 21787 12297
rect 21729 12257 21741 12291
rect 21775 12288 21787 12291
rect 21818 12288 21824 12300
rect 21775 12260 21824 12288
rect 21775 12257 21787 12260
rect 21729 12251 21787 12257
rect 21818 12248 21824 12260
rect 21876 12248 21882 12300
rect 5166 12180 5172 12232
rect 5224 12220 5230 12232
rect 5997 12223 6055 12229
rect 5997 12220 6009 12223
rect 5224 12192 6009 12220
rect 5224 12180 5230 12192
rect 5997 12189 6009 12192
rect 6043 12189 6055 12223
rect 5997 12183 6055 12189
rect 7466 12180 7472 12232
rect 7524 12220 7530 12232
rect 12342 12220 12348 12232
rect 7524 12192 12348 12220
rect 7524 12180 7530 12192
rect 12342 12180 12348 12192
rect 12400 12180 12406 12232
rect 15657 12223 15715 12229
rect 15657 12189 15669 12223
rect 15703 12220 15715 12223
rect 16114 12220 16120 12232
rect 15703 12192 16120 12220
rect 15703 12189 15715 12192
rect 15657 12183 15715 12189
rect 16114 12180 16120 12192
rect 16172 12220 16178 12232
rect 17405 12223 17463 12229
rect 17405 12220 17417 12223
rect 16172 12192 17417 12220
rect 16172 12180 16178 12192
rect 17405 12189 17417 12192
rect 17451 12189 17463 12223
rect 17405 12183 17463 12189
rect 5166 12044 5172 12096
rect 5224 12084 5230 12096
rect 5813 12087 5871 12093
rect 5813 12084 5825 12087
rect 5224 12056 5825 12084
rect 5224 12044 5230 12056
rect 5813 12053 5825 12056
rect 5859 12053 5871 12087
rect 5813 12047 5871 12053
rect 7193 12087 7251 12093
rect 7193 12053 7205 12087
rect 7239 12084 7251 12087
rect 7282 12084 7288 12096
rect 7239 12056 7288 12084
rect 7239 12053 7251 12056
rect 7193 12047 7251 12053
rect 7282 12044 7288 12056
rect 7340 12044 7346 12096
rect 8294 12084 8300 12096
rect 8255 12056 8300 12084
rect 8294 12044 8300 12056
rect 8352 12044 8358 12096
rect 16390 12044 16396 12096
rect 16448 12084 16454 12096
rect 18141 12087 18199 12093
rect 18141 12084 18153 12087
rect 16448 12056 18153 12084
rect 16448 12044 16454 12056
rect 18141 12053 18153 12056
rect 18187 12084 18199 12087
rect 19334 12084 19340 12096
rect 18187 12056 19340 12084
rect 18187 12053 18199 12056
rect 18141 12047 18199 12053
rect 19334 12044 19340 12056
rect 19392 12044 19398 12096
rect 1104 11994 24656 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 24656 11994
rect 1104 11920 24656 11942
rect 4341 11883 4399 11889
rect 4341 11849 4353 11883
rect 4387 11880 4399 11883
rect 7374 11880 7380 11892
rect 4387 11852 7380 11880
rect 4387 11849 4399 11852
rect 4341 11843 4399 11849
rect 2777 11747 2835 11753
rect 2777 11713 2789 11747
rect 2823 11744 2835 11747
rect 4356 11744 4384 11843
rect 7374 11840 7380 11852
rect 7432 11840 7438 11892
rect 8386 11880 8392 11892
rect 8347 11852 8392 11880
rect 8386 11840 8392 11852
rect 8444 11840 8450 11892
rect 16574 11880 16580 11892
rect 16535 11852 16580 11880
rect 16574 11840 16580 11852
rect 16632 11840 16638 11892
rect 16853 11883 16911 11889
rect 16853 11849 16865 11883
rect 16899 11880 16911 11883
rect 17310 11880 17316 11892
rect 16899 11852 17316 11880
rect 16899 11849 16911 11852
rect 16853 11843 16911 11849
rect 4525 11815 4583 11821
rect 4525 11781 4537 11815
rect 4571 11812 4583 11815
rect 4614 11812 4620 11824
rect 4571 11784 4620 11812
rect 4571 11781 4583 11784
rect 4525 11775 4583 11781
rect 2823 11716 4384 11744
rect 4540 11744 4568 11775
rect 4614 11772 4620 11784
rect 4672 11772 4678 11824
rect 7009 11747 7067 11753
rect 7009 11744 7021 11747
rect 4540 11716 7021 11744
rect 2823 11713 2835 11716
rect 2777 11707 2835 11713
rect 2498 11676 2504 11688
rect 2411 11648 2504 11676
rect 2498 11636 2504 11648
rect 2556 11676 2562 11688
rect 4540 11676 4568 11716
rect 7009 11713 7021 11716
rect 7055 11713 7067 11747
rect 7282 11744 7288 11756
rect 7243 11716 7288 11744
rect 7009 11707 7067 11713
rect 2556 11648 4568 11676
rect 7024 11676 7052 11707
rect 7282 11704 7288 11716
rect 7340 11704 7346 11756
rect 7098 11676 7104 11688
rect 7024 11648 7104 11676
rect 2556 11636 2562 11648
rect 7098 11636 7104 11648
rect 7156 11676 7162 11688
rect 8757 11679 8815 11685
rect 8757 11676 8769 11679
rect 7156 11648 8769 11676
rect 7156 11636 7162 11648
rect 8757 11645 8769 11648
rect 8803 11676 8815 11679
rect 8846 11676 8852 11688
rect 8803 11648 8852 11676
rect 8803 11645 8815 11648
rect 8757 11639 8815 11645
rect 8846 11636 8852 11648
rect 8904 11636 8910 11688
rect 16485 11679 16543 11685
rect 16485 11645 16497 11679
rect 16531 11676 16543 11679
rect 16868 11676 16896 11843
rect 17310 11840 17316 11852
rect 17368 11840 17374 11892
rect 19886 11880 19892 11892
rect 19536 11852 19892 11880
rect 19536 11753 19564 11852
rect 19886 11840 19892 11852
rect 19944 11880 19950 11892
rect 21358 11880 21364 11892
rect 19944 11852 21364 11880
rect 19944 11840 19950 11852
rect 21358 11840 21364 11852
rect 21416 11840 21422 11892
rect 22278 11880 22284 11892
rect 22239 11852 22284 11880
rect 22278 11840 22284 11852
rect 22336 11840 22342 11892
rect 19521 11747 19579 11753
rect 19521 11713 19533 11747
rect 19567 11713 19579 11747
rect 19521 11707 19579 11713
rect 19797 11747 19855 11753
rect 19797 11713 19809 11747
rect 19843 11744 19855 11747
rect 20806 11744 20812 11756
rect 19843 11716 20812 11744
rect 19843 11713 19855 11716
rect 19797 11707 19855 11713
rect 20806 11704 20812 11716
rect 20864 11704 20870 11756
rect 16531 11648 16896 11676
rect 22189 11679 22247 11685
rect 16531 11645 16543 11648
rect 16485 11639 16543 11645
rect 22189 11645 22201 11679
rect 22235 11676 22247 11679
rect 23382 11676 23388 11688
rect 22235 11648 23388 11676
rect 22235 11645 22247 11648
rect 22189 11639 22247 11645
rect 23382 11636 23388 11648
rect 23440 11636 23446 11688
rect 3878 11540 3884 11552
rect 3839 11512 3884 11540
rect 3878 11500 3884 11512
rect 3936 11500 3942 11552
rect 20898 11540 20904 11552
rect 20859 11512 20904 11540
rect 20898 11500 20904 11512
rect 20956 11500 20962 11552
rect 1104 11450 24656 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 24656 11450
rect 1104 11376 24656 11398
rect 8478 11336 8484 11348
rect 8439 11308 8484 11336
rect 8478 11296 8484 11308
rect 8536 11296 8542 11348
rect 8846 11336 8852 11348
rect 8807 11308 8852 11336
rect 8846 11296 8852 11308
rect 8904 11296 8910 11348
rect 19061 11339 19119 11345
rect 19061 11305 19073 11339
rect 19107 11336 19119 11339
rect 19426 11336 19432 11348
rect 19107 11308 19432 11336
rect 19107 11305 19119 11308
rect 19061 11299 19119 11305
rect 7098 11200 7104 11212
rect 7059 11172 7104 11200
rect 7098 11160 7104 11172
rect 7156 11160 7162 11212
rect 12894 11160 12900 11212
rect 12952 11200 12958 11212
rect 13265 11203 13323 11209
rect 13265 11200 13277 11203
rect 12952 11172 13277 11200
rect 12952 11160 12958 11172
rect 13265 11169 13277 11172
rect 13311 11169 13323 11203
rect 13265 11163 13323 11169
rect 13633 11203 13691 11209
rect 13633 11169 13645 11203
rect 13679 11200 13691 11203
rect 13998 11200 14004 11212
rect 13679 11172 14004 11200
rect 13679 11169 13691 11172
rect 13633 11163 13691 11169
rect 13998 11160 14004 11172
rect 14056 11160 14062 11212
rect 16390 11200 16396 11212
rect 16351 11172 16396 11200
rect 16390 11160 16396 11172
rect 16448 11160 16454 11212
rect 7374 11132 7380 11144
rect 7335 11104 7380 11132
rect 7374 11092 7380 11104
rect 7432 11092 7438 11144
rect 12710 11132 12716 11144
rect 12671 11104 12716 11132
rect 12710 11092 12716 11104
rect 12768 11092 12774 11144
rect 13357 11135 13415 11141
rect 13357 11101 13369 11135
rect 13403 11101 13415 11135
rect 13357 11095 13415 11101
rect 13541 11135 13599 11141
rect 13541 11101 13553 11135
rect 13587 11132 13599 11135
rect 13814 11132 13820 11144
rect 13587 11104 13820 11132
rect 13587 11101 13599 11104
rect 13541 11095 13599 11101
rect 13372 11064 13400 11095
rect 13814 11092 13820 11104
rect 13872 11092 13878 11144
rect 17221 11135 17279 11141
rect 17221 11101 17233 11135
rect 17267 11101 17279 11135
rect 17221 11095 17279 11101
rect 17497 11135 17555 11141
rect 17497 11101 17509 11135
rect 17543 11132 17555 11135
rect 19076 11132 19104 11299
rect 19426 11296 19432 11308
rect 19484 11336 19490 11348
rect 24210 11336 24216 11348
rect 19484 11308 24216 11336
rect 19484 11296 19490 11308
rect 24210 11296 24216 11308
rect 24268 11296 24274 11348
rect 19334 11160 19340 11212
rect 19392 11200 19398 11212
rect 19889 11203 19947 11209
rect 19889 11200 19901 11203
rect 19392 11172 19901 11200
rect 19392 11160 19398 11172
rect 19889 11169 19901 11172
rect 19935 11169 19947 11203
rect 19889 11163 19947 11169
rect 17543 11104 19104 11132
rect 17543 11101 17555 11104
rect 17497 11095 17555 11101
rect 13722 11064 13728 11076
rect 13372 11036 13728 11064
rect 13722 11024 13728 11036
rect 13780 11064 13786 11076
rect 13909 11067 13967 11073
rect 13909 11064 13921 11067
rect 13780 11036 13921 11064
rect 13780 11024 13786 11036
rect 13909 11033 13921 11036
rect 13955 11033 13967 11067
rect 16206 11064 16212 11076
rect 16167 11036 16212 11064
rect 13909 11027 13967 11033
rect 16206 11024 16212 11036
rect 16264 11024 16270 11076
rect 12802 10956 12808 11008
rect 12860 10996 12866 11008
rect 16574 10996 16580 11008
rect 12860 10968 16580 10996
rect 12860 10956 12866 10968
rect 16574 10956 16580 10968
rect 16632 10956 16638 11008
rect 17236 10996 17264 11095
rect 19245 11067 19303 11073
rect 19245 11064 19257 11067
rect 18156 11036 19257 11064
rect 18156 10996 18184 11036
rect 19245 11033 19257 11036
rect 19291 11064 19303 11067
rect 19705 11067 19763 11073
rect 19705 11064 19717 11067
rect 19291 11036 19717 11064
rect 19291 11033 19303 11036
rect 19245 11027 19303 11033
rect 19705 11033 19717 11036
rect 19751 11064 19763 11067
rect 19886 11064 19892 11076
rect 19751 11036 19892 11064
rect 19751 11033 19763 11036
rect 19705 11027 19763 11033
rect 19886 11024 19892 11036
rect 19944 11024 19950 11076
rect 17236 10968 18184 10996
rect 18322 10956 18328 11008
rect 18380 10996 18386 11008
rect 18601 10999 18659 11005
rect 18601 10996 18613 10999
rect 18380 10968 18613 10996
rect 18380 10956 18386 10968
rect 18601 10965 18613 10968
rect 18647 10965 18659 10999
rect 18601 10959 18659 10965
rect 1104 10906 24656 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 24656 10906
rect 1104 10832 24656 10854
rect 4341 10795 4399 10801
rect 4341 10761 4353 10795
rect 4387 10792 4399 10795
rect 4614 10792 4620 10804
rect 4387 10764 4620 10792
rect 4387 10761 4399 10764
rect 4341 10755 4399 10761
rect 4614 10752 4620 10764
rect 4672 10752 4678 10804
rect 7374 10752 7380 10804
rect 7432 10792 7438 10804
rect 8021 10795 8079 10801
rect 8021 10792 8033 10795
rect 7432 10764 8033 10792
rect 7432 10752 7438 10764
rect 8021 10761 8033 10764
rect 8067 10761 8079 10795
rect 8021 10755 8079 10761
rect 8110 10752 8116 10804
rect 8168 10792 8174 10804
rect 12802 10792 12808 10804
rect 8168 10764 12808 10792
rect 8168 10752 8174 10764
rect 12802 10752 12808 10764
rect 12860 10752 12866 10804
rect 12894 10752 12900 10804
rect 12952 10792 12958 10804
rect 13817 10795 13875 10801
rect 13817 10792 13829 10795
rect 12952 10764 13829 10792
rect 12952 10752 12958 10764
rect 13817 10761 13829 10764
rect 13863 10761 13875 10795
rect 13817 10755 13875 10761
rect 13998 10752 14004 10804
rect 14056 10792 14062 10804
rect 19429 10795 19487 10801
rect 19429 10792 19441 10795
rect 14056 10764 19441 10792
rect 14056 10752 14062 10764
rect 19429 10761 19441 10764
rect 19475 10761 19487 10795
rect 19429 10755 19487 10761
rect 19886 10752 19892 10804
rect 19944 10792 19950 10804
rect 20349 10795 20407 10801
rect 20349 10792 20361 10795
rect 19944 10764 20361 10792
rect 19944 10752 19950 10764
rect 20349 10761 20361 10764
rect 20395 10761 20407 10795
rect 20349 10755 20407 10761
rect 14277 10727 14335 10733
rect 14277 10693 14289 10727
rect 14323 10724 14335 10727
rect 15378 10724 15384 10736
rect 14323 10696 15384 10724
rect 14323 10693 14335 10696
rect 14277 10687 14335 10693
rect 2498 10656 2504 10668
rect 2459 10628 2504 10656
rect 2498 10616 2504 10628
rect 2556 10616 2562 10668
rect 6730 10616 6736 10668
rect 6788 10656 6794 10668
rect 6788 10628 7236 10656
rect 6788 10616 6794 10628
rect 2774 10548 2780 10600
rect 2832 10588 2838 10600
rect 2832 10560 2877 10588
rect 2832 10548 2838 10560
rect 6546 10548 6552 10600
rect 6604 10588 6610 10600
rect 6822 10588 6828 10600
rect 6604 10560 6828 10588
rect 6604 10548 6610 10560
rect 6822 10548 6828 10560
rect 6880 10548 6886 10600
rect 7024 10597 7052 10628
rect 7009 10591 7067 10597
rect 7009 10557 7021 10591
rect 7055 10557 7067 10591
rect 7208 10588 7236 10628
rect 8018 10616 8024 10668
rect 8076 10656 8082 10668
rect 12158 10656 12164 10668
rect 8076 10628 12164 10656
rect 8076 10616 8082 10628
rect 12158 10616 12164 10628
rect 12216 10616 12222 10668
rect 12710 10656 12716 10668
rect 12671 10628 12716 10656
rect 12710 10616 12716 10628
rect 12768 10616 12774 10668
rect 14292 10656 14320 10687
rect 15378 10684 15384 10696
rect 15436 10684 15442 10736
rect 16574 10684 16580 10736
rect 16632 10724 16638 10736
rect 17770 10724 17776 10736
rect 16632 10696 17776 10724
rect 16632 10684 16638 10696
rect 17770 10684 17776 10696
rect 17828 10684 17834 10736
rect 18322 10656 18328 10668
rect 13280 10628 14320 10656
rect 18283 10628 18328 10656
rect 7561 10591 7619 10597
rect 7561 10588 7573 10591
rect 7208 10560 7573 10588
rect 7009 10551 7067 10557
rect 7561 10557 7573 10560
rect 7607 10557 7619 10591
rect 7561 10551 7619 10557
rect 7745 10591 7803 10597
rect 7745 10557 7757 10591
rect 7791 10588 7803 10591
rect 8294 10588 8300 10600
rect 7791 10560 8300 10588
rect 7791 10557 7803 10560
rect 7745 10551 7803 10557
rect 8294 10548 8300 10560
rect 8352 10548 8358 10600
rect 12437 10591 12495 10597
rect 12437 10557 12449 10591
rect 12483 10588 12495 10591
rect 13280 10588 13308 10628
rect 18322 10616 18328 10628
rect 18380 10616 18386 10668
rect 20364 10656 20392 10755
rect 20530 10656 20536 10668
rect 20364 10628 20536 10656
rect 20530 10616 20536 10628
rect 20588 10616 20594 10668
rect 20809 10659 20867 10665
rect 20809 10625 20821 10659
rect 20855 10656 20867 10659
rect 20898 10656 20904 10668
rect 20855 10628 20904 10656
rect 20855 10625 20867 10628
rect 20809 10619 20867 10625
rect 20898 10616 20904 10628
rect 20956 10616 20962 10668
rect 12483 10560 13308 10588
rect 18049 10591 18107 10597
rect 12483 10557 12495 10560
rect 12437 10551 12495 10557
rect 18049 10557 18061 10591
rect 18095 10557 18107 10591
rect 18049 10551 18107 10557
rect 18064 10520 18092 10551
rect 17788 10492 18092 10520
rect 3878 10452 3884 10464
rect 3839 10424 3884 10452
rect 3878 10412 3884 10424
rect 3936 10412 3942 10464
rect 6546 10452 6552 10464
rect 6507 10424 6552 10452
rect 6546 10412 6552 10424
rect 6604 10412 6610 10464
rect 16206 10412 16212 10464
rect 16264 10452 16270 10464
rect 17788 10461 17816 10492
rect 17773 10455 17831 10461
rect 17773 10452 17785 10455
rect 16264 10424 17785 10452
rect 16264 10412 16270 10424
rect 17773 10421 17785 10424
rect 17819 10421 17831 10455
rect 17773 10415 17831 10421
rect 21450 10412 21456 10464
rect 21508 10452 21514 10464
rect 21913 10455 21971 10461
rect 21913 10452 21925 10455
rect 21508 10424 21925 10452
rect 21508 10412 21514 10424
rect 21913 10421 21925 10424
rect 21959 10421 21971 10455
rect 21913 10415 21971 10421
rect 1104 10362 24656 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 24656 10362
rect 1104 10288 24656 10310
rect 13630 10208 13636 10260
rect 13688 10248 13694 10260
rect 13817 10251 13875 10257
rect 13817 10248 13829 10251
rect 13688 10220 13829 10248
rect 13688 10208 13694 10220
rect 13817 10217 13829 10220
rect 13863 10217 13875 10251
rect 13817 10211 13875 10217
rect 20530 10208 20536 10260
rect 20588 10248 20594 10260
rect 20901 10251 20959 10257
rect 20901 10248 20913 10251
rect 20588 10220 20913 10248
rect 20588 10208 20594 10220
rect 20901 10217 20913 10220
rect 20947 10217 20959 10251
rect 20901 10211 20959 10217
rect 2774 10140 2780 10192
rect 2832 10180 2838 10192
rect 8205 10183 8263 10189
rect 8205 10180 8217 10183
rect 2832 10152 8217 10180
rect 2832 10140 2838 10152
rect 8205 10149 8217 10152
rect 8251 10149 8263 10183
rect 8205 10143 8263 10149
rect 6549 10115 6607 10121
rect 6549 10081 6561 10115
rect 6595 10112 6607 10115
rect 7006 10112 7012 10124
rect 6595 10084 7012 10112
rect 6595 10081 6607 10084
rect 6549 10075 6607 10081
rect 7006 10072 7012 10084
rect 7064 10072 7070 10124
rect 7745 10115 7803 10121
rect 7745 10081 7757 10115
rect 7791 10112 7803 10115
rect 13538 10112 13544 10124
rect 7791 10084 13544 10112
rect 7791 10081 7803 10084
rect 7745 10075 7803 10081
rect 13538 10072 13544 10084
rect 13596 10072 13602 10124
rect 13906 10072 13912 10124
rect 13964 10112 13970 10124
rect 15289 10115 15347 10121
rect 15289 10112 15301 10115
rect 13964 10084 15301 10112
rect 13964 10072 13970 10084
rect 15289 10081 15301 10084
rect 15335 10081 15347 10115
rect 20916 10112 20944 10211
rect 21085 10115 21143 10121
rect 21085 10112 21097 10115
rect 20916 10084 21097 10112
rect 15289 10075 15347 10081
rect 21085 10081 21097 10084
rect 21131 10081 21143 10115
rect 21085 10075 21143 10081
rect 21361 10115 21419 10121
rect 21361 10081 21373 10115
rect 21407 10112 21419 10115
rect 21450 10112 21456 10124
rect 21407 10084 21456 10112
rect 21407 10081 21419 10084
rect 21361 10075 21419 10081
rect 21450 10072 21456 10084
rect 21508 10072 21514 10124
rect 7653 10047 7711 10053
rect 7653 10013 7665 10047
rect 7699 10013 7711 10047
rect 12250 10044 12256 10056
rect 12211 10016 12256 10044
rect 7653 10007 7711 10013
rect 6733 9979 6791 9985
rect 6733 9945 6745 9979
rect 6779 9976 6791 9979
rect 7668 9976 7696 10007
rect 12250 10004 12256 10016
rect 12308 10004 12314 10056
rect 12526 10044 12532 10056
rect 12487 10016 12532 10044
rect 12526 10004 12532 10016
rect 12584 10004 12590 10056
rect 7742 9976 7748 9988
rect 6779 9948 7748 9976
rect 6779 9945 6791 9948
rect 6733 9939 6791 9945
rect 7742 9936 7748 9948
rect 7800 9936 7806 9988
rect 13906 9936 13912 9988
rect 13964 9976 13970 9988
rect 15381 9979 15439 9985
rect 15381 9976 15393 9979
rect 13964 9948 15393 9976
rect 13964 9936 13970 9948
rect 15381 9945 15393 9948
rect 15427 9945 15439 9979
rect 15381 9939 15439 9945
rect 7006 9908 7012 9920
rect 6967 9880 7012 9908
rect 7006 9868 7012 9880
rect 7064 9868 7070 9920
rect 13998 9908 14004 9920
rect 13959 9880 14004 9908
rect 13998 9868 14004 9880
rect 14056 9908 14062 9920
rect 16206 9908 16212 9920
rect 14056 9880 16212 9908
rect 14056 9868 14062 9880
rect 16206 9868 16212 9880
rect 16264 9868 16270 9920
rect 22462 9908 22468 9920
rect 22423 9880 22468 9908
rect 22462 9868 22468 9880
rect 22520 9868 22526 9920
rect 1104 9818 24656 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 24656 9818
rect 1104 9744 24656 9766
rect 20530 9664 20536 9716
rect 20588 9704 20594 9716
rect 20717 9707 20775 9713
rect 20717 9704 20729 9707
rect 20588 9676 20729 9704
rect 20588 9664 20594 9676
rect 20717 9673 20729 9676
rect 20763 9673 20775 9707
rect 20717 9667 20775 9673
rect 7742 9636 7748 9648
rect 7655 9608 7748 9636
rect 7742 9596 7748 9608
rect 7800 9636 7806 9648
rect 7800 9608 9352 9636
rect 7800 9596 7806 9608
rect 2774 9528 2780 9580
rect 2832 9568 2838 9580
rect 9324 9577 9352 9608
rect 12342 9596 12348 9648
rect 12400 9636 12406 9648
rect 13998 9636 14004 9648
rect 12400 9608 14004 9636
rect 12400 9596 12406 9608
rect 13998 9596 14004 9608
rect 14056 9596 14062 9648
rect 4249 9571 4307 9577
rect 4249 9568 4261 9571
rect 2832 9540 2877 9568
rect 2976 9540 4261 9568
rect 2832 9528 2838 9540
rect 2498 9500 2504 9512
rect 2411 9472 2504 9500
rect 2498 9460 2504 9472
rect 2556 9500 2562 9512
rect 2976 9500 3004 9540
rect 4249 9537 4261 9540
rect 4295 9537 4307 9571
rect 8481 9571 8539 9577
rect 8481 9568 8493 9571
rect 4249 9531 4307 9537
rect 5644 9540 8493 9568
rect 5644 9500 5672 9540
rect 8481 9537 8493 9540
rect 8527 9537 8539 9571
rect 8481 9531 8539 9537
rect 9309 9571 9367 9577
rect 9309 9537 9321 9571
rect 9355 9537 9367 9571
rect 9309 9531 9367 9537
rect 12526 9528 12532 9580
rect 12584 9568 12590 9580
rect 12897 9571 12955 9577
rect 12897 9568 12909 9571
rect 12584 9540 12909 9568
rect 12584 9528 12590 9540
rect 12897 9537 12909 9540
rect 12943 9537 12955 9571
rect 13814 9568 13820 9580
rect 13775 9540 13820 9568
rect 12897 9531 12955 9537
rect 13814 9528 13820 9540
rect 13872 9528 13878 9580
rect 20349 9571 20407 9577
rect 20349 9568 20361 9571
rect 13924 9540 20361 9568
rect 2556 9472 3004 9500
rect 3712 9472 5672 9500
rect 8021 9503 8079 9509
rect 2556 9460 2562 9472
rect 2774 9324 2780 9376
rect 2832 9364 2838 9376
rect 3712 9364 3740 9472
rect 8021 9469 8033 9503
rect 8067 9469 8079 9503
rect 9398 9500 9404 9512
rect 9359 9472 9404 9500
rect 8021 9463 8079 9469
rect 7926 9432 7932 9444
rect 7887 9404 7932 9432
rect 7926 9392 7932 9404
rect 7984 9392 7990 9444
rect 3878 9364 3884 9376
rect 2832 9336 3740 9364
rect 3839 9336 3884 9364
rect 2832 9324 2838 9336
rect 3878 9324 3884 9336
rect 3936 9324 3942 9376
rect 8036 9364 8064 9463
rect 9398 9460 9404 9472
rect 9456 9460 9462 9512
rect 10134 9460 10140 9512
rect 10192 9500 10198 9512
rect 13357 9503 13415 9509
rect 13357 9500 13369 9503
rect 10192 9472 13369 9500
rect 10192 9460 10198 9472
rect 13357 9469 13369 9472
rect 13403 9469 13415 9503
rect 13357 9463 13415 9469
rect 13541 9503 13599 9509
rect 13541 9469 13553 9503
rect 13587 9500 13599 9503
rect 13630 9500 13636 9512
rect 13587 9472 13636 9500
rect 13587 9469 13599 9472
rect 13541 9463 13599 9469
rect 8110 9392 8116 9444
rect 8168 9432 8174 9444
rect 9861 9435 9919 9441
rect 9861 9432 9873 9435
rect 8168 9404 9873 9432
rect 8168 9392 8174 9404
rect 9861 9401 9873 9404
rect 9907 9401 9919 9435
rect 9861 9395 9919 9401
rect 8665 9367 8723 9373
rect 8665 9364 8677 9367
rect 8036 9336 8677 9364
rect 8665 9333 8677 9336
rect 8711 9364 8723 9367
rect 11974 9364 11980 9376
rect 8711 9336 11980 9364
rect 8711 9333 8723 9336
rect 8665 9327 8723 9333
rect 11974 9324 11980 9336
rect 12032 9324 12038 9376
rect 13372 9364 13400 9463
rect 13630 9460 13636 9472
rect 13688 9460 13694 9512
rect 13924 9509 13952 9540
rect 20349 9537 20361 9540
rect 20395 9537 20407 9571
rect 20349 9531 20407 9537
rect 13909 9503 13967 9509
rect 13909 9469 13921 9503
rect 13955 9469 13967 9503
rect 13909 9463 13967 9469
rect 18969 9503 19027 9509
rect 18969 9469 18981 9503
rect 19015 9500 19027 9503
rect 19245 9503 19303 9509
rect 19015 9472 19104 9500
rect 19015 9469 19027 9472
rect 18969 9463 19027 9469
rect 13722 9364 13728 9376
rect 13372 9336 13728 9364
rect 13722 9324 13728 9336
rect 13780 9364 13786 9376
rect 14277 9367 14335 9373
rect 14277 9364 14289 9367
rect 13780 9336 14289 9364
rect 13780 9324 13786 9336
rect 14277 9333 14289 9336
rect 14323 9364 14335 9367
rect 15286 9364 15292 9376
rect 14323 9336 15292 9364
rect 14323 9333 14335 9336
rect 14277 9327 14335 9333
rect 15286 9324 15292 9336
rect 15344 9324 15350 9376
rect 19076 9364 19104 9472
rect 19245 9469 19257 9503
rect 19291 9500 19303 9503
rect 20070 9500 20076 9512
rect 19291 9472 20076 9500
rect 19291 9469 19303 9472
rect 19245 9463 19303 9469
rect 20070 9460 20076 9472
rect 20128 9460 20134 9512
rect 20530 9364 20536 9376
rect 19076 9336 20536 9364
rect 20530 9324 20536 9336
rect 20588 9324 20594 9376
rect 1104 9274 24656 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 24656 9274
rect 1104 9200 24656 9222
rect 7926 9120 7932 9172
rect 7984 9160 7990 9172
rect 9953 9163 10011 9169
rect 9953 9160 9965 9163
rect 7984 9132 9965 9160
rect 7984 9120 7990 9132
rect 9953 9129 9965 9132
rect 9999 9129 10011 9163
rect 14090 9160 14096 9172
rect 14051 9132 14096 9160
rect 9953 9123 10011 9129
rect 14090 9120 14096 9132
rect 14148 9120 14154 9172
rect 19426 9160 19432 9172
rect 19387 9132 19432 9160
rect 19426 9120 19432 9132
rect 19484 9120 19490 9172
rect 20530 9120 20536 9172
rect 20588 9160 20594 9172
rect 21361 9163 21419 9169
rect 21361 9160 21373 9163
rect 20588 9132 21373 9160
rect 20588 9120 20594 9132
rect 21361 9129 21373 9132
rect 21407 9129 21419 9163
rect 21361 9123 21419 9129
rect 7834 9092 7840 9104
rect 6472 9064 7840 9092
rect 6472 9033 6500 9064
rect 7834 9052 7840 9064
rect 7892 9052 7898 9104
rect 8665 9095 8723 9101
rect 8665 9092 8677 9095
rect 8036 9064 8677 9092
rect 6457 9027 6515 9033
rect 6457 8993 6469 9027
rect 6503 8993 6515 9027
rect 7742 9024 7748 9036
rect 7703 8996 7748 9024
rect 6457 8987 6515 8993
rect 7742 8984 7748 8996
rect 7800 8984 7806 9036
rect 8036 9033 8064 9064
rect 8665 9061 8677 9064
rect 8711 9092 8723 9095
rect 12066 9092 12072 9104
rect 8711 9064 12072 9092
rect 8711 9061 8723 9064
rect 8665 9055 8723 9061
rect 12066 9052 12072 9064
rect 12124 9052 12130 9104
rect 13814 9052 13820 9104
rect 13872 9092 13878 9104
rect 15381 9095 15439 9101
rect 15381 9092 15393 9095
rect 13872 9064 15393 9092
rect 13872 9052 13878 9064
rect 15381 9061 15393 9064
rect 15427 9061 15439 9095
rect 15381 9055 15439 9061
rect 7929 9027 7987 9033
rect 7929 8993 7941 9027
rect 7975 8993 7987 9027
rect 7929 8987 7987 8993
rect 8021 9027 8079 9033
rect 8021 8993 8033 9027
rect 8067 8993 8079 9027
rect 9674 9024 9680 9036
rect 9635 8996 9680 9024
rect 8021 8987 8079 8993
rect 6365 8959 6423 8965
rect 6365 8925 6377 8959
rect 6411 8956 6423 8959
rect 7760 8956 7788 8984
rect 6411 8928 7788 8956
rect 7944 8956 7972 8987
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 9861 9027 9919 9033
rect 9861 8993 9873 9027
rect 9907 8993 9919 9027
rect 9861 8987 9919 8993
rect 8294 8956 8300 8968
rect 7944 8928 8300 8956
rect 6411 8925 6423 8928
rect 6365 8919 6423 8925
rect 8294 8916 8300 8928
rect 8352 8916 8358 8968
rect 8386 8916 8392 8968
rect 8444 8956 8450 8968
rect 9876 8956 9904 8987
rect 13998 8984 14004 9036
rect 14056 9024 14062 9036
rect 14461 9027 14519 9033
rect 14461 9024 14473 9027
rect 14056 8996 14473 9024
rect 14056 8984 14062 8996
rect 14461 8993 14473 8996
rect 14507 8993 14519 9027
rect 15286 9024 15292 9036
rect 15199 8996 15292 9024
rect 14461 8987 14519 8993
rect 15286 8984 15292 8996
rect 15344 9024 15350 9036
rect 18601 9027 18659 9033
rect 15344 8996 15700 9024
rect 15344 8984 15350 8996
rect 8444 8928 9904 8956
rect 8444 8916 8450 8928
rect 10962 8916 10968 8968
rect 11020 8956 11026 8968
rect 12342 8956 12348 8968
rect 11020 8928 12348 8956
rect 11020 8916 11026 8928
rect 12342 8916 12348 8928
rect 12400 8956 12406 8968
rect 12713 8959 12771 8965
rect 12713 8956 12725 8959
rect 12400 8928 12725 8956
rect 12400 8916 12406 8928
rect 12713 8925 12725 8928
rect 12759 8925 12771 8959
rect 12986 8956 12992 8968
rect 12947 8928 12992 8956
rect 12713 8919 12771 8925
rect 12986 8916 12992 8928
rect 13044 8916 13050 8968
rect 4062 8848 4068 8900
rect 4120 8888 4126 8900
rect 12618 8888 12624 8900
rect 4120 8860 12624 8888
rect 4120 8848 4126 8860
rect 12618 8848 12624 8860
rect 12676 8848 12682 8900
rect 15672 8897 15700 8996
rect 18601 8993 18613 9027
rect 18647 9024 18659 9027
rect 19444 9024 19472 9120
rect 18647 8996 19472 9024
rect 21376 9024 21404 9123
rect 21545 9027 21603 9033
rect 21545 9024 21557 9027
rect 21376 8996 21557 9024
rect 18647 8993 18659 8996
rect 18601 8987 18659 8993
rect 21545 8993 21557 8996
rect 21591 8993 21603 9027
rect 21545 8987 21603 8993
rect 21821 9027 21879 9033
rect 21821 8993 21833 9027
rect 21867 9024 21879 9027
rect 22462 9024 22468 9036
rect 21867 8996 22468 9024
rect 21867 8993 21879 8996
rect 21821 8987 21879 8993
rect 22462 8984 22468 8996
rect 22520 8984 22526 9036
rect 15657 8891 15715 8897
rect 15657 8857 15669 8891
rect 15703 8888 15715 8891
rect 15703 8860 21496 8888
rect 15703 8857 15715 8860
rect 15657 8851 15715 8857
rect 2774 8780 2780 8832
rect 2832 8820 2838 8832
rect 6641 8823 6699 8829
rect 6641 8820 6653 8823
rect 2832 8792 6653 8820
rect 2832 8780 2838 8792
rect 6641 8789 6653 8792
rect 6687 8789 6699 8823
rect 8202 8820 8208 8832
rect 8163 8792 8208 8820
rect 6641 8783 6699 8789
rect 8202 8780 8208 8792
rect 8260 8780 8266 8832
rect 19245 8823 19303 8829
rect 19245 8789 19257 8823
rect 19291 8820 19303 8823
rect 19334 8820 19340 8832
rect 19291 8792 19340 8820
rect 19291 8789 19303 8792
rect 19245 8783 19303 8789
rect 19334 8780 19340 8792
rect 19392 8780 19398 8832
rect 21468 8820 21496 8860
rect 22925 8823 22983 8829
rect 22925 8820 22937 8823
rect 21468 8792 22937 8820
rect 22925 8789 22937 8792
rect 22971 8789 22983 8823
rect 22925 8783 22983 8789
rect 1104 8730 24656 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 24656 8730
rect 1104 8656 24656 8678
rect 8386 8616 8392 8628
rect 8347 8588 8392 8616
rect 8386 8576 8392 8588
rect 8444 8576 8450 8628
rect 10134 8616 10140 8628
rect 10095 8588 10140 8616
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 18601 8619 18659 8625
rect 18601 8585 18613 8619
rect 18647 8616 18659 8619
rect 20070 8616 20076 8628
rect 18647 8588 19656 8616
rect 20031 8588 20076 8616
rect 18647 8585 18659 8588
rect 18601 8579 18659 8585
rect 15749 8551 15807 8557
rect 15749 8517 15761 8551
rect 15795 8548 15807 8551
rect 16206 8548 16212 8560
rect 15795 8520 16212 8548
rect 15795 8517 15807 8520
rect 15749 8511 15807 8517
rect 16206 8508 16212 8520
rect 16264 8508 16270 8560
rect 19628 8548 19656 8588
rect 20070 8576 20076 8588
rect 20128 8576 20134 8628
rect 20530 8616 20536 8628
rect 20491 8588 20536 8616
rect 20530 8576 20536 8588
rect 20588 8576 20594 8628
rect 20548 8548 20576 8576
rect 20714 8548 20720 8560
rect 19628 8520 20720 8548
rect 20714 8508 20720 8520
rect 20772 8508 20778 8560
rect 2777 8483 2835 8489
rect 2777 8449 2789 8483
rect 2823 8480 2835 8483
rect 8202 8480 8208 8492
rect 2823 8452 8208 8480
rect 2823 8449 2835 8452
rect 2777 8443 2835 8449
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 12986 8440 12992 8492
rect 13044 8480 13050 8492
rect 13541 8483 13599 8489
rect 13541 8480 13553 8483
rect 13044 8452 13553 8480
rect 13044 8440 13050 8452
rect 13541 8449 13553 8452
rect 13587 8449 13599 8483
rect 13541 8443 13599 8449
rect 13814 8440 13820 8492
rect 13872 8480 13878 8492
rect 14461 8483 14519 8489
rect 14461 8480 14473 8483
rect 13872 8452 14473 8480
rect 13872 8440 13878 8452
rect 14461 8449 14473 8452
rect 14507 8449 14519 8483
rect 22278 8480 22284 8492
rect 14461 8443 14519 8449
rect 14568 8452 22284 8480
rect 2501 8415 2559 8421
rect 2501 8381 2513 8415
rect 2547 8412 2559 8415
rect 6822 8412 6828 8424
rect 2547 8384 4384 8412
rect 6783 8384 6828 8412
rect 2547 8381 2559 8384
rect 2501 8375 2559 8381
rect 4356 8353 4384 8384
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 7098 8412 7104 8424
rect 7059 8384 7104 8412
rect 7098 8372 7104 8384
rect 7156 8372 7162 8424
rect 9677 8415 9735 8421
rect 9677 8381 9689 8415
rect 9723 8412 9735 8415
rect 9766 8412 9772 8424
rect 9723 8384 9772 8412
rect 9723 8381 9735 8384
rect 9677 8375 9735 8381
rect 9766 8372 9772 8384
rect 9824 8412 9830 8424
rect 10134 8412 10140 8424
rect 9824 8384 10140 8412
rect 9824 8372 9830 8384
rect 10134 8372 10140 8384
rect 10192 8372 10198 8424
rect 13998 8412 14004 8424
rect 13959 8384 14004 8412
rect 13998 8372 14004 8384
rect 14056 8372 14062 8424
rect 14090 8372 14096 8424
rect 14148 8412 14154 8424
rect 14185 8415 14243 8421
rect 14185 8412 14197 8415
rect 14148 8384 14197 8412
rect 14148 8372 14154 8384
rect 14185 8381 14197 8384
rect 14231 8381 14243 8415
rect 14185 8375 14243 8381
rect 4341 8347 4399 8353
rect 4341 8313 4353 8347
rect 4387 8344 4399 8347
rect 4614 8344 4620 8356
rect 4387 8316 4620 8344
rect 4387 8313 4399 8316
rect 4341 8307 4399 8313
rect 4614 8304 4620 8316
rect 4672 8344 4678 8356
rect 5442 8344 5448 8356
rect 4672 8316 5448 8344
rect 4672 8304 4678 8316
rect 5442 8304 5448 8316
rect 5500 8304 5506 8356
rect 14476 8344 14504 8443
rect 14568 8421 14596 8452
rect 22278 8440 22284 8452
rect 22336 8440 22342 8492
rect 14553 8415 14611 8421
rect 14553 8381 14565 8415
rect 14599 8381 14611 8415
rect 14553 8375 14611 8381
rect 15565 8415 15623 8421
rect 15565 8381 15577 8415
rect 15611 8381 15623 8415
rect 15565 8375 15623 8381
rect 18601 8415 18659 8421
rect 18601 8381 18613 8415
rect 18647 8412 18659 8415
rect 18693 8415 18751 8421
rect 18693 8412 18705 8415
rect 18647 8384 18705 8412
rect 18647 8381 18659 8384
rect 18601 8375 18659 8381
rect 18693 8381 18705 8384
rect 18739 8381 18751 8415
rect 18693 8375 18751 8381
rect 18969 8415 19027 8421
rect 18969 8381 18981 8415
rect 19015 8412 19027 8415
rect 19334 8412 19340 8424
rect 19015 8384 19340 8412
rect 19015 8381 19027 8384
rect 18969 8375 19027 8381
rect 15580 8344 15608 8375
rect 19334 8372 19340 8384
rect 19392 8372 19398 8424
rect 14476 8316 15608 8344
rect 3878 8276 3884 8288
rect 3839 8248 3884 8276
rect 3878 8236 3884 8248
rect 3936 8236 3942 8288
rect 4062 8236 4068 8288
rect 4120 8276 4126 8288
rect 6546 8276 6552 8288
rect 4120 8248 6552 8276
rect 4120 8236 4126 8248
rect 6546 8236 6552 8248
rect 6604 8236 6610 8288
rect 6822 8236 6828 8288
rect 6880 8276 6886 8288
rect 8202 8276 8208 8288
rect 6880 8248 8208 8276
rect 6880 8236 6886 8248
rect 8202 8236 8208 8248
rect 8260 8276 8266 8288
rect 8573 8279 8631 8285
rect 8573 8276 8585 8279
rect 8260 8248 8585 8276
rect 8260 8236 8266 8248
rect 8573 8245 8585 8248
rect 8619 8245 8631 8279
rect 9858 8276 9864 8288
rect 9819 8248 9864 8276
rect 8573 8239 8631 8245
rect 9858 8236 9864 8248
rect 9916 8236 9922 8288
rect 12894 8236 12900 8288
rect 12952 8276 12958 8288
rect 13906 8276 13912 8288
rect 12952 8248 13912 8276
rect 12952 8236 12958 8248
rect 13906 8236 13912 8248
rect 13964 8236 13970 8288
rect 1104 8186 24656 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 24656 8186
rect 1104 8112 24656 8134
rect 8294 8032 8300 8084
rect 8352 8072 8358 8084
rect 9953 8075 10011 8081
rect 9953 8072 9965 8075
rect 8352 8044 9965 8072
rect 8352 8032 8358 8044
rect 9953 8041 9965 8044
rect 9999 8041 10011 8075
rect 14093 8075 14151 8081
rect 9953 8035 10011 8041
rect 12452 8044 13400 8072
rect 7098 7964 7104 8016
rect 7156 8004 7162 8016
rect 7377 8007 7435 8013
rect 7377 8004 7389 8007
rect 7156 7976 7389 8004
rect 7156 7964 7162 7976
rect 7377 7973 7389 7976
rect 7423 7973 7435 8007
rect 9674 8004 9680 8016
rect 7377 7967 7435 7973
rect 8404 7976 8800 8004
rect 9635 7976 9680 8004
rect 8404 7945 8432 7976
rect 8021 7939 8079 7945
rect 8021 7905 8033 7939
rect 8067 7936 8079 7939
rect 8389 7939 8447 7945
rect 8067 7908 8340 7936
rect 8067 7905 8079 7908
rect 8021 7899 8079 7905
rect 7098 7828 7104 7880
rect 7156 7868 7162 7880
rect 7837 7871 7895 7877
rect 7837 7868 7849 7871
rect 7156 7840 7849 7868
rect 7156 7828 7162 7840
rect 7837 7837 7849 7840
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 8312 7800 8340 7908
rect 8389 7905 8401 7939
rect 8435 7905 8447 7939
rect 8389 7899 8447 7905
rect 8478 7896 8484 7948
rect 8536 7936 8542 7948
rect 8772 7945 8800 7976
rect 9674 7964 9680 7976
rect 9732 8004 9738 8016
rect 11793 8007 11851 8013
rect 11793 8004 11805 8007
rect 9732 7976 11805 8004
rect 9732 7964 9738 7976
rect 11793 7973 11805 7976
rect 11839 7973 11851 8007
rect 11793 7967 11851 7973
rect 8757 7939 8815 7945
rect 8536 7908 8581 7936
rect 8536 7896 8542 7908
rect 8757 7905 8769 7939
rect 8803 7936 8815 7939
rect 9766 7936 9772 7948
rect 8803 7908 9772 7936
rect 8803 7905 8815 7908
rect 8757 7899 8815 7905
rect 9766 7896 9772 7908
rect 9824 7896 9830 7948
rect 9861 7939 9919 7945
rect 9861 7905 9873 7939
rect 9907 7905 9919 7939
rect 9861 7899 9919 7905
rect 8570 7828 8576 7880
rect 8628 7868 8634 7880
rect 9876 7868 9904 7899
rect 8628 7840 9904 7868
rect 11808 7868 11836 7967
rect 11977 7939 12035 7945
rect 11977 7905 11989 7939
rect 12023 7936 12035 7939
rect 12158 7936 12164 7948
rect 12023 7908 12164 7936
rect 12023 7905 12035 7908
rect 11977 7899 12035 7905
rect 12158 7896 12164 7908
rect 12216 7896 12222 7948
rect 12345 7939 12403 7945
rect 12345 7905 12357 7939
rect 12391 7936 12403 7939
rect 12452 7936 12480 8044
rect 13372 7945 13400 8044
rect 14093 8041 14105 8075
rect 14139 8072 14151 8075
rect 17862 8072 17868 8084
rect 14139 8044 17868 8072
rect 14139 8041 14151 8044
rect 14093 8035 14151 8041
rect 12391 7908 12480 7936
rect 13357 7939 13415 7945
rect 12391 7905 12403 7908
rect 12345 7899 12403 7905
rect 13357 7905 13369 7939
rect 13403 7905 13415 7939
rect 13357 7899 13415 7905
rect 13449 7939 13507 7945
rect 13449 7905 13461 7939
rect 13495 7936 13507 7939
rect 14108 7936 14136 8035
rect 17862 8032 17868 8044
rect 17920 8032 17926 8084
rect 15470 7936 15476 7948
rect 13495 7908 14136 7936
rect 15431 7908 15476 7936
rect 13495 7905 13507 7908
rect 13449 7899 13507 7905
rect 15470 7896 15476 7908
rect 15528 7896 15534 7948
rect 15562 7896 15568 7948
rect 15620 7936 15626 7948
rect 15620 7908 15665 7936
rect 15620 7896 15626 7908
rect 12894 7868 12900 7880
rect 11808 7840 12900 7868
rect 8628 7828 8634 7840
rect 12894 7828 12900 7840
rect 12952 7828 12958 7880
rect 16025 7871 16083 7877
rect 16025 7868 16037 7871
rect 13004 7840 16037 7868
rect 9030 7800 9036 7812
rect 8312 7772 9036 7800
rect 9030 7760 9036 7772
rect 9088 7760 9094 7812
rect 9674 7760 9680 7812
rect 9732 7800 9738 7812
rect 13004 7800 13032 7840
rect 16025 7837 16037 7840
rect 16071 7837 16083 7871
rect 16025 7831 16083 7837
rect 9732 7772 13032 7800
rect 13081 7803 13139 7809
rect 9732 7760 9738 7772
rect 13081 7769 13093 7803
rect 13127 7800 13139 7803
rect 13173 7803 13231 7809
rect 13173 7800 13185 7803
rect 13127 7772 13185 7800
rect 13127 7769 13139 7772
rect 13081 7763 13139 7769
rect 13173 7769 13185 7772
rect 13219 7800 13231 7803
rect 13219 7772 15148 7800
rect 13219 7769 13231 7772
rect 13173 7763 13231 7769
rect 7006 7692 7012 7744
rect 7064 7732 7070 7744
rect 13096 7732 13124 7763
rect 13630 7732 13636 7744
rect 7064 7704 13124 7732
rect 13591 7704 13636 7732
rect 7064 7692 7070 7704
rect 13630 7692 13636 7704
rect 13688 7692 13694 7744
rect 15120 7741 15148 7772
rect 15105 7735 15163 7741
rect 15105 7701 15117 7735
rect 15151 7732 15163 7735
rect 15289 7735 15347 7741
rect 15289 7732 15301 7735
rect 15151 7704 15301 7732
rect 15151 7701 15163 7704
rect 15105 7695 15163 7701
rect 15289 7701 15301 7704
rect 15335 7701 15347 7735
rect 15289 7695 15347 7701
rect 1104 7642 24656 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 24656 7642
rect 1104 7568 24656 7590
rect 8570 7528 8576 7540
rect 8531 7500 8576 7528
rect 8570 7488 8576 7500
rect 8628 7488 8634 7540
rect 14366 7488 14372 7540
rect 14424 7528 14430 7540
rect 15102 7528 15108 7540
rect 14424 7500 15108 7528
rect 14424 7488 14430 7500
rect 15102 7488 15108 7500
rect 15160 7528 15166 7540
rect 15289 7531 15347 7537
rect 15289 7528 15301 7531
rect 15160 7500 15301 7528
rect 15160 7488 15166 7500
rect 15289 7497 15301 7500
rect 15335 7497 15347 7531
rect 15289 7491 15347 7497
rect 15378 7488 15384 7540
rect 15436 7528 15442 7540
rect 15473 7531 15531 7537
rect 15473 7528 15485 7531
rect 15436 7500 15485 7528
rect 15436 7488 15442 7500
rect 15473 7497 15485 7500
rect 15519 7497 15531 7531
rect 20714 7528 20720 7540
rect 20675 7500 20720 7528
rect 15473 7491 15531 7497
rect 20714 7488 20720 7500
rect 20772 7488 20778 7540
rect 22278 7528 22284 7540
rect 22239 7500 22284 7528
rect 22278 7488 22284 7500
rect 22336 7488 22342 7540
rect 2777 7395 2835 7401
rect 2777 7361 2789 7395
rect 2823 7392 2835 7395
rect 9766 7392 9772 7404
rect 2823 7364 9772 7392
rect 2823 7361 2835 7364
rect 2777 7355 2835 7361
rect 9766 7352 9772 7364
rect 9824 7352 9830 7404
rect 12802 7352 12808 7404
rect 12860 7392 12866 7404
rect 13725 7395 13783 7401
rect 13725 7392 13737 7395
rect 12860 7364 13737 7392
rect 12860 7352 12866 7364
rect 13725 7361 13737 7364
rect 13771 7392 13783 7395
rect 15396 7392 15424 7488
rect 19334 7392 19340 7404
rect 13771 7364 15424 7392
rect 19295 7364 19340 7392
rect 13771 7361 13783 7364
rect 13725 7355 13783 7361
rect 19334 7352 19340 7364
rect 19392 7352 19398 7404
rect 20732 7392 20760 7488
rect 20901 7395 20959 7401
rect 20901 7392 20913 7395
rect 20732 7364 20913 7392
rect 20901 7361 20913 7364
rect 20947 7361 20959 7395
rect 20901 7355 20959 7361
rect 2498 7324 2504 7336
rect 2459 7296 2504 7324
rect 2498 7284 2504 7296
rect 2556 7284 2562 7336
rect 6822 7284 6828 7336
rect 6880 7324 6886 7336
rect 7009 7327 7067 7333
rect 7009 7324 7021 7327
rect 6880 7296 7021 7324
rect 6880 7284 6886 7296
rect 7009 7293 7021 7296
rect 7055 7293 7067 7327
rect 7282 7324 7288 7336
rect 7243 7296 7288 7324
rect 7009 7287 7067 7293
rect 7282 7284 7288 7296
rect 7340 7284 7346 7336
rect 14001 7327 14059 7333
rect 14001 7293 14013 7327
rect 14047 7324 14059 7327
rect 15286 7324 15292 7336
rect 14047 7296 15292 7324
rect 14047 7293 14059 7296
rect 14001 7287 14059 7293
rect 15286 7284 15292 7296
rect 15344 7284 15350 7336
rect 21177 7327 21235 7333
rect 21177 7293 21189 7327
rect 21223 7324 21235 7327
rect 22278 7324 22284 7336
rect 21223 7296 22284 7324
rect 21223 7293 21235 7296
rect 21177 7287 21235 7293
rect 22278 7284 22284 7296
rect 22336 7284 22342 7336
rect 3878 7188 3884 7200
rect 3839 7160 3884 7188
rect 3878 7148 3884 7160
rect 3936 7148 3942 7200
rect 4341 7191 4399 7197
rect 4341 7157 4353 7191
rect 4387 7188 4399 7191
rect 4614 7188 4620 7200
rect 4387 7160 4620 7188
rect 4387 7157 4399 7160
rect 4341 7151 4399 7157
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 8202 7148 8208 7200
rect 8260 7188 8266 7200
rect 8757 7191 8815 7197
rect 8757 7188 8769 7191
rect 8260 7160 8769 7188
rect 8260 7148 8266 7160
rect 8757 7157 8769 7160
rect 8803 7188 8815 7191
rect 10962 7188 10968 7200
rect 8803 7160 10968 7188
rect 8803 7157 8815 7160
rect 8757 7151 8815 7157
rect 10962 7148 10968 7160
rect 11020 7148 11026 7200
rect 19978 7188 19984 7200
rect 19939 7160 19984 7188
rect 19978 7148 19984 7160
rect 20036 7148 20042 7200
rect 1104 7098 24656 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 24656 7098
rect 1104 7024 24656 7046
rect 15102 6984 15108 6996
rect 15063 6956 15108 6984
rect 15102 6944 15108 6956
rect 15160 6984 15166 6996
rect 20714 6984 20720 6996
rect 15160 6956 15976 6984
rect 20675 6956 20720 6984
rect 15160 6944 15166 6956
rect 7098 6916 7104 6928
rect 7059 6888 7104 6916
rect 7098 6876 7104 6888
rect 7156 6876 7162 6928
rect 15286 6916 15292 6928
rect 15247 6888 15292 6916
rect 15286 6876 15292 6888
rect 15344 6876 15350 6928
rect 4062 6808 4068 6860
rect 4120 6848 4126 6860
rect 5166 6848 5172 6860
rect 4120 6820 5172 6848
rect 4120 6808 4126 6820
rect 5166 6808 5172 6820
rect 5224 6808 5230 6860
rect 10962 6808 10968 6860
rect 11020 6848 11026 6860
rect 11149 6851 11207 6857
rect 11149 6848 11161 6851
rect 11020 6820 11161 6848
rect 11020 6808 11026 6820
rect 11149 6817 11161 6820
rect 11195 6848 11207 6851
rect 12986 6848 12992 6860
rect 11195 6820 12992 6848
rect 11195 6817 11207 6820
rect 11149 6811 11207 6817
rect 12986 6808 12992 6820
rect 13044 6808 13050 6860
rect 13817 6851 13875 6857
rect 13817 6817 13829 6851
rect 13863 6848 13875 6851
rect 13906 6848 13912 6860
rect 13863 6820 13912 6848
rect 13863 6817 13875 6820
rect 13817 6811 13875 6817
rect 13906 6808 13912 6820
rect 13964 6808 13970 6860
rect 14001 6851 14059 6857
rect 14001 6817 14013 6851
rect 14047 6817 14059 6851
rect 14001 6811 14059 6817
rect 14369 6851 14427 6857
rect 14369 6817 14381 6851
rect 14415 6848 14427 6851
rect 15470 6848 15476 6860
rect 14415 6820 15476 6848
rect 14415 6817 14427 6820
rect 14369 6811 14427 6817
rect 5442 6780 5448 6792
rect 5355 6752 5448 6780
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 5718 6780 5724 6792
rect 5679 6752 5724 6780
rect 5718 6740 5724 6752
rect 5776 6740 5782 6792
rect 11422 6780 11428 6792
rect 11383 6752 11428 6780
rect 11422 6740 11428 6752
rect 11480 6740 11486 6792
rect 12158 6740 12164 6792
rect 12216 6780 12222 6792
rect 12529 6783 12587 6789
rect 12529 6780 12541 6783
rect 12216 6752 12541 6780
rect 12216 6740 12222 6752
rect 12529 6749 12541 6752
rect 12575 6749 12587 6783
rect 14016 6780 14044 6811
rect 15470 6808 15476 6820
rect 15528 6808 15534 6860
rect 15948 6857 15976 6956
rect 20714 6944 20720 6956
rect 20772 6944 20778 6996
rect 22278 6984 22284 6996
rect 22239 6956 22284 6984
rect 22278 6944 22284 6956
rect 22336 6944 22342 6996
rect 15933 6851 15991 6857
rect 15933 6817 15945 6851
rect 15979 6817 15991 6851
rect 16298 6848 16304 6860
rect 16259 6820 16304 6848
rect 15933 6811 15991 6817
rect 16298 6808 16304 6820
rect 16356 6808 16362 6860
rect 19245 6851 19303 6857
rect 19245 6817 19257 6851
rect 19291 6848 19303 6851
rect 19978 6848 19984 6860
rect 19291 6820 19984 6848
rect 19291 6817 19303 6820
rect 19245 6811 19303 6817
rect 19978 6808 19984 6820
rect 20036 6848 20042 6860
rect 21177 6851 21235 6857
rect 21177 6848 21189 6851
rect 20036 6820 21189 6848
rect 20036 6808 20042 6820
rect 21177 6817 21189 6820
rect 21223 6817 21235 6851
rect 21177 6811 21235 6817
rect 15654 6780 15660 6792
rect 14016 6752 15660 6780
rect 12529 6743 12587 6749
rect 15654 6740 15660 6752
rect 15712 6740 15718 6792
rect 15749 6783 15807 6789
rect 15749 6749 15761 6783
rect 15795 6749 15807 6783
rect 16206 6780 16212 6792
rect 16167 6752 16212 6780
rect 15749 6743 15807 6749
rect 5460 6644 5488 6740
rect 15102 6672 15108 6724
rect 15160 6712 15166 6724
rect 15764 6712 15792 6743
rect 16206 6740 16212 6752
rect 16264 6740 16270 6792
rect 20714 6740 20720 6792
rect 20772 6780 20778 6792
rect 20901 6783 20959 6789
rect 20901 6780 20913 6783
rect 20772 6752 20913 6780
rect 20772 6740 20778 6752
rect 20901 6749 20913 6752
rect 20947 6749 20959 6783
rect 20901 6743 20959 6749
rect 15160 6684 15792 6712
rect 15160 6672 15166 6684
rect 7285 6647 7343 6653
rect 7285 6644 7297 6647
rect 5460 6616 7297 6644
rect 7285 6613 7297 6616
rect 7331 6644 7343 6647
rect 11330 6644 11336 6656
rect 7331 6616 11336 6644
rect 7331 6613 7343 6616
rect 7285 6607 7343 6613
rect 11330 6604 11336 6616
rect 11388 6644 11394 6656
rect 12802 6644 12808 6656
rect 11388 6616 12808 6644
rect 11388 6604 11394 6616
rect 12802 6604 12808 6616
rect 12860 6604 12866 6656
rect 12986 6644 12992 6656
rect 12947 6616 12992 6644
rect 12986 6604 12992 6616
rect 13044 6604 13050 6656
rect 19886 6644 19892 6656
rect 19847 6616 19892 6644
rect 19886 6604 19892 6616
rect 19944 6604 19950 6656
rect 1104 6554 24656 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 24656 6554
rect 1104 6480 24656 6502
rect 4341 6443 4399 6449
rect 4341 6409 4353 6443
rect 4387 6440 4399 6443
rect 9674 6440 9680 6452
rect 4387 6412 9680 6440
rect 4387 6409 4399 6412
rect 4341 6403 4399 6409
rect 2498 6236 2504 6248
rect 2459 6208 2504 6236
rect 2498 6196 2504 6208
rect 2556 6196 2562 6248
rect 2777 6239 2835 6245
rect 2777 6205 2789 6239
rect 2823 6236 2835 6239
rect 4540 6236 4568 6412
rect 9674 6400 9680 6412
rect 9732 6400 9738 6452
rect 16298 6400 16304 6452
rect 16356 6440 16362 6452
rect 21637 6443 21695 6449
rect 21637 6440 21649 6443
rect 16356 6412 21649 6440
rect 16356 6400 16362 6412
rect 21637 6409 21649 6412
rect 21683 6409 21695 6443
rect 21637 6403 21695 6409
rect 7282 6264 7288 6316
rect 7340 6304 7346 6316
rect 7837 6307 7895 6313
rect 7837 6304 7849 6307
rect 7340 6276 7849 6304
rect 7340 6264 7346 6276
rect 7837 6273 7849 6276
rect 7883 6273 7895 6307
rect 7837 6267 7895 6273
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6304 8447 6307
rect 9858 6304 9864 6316
rect 8435 6276 9864 6304
rect 8435 6273 8447 6276
rect 8389 6267 8447 6273
rect 9858 6264 9864 6276
rect 9916 6264 9922 6316
rect 20165 6307 20223 6313
rect 20165 6273 20177 6307
rect 20211 6304 20223 6307
rect 20257 6307 20315 6313
rect 20257 6304 20269 6307
rect 20211 6276 20269 6304
rect 20211 6273 20223 6276
rect 20165 6267 20223 6273
rect 20257 6273 20269 6276
rect 20303 6304 20315 6307
rect 20714 6304 20720 6316
rect 20303 6276 20720 6304
rect 20303 6273 20315 6276
rect 20257 6267 20315 6273
rect 20714 6264 20720 6276
rect 20772 6264 20778 6316
rect 2823 6208 4568 6236
rect 8481 6239 8539 6245
rect 2823 6205 2835 6208
rect 2777 6199 2835 6205
rect 8481 6205 8493 6239
rect 8527 6236 8539 6239
rect 8570 6236 8576 6248
rect 8527 6208 8576 6236
rect 8527 6205 8539 6208
rect 8481 6199 8539 6205
rect 8570 6196 8576 6208
rect 8628 6196 8634 6248
rect 8846 6236 8852 6248
rect 8807 6208 8852 6236
rect 8846 6196 8852 6208
rect 8904 6196 8910 6248
rect 9030 6236 9036 6248
rect 8991 6208 9036 6236
rect 9030 6196 9036 6208
rect 9088 6196 9094 6248
rect 15102 6196 15108 6248
rect 15160 6236 15166 6248
rect 15381 6239 15439 6245
rect 15381 6236 15393 6239
rect 15160 6208 15393 6236
rect 15160 6196 15166 6208
rect 15381 6205 15393 6208
rect 15427 6205 15439 6239
rect 15381 6199 15439 6205
rect 15565 6239 15623 6245
rect 15565 6205 15577 6239
rect 15611 6236 15623 6239
rect 15654 6236 15660 6248
rect 15611 6208 15660 6236
rect 15611 6205 15623 6208
rect 15565 6199 15623 6205
rect 15654 6196 15660 6208
rect 15712 6196 15718 6248
rect 15933 6239 15991 6245
rect 15933 6205 15945 6239
rect 15979 6205 15991 6239
rect 15933 6199 15991 6205
rect 16117 6239 16175 6245
rect 16117 6205 16129 6239
rect 16163 6236 16175 6239
rect 16206 6236 16212 6248
rect 16163 6208 16212 6236
rect 16163 6205 16175 6208
rect 16117 6199 16175 6205
rect 15948 6168 15976 6199
rect 16206 6196 16212 6208
rect 16264 6196 16270 6248
rect 20533 6239 20591 6245
rect 20533 6205 20545 6239
rect 20579 6236 20591 6239
rect 20898 6236 20904 6248
rect 20579 6208 20904 6236
rect 20579 6205 20591 6208
rect 20533 6199 20591 6205
rect 20898 6196 20904 6208
rect 20956 6196 20962 6248
rect 16850 6168 16856 6180
rect 15948 6140 16856 6168
rect 16850 6128 16856 6140
rect 16908 6128 16914 6180
rect 3878 6100 3884 6112
rect 3839 6072 3884 6100
rect 3878 6060 3884 6072
rect 3936 6060 3942 6112
rect 4062 6060 4068 6112
rect 4120 6100 4126 6112
rect 4525 6103 4583 6109
rect 4525 6100 4537 6103
rect 4120 6072 4537 6100
rect 4120 6060 4126 6072
rect 4525 6069 4537 6072
rect 4571 6100 4583 6103
rect 4614 6100 4620 6112
rect 4571 6072 4620 6100
rect 4571 6069 4583 6072
rect 4525 6063 4583 6069
rect 4614 6060 4620 6072
rect 4672 6100 4678 6112
rect 5902 6100 5908 6112
rect 4672 6072 5908 6100
rect 4672 6060 4678 6072
rect 5902 6060 5908 6072
rect 5960 6060 5966 6112
rect 15197 6103 15255 6109
rect 15197 6069 15209 6103
rect 15243 6100 15255 6103
rect 15562 6100 15568 6112
rect 15243 6072 15568 6100
rect 15243 6069 15255 6072
rect 15197 6063 15255 6069
rect 15562 6060 15568 6072
rect 15620 6060 15626 6112
rect 1104 6010 24656 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 24656 6010
rect 1104 5936 24656 5958
rect 5902 5896 5908 5908
rect 5815 5868 5908 5896
rect 5902 5856 5908 5868
rect 5960 5896 5966 5908
rect 6822 5896 6828 5908
rect 5960 5868 6828 5896
rect 5960 5856 5966 5868
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 15013 5899 15071 5905
rect 15013 5865 15025 5899
rect 15059 5896 15071 5899
rect 15194 5896 15200 5908
rect 15059 5868 15200 5896
rect 15059 5865 15071 5868
rect 15013 5859 15071 5865
rect 15194 5856 15200 5868
rect 15252 5896 15258 5908
rect 15378 5896 15384 5908
rect 15252 5868 15384 5896
rect 15252 5856 15258 5868
rect 15378 5856 15384 5868
rect 15436 5856 15442 5908
rect 15654 5856 15660 5908
rect 15712 5896 15718 5908
rect 16669 5899 16727 5905
rect 16669 5896 16681 5899
rect 15712 5868 16681 5896
rect 15712 5856 15718 5868
rect 16669 5865 16681 5868
rect 16715 5865 16727 5899
rect 16669 5859 16727 5865
rect 20714 5856 20720 5908
rect 20772 5896 20778 5908
rect 21545 5899 21603 5905
rect 21545 5896 21557 5899
rect 20772 5868 21557 5896
rect 20772 5856 20778 5868
rect 21545 5865 21557 5868
rect 21591 5865 21603 5899
rect 21726 5896 21732 5908
rect 21687 5868 21732 5896
rect 21545 5859 21603 5865
rect 5718 5828 5724 5840
rect 5679 5800 5724 5828
rect 5718 5788 5724 5800
rect 5776 5788 5782 5840
rect 11422 5788 11428 5840
rect 11480 5828 11486 5840
rect 11517 5831 11575 5837
rect 11517 5828 11529 5831
rect 11480 5800 11529 5828
rect 11480 5788 11486 5800
rect 11517 5797 11529 5800
rect 11563 5797 11575 5831
rect 13998 5828 14004 5840
rect 11517 5791 11575 5797
rect 11992 5800 14004 5828
rect 9858 5720 9864 5772
rect 9916 5760 9922 5772
rect 11992 5769 12020 5800
rect 13998 5788 14004 5800
rect 14056 5828 14062 5840
rect 15102 5828 15108 5840
rect 14056 5800 15108 5828
rect 14056 5788 14062 5800
rect 15102 5788 15108 5800
rect 15160 5788 15166 5840
rect 11977 5763 12035 5769
rect 11977 5760 11989 5763
rect 9916 5732 11989 5760
rect 9916 5720 9922 5732
rect 11977 5729 11989 5732
rect 12023 5729 12035 5763
rect 12158 5760 12164 5772
rect 12119 5732 12164 5760
rect 11977 5723 12035 5729
rect 12158 5720 12164 5732
rect 12216 5720 12222 5772
rect 12526 5760 12532 5772
rect 12487 5732 12532 5760
rect 12526 5720 12532 5732
rect 12584 5720 12590 5772
rect 12713 5763 12771 5769
rect 12713 5729 12725 5763
rect 12759 5760 12771 5763
rect 15562 5760 15568 5772
rect 12759 5732 15424 5760
rect 15523 5732 15568 5760
rect 12759 5729 12771 5732
rect 12713 5723 12771 5729
rect 4062 5692 4068 5704
rect 4023 5664 4068 5692
rect 4062 5652 4068 5664
rect 4120 5652 4126 5704
rect 4341 5695 4399 5701
rect 4341 5661 4353 5695
rect 4387 5692 4399 5695
rect 5626 5692 5632 5704
rect 4387 5664 5632 5692
rect 4387 5661 4399 5664
rect 4341 5655 4399 5661
rect 5626 5652 5632 5664
rect 5684 5652 5690 5704
rect 9030 5652 9036 5704
rect 9088 5692 9094 5704
rect 12728 5692 12756 5723
rect 9088 5664 12756 5692
rect 9088 5652 9094 5664
rect 15194 5652 15200 5704
rect 15252 5692 15258 5704
rect 15289 5695 15347 5701
rect 15289 5692 15301 5695
rect 15252 5664 15301 5692
rect 15252 5652 15258 5664
rect 15289 5661 15301 5664
rect 15335 5661 15347 5695
rect 15396 5692 15424 5732
rect 15562 5720 15568 5732
rect 15620 5720 15626 5772
rect 19153 5763 19211 5769
rect 19153 5729 19165 5763
rect 19199 5760 19211 5763
rect 19886 5760 19892 5772
rect 19199 5732 19892 5760
rect 19199 5729 19211 5732
rect 19153 5723 19211 5729
rect 19886 5720 19892 5732
rect 19944 5720 19950 5772
rect 16206 5692 16212 5704
rect 15396 5664 16212 5692
rect 15289 5655 15347 5661
rect 16206 5652 16212 5664
rect 16264 5652 16270 5704
rect 21358 5652 21364 5704
rect 21416 5692 21422 5704
rect 21560 5692 21588 5859
rect 21726 5856 21732 5868
rect 21784 5856 21790 5908
rect 21744 5760 21772 5856
rect 22189 5763 22247 5769
rect 22189 5760 22201 5763
rect 21744 5732 22201 5760
rect 22189 5729 22201 5732
rect 22235 5729 22247 5763
rect 22189 5723 22247 5729
rect 21913 5695 21971 5701
rect 21913 5692 21925 5695
rect 21416 5664 21925 5692
rect 21416 5652 21422 5664
rect 21913 5661 21925 5664
rect 21959 5661 21971 5695
rect 21913 5655 21971 5661
rect 19334 5516 19340 5568
rect 19392 5556 19398 5568
rect 19797 5559 19855 5565
rect 19797 5556 19809 5559
rect 19392 5528 19809 5556
rect 19392 5516 19398 5528
rect 19797 5525 19809 5528
rect 19843 5525 19855 5559
rect 23474 5556 23480 5568
rect 23435 5528 23480 5556
rect 19797 5519 19855 5525
rect 23474 5516 23480 5528
rect 23532 5516 23538 5568
rect 1104 5466 24656 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 24656 5466
rect 1104 5392 24656 5414
rect 4062 5312 4068 5364
rect 4120 5352 4126 5364
rect 4249 5355 4307 5361
rect 4249 5352 4261 5355
rect 4120 5324 4261 5352
rect 4120 5312 4126 5324
rect 4249 5321 4261 5324
rect 4295 5321 4307 5355
rect 5626 5352 5632 5364
rect 5587 5324 5632 5352
rect 4249 5315 4307 5321
rect 5626 5312 5632 5324
rect 5684 5312 5690 5364
rect 8481 5355 8539 5361
rect 8481 5321 8493 5355
rect 8527 5352 8539 5355
rect 8846 5352 8852 5364
rect 8527 5324 8852 5352
rect 8527 5321 8539 5324
rect 8481 5315 8539 5321
rect 8846 5312 8852 5324
rect 8904 5312 8910 5364
rect 15194 5312 15200 5364
rect 15252 5352 15258 5364
rect 15289 5355 15347 5361
rect 15289 5352 15301 5355
rect 15252 5324 15301 5352
rect 15252 5312 15258 5324
rect 15289 5321 15301 5324
rect 15335 5321 15347 5355
rect 16850 5352 16856 5364
rect 16811 5324 16856 5352
rect 15289 5315 15347 5321
rect 2774 5176 2780 5228
rect 2832 5216 2838 5228
rect 2832 5188 2877 5216
rect 2832 5176 2838 5188
rect 4062 5176 4068 5228
rect 4120 5216 4126 5228
rect 5534 5216 5540 5228
rect 4120 5188 5540 5216
rect 4120 5176 4126 5188
rect 5534 5176 5540 5188
rect 5592 5176 5598 5228
rect 15304 5216 15332 5315
rect 16850 5312 16856 5324
rect 16908 5312 16914 5364
rect 20898 5352 20904 5364
rect 20859 5324 20904 5352
rect 20898 5312 20904 5324
rect 20956 5312 20962 5364
rect 21358 5352 21364 5364
rect 21319 5324 21364 5352
rect 21358 5312 21364 5324
rect 21416 5312 21422 5364
rect 15473 5219 15531 5225
rect 15473 5216 15485 5219
rect 15304 5188 15485 5216
rect 15473 5185 15485 5188
rect 15519 5185 15531 5219
rect 15473 5179 15531 5185
rect 19797 5219 19855 5225
rect 19797 5185 19809 5219
rect 19843 5216 19855 5219
rect 19886 5216 19892 5228
rect 19843 5188 19892 5216
rect 19843 5185 19855 5188
rect 19797 5179 19855 5185
rect 19886 5176 19892 5188
rect 19944 5176 19950 5228
rect 2498 5148 2504 5160
rect 2459 5120 2504 5148
rect 2498 5108 2504 5120
rect 2556 5108 2562 5160
rect 4985 5151 5043 5157
rect 4985 5117 4997 5151
rect 5031 5148 5043 5151
rect 5810 5148 5816 5160
rect 5031 5120 5816 5148
rect 5031 5117 5043 5120
rect 4985 5111 5043 5117
rect 5810 5108 5816 5120
rect 5868 5108 5874 5160
rect 6914 5148 6920 5160
rect 6875 5120 6920 5148
rect 6914 5108 6920 5120
rect 6972 5108 6978 5160
rect 7190 5148 7196 5160
rect 7151 5120 7196 5148
rect 7190 5108 7196 5120
rect 7248 5108 7254 5160
rect 15749 5151 15807 5157
rect 15749 5117 15761 5151
rect 15795 5148 15807 5151
rect 16666 5148 16672 5160
rect 15795 5120 16672 5148
rect 15795 5117 15807 5120
rect 15749 5111 15807 5117
rect 16666 5108 16672 5120
rect 16724 5108 16730 5160
rect 19521 5151 19579 5157
rect 19521 5117 19533 5151
rect 19567 5148 19579 5151
rect 20714 5148 20720 5160
rect 19567 5120 20720 5148
rect 19567 5117 19579 5120
rect 19521 5111 19579 5117
rect 20714 5108 20720 5120
rect 20772 5108 20778 5160
rect 3878 5012 3884 5024
rect 3839 4984 3884 5012
rect 3878 4972 3884 4984
rect 3936 4972 3942 5024
rect 8754 5012 8760 5024
rect 8667 4984 8760 5012
rect 8754 4972 8760 4984
rect 8812 5012 8818 5024
rect 10502 5012 10508 5024
rect 8812 4984 10508 5012
rect 8812 4972 8818 4984
rect 10502 4972 10508 4984
rect 10560 4972 10566 5024
rect 1104 4922 24656 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 24656 4922
rect 1104 4848 24656 4870
rect 6914 4768 6920 4820
rect 6972 4808 6978 4820
rect 7285 4811 7343 4817
rect 7285 4808 7297 4811
rect 6972 4780 7297 4808
rect 6972 4768 6978 4780
rect 7285 4777 7297 4780
rect 7331 4808 7343 4811
rect 8754 4808 8760 4820
rect 7331 4780 8760 4808
rect 7331 4777 7343 4780
rect 7285 4771 7343 4777
rect 8754 4768 8760 4780
rect 8812 4768 8818 4820
rect 16666 4808 16672 4820
rect 16627 4780 16672 4808
rect 16666 4768 16672 4780
rect 16724 4768 16730 4820
rect 7190 4740 7196 4752
rect 7151 4712 7196 4740
rect 7190 4700 7196 4712
rect 7248 4700 7254 4752
rect 12437 4743 12495 4749
rect 12437 4709 12449 4743
rect 12483 4740 12495 4743
rect 12526 4740 12532 4752
rect 12483 4712 12532 4740
rect 12483 4709 12495 4712
rect 12437 4703 12495 4709
rect 12526 4700 12532 4712
rect 12584 4700 12590 4752
rect 5258 4632 5264 4684
rect 5316 4672 5322 4684
rect 5537 4675 5595 4681
rect 5537 4672 5549 4675
rect 5316 4644 5549 4672
rect 5316 4632 5322 4644
rect 5537 4641 5549 4644
rect 5583 4672 5595 4675
rect 5902 4672 5908 4684
rect 5583 4644 5908 4672
rect 5583 4641 5595 4644
rect 5537 4635 5595 4641
rect 5902 4632 5908 4644
rect 5960 4632 5966 4684
rect 10502 4632 10508 4684
rect 10560 4672 10566 4684
rect 10781 4675 10839 4681
rect 10781 4672 10793 4675
rect 10560 4644 10793 4672
rect 10560 4632 10566 4644
rect 10781 4641 10793 4644
rect 10827 4672 10839 4675
rect 13265 4675 13323 4681
rect 10827 4644 12664 4672
rect 10827 4641 10839 4644
rect 10781 4635 10839 4641
rect 5810 4604 5816 4616
rect 5771 4576 5816 4604
rect 5810 4564 5816 4576
rect 5868 4564 5874 4616
rect 11054 4604 11060 4616
rect 11015 4576 11060 4604
rect 11054 4564 11060 4576
rect 11112 4564 11118 4616
rect 12636 4545 12664 4644
rect 13265 4641 13277 4675
rect 13311 4672 13323 4675
rect 15565 4675 15623 4681
rect 15565 4672 15577 4675
rect 13311 4644 15577 4672
rect 13311 4641 13323 4644
rect 13265 4635 13323 4641
rect 15565 4641 15577 4644
rect 15611 4672 15623 4675
rect 19334 4672 19340 4684
rect 15611 4644 19340 4672
rect 15611 4641 15623 4644
rect 15565 4635 15623 4641
rect 19334 4632 19340 4644
rect 19392 4632 19398 4684
rect 15289 4607 15347 4613
rect 15289 4573 15301 4607
rect 15335 4573 15347 4607
rect 15289 4567 15347 4573
rect 12621 4539 12679 4545
rect 12621 4505 12633 4539
rect 12667 4536 12679 4539
rect 12986 4536 12992 4548
rect 12667 4508 12992 4536
rect 12667 4505 12679 4508
rect 12621 4499 12679 4505
rect 12986 4496 12992 4508
rect 13044 4536 13050 4548
rect 15304 4536 15332 4567
rect 13044 4508 15332 4536
rect 13044 4496 13050 4508
rect 13170 4428 13176 4480
rect 13228 4468 13234 4480
rect 13909 4471 13967 4477
rect 13909 4468 13921 4471
rect 13228 4440 13921 4468
rect 13228 4428 13234 4440
rect 13909 4437 13921 4440
rect 13955 4437 13967 4471
rect 15304 4468 15332 4508
rect 17037 4471 17095 4477
rect 17037 4468 17049 4471
rect 15304 4440 17049 4468
rect 13909 4431 13967 4437
rect 17037 4437 17049 4440
rect 17083 4437 17095 4471
rect 17037 4431 17095 4437
rect 1104 4378 24656 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 24656 4378
rect 1104 4304 24656 4326
rect 3970 4224 3976 4276
rect 4028 4264 4034 4276
rect 4249 4267 4307 4273
rect 4249 4264 4261 4267
rect 4028 4236 4261 4264
rect 4028 4224 4034 4236
rect 4249 4233 4261 4236
rect 4295 4233 4307 4267
rect 4249 4227 4307 4233
rect 11054 4224 11060 4276
rect 11112 4264 11118 4276
rect 11149 4267 11207 4273
rect 11149 4264 11161 4267
rect 11112 4236 11161 4264
rect 11112 4224 11118 4236
rect 11149 4233 11161 4236
rect 11195 4233 11207 4267
rect 11149 4227 11207 4233
rect 2498 4128 2504 4140
rect 2411 4100 2504 4128
rect 2498 4088 2504 4100
rect 2556 4128 2562 4140
rect 3970 4128 3976 4140
rect 2556 4100 3976 4128
rect 2556 4088 2562 4100
rect 3970 4088 3976 4100
rect 4028 4088 4034 4140
rect 6825 4131 6883 4137
rect 6825 4097 6837 4131
rect 6871 4128 6883 4131
rect 9861 4131 9919 4137
rect 9861 4128 9873 4131
rect 6871 4100 9873 4128
rect 6871 4097 6883 4100
rect 6825 4091 6883 4097
rect 9861 4097 9873 4100
rect 9907 4128 9919 4131
rect 13170 4128 13176 4140
rect 9907 4100 13176 4128
rect 9907 4097 9919 4100
rect 9861 4091 9919 4097
rect 13170 4088 13176 4100
rect 13228 4088 13234 4140
rect 2777 4063 2835 4069
rect 2777 4029 2789 4063
rect 2823 4060 2835 4063
rect 2823 4032 4292 4060
rect 2823 4029 2835 4032
rect 2777 4023 2835 4029
rect 4264 3992 4292 4032
rect 5810 4020 5816 4072
rect 5868 4060 5874 4072
rect 7469 4063 7527 4069
rect 7469 4060 7481 4063
rect 5868 4032 7481 4060
rect 5868 4020 5874 4032
rect 7469 4029 7481 4032
rect 7515 4029 7527 4063
rect 7469 4023 7527 4029
rect 9585 4063 9643 4069
rect 9585 4029 9597 4063
rect 9631 4060 9643 4063
rect 11330 4060 11336 4072
rect 9631 4032 11336 4060
rect 9631 4029 9643 4032
rect 9585 4023 9643 4029
rect 11330 4020 11336 4032
rect 11388 4020 11394 4072
rect 8110 3992 8116 4004
rect 4264 3964 8116 3992
rect 8110 3952 8116 3964
rect 8168 3952 8174 4004
rect 3878 3924 3884 3936
rect 3839 3896 3884 3924
rect 3878 3884 3884 3896
rect 3936 3884 3942 3936
rect 1104 3834 24656 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 24656 3834
rect 1104 3760 24656 3782
rect 4062 3680 4068 3732
rect 4120 3720 4126 3732
rect 7098 3720 7104 3732
rect 4120 3692 7104 3720
rect 4120 3680 4126 3692
rect 7098 3680 7104 3692
rect 7156 3680 7162 3732
rect 1104 3290 24656 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 24656 3290
rect 1104 3216 24656 3238
rect 5258 3176 5264 3188
rect 5219 3148 5264 3176
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 10502 3176 10508 3188
rect 8680 3148 10508 3176
rect 3237 3043 3295 3049
rect 3237 3009 3249 3043
rect 3283 3040 3295 3043
rect 3970 3040 3976 3052
rect 3283 3012 3976 3040
rect 3283 3009 3295 3012
rect 3237 3003 3295 3009
rect 3970 3000 3976 3012
rect 4028 3000 4034 3052
rect 8680 3049 8708 3148
rect 10502 3136 10508 3148
rect 10560 3136 10566 3188
rect 8665 3043 8723 3049
rect 8665 3009 8677 3043
rect 8711 3009 8723 3043
rect 8665 3003 8723 3009
rect 8941 3043 8999 3049
rect 8941 3009 8953 3043
rect 8987 3040 8999 3043
rect 10318 3040 10324 3052
rect 8987 3012 10324 3040
rect 8987 3009 8999 3012
rect 8941 3003 8999 3009
rect 10318 3000 10324 3012
rect 10376 3000 10382 3052
rect 3513 2975 3571 2981
rect 3513 2941 3525 2975
rect 3559 2972 3571 2975
rect 5077 2975 5135 2981
rect 5077 2972 5089 2975
rect 3559 2944 5089 2972
rect 3559 2941 3571 2944
rect 3513 2935 3571 2941
rect 5077 2941 5089 2944
rect 5123 2972 5135 2975
rect 7558 2972 7564 2984
rect 5123 2944 7564 2972
rect 5123 2941 5135 2944
rect 5077 2935 5135 2941
rect 7558 2932 7564 2944
rect 7616 2932 7622 2984
rect 2774 2796 2780 2848
rect 2832 2836 2838 2848
rect 4617 2839 4675 2845
rect 4617 2836 4629 2839
rect 2832 2808 4629 2836
rect 2832 2796 2838 2808
rect 4617 2805 4629 2808
rect 4663 2805 4675 2839
rect 10042 2836 10048 2848
rect 10003 2808 10048 2836
rect 4617 2799 4675 2805
rect 10042 2796 10048 2808
rect 10100 2796 10106 2848
rect 1104 2746 24656 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 24656 2746
rect 1104 2672 24656 2694
rect 3510 2592 3516 2644
rect 3568 2632 3574 2644
rect 10042 2632 10048 2644
rect 3568 2604 10048 2632
rect 3568 2592 3574 2604
rect 10042 2592 10048 2604
rect 10100 2592 10106 2644
rect 2866 2524 2872 2576
rect 2924 2564 2930 2576
rect 4982 2564 4988 2576
rect 2924 2536 4988 2564
rect 2924 2524 2930 2536
rect 4982 2524 4988 2536
rect 5040 2524 5046 2576
rect 1104 2202 24656 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 24656 2202
rect 1104 2128 24656 2150
rect 52546 892 52552 944
rect 52604 932 52610 944
rect 53374 932 53380 944
rect 52604 904 53380 932
rect 52604 892 52610 904
rect 53374 892 53380 904
rect 53432 892 53438 944
rect 2774 416 2780 468
rect 2832 456 2838 468
rect 5350 456 5356 468
rect 2832 428 5356 456
rect 2832 416 2838 428
rect 5350 416 5356 428
rect 5408 416 5414 468
<< via1 >>
rect 4068 44140 4120 44192
rect 75552 44140 75604 44192
rect 19606 44038 19658 44090
rect 19670 44038 19722 44090
rect 19734 44038 19786 44090
rect 19798 44038 19850 44090
rect 50326 44038 50378 44090
rect 50390 44038 50442 44090
rect 50454 44038 50506 44090
rect 50518 44038 50570 44090
rect 81046 44038 81098 44090
rect 81110 44038 81162 44090
rect 81174 44038 81226 44090
rect 81238 44038 81290 44090
rect 17868 43868 17920 43920
rect 28264 43843 28316 43852
rect 15660 43775 15712 43784
rect 15660 43741 15669 43775
rect 15669 43741 15703 43775
rect 15703 43741 15712 43775
rect 15660 43732 15712 43741
rect 17040 43596 17092 43648
rect 28264 43809 28273 43843
rect 28273 43809 28307 43843
rect 28307 43809 28316 43843
rect 28264 43800 28316 43809
rect 45928 43868 45980 43920
rect 43628 43732 43680 43784
rect 44456 43775 44508 43784
rect 44456 43741 44465 43775
rect 44465 43741 44499 43775
rect 44499 43741 44508 43775
rect 44456 43732 44508 43741
rect 48780 43800 48832 43852
rect 54576 43800 54628 43852
rect 58532 43843 58584 43852
rect 58532 43809 58541 43843
rect 58541 43809 58575 43843
rect 58575 43809 58584 43843
rect 58532 43800 58584 43809
rect 59544 43843 59596 43852
rect 59544 43809 59553 43843
rect 59553 43809 59587 43843
rect 59587 43809 59596 43843
rect 59544 43800 59596 43809
rect 60004 43800 60056 43852
rect 74080 43800 74132 43852
rect 78588 43800 78640 43852
rect 78864 43800 78916 43852
rect 49608 43732 49660 43784
rect 61016 43732 61068 43784
rect 78680 43732 78732 43784
rect 81440 43800 81492 43852
rect 82360 43843 82412 43852
rect 82360 43809 82369 43843
rect 82369 43809 82403 43843
rect 82403 43809 82412 43843
rect 82360 43800 82412 43809
rect 82820 43775 82872 43784
rect 82820 43741 82829 43775
rect 82829 43741 82863 43775
rect 82863 43741 82872 43775
rect 82820 43732 82872 43741
rect 26240 43664 26292 43716
rect 48320 43664 48372 43716
rect 74264 43664 74316 43716
rect 78496 43664 78548 43716
rect 18420 43596 18472 43648
rect 44548 43596 44600 43648
rect 45652 43639 45704 43648
rect 45652 43605 45661 43639
rect 45661 43605 45695 43639
rect 45695 43605 45704 43639
rect 45652 43596 45704 43605
rect 45928 43639 45980 43648
rect 45928 43605 45937 43639
rect 45937 43605 45971 43639
rect 45971 43605 45980 43639
rect 45928 43596 45980 43605
rect 53840 43639 53892 43648
rect 53840 43605 53849 43639
rect 53849 43605 53883 43639
rect 53883 43605 53892 43639
rect 53840 43596 53892 43605
rect 59084 43596 59136 43648
rect 74080 43639 74132 43648
rect 74080 43605 74089 43639
rect 74089 43605 74123 43639
rect 74123 43605 74132 43639
rect 74080 43596 74132 43605
rect 78772 43596 78824 43648
rect 82084 43639 82136 43648
rect 82084 43605 82093 43639
rect 82093 43605 82127 43639
rect 82127 43605 82136 43639
rect 82084 43596 82136 43605
rect 4246 43494 4298 43546
rect 4310 43494 4362 43546
rect 4374 43494 4426 43546
rect 4438 43494 4490 43546
rect 34966 43494 35018 43546
rect 35030 43494 35082 43546
rect 35094 43494 35146 43546
rect 35158 43494 35210 43546
rect 65686 43494 65738 43546
rect 65750 43494 65802 43546
rect 65814 43494 65866 43546
rect 65878 43494 65930 43546
rect 96406 43494 96458 43546
rect 96470 43494 96522 43546
rect 96534 43494 96586 43546
rect 96598 43494 96650 43546
rect 18420 43392 18472 43444
rect 48320 43435 48372 43444
rect 2780 43299 2832 43308
rect 2780 43265 2789 43299
rect 2789 43265 2823 43299
rect 2823 43265 2832 43299
rect 2780 43256 2832 43265
rect 3148 43256 3200 43308
rect 8576 43256 8628 43308
rect 27160 43256 27212 43308
rect 48320 43401 48329 43435
rect 48329 43401 48363 43435
rect 48363 43401 48372 43435
rect 48320 43392 48372 43401
rect 7840 43231 7892 43240
rect 7840 43197 7849 43231
rect 7849 43197 7883 43231
rect 7883 43197 7892 43231
rect 7840 43188 7892 43197
rect 12348 43188 12400 43240
rect 15476 43231 15528 43240
rect 15476 43197 15485 43231
rect 15485 43197 15519 43231
rect 15519 43197 15528 43231
rect 15476 43188 15528 43197
rect 16672 43188 16724 43240
rect 3884 43095 3936 43104
rect 3884 43061 3893 43095
rect 3893 43061 3927 43095
rect 3927 43061 3936 43095
rect 3884 43052 3936 43061
rect 4804 43052 4856 43104
rect 8944 43095 8996 43104
rect 8944 43061 8953 43095
rect 8953 43061 8987 43095
rect 8987 43061 8996 43095
rect 8944 43052 8996 43061
rect 12532 43095 12584 43104
rect 12532 43061 12541 43095
rect 12541 43061 12575 43095
rect 12575 43061 12584 43095
rect 12532 43052 12584 43061
rect 16488 43052 16540 43104
rect 18144 43095 18196 43104
rect 18144 43061 18153 43095
rect 18153 43061 18187 43095
rect 18187 43061 18196 43095
rect 18144 43052 18196 43061
rect 20168 43052 20220 43104
rect 21180 43231 21232 43240
rect 21180 43197 21189 43231
rect 21189 43197 21223 43231
rect 21223 43197 21232 43231
rect 21180 43188 21232 43197
rect 21456 43052 21508 43104
rect 29184 43120 29236 43172
rect 22100 43052 22152 43104
rect 26700 43052 26752 43104
rect 28448 43095 28500 43104
rect 28448 43061 28457 43095
rect 28457 43061 28491 43095
rect 28491 43061 28500 43095
rect 28448 43052 28500 43061
rect 31944 43052 31996 43104
rect 32312 43052 32364 43104
rect 33232 43231 33284 43240
rect 33232 43197 33241 43231
rect 33241 43197 33275 43231
rect 33275 43197 33284 43231
rect 33232 43188 33284 43197
rect 33968 43188 34020 43240
rect 38844 43256 38896 43308
rect 40040 43256 40092 43308
rect 35256 43120 35308 43172
rect 33232 43052 33284 43104
rect 34152 43095 34204 43104
rect 34152 43061 34161 43095
rect 34161 43061 34195 43095
rect 34195 43061 34204 43095
rect 34152 43052 34204 43061
rect 48780 43231 48832 43240
rect 48780 43197 48789 43231
rect 48789 43197 48823 43231
rect 48823 43197 48832 43231
rect 48780 43188 48832 43197
rect 53840 43392 53892 43444
rect 54576 43435 54628 43444
rect 54576 43401 54585 43435
rect 54585 43401 54619 43435
rect 54619 43401 54628 43435
rect 54576 43392 54628 43401
rect 54668 43392 54720 43444
rect 53380 43256 53432 43308
rect 61108 43392 61160 43444
rect 74632 43435 74684 43444
rect 74632 43401 74641 43435
rect 74641 43401 74675 43435
rect 74675 43401 74684 43435
rect 74632 43392 74684 43401
rect 75552 43435 75604 43444
rect 75552 43401 75561 43435
rect 75561 43401 75595 43435
rect 75595 43401 75604 43435
rect 75552 43392 75604 43401
rect 46572 43120 46624 43172
rect 54668 43188 54720 43240
rect 59084 43299 59136 43308
rect 59084 43265 59093 43299
rect 59093 43265 59127 43299
rect 59127 43265 59136 43299
rect 59084 43256 59136 43265
rect 73896 43256 73948 43308
rect 78496 43256 78548 43308
rect 82360 43299 82412 43308
rect 82360 43265 82369 43299
rect 82369 43265 82403 43299
rect 82403 43265 82412 43299
rect 82360 43256 82412 43265
rect 59360 43188 59412 43240
rect 63868 43188 63920 43240
rect 66904 43231 66956 43240
rect 66904 43197 66913 43231
rect 66913 43197 66947 43231
rect 66947 43197 66956 43231
rect 66904 43188 66956 43197
rect 67364 43231 67416 43240
rect 66260 43120 66312 43172
rect 67364 43197 67373 43231
rect 67373 43197 67407 43231
rect 67407 43197 67416 43231
rect 67364 43188 67416 43197
rect 70584 43231 70636 43240
rect 70584 43197 70593 43231
rect 70593 43197 70627 43231
rect 70627 43197 70636 43231
rect 70584 43188 70636 43197
rect 74172 43231 74224 43240
rect 74172 43197 74181 43231
rect 74181 43197 74215 43231
rect 74215 43197 74224 43231
rect 74172 43188 74224 43197
rect 74540 43188 74592 43240
rect 75552 43188 75604 43240
rect 78680 43231 78732 43240
rect 78680 43197 78689 43231
rect 78689 43197 78723 43231
rect 78723 43197 78732 43231
rect 78680 43188 78732 43197
rect 78864 43231 78916 43240
rect 78864 43197 78873 43231
rect 78873 43197 78907 43231
rect 78907 43197 78916 43231
rect 78864 43188 78916 43197
rect 81992 43231 82044 43240
rect 81992 43197 82001 43231
rect 82001 43197 82035 43231
rect 82035 43197 82044 43231
rect 81992 43188 82044 43197
rect 67916 43120 67968 43172
rect 69204 43120 69256 43172
rect 73252 43120 73304 43172
rect 78772 43120 78824 43172
rect 81532 43120 81584 43172
rect 39028 43052 39080 43104
rect 40960 43095 41012 43104
rect 40960 43061 40969 43095
rect 40969 43061 41003 43095
rect 41003 43061 41012 43095
rect 40960 43052 41012 43061
rect 42616 43095 42668 43104
rect 42616 43061 42625 43095
rect 42625 43061 42659 43095
rect 42659 43061 42668 43095
rect 42616 43052 42668 43061
rect 49792 43095 49844 43104
rect 49792 43061 49801 43095
rect 49801 43061 49835 43095
rect 49835 43061 49844 43095
rect 49792 43052 49844 43061
rect 52276 43095 52328 43104
rect 52276 43061 52285 43095
rect 52285 43061 52319 43095
rect 52319 43061 52328 43095
rect 52276 43052 52328 43061
rect 58440 43052 58492 43104
rect 59912 43052 59964 43104
rect 63776 43095 63828 43104
rect 63776 43061 63785 43095
rect 63785 43061 63819 43095
rect 63819 43061 63828 43095
rect 63776 43052 63828 43061
rect 71780 43052 71832 43104
rect 75920 43095 75972 43104
rect 75920 43061 75929 43095
rect 75929 43061 75963 43095
rect 75963 43061 75972 43095
rect 75920 43052 75972 43061
rect 83832 43095 83884 43104
rect 83832 43061 83841 43095
rect 83841 43061 83875 43095
rect 83875 43061 83884 43095
rect 83832 43052 83884 43061
rect 19606 42950 19658 43002
rect 19670 42950 19722 43002
rect 19734 42950 19786 43002
rect 19798 42950 19850 43002
rect 50326 42950 50378 43002
rect 50390 42950 50442 43002
rect 50454 42950 50506 43002
rect 50518 42950 50570 43002
rect 81046 42950 81098 43002
rect 81110 42950 81162 43002
rect 81174 42950 81226 43002
rect 81238 42950 81290 43002
rect 3516 42848 3568 42900
rect 7564 42848 7616 42900
rect 12348 42891 12400 42900
rect 12348 42857 12357 42891
rect 12357 42857 12391 42891
rect 12391 42857 12400 42891
rect 12348 42848 12400 42857
rect 21180 42848 21232 42900
rect 26056 42848 26108 42900
rect 28264 42891 28316 42900
rect 28264 42857 28273 42891
rect 28273 42857 28307 42891
rect 28307 42857 28316 42891
rect 28264 42848 28316 42857
rect 29368 42848 29420 42900
rect 2688 42755 2740 42764
rect 2688 42721 2697 42755
rect 2697 42721 2731 42755
rect 2731 42721 2740 42755
rect 2688 42712 2740 42721
rect 23848 42780 23900 42832
rect 4068 42712 4120 42764
rect 8116 42755 8168 42764
rect 8116 42721 8125 42755
rect 8125 42721 8159 42755
rect 8159 42721 8168 42755
rect 8116 42712 8168 42721
rect 2688 42576 2740 42628
rect 2780 42508 2832 42560
rect 3056 42508 3108 42560
rect 6552 42508 6604 42560
rect 6920 42508 6972 42560
rect 8024 42576 8076 42628
rect 15476 42712 15528 42764
rect 16488 42712 16540 42764
rect 17040 42755 17092 42764
rect 10784 42687 10836 42696
rect 10784 42653 10793 42687
rect 10793 42653 10827 42687
rect 10827 42653 10836 42687
rect 10784 42644 10836 42653
rect 11520 42644 11572 42696
rect 17040 42721 17049 42755
rect 17049 42721 17083 42755
rect 17083 42721 17092 42755
rect 17040 42712 17092 42721
rect 20904 42644 20956 42696
rect 21456 42644 21508 42696
rect 22008 42712 22060 42764
rect 24768 42712 24820 42764
rect 8852 42508 8904 42560
rect 10048 42551 10100 42560
rect 10048 42517 10057 42551
rect 10057 42517 10091 42551
rect 10091 42517 10100 42551
rect 10048 42508 10100 42517
rect 13728 42508 13780 42560
rect 18328 42551 18380 42560
rect 18328 42517 18337 42551
rect 18337 42517 18371 42551
rect 18371 42517 18380 42551
rect 18328 42508 18380 42517
rect 21916 42508 21968 42560
rect 22560 42508 22612 42560
rect 23112 42551 23164 42560
rect 23112 42517 23121 42551
rect 23121 42517 23155 42551
rect 23155 42517 23164 42551
rect 23112 42508 23164 42517
rect 24032 42551 24084 42560
rect 24032 42517 24041 42551
rect 24041 42517 24075 42551
rect 24075 42517 24084 42551
rect 29184 42755 29236 42764
rect 26240 42644 26292 42696
rect 26700 42687 26752 42696
rect 26700 42653 26709 42687
rect 26709 42653 26743 42687
rect 26743 42653 26752 42687
rect 26700 42644 26752 42653
rect 24032 42508 24084 42517
rect 24768 42508 24820 42560
rect 29184 42721 29193 42755
rect 29193 42721 29227 42755
rect 29227 42721 29236 42755
rect 29184 42712 29236 42721
rect 29276 42712 29328 42764
rect 33232 42780 33284 42832
rect 32220 42755 32272 42764
rect 32220 42721 32229 42755
rect 32229 42721 32263 42755
rect 32263 42721 32272 42755
rect 32220 42712 32272 42721
rect 35256 42755 35308 42764
rect 31944 42644 31996 42696
rect 32312 42644 32364 42696
rect 27896 42576 27948 42628
rect 34980 42687 35032 42696
rect 34980 42653 34989 42687
rect 34989 42653 35023 42687
rect 35023 42653 35032 42687
rect 34980 42644 35032 42653
rect 35256 42721 35265 42755
rect 35265 42721 35299 42755
rect 35299 42721 35308 42755
rect 35256 42712 35308 42721
rect 66904 42848 66956 42900
rect 78588 42848 78640 42900
rect 81440 42891 81492 42900
rect 40132 42712 40184 42764
rect 40500 42712 40552 42764
rect 44916 42712 44968 42764
rect 53840 42780 53892 42832
rect 37740 42644 37792 42696
rect 38200 42644 38252 42696
rect 46572 42755 46624 42764
rect 46572 42721 46581 42755
rect 46581 42721 46615 42755
rect 46615 42721 46624 42755
rect 46572 42712 46624 42721
rect 46020 42687 46072 42696
rect 46020 42653 46029 42687
rect 46029 42653 46063 42687
rect 46063 42653 46072 42687
rect 46020 42644 46072 42653
rect 46112 42644 46164 42696
rect 51356 42712 51408 42764
rect 53748 42712 53800 42764
rect 28448 42551 28500 42560
rect 28448 42517 28457 42551
rect 28457 42517 28491 42551
rect 28491 42517 28500 42551
rect 28448 42508 28500 42517
rect 33876 42508 33928 42560
rect 39028 42576 39080 42628
rect 43536 42576 43588 42628
rect 39304 42508 39356 42560
rect 39580 42551 39632 42560
rect 39580 42517 39589 42551
rect 39589 42517 39623 42551
rect 39623 42517 39632 42551
rect 39580 42508 39632 42517
rect 39672 42508 39724 42560
rect 50804 42576 50856 42628
rect 54668 42712 54720 42764
rect 57152 42755 57204 42764
rect 57152 42721 57161 42755
rect 57161 42721 57195 42755
rect 57195 42721 57204 42755
rect 57152 42712 57204 42721
rect 57336 42755 57388 42764
rect 57336 42721 57345 42755
rect 57345 42721 57379 42755
rect 57379 42721 57388 42755
rect 57336 42712 57388 42721
rect 58348 42712 58400 42764
rect 60004 42780 60056 42832
rect 54852 42644 54904 42696
rect 60464 42755 60516 42764
rect 60464 42721 60473 42755
rect 60473 42721 60507 42755
rect 60507 42721 60516 42755
rect 60464 42712 60516 42721
rect 61016 42712 61068 42764
rect 63776 42712 63828 42764
rect 66260 42712 66312 42764
rect 67364 42712 67416 42764
rect 69204 42755 69256 42764
rect 43720 42508 43772 42560
rect 50988 42508 51040 42560
rect 58440 42576 58492 42628
rect 58900 42576 58952 42628
rect 52368 42551 52420 42560
rect 52368 42517 52377 42551
rect 52377 42517 52411 42551
rect 52411 42517 52420 42551
rect 52368 42508 52420 42517
rect 53104 42508 53156 42560
rect 55680 42508 55732 42560
rect 59360 42644 59412 42696
rect 61108 42644 61160 42696
rect 59636 42576 59688 42628
rect 69204 42721 69213 42755
rect 69213 42721 69247 42755
rect 69247 42721 69256 42755
rect 69204 42712 69256 42721
rect 71228 42712 71280 42764
rect 75552 42780 75604 42832
rect 81440 42857 81449 42891
rect 81449 42857 81483 42891
rect 81483 42857 81492 42891
rect 81440 42848 81492 42857
rect 85212 42848 85264 42900
rect 73896 42755 73948 42764
rect 73896 42721 73905 42755
rect 73905 42721 73939 42755
rect 73939 42721 73948 42755
rect 73896 42712 73948 42721
rect 74632 42712 74684 42764
rect 60096 42508 60148 42560
rect 63592 42508 63644 42560
rect 64236 42508 64288 42560
rect 65524 42551 65576 42560
rect 65524 42517 65533 42551
rect 65533 42517 65567 42551
rect 65567 42517 65576 42551
rect 65524 42508 65576 42517
rect 67272 42551 67324 42560
rect 67272 42517 67281 42551
rect 67281 42517 67315 42551
rect 67315 42517 67324 42551
rect 67272 42508 67324 42517
rect 71504 42619 71556 42628
rect 71504 42585 71513 42619
rect 71513 42585 71547 42619
rect 71547 42585 71556 42619
rect 71504 42576 71556 42585
rect 71228 42551 71280 42560
rect 71228 42517 71237 42551
rect 71237 42517 71271 42551
rect 71271 42517 71280 42551
rect 71228 42508 71280 42517
rect 73252 42644 73304 42696
rect 77668 42576 77720 42628
rect 72700 42551 72752 42560
rect 72700 42517 72709 42551
rect 72709 42517 72743 42551
rect 72743 42517 72752 42551
rect 72700 42508 72752 42517
rect 73436 42508 73488 42560
rect 74080 42508 74132 42560
rect 78312 42508 78364 42560
rect 78772 42644 78824 42696
rect 81440 42712 81492 42764
rect 82820 42712 82872 42764
rect 81992 42644 82044 42696
rect 82728 42687 82780 42696
rect 82728 42653 82737 42687
rect 82737 42653 82771 42687
rect 82771 42653 82780 42687
rect 82728 42644 82780 42653
rect 79876 42508 79928 42560
rect 83004 42508 83056 42560
rect 83832 42508 83884 42560
rect 4246 42406 4298 42458
rect 4310 42406 4362 42458
rect 4374 42406 4426 42458
rect 4438 42406 4490 42458
rect 34966 42406 35018 42458
rect 35030 42406 35082 42458
rect 35094 42406 35146 42458
rect 35158 42406 35210 42458
rect 65686 42406 65738 42458
rect 65750 42406 65802 42458
rect 65814 42406 65866 42458
rect 65878 42406 65930 42458
rect 96406 42406 96458 42458
rect 96470 42406 96522 42458
rect 96534 42406 96586 42458
rect 96598 42406 96650 42458
rect 4068 42304 4120 42356
rect 3056 42211 3108 42220
rect 3056 42177 3065 42211
rect 3065 42177 3099 42211
rect 3099 42177 3108 42211
rect 3056 42168 3108 42177
rect 3700 42168 3752 42220
rect 11796 42304 11848 42356
rect 8576 42211 8628 42220
rect 8576 42177 8585 42211
rect 8585 42177 8619 42211
rect 8619 42177 8628 42211
rect 8576 42168 8628 42177
rect 8852 42211 8904 42220
rect 8852 42177 8861 42211
rect 8861 42177 8895 42211
rect 8895 42177 8904 42211
rect 8852 42168 8904 42177
rect 10048 42168 10100 42220
rect 21824 42304 21876 42356
rect 21916 42304 21968 42356
rect 38660 42304 38712 42356
rect 16672 42279 16724 42288
rect 16672 42245 16681 42279
rect 16681 42245 16715 42279
rect 16715 42245 16724 42279
rect 16672 42236 16724 42245
rect 15660 42211 15712 42220
rect 15660 42177 15669 42211
rect 15669 42177 15703 42211
rect 15703 42177 15712 42211
rect 15660 42168 15712 42177
rect 16764 42168 16816 42220
rect 18052 42168 18104 42220
rect 10784 42100 10836 42152
rect 16212 42143 16264 42152
rect 16212 42109 16221 42143
rect 16221 42109 16255 42143
rect 16255 42109 16264 42143
rect 16212 42100 16264 42109
rect 21180 42236 21232 42288
rect 21364 42236 21416 42288
rect 18420 42211 18472 42220
rect 18420 42177 18429 42211
rect 18429 42177 18463 42211
rect 18463 42177 18472 42211
rect 18420 42168 18472 42177
rect 27160 42211 27212 42220
rect 18328 42143 18380 42152
rect 18328 42109 18337 42143
rect 18337 42109 18371 42143
rect 18371 42109 18380 42143
rect 18328 42100 18380 42109
rect 16948 42032 17000 42084
rect 4804 41964 4856 42016
rect 10508 41964 10560 42016
rect 11428 42007 11480 42016
rect 11428 41973 11437 42007
rect 11437 41973 11471 42007
rect 11471 41973 11480 42007
rect 11428 41964 11480 41973
rect 16212 41964 16264 42016
rect 16764 41964 16816 42016
rect 17868 41964 17920 42016
rect 27160 42177 27169 42211
rect 27169 42177 27203 42211
rect 27203 42177 27212 42211
rect 27160 42168 27212 42177
rect 32220 42211 32272 42220
rect 32220 42177 32229 42211
rect 32229 42177 32263 42211
rect 32263 42177 32272 42211
rect 32220 42168 32272 42177
rect 32588 42211 32640 42220
rect 32588 42177 32597 42211
rect 32597 42177 32631 42211
rect 32631 42177 32640 42211
rect 32588 42168 32640 42177
rect 22560 42143 22612 42152
rect 21548 42032 21600 42084
rect 20168 41964 20220 42016
rect 21180 41964 21232 42016
rect 22560 42109 22569 42143
rect 22569 42109 22603 42143
rect 22603 42109 22612 42143
rect 22560 42100 22612 42109
rect 24032 42100 24084 42152
rect 26056 42100 26108 42152
rect 26608 42143 26660 42152
rect 26608 42109 26617 42143
rect 26617 42109 26651 42143
rect 26651 42109 26660 42143
rect 26608 42100 26660 42109
rect 26700 42143 26752 42152
rect 26700 42109 26709 42143
rect 26709 42109 26743 42143
rect 26743 42109 26752 42143
rect 26700 42100 26752 42109
rect 34152 42168 34204 42220
rect 37096 42168 37148 42220
rect 37372 42236 37424 42288
rect 39028 42304 39080 42356
rect 39120 42304 39172 42356
rect 33508 42143 33560 42152
rect 33508 42109 33517 42143
rect 33517 42109 33551 42143
rect 33551 42109 33560 42143
rect 33508 42100 33560 42109
rect 34428 42100 34480 42152
rect 37372 42143 37424 42152
rect 37372 42109 37381 42143
rect 37381 42109 37415 42143
rect 37415 42109 37424 42143
rect 37372 42100 37424 42109
rect 39396 42236 39448 42288
rect 40960 42304 41012 42356
rect 40408 42168 40460 42220
rect 41880 42236 41932 42288
rect 41972 42168 42024 42220
rect 43536 42304 43588 42356
rect 48872 42304 48924 42356
rect 53748 42347 53800 42356
rect 53748 42313 53757 42347
rect 53757 42313 53791 42347
rect 53791 42313 53800 42347
rect 53748 42304 53800 42313
rect 46112 42236 46164 42288
rect 42248 42168 42300 42220
rect 58532 42236 58584 42288
rect 59176 42236 59228 42288
rect 61200 42236 61252 42288
rect 66720 42279 66772 42288
rect 49148 42168 49200 42220
rect 63868 42211 63920 42220
rect 63868 42177 63877 42211
rect 63877 42177 63911 42211
rect 63911 42177 63920 42211
rect 63868 42168 63920 42177
rect 64420 42168 64472 42220
rect 39304 42100 39356 42152
rect 39580 42100 39632 42152
rect 39856 42100 39908 42152
rect 30748 42032 30800 42084
rect 33140 42032 33192 42084
rect 43904 42100 43956 42152
rect 44916 42100 44968 42152
rect 48320 42100 48372 42152
rect 48596 42143 48648 42152
rect 21732 41964 21784 42016
rect 22100 41964 22152 42016
rect 22836 41964 22888 42016
rect 25688 42007 25740 42016
rect 25688 41973 25697 42007
rect 25697 41973 25731 42007
rect 25731 41973 25740 42007
rect 25688 41964 25740 41973
rect 25780 41964 25832 42016
rect 26608 41964 26660 42016
rect 29368 41964 29420 42016
rect 32128 41964 32180 42016
rect 32588 41964 32640 42016
rect 34336 41964 34388 42016
rect 35532 41964 35584 42016
rect 40040 41964 40092 42016
rect 40132 41964 40184 42016
rect 40592 42007 40644 42016
rect 40592 41973 40601 42007
rect 40601 41973 40635 42007
rect 40635 41973 40644 42007
rect 40592 41964 40644 41973
rect 41880 41964 41932 42016
rect 47768 42032 47820 42084
rect 48596 42109 48605 42143
rect 48605 42109 48639 42143
rect 48639 42109 48648 42143
rect 48596 42100 48648 42109
rect 44180 41964 44232 42016
rect 45192 41964 45244 42016
rect 48504 41964 48556 42016
rect 50068 42100 50120 42152
rect 49700 42032 49752 42084
rect 49516 42007 49568 42016
rect 49516 41973 49525 42007
rect 49525 41973 49559 42007
rect 49559 41973 49568 42007
rect 49516 41964 49568 41973
rect 49608 41964 49660 42016
rect 52368 42100 52420 42152
rect 51080 41964 51132 42016
rect 54208 41964 54260 42016
rect 54484 42100 54536 42152
rect 54668 42143 54720 42152
rect 54668 42109 54677 42143
rect 54677 42109 54711 42143
rect 54711 42109 54720 42143
rect 54668 42100 54720 42109
rect 54852 42143 54904 42152
rect 54852 42109 54861 42143
rect 54861 42109 54895 42143
rect 54895 42109 54904 42143
rect 54852 42100 54904 42109
rect 55680 42143 55732 42152
rect 55680 42109 55689 42143
rect 55689 42109 55723 42143
rect 55723 42109 55732 42143
rect 55680 42100 55732 42109
rect 57152 42100 57204 42152
rect 59636 42143 59688 42152
rect 59636 42109 59645 42143
rect 59645 42109 59679 42143
rect 59679 42109 59688 42143
rect 59636 42100 59688 42109
rect 60004 42143 60056 42152
rect 60004 42109 60013 42143
rect 60013 42109 60047 42143
rect 60047 42109 60056 42143
rect 60004 42100 60056 42109
rect 60188 42143 60240 42152
rect 60188 42109 60197 42143
rect 60197 42109 60231 42143
rect 60231 42109 60240 42143
rect 60188 42100 60240 42109
rect 60648 42100 60700 42152
rect 61016 42143 61068 42152
rect 61016 42109 61025 42143
rect 61025 42109 61059 42143
rect 61059 42109 61068 42143
rect 61016 42100 61068 42109
rect 61200 42143 61252 42152
rect 61200 42109 61209 42143
rect 61209 42109 61243 42143
rect 61243 42109 61252 42143
rect 61200 42100 61252 42109
rect 64512 42143 64564 42152
rect 64512 42109 64521 42143
rect 64521 42109 64555 42143
rect 64555 42109 64564 42143
rect 64512 42100 64564 42109
rect 64880 42143 64932 42152
rect 64880 42109 64889 42143
rect 64889 42109 64923 42143
rect 64923 42109 64932 42143
rect 64880 42100 64932 42109
rect 65064 42143 65116 42152
rect 65064 42109 65073 42143
rect 65073 42109 65107 42143
rect 65107 42109 65116 42143
rect 65064 42100 65116 42109
rect 66720 42245 66729 42279
rect 66729 42245 66763 42279
rect 66763 42245 66772 42279
rect 66720 42236 66772 42245
rect 67364 42236 67416 42288
rect 72700 42236 72752 42288
rect 78588 42236 78640 42288
rect 70584 42211 70636 42220
rect 70584 42177 70593 42211
rect 70593 42177 70627 42211
rect 70627 42177 70636 42211
rect 70584 42168 70636 42177
rect 71504 42168 71556 42220
rect 73252 42211 73304 42220
rect 67272 42100 67324 42152
rect 69848 42075 69900 42084
rect 54668 41964 54720 42016
rect 55956 41964 56008 42016
rect 60096 41964 60148 42016
rect 60464 41964 60516 42016
rect 69848 42041 69857 42075
rect 69857 42041 69891 42075
rect 69891 42041 69900 42075
rect 69848 42032 69900 42041
rect 66352 41964 66404 42016
rect 69664 42007 69716 42016
rect 69664 41973 69673 42007
rect 69673 41973 69707 42007
rect 69707 41973 69716 42007
rect 71228 42100 71280 42152
rect 73252 42177 73261 42211
rect 73261 42177 73295 42211
rect 73295 42177 73304 42211
rect 73252 42168 73304 42177
rect 74356 42168 74408 42220
rect 74540 42211 74592 42220
rect 74540 42177 74549 42211
rect 74549 42177 74583 42211
rect 74583 42177 74592 42211
rect 74540 42168 74592 42177
rect 75920 42168 75972 42220
rect 82084 42304 82136 42356
rect 82360 42304 82412 42356
rect 74264 42100 74316 42152
rect 77668 42143 77720 42152
rect 77668 42109 77677 42143
rect 77677 42109 77711 42143
rect 77711 42109 77720 42143
rect 77668 42100 77720 42109
rect 78404 42100 78456 42152
rect 79876 42143 79928 42152
rect 79876 42109 79885 42143
rect 79885 42109 79919 42143
rect 79919 42109 79928 42143
rect 79876 42100 79928 42109
rect 85764 42168 85816 42220
rect 82728 42100 82780 42152
rect 83096 42143 83148 42152
rect 69664 41964 69716 41973
rect 73252 42032 73304 42084
rect 74356 41964 74408 42016
rect 76748 42007 76800 42016
rect 76748 41973 76757 42007
rect 76757 41973 76791 42007
rect 76791 41973 76800 42007
rect 76748 41964 76800 41973
rect 79968 42007 80020 42016
rect 79968 41973 79977 42007
rect 79977 41973 80011 42007
rect 80011 41973 80020 42007
rect 79968 41964 80020 41973
rect 83096 42109 83105 42143
rect 83105 42109 83139 42143
rect 83139 42109 83148 42143
rect 83096 42100 83148 42109
rect 87144 42032 87196 42084
rect 84108 41964 84160 42016
rect 19606 41862 19658 41914
rect 19670 41862 19722 41914
rect 19734 41862 19786 41914
rect 19798 41862 19850 41914
rect 50326 41862 50378 41914
rect 50390 41862 50442 41914
rect 50454 41862 50506 41914
rect 50518 41862 50570 41914
rect 81046 41862 81098 41914
rect 81110 41862 81162 41914
rect 81174 41862 81226 41914
rect 81238 41862 81290 41914
rect 7840 41760 7892 41812
rect 11520 41803 11572 41812
rect 11520 41769 11529 41803
rect 11529 41769 11563 41803
rect 11563 41769 11572 41803
rect 11520 41760 11572 41769
rect 7472 41667 7524 41676
rect 7472 41633 7481 41667
rect 7481 41633 7515 41667
rect 7515 41633 7524 41667
rect 7472 41624 7524 41633
rect 9128 41692 9180 41744
rect 12532 41760 12584 41812
rect 13728 41760 13780 41812
rect 16764 41803 16816 41812
rect 16764 41769 16773 41803
rect 16773 41769 16807 41803
rect 16807 41769 16816 41803
rect 16764 41760 16816 41769
rect 16948 41803 17000 41812
rect 16948 41769 16957 41803
rect 16957 41769 16991 41803
rect 16991 41769 17000 41803
rect 16948 41760 17000 41769
rect 7932 41624 7984 41676
rect 8116 41624 8168 41676
rect 10508 41667 10560 41676
rect 10508 41633 10517 41667
rect 10517 41633 10551 41667
rect 10551 41633 10560 41667
rect 10508 41624 10560 41633
rect 11796 41692 11848 41744
rect 27896 41803 27948 41812
rect 27896 41769 27905 41803
rect 27905 41769 27939 41803
rect 27939 41769 27948 41803
rect 27896 41760 27948 41769
rect 25780 41735 25832 41744
rect 11060 41667 11112 41676
rect 11060 41633 11069 41667
rect 11069 41633 11103 41667
rect 11103 41633 11112 41667
rect 14188 41667 14240 41676
rect 11060 41624 11112 41633
rect 14188 41633 14197 41667
rect 14197 41633 14231 41667
rect 14231 41633 14240 41667
rect 14188 41624 14240 41633
rect 16028 41667 16080 41676
rect 16028 41633 16037 41667
rect 16037 41633 16071 41667
rect 16071 41633 16080 41667
rect 16028 41624 16080 41633
rect 16488 41624 16540 41676
rect 16764 41624 16816 41676
rect 21180 41667 21232 41676
rect 6920 41599 6972 41608
rect 6920 41565 6929 41599
rect 6929 41565 6963 41599
rect 6963 41565 6972 41599
rect 6920 41556 6972 41565
rect 10324 41599 10376 41608
rect 10324 41565 10333 41599
rect 10333 41565 10367 41599
rect 10367 41565 10376 41599
rect 10324 41556 10376 41565
rect 12532 41556 12584 41608
rect 16948 41556 17000 41608
rect 5080 41488 5132 41540
rect 20904 41599 20956 41608
rect 20904 41565 20913 41599
rect 20913 41565 20947 41599
rect 20947 41565 20956 41599
rect 20904 41556 20956 41565
rect 21180 41633 21189 41667
rect 21189 41633 21223 41667
rect 21223 41633 21232 41667
rect 21180 41624 21232 41633
rect 25044 41667 25096 41676
rect 25044 41633 25053 41667
rect 25053 41633 25087 41667
rect 25087 41633 25096 41667
rect 25044 41624 25096 41633
rect 18144 41488 18196 41540
rect 2964 41420 3016 41472
rect 6920 41420 6972 41472
rect 11060 41420 11112 41472
rect 13084 41420 13136 41472
rect 14280 41463 14332 41472
rect 14280 41429 14289 41463
rect 14289 41429 14323 41463
rect 14323 41429 14332 41463
rect 14280 41420 14332 41429
rect 16488 41420 16540 41472
rect 20720 41420 20772 41472
rect 21916 41488 21968 41540
rect 25780 41701 25789 41735
rect 25789 41701 25823 41735
rect 25823 41701 25832 41735
rect 25780 41692 25832 41701
rect 25688 41624 25740 41676
rect 26700 41692 26752 41744
rect 26148 41624 26200 41676
rect 27344 41624 27396 41676
rect 27896 41624 27948 41676
rect 26332 41556 26384 41608
rect 29276 41760 29328 41812
rect 31576 41760 31628 41812
rect 35532 41803 35584 41812
rect 28172 41692 28224 41744
rect 34060 41692 34112 41744
rect 34704 41692 34756 41744
rect 35532 41769 35541 41803
rect 35541 41769 35575 41803
rect 35575 41769 35584 41803
rect 35532 41760 35584 41769
rect 38016 41760 38068 41812
rect 39396 41803 39448 41812
rect 39396 41769 39405 41803
rect 39405 41769 39439 41803
rect 39439 41769 39448 41803
rect 39396 41760 39448 41769
rect 39672 41760 39724 41812
rect 30932 41667 30984 41676
rect 30932 41633 30941 41667
rect 30941 41633 30975 41667
rect 30975 41633 30984 41667
rect 30932 41624 30984 41633
rect 32404 41624 32456 41676
rect 32680 41624 32732 41676
rect 33876 41624 33928 41676
rect 33968 41667 34020 41676
rect 33968 41633 33977 41667
rect 33977 41633 34011 41667
rect 34011 41633 34020 41667
rect 33968 41624 34020 41633
rect 34336 41667 34388 41676
rect 31760 41556 31812 41608
rect 34336 41633 34345 41667
rect 34345 41633 34379 41667
rect 34379 41633 34388 41667
rect 34336 41624 34388 41633
rect 38016 41667 38068 41676
rect 26240 41531 26292 41540
rect 26240 41497 26249 41531
rect 26249 41497 26283 41531
rect 26283 41497 26292 41531
rect 26240 41488 26292 41497
rect 27160 41488 27212 41540
rect 30748 41531 30800 41540
rect 30748 41497 30757 41531
rect 30757 41497 30791 41531
rect 30791 41497 30800 41531
rect 30748 41488 30800 41497
rect 32220 41488 32272 41540
rect 21364 41420 21416 41472
rect 22284 41463 22336 41472
rect 22284 41429 22293 41463
rect 22293 41429 22327 41463
rect 22327 41429 22336 41463
rect 22284 41420 22336 41429
rect 23112 41420 23164 41472
rect 31484 41420 31536 41472
rect 32680 41420 32732 41472
rect 32864 41488 32916 41540
rect 33692 41531 33744 41540
rect 33692 41497 33701 41531
rect 33701 41497 33735 41531
rect 33735 41497 33744 41531
rect 33692 41488 33744 41497
rect 38016 41633 38025 41667
rect 38025 41633 38059 41667
rect 38059 41633 38068 41667
rect 38016 41624 38068 41633
rect 38660 41692 38712 41744
rect 43168 41760 43220 41812
rect 40592 41692 40644 41744
rect 43628 41692 43680 41744
rect 38568 41667 38620 41676
rect 38568 41633 38577 41667
rect 38577 41633 38611 41667
rect 38611 41633 38620 41667
rect 38568 41624 38620 41633
rect 39672 41624 39724 41676
rect 42616 41624 42668 41676
rect 43536 41624 43588 41676
rect 44824 41760 44876 41812
rect 45928 41760 45980 41812
rect 48228 41760 48280 41812
rect 45652 41692 45704 41744
rect 47768 41692 47820 41744
rect 48596 41760 48648 41812
rect 44548 41667 44600 41676
rect 44548 41633 44557 41667
rect 44557 41633 44591 41667
rect 44591 41633 44600 41667
rect 44548 41624 44600 41633
rect 44824 41624 44876 41676
rect 45560 41667 45612 41676
rect 45560 41633 45569 41667
rect 45569 41633 45603 41667
rect 45603 41633 45612 41667
rect 45560 41624 45612 41633
rect 48504 41624 48556 41676
rect 51264 41760 51316 41812
rect 69664 41760 69716 41812
rect 64420 41692 64472 41744
rect 49608 41624 49660 41676
rect 49884 41667 49936 41676
rect 49884 41633 49893 41667
rect 49893 41633 49927 41667
rect 49927 41633 49936 41667
rect 49884 41624 49936 41633
rect 53104 41667 53156 41676
rect 53104 41633 53113 41667
rect 53113 41633 53147 41667
rect 53147 41633 53156 41667
rect 53104 41624 53156 41633
rect 53288 41667 53340 41676
rect 53288 41633 53297 41667
rect 53297 41633 53331 41667
rect 53331 41633 53340 41667
rect 53288 41624 53340 41633
rect 55036 41667 55088 41676
rect 55036 41633 55045 41667
rect 55045 41633 55079 41667
rect 55079 41633 55088 41667
rect 55036 41624 55088 41633
rect 55128 41667 55180 41676
rect 55128 41633 55149 41667
rect 55149 41633 55180 41667
rect 55128 41624 55180 41633
rect 37924 41599 37976 41608
rect 37924 41565 37933 41599
rect 37933 41565 37967 41599
rect 37967 41565 37976 41599
rect 37924 41556 37976 41565
rect 39028 41599 39080 41608
rect 39028 41565 39037 41599
rect 39037 41565 39071 41599
rect 39071 41565 39080 41599
rect 42340 41599 42392 41608
rect 39028 41556 39080 41565
rect 42340 41565 42349 41599
rect 42349 41565 42383 41599
rect 42383 41565 42392 41599
rect 42340 41556 42392 41565
rect 43720 41556 43772 41608
rect 45836 41556 45888 41608
rect 46020 41556 46072 41608
rect 48964 41599 49016 41608
rect 48964 41565 48973 41599
rect 48973 41565 49007 41599
rect 49007 41565 49016 41599
rect 48964 41556 49016 41565
rect 55956 41624 56008 41676
rect 57336 41624 57388 41676
rect 59176 41624 59228 41676
rect 59912 41624 59964 41676
rect 64328 41667 64380 41676
rect 64328 41633 64337 41667
rect 64337 41633 64371 41667
rect 64371 41633 64380 41667
rect 64328 41624 64380 41633
rect 64880 41692 64932 41744
rect 66352 41692 66404 41744
rect 71688 41760 71740 41812
rect 74356 41760 74408 41812
rect 69848 41692 69900 41744
rect 55864 41556 55916 41608
rect 60096 41556 60148 41608
rect 65064 41624 65116 41676
rect 67548 41624 67600 41676
rect 71780 41667 71832 41676
rect 71780 41633 71789 41667
rect 71789 41633 71823 41667
rect 71823 41633 71832 41667
rect 71780 41624 71832 41633
rect 73252 41692 73304 41744
rect 74172 41692 74224 41744
rect 73160 41624 73212 41676
rect 65432 41556 65484 41608
rect 66352 41599 66404 41608
rect 66352 41565 66361 41599
rect 66361 41565 66395 41599
rect 66395 41565 66404 41599
rect 66352 41556 66404 41565
rect 73252 41599 73304 41608
rect 73252 41565 73261 41599
rect 73261 41565 73295 41599
rect 73295 41565 73304 41599
rect 73252 41556 73304 41565
rect 73344 41556 73396 41608
rect 78680 41624 78732 41676
rect 81164 41667 81216 41676
rect 81164 41633 81173 41667
rect 81173 41633 81207 41667
rect 81207 41633 81216 41667
rect 81164 41624 81216 41633
rect 81992 41692 82044 41744
rect 80888 41556 80940 41608
rect 82360 41624 82412 41676
rect 82912 41667 82964 41676
rect 82912 41633 82921 41667
rect 82921 41633 82955 41667
rect 82955 41633 82964 41667
rect 82912 41624 82964 41633
rect 83648 41624 83700 41676
rect 84108 41624 84160 41676
rect 33508 41420 33560 41472
rect 33876 41463 33928 41472
rect 33876 41429 33885 41463
rect 33885 41429 33919 41463
rect 33919 41429 33928 41463
rect 33876 41420 33928 41429
rect 34060 41420 34112 41472
rect 38936 41420 38988 41472
rect 39120 41488 39172 41540
rect 78864 41488 78916 41540
rect 42340 41420 42392 41472
rect 43444 41420 43496 41472
rect 44548 41420 44600 41472
rect 45928 41420 45980 41472
rect 46388 41463 46440 41472
rect 46388 41429 46397 41463
rect 46397 41429 46431 41463
rect 46431 41429 46440 41463
rect 46388 41420 46440 41429
rect 46572 41463 46624 41472
rect 46572 41429 46581 41463
rect 46581 41429 46615 41463
rect 46615 41429 46624 41463
rect 46572 41420 46624 41429
rect 50160 41463 50212 41472
rect 50160 41429 50169 41463
rect 50169 41429 50203 41463
rect 50203 41429 50212 41463
rect 50160 41420 50212 41429
rect 55036 41420 55088 41472
rect 64236 41420 64288 41472
rect 66720 41420 66772 41472
rect 72608 41420 72660 41472
rect 73344 41420 73396 41472
rect 73528 41463 73580 41472
rect 73528 41429 73537 41463
rect 73537 41429 73571 41463
rect 73571 41429 73580 41463
rect 73528 41420 73580 41429
rect 83096 41463 83148 41472
rect 83096 41429 83105 41463
rect 83105 41429 83139 41463
rect 83139 41429 83148 41463
rect 83096 41420 83148 41429
rect 4246 41318 4298 41370
rect 4310 41318 4362 41370
rect 4374 41318 4426 41370
rect 4438 41318 4490 41370
rect 34966 41318 35018 41370
rect 35030 41318 35082 41370
rect 35094 41318 35146 41370
rect 35158 41318 35210 41370
rect 65686 41318 65738 41370
rect 65750 41318 65802 41370
rect 65814 41318 65866 41370
rect 65878 41318 65930 41370
rect 96406 41318 96458 41370
rect 96470 41318 96522 41370
rect 96534 41318 96586 41370
rect 96598 41318 96650 41370
rect 4804 41216 4856 41268
rect 8392 41216 8444 41268
rect 8944 41216 8996 41268
rect 14188 41148 14240 41200
rect 26056 41148 26108 41200
rect 26240 41148 26292 41200
rect 9680 41080 9732 41132
rect 26700 41080 26752 41132
rect 27804 41148 27856 41200
rect 30932 41148 30984 41200
rect 34428 41148 34480 41200
rect 26976 41080 27028 41132
rect 32128 41080 32180 41132
rect 33416 41080 33468 41132
rect 3792 41012 3844 41064
rect 8392 41055 8444 41064
rect 8392 41021 8401 41055
rect 8401 41021 8435 41055
rect 8435 41021 8444 41055
rect 8392 41012 8444 41021
rect 12992 41055 13044 41064
rect 5632 40944 5684 40996
rect 7472 40876 7524 40928
rect 12992 41021 13001 41055
rect 13001 41021 13035 41055
rect 13035 41021 13044 41055
rect 12992 41012 13044 41021
rect 13728 41012 13780 41064
rect 19340 41012 19392 41064
rect 19984 41055 20036 41064
rect 19984 41021 19993 41055
rect 19993 41021 20027 41055
rect 20027 41021 20036 41055
rect 19984 41012 20036 41021
rect 22284 41055 22336 41064
rect 14280 40944 14332 40996
rect 13636 40876 13688 40928
rect 15384 40919 15436 40928
rect 15384 40885 15393 40919
rect 15393 40885 15427 40919
rect 15427 40885 15436 40919
rect 15384 40876 15436 40885
rect 21640 40944 21692 40996
rect 22284 41021 22293 41055
rect 22293 41021 22327 41055
rect 22327 41021 22336 41055
rect 22284 41012 22336 41021
rect 24860 41012 24912 41064
rect 26148 41012 26200 41064
rect 27252 41055 27304 41064
rect 27252 41021 27261 41055
rect 27261 41021 27295 41055
rect 27295 41021 27304 41055
rect 27252 41012 27304 41021
rect 27620 41012 27672 41064
rect 27712 41012 27764 41064
rect 31484 41012 31536 41064
rect 31576 41055 31628 41064
rect 31576 41021 31585 41055
rect 31585 41021 31619 41055
rect 31619 41021 31628 41055
rect 31576 41012 31628 41021
rect 31944 41055 31996 41064
rect 31944 41021 31953 41055
rect 31953 41021 31987 41055
rect 31987 41021 31996 41055
rect 31944 41012 31996 41021
rect 32404 41055 32456 41064
rect 32404 41021 32413 41055
rect 32413 41021 32447 41055
rect 32447 41021 32456 41055
rect 32404 41012 32456 41021
rect 32496 41055 32548 41064
rect 32496 41021 32505 41055
rect 32505 41021 32539 41055
rect 32539 41021 32548 41055
rect 32496 41012 32548 41021
rect 32680 41012 32732 41064
rect 33416 40944 33468 40996
rect 34796 41012 34848 41064
rect 21456 40919 21508 40928
rect 21456 40885 21465 40919
rect 21465 40885 21499 40919
rect 21499 40885 21508 40919
rect 21456 40876 21508 40885
rect 22376 40919 22428 40928
rect 22376 40885 22385 40919
rect 22385 40885 22419 40919
rect 22419 40885 22428 40919
rect 22376 40876 22428 40885
rect 24860 40876 24912 40928
rect 25044 40876 25096 40928
rect 26148 40876 26200 40928
rect 26332 40919 26384 40928
rect 26332 40885 26341 40919
rect 26341 40885 26375 40919
rect 26375 40885 26384 40919
rect 26332 40876 26384 40885
rect 26424 40876 26476 40928
rect 27436 40876 27488 40928
rect 27620 40919 27672 40928
rect 27620 40885 27629 40919
rect 27629 40885 27663 40919
rect 27663 40885 27672 40919
rect 27620 40876 27672 40885
rect 27804 40919 27856 40928
rect 27804 40885 27813 40919
rect 27813 40885 27847 40919
rect 27847 40885 27856 40919
rect 27804 40876 27856 40885
rect 30288 40876 30340 40928
rect 31760 40876 31812 40928
rect 32404 40876 32456 40928
rect 33140 40876 33192 40928
rect 33324 40919 33376 40928
rect 33324 40885 33333 40919
rect 33333 40885 33367 40919
rect 33367 40885 33376 40919
rect 33324 40876 33376 40885
rect 33508 40919 33560 40928
rect 33508 40885 33517 40919
rect 33517 40885 33551 40919
rect 33551 40885 33560 40919
rect 33508 40876 33560 40885
rect 38752 41080 38804 41132
rect 44180 41148 44232 41200
rect 45928 41216 45980 41268
rect 48964 41216 49016 41268
rect 49056 41216 49108 41268
rect 51264 41216 51316 41268
rect 53288 41216 53340 41268
rect 50068 41191 50120 41200
rect 50068 41157 50077 41191
rect 50077 41157 50111 41191
rect 50111 41157 50120 41191
rect 55864 41216 55916 41268
rect 63776 41259 63828 41268
rect 63776 41225 63785 41259
rect 63785 41225 63819 41259
rect 63819 41225 63828 41259
rect 63776 41216 63828 41225
rect 64512 41216 64564 41268
rect 67548 41216 67600 41268
rect 71228 41216 71280 41268
rect 76748 41216 76800 41268
rect 78680 41216 78732 41268
rect 79968 41216 80020 41268
rect 80888 41259 80940 41268
rect 50068 41148 50120 41157
rect 43904 41123 43956 41132
rect 43904 41089 43913 41123
rect 43913 41089 43947 41123
rect 43947 41089 43956 41123
rect 43904 41080 43956 41089
rect 45100 41080 45152 41132
rect 37372 41012 37424 41064
rect 37648 41055 37700 41064
rect 37648 41021 37657 41055
rect 37657 41021 37691 41055
rect 37691 41021 37700 41055
rect 37648 41012 37700 41021
rect 38108 41012 38160 41064
rect 43996 41055 44048 41064
rect 43996 41021 44005 41055
rect 44005 41021 44039 41055
rect 44039 41021 44048 41055
rect 43996 41012 44048 41021
rect 44088 41012 44140 41064
rect 45192 41012 45244 41064
rect 45468 41012 45520 41064
rect 48688 41080 48740 41132
rect 49516 41080 49568 41132
rect 48504 41055 48556 41064
rect 48504 41021 48513 41055
rect 48513 41021 48547 41055
rect 48547 41021 48556 41055
rect 48504 41012 48556 41021
rect 48964 41055 49016 41064
rect 48964 41021 48973 41055
rect 48973 41021 49007 41055
rect 49007 41021 49016 41055
rect 48964 41012 49016 41021
rect 49056 41055 49108 41064
rect 49056 41021 49065 41055
rect 49065 41021 49099 41055
rect 49099 41021 49108 41055
rect 52644 41055 52696 41064
rect 49056 41012 49108 41021
rect 52644 41021 52653 41055
rect 52653 41021 52687 41055
rect 52687 41021 52696 41055
rect 52644 41012 52696 41021
rect 48320 40944 48372 40996
rect 38936 40876 38988 40928
rect 45192 40876 45244 40928
rect 45376 40876 45428 40928
rect 55036 41055 55088 41064
rect 55036 41021 55045 41055
rect 55045 41021 55079 41055
rect 55079 41021 55088 41055
rect 55036 41012 55088 41021
rect 64880 41055 64932 41064
rect 64880 41021 64889 41055
rect 64889 41021 64923 41055
rect 64923 41021 64932 41055
rect 64880 41012 64932 41021
rect 65064 40944 65116 40996
rect 49332 40876 49384 40928
rect 54576 40919 54628 40928
rect 54576 40885 54585 40919
rect 54585 40885 54619 40919
rect 54619 40885 54628 40919
rect 54576 40876 54628 40885
rect 54852 40876 54904 40928
rect 63500 40876 63552 40928
rect 64328 40876 64380 40928
rect 71688 41148 71740 41200
rect 73068 41148 73120 41200
rect 73528 41148 73580 41200
rect 73252 41012 73304 41064
rect 73436 41012 73488 41064
rect 66260 40876 66312 40928
rect 67364 40876 67416 40928
rect 73528 40944 73580 40996
rect 74724 41012 74776 41064
rect 78404 41055 78456 41064
rect 78404 41021 78413 41055
rect 78413 41021 78447 41055
rect 78447 41021 78456 41055
rect 78404 41012 78456 41021
rect 80888 41225 80897 41259
rect 80897 41225 80931 41259
rect 80931 41225 80940 41259
rect 80888 41216 80940 41225
rect 87144 41259 87196 41268
rect 87144 41225 87153 41259
rect 87153 41225 87187 41259
rect 87187 41225 87196 41259
rect 87144 41216 87196 41225
rect 81440 41148 81492 41200
rect 74908 40944 74960 40996
rect 80796 41012 80848 41064
rect 88984 41080 89036 41132
rect 83648 41012 83700 41064
rect 87604 41055 87656 41064
rect 87604 41021 87613 41055
rect 87613 41021 87647 41055
rect 87647 41021 87656 41055
rect 87604 41012 87656 41021
rect 72148 40876 72200 40928
rect 72976 40919 73028 40928
rect 72976 40885 72985 40919
rect 72985 40885 73019 40919
rect 73019 40885 73028 40919
rect 72976 40876 73028 40885
rect 73160 40876 73212 40928
rect 74816 40919 74868 40928
rect 74816 40885 74825 40919
rect 74825 40885 74859 40919
rect 74859 40885 74868 40919
rect 74816 40876 74868 40885
rect 79416 40876 79468 40928
rect 80796 40876 80848 40928
rect 82728 40876 82780 40928
rect 88524 40876 88576 40928
rect 19606 40774 19658 40826
rect 19670 40774 19722 40826
rect 19734 40774 19786 40826
rect 19798 40774 19850 40826
rect 50326 40774 50378 40826
rect 50390 40774 50442 40826
rect 50454 40774 50506 40826
rect 50518 40774 50570 40826
rect 81046 40774 81098 40826
rect 81110 40774 81162 40826
rect 81174 40774 81226 40826
rect 81238 40774 81290 40826
rect 2872 40672 2924 40724
rect 4988 40672 5040 40724
rect 5632 40579 5684 40588
rect 4804 40468 4856 40520
rect 5632 40545 5641 40579
rect 5641 40545 5675 40579
rect 5675 40545 5684 40579
rect 5632 40536 5684 40545
rect 7472 40536 7524 40588
rect 8208 40604 8260 40656
rect 12992 40672 13044 40724
rect 17868 40672 17920 40724
rect 20720 40715 20772 40724
rect 20720 40681 20729 40715
rect 20729 40681 20763 40715
rect 20763 40681 20772 40715
rect 20720 40672 20772 40681
rect 21916 40672 21968 40724
rect 24952 40672 25004 40724
rect 26424 40672 26476 40724
rect 27804 40672 27856 40724
rect 31760 40672 31812 40724
rect 26332 40604 26384 40656
rect 27528 40604 27580 40656
rect 8484 40536 8536 40588
rect 11980 40536 12032 40588
rect 12072 40579 12124 40588
rect 12072 40545 12081 40579
rect 12081 40545 12115 40579
rect 12115 40545 12124 40579
rect 12072 40536 12124 40545
rect 12716 40536 12768 40588
rect 13544 40579 13596 40588
rect 8024 40511 8076 40520
rect 8024 40477 8033 40511
rect 8033 40477 8067 40511
rect 8067 40477 8076 40511
rect 8024 40468 8076 40477
rect 10968 40468 11020 40520
rect 13544 40545 13553 40579
rect 13553 40545 13587 40579
rect 13587 40545 13596 40579
rect 13544 40536 13596 40545
rect 13728 40536 13780 40588
rect 16580 40536 16632 40588
rect 14280 40468 14332 40520
rect 16028 40468 16080 40520
rect 21916 40579 21968 40588
rect 21916 40545 21925 40579
rect 21925 40545 21959 40579
rect 21959 40545 21968 40579
rect 21916 40536 21968 40545
rect 22100 40579 22152 40588
rect 22100 40545 22109 40579
rect 22109 40545 22143 40579
rect 22143 40545 22152 40579
rect 22100 40536 22152 40545
rect 22376 40536 22428 40588
rect 21732 40468 21784 40520
rect 26516 40511 26568 40520
rect 26516 40477 26525 40511
rect 26525 40477 26559 40511
rect 26559 40477 26568 40511
rect 26516 40468 26568 40477
rect 26792 40511 26844 40520
rect 26792 40477 26801 40511
rect 26801 40477 26835 40511
rect 26835 40477 26844 40511
rect 26792 40468 26844 40477
rect 30932 40536 30984 40588
rect 32036 40604 32088 40656
rect 33692 40647 33744 40656
rect 32772 40579 32824 40588
rect 31576 40468 31628 40520
rect 31944 40468 31996 40520
rect 32772 40545 32781 40579
rect 32781 40545 32815 40579
rect 32815 40545 32824 40579
rect 32772 40536 32824 40545
rect 33692 40613 33701 40647
rect 33701 40613 33735 40647
rect 33735 40613 33744 40647
rect 33692 40604 33744 40613
rect 37648 40672 37700 40724
rect 38476 40672 38528 40724
rect 43168 40715 43220 40724
rect 43168 40681 43177 40715
rect 43177 40681 43211 40715
rect 43211 40681 43220 40715
rect 43168 40672 43220 40681
rect 43444 40672 43496 40724
rect 44180 40672 44232 40724
rect 45560 40672 45612 40724
rect 45928 40672 45980 40724
rect 82728 40672 82780 40724
rect 82912 40715 82964 40724
rect 82912 40681 82921 40715
rect 82921 40681 82955 40715
rect 82955 40681 82964 40715
rect 82912 40672 82964 40681
rect 88984 40715 89036 40724
rect 88984 40681 88993 40715
rect 88993 40681 89027 40715
rect 89027 40681 89036 40715
rect 88984 40672 89036 40681
rect 38108 40536 38160 40588
rect 42708 40536 42760 40588
rect 25044 40400 25096 40452
rect 27620 40400 27672 40452
rect 32220 40400 32272 40452
rect 34612 40468 34664 40520
rect 38016 40468 38068 40520
rect 40592 40468 40644 40520
rect 42892 40468 42944 40520
rect 43444 40468 43496 40520
rect 44180 40536 44232 40588
rect 46388 40604 46440 40656
rect 50160 40604 50212 40656
rect 54668 40647 54720 40656
rect 54668 40613 54677 40647
rect 54677 40613 54711 40647
rect 54711 40613 54720 40647
rect 54668 40604 54720 40613
rect 81348 40647 81400 40656
rect 45192 40536 45244 40588
rect 54852 40579 54904 40588
rect 54852 40545 54861 40579
rect 54861 40545 54895 40579
rect 54895 40545 54904 40579
rect 57796 40579 57848 40588
rect 54852 40536 54904 40545
rect 57796 40545 57805 40579
rect 57805 40545 57839 40579
rect 57839 40545 57848 40579
rect 57796 40536 57848 40545
rect 58808 40579 58860 40588
rect 58808 40545 58817 40579
rect 58817 40545 58851 40579
rect 58851 40545 58860 40579
rect 58808 40536 58860 40545
rect 62948 40579 63000 40588
rect 49516 40468 49568 40520
rect 49792 40511 49844 40520
rect 49792 40477 49801 40511
rect 49801 40477 49835 40511
rect 49835 40477 49844 40511
rect 49792 40468 49844 40477
rect 52644 40468 52696 40520
rect 52920 40468 52972 40520
rect 55128 40511 55180 40520
rect 55128 40477 55137 40511
rect 55137 40477 55171 40511
rect 55171 40477 55180 40511
rect 55128 40468 55180 40477
rect 62948 40545 62957 40579
rect 62957 40545 62991 40579
rect 62991 40545 63000 40579
rect 62948 40536 63000 40545
rect 63776 40536 63828 40588
rect 64328 40579 64380 40588
rect 64328 40545 64337 40579
rect 64337 40545 64371 40579
rect 64371 40545 64380 40579
rect 64328 40536 64380 40545
rect 64696 40536 64748 40588
rect 66076 40536 66128 40588
rect 66260 40536 66312 40588
rect 66352 40579 66404 40588
rect 66352 40545 66361 40579
rect 66361 40545 66395 40579
rect 66395 40545 66404 40579
rect 67364 40579 67416 40588
rect 66352 40536 66404 40545
rect 67364 40545 67373 40579
rect 67373 40545 67407 40579
rect 67407 40545 67416 40579
rect 67364 40536 67416 40545
rect 67456 40536 67508 40588
rect 67916 40579 67968 40588
rect 67916 40545 67925 40579
rect 67925 40545 67959 40579
rect 67959 40545 67968 40579
rect 67916 40536 67968 40545
rect 72976 40536 73028 40588
rect 73068 40579 73120 40588
rect 73068 40545 73077 40579
rect 73077 40545 73111 40579
rect 73111 40545 73120 40579
rect 73436 40579 73488 40588
rect 73068 40536 73120 40545
rect 73436 40545 73445 40579
rect 73445 40545 73479 40579
rect 73479 40545 73488 40579
rect 73436 40536 73488 40545
rect 74724 40579 74776 40588
rect 74724 40545 74733 40579
rect 74733 40545 74767 40579
rect 74767 40545 74776 40579
rect 74724 40536 74776 40545
rect 74908 40579 74960 40588
rect 74908 40545 74917 40579
rect 74917 40545 74951 40579
rect 74951 40545 74960 40579
rect 74908 40536 74960 40545
rect 64604 40468 64656 40520
rect 64972 40468 65024 40520
rect 71044 40468 71096 40520
rect 73160 40511 73212 40520
rect 73160 40477 73169 40511
rect 73169 40477 73203 40511
rect 73203 40477 73212 40511
rect 73528 40511 73580 40520
rect 73160 40468 73212 40477
rect 73528 40477 73537 40511
rect 73537 40477 73571 40511
rect 73571 40477 73580 40511
rect 73528 40468 73580 40477
rect 80888 40536 80940 40588
rect 81348 40613 81357 40647
rect 81357 40613 81391 40647
rect 81391 40613 81400 40647
rect 81348 40604 81400 40613
rect 81440 40536 81492 40588
rect 87604 40604 87656 40656
rect 86500 40579 86552 40588
rect 86500 40545 86509 40579
rect 86509 40545 86543 40579
rect 86543 40545 86552 40579
rect 86500 40536 86552 40545
rect 33232 40400 33284 40452
rect 33324 40400 33376 40452
rect 67272 40400 67324 40452
rect 75828 40400 75880 40452
rect 78680 40400 78732 40452
rect 83004 40468 83056 40520
rect 86224 40511 86276 40520
rect 86224 40477 86233 40511
rect 86233 40477 86267 40511
rect 86267 40477 86276 40511
rect 86224 40468 86276 40477
rect 86684 40511 86736 40520
rect 86684 40477 86693 40511
rect 86693 40477 86727 40511
rect 86727 40477 86736 40511
rect 86684 40468 86736 40477
rect 89444 40511 89496 40520
rect 89444 40477 89453 40511
rect 89453 40477 89487 40511
rect 89487 40477 89496 40511
rect 89444 40468 89496 40477
rect 5724 40375 5776 40384
rect 5724 40341 5733 40375
rect 5733 40341 5767 40375
rect 5767 40341 5776 40375
rect 5724 40332 5776 40341
rect 6368 40332 6420 40384
rect 7288 40332 7340 40384
rect 10324 40332 10376 40384
rect 10968 40332 11020 40384
rect 13728 40375 13780 40384
rect 13728 40341 13737 40375
rect 13737 40341 13771 40375
rect 13771 40341 13780 40375
rect 13728 40332 13780 40341
rect 22100 40332 22152 40384
rect 27528 40332 27580 40384
rect 27896 40375 27948 40384
rect 27896 40341 27905 40375
rect 27905 40341 27939 40375
rect 27939 40341 27948 40375
rect 27896 40332 27948 40341
rect 28264 40375 28316 40384
rect 28264 40341 28273 40375
rect 28273 40341 28307 40375
rect 28307 40341 28316 40375
rect 28264 40332 28316 40341
rect 33508 40332 33560 40384
rect 37648 40332 37700 40384
rect 39304 40375 39356 40384
rect 39304 40341 39313 40375
rect 39313 40341 39347 40375
rect 39347 40341 39356 40375
rect 39304 40332 39356 40341
rect 42892 40375 42944 40384
rect 42892 40341 42901 40375
rect 42901 40341 42935 40375
rect 42935 40341 42944 40375
rect 42892 40332 42944 40341
rect 43996 40332 44048 40384
rect 45376 40332 45428 40384
rect 48320 40332 48372 40384
rect 49700 40375 49752 40384
rect 49700 40341 49709 40375
rect 49709 40341 49743 40375
rect 49743 40341 49752 40375
rect 49700 40332 49752 40341
rect 51448 40332 51500 40384
rect 57704 40332 57756 40384
rect 59176 40332 59228 40384
rect 63592 40332 63644 40384
rect 64972 40375 65024 40384
rect 64972 40341 64981 40375
rect 64981 40341 65015 40375
rect 65015 40341 65024 40375
rect 64972 40332 65024 40341
rect 65432 40332 65484 40384
rect 66352 40332 66404 40384
rect 67364 40332 67416 40384
rect 71964 40332 72016 40384
rect 73160 40332 73212 40384
rect 80796 40332 80848 40384
rect 80888 40332 80940 40384
rect 89904 40332 89956 40384
rect 4246 40230 4298 40282
rect 4310 40230 4362 40282
rect 4374 40230 4426 40282
rect 4438 40230 4490 40282
rect 34966 40230 35018 40282
rect 35030 40230 35082 40282
rect 35094 40230 35146 40282
rect 35158 40230 35210 40282
rect 65686 40230 65738 40282
rect 65750 40230 65802 40282
rect 65814 40230 65866 40282
rect 65878 40230 65930 40282
rect 96406 40230 96458 40282
rect 96470 40230 96522 40282
rect 96534 40230 96586 40282
rect 96598 40230 96650 40282
rect 1492 40128 1544 40180
rect 9680 40128 9732 40180
rect 12440 40128 12492 40180
rect 13544 40128 13596 40180
rect 15384 40128 15436 40180
rect 23848 40128 23900 40180
rect 26792 40128 26844 40180
rect 27344 40128 27396 40180
rect 27988 40128 28040 40180
rect 31760 40128 31812 40180
rect 34704 40128 34756 40180
rect 38108 40128 38160 40180
rect 39304 40128 39356 40180
rect 3792 40103 3844 40112
rect 3792 40069 3801 40103
rect 3801 40069 3835 40103
rect 3835 40069 3844 40103
rect 3792 40060 3844 40069
rect 2780 39992 2832 40044
rect 2964 39967 3016 39976
rect 2964 39933 2973 39967
rect 2973 39933 3007 39967
rect 3007 39933 3016 39967
rect 3424 39967 3476 39976
rect 2964 39924 3016 39933
rect 3424 39933 3433 39967
rect 3433 39933 3467 39967
rect 3467 39933 3476 39967
rect 3424 39924 3476 39933
rect 5724 40060 5776 40112
rect 9128 40103 9180 40112
rect 8576 39992 8628 40044
rect 4804 39924 4856 39976
rect 3240 39856 3292 39908
rect 8208 39924 8260 39976
rect 8484 39924 8536 39976
rect 9128 40069 9137 40103
rect 9137 40069 9171 40103
rect 9171 40069 9180 40103
rect 9128 40060 9180 40069
rect 8944 39992 8996 40044
rect 12716 40060 12768 40112
rect 12808 39992 12860 40044
rect 12072 39924 12124 39976
rect 13728 40060 13780 40112
rect 26516 40060 26568 40112
rect 28264 40060 28316 40112
rect 31668 40060 31720 40112
rect 13728 39967 13780 39976
rect 13728 39933 13737 39967
rect 13737 39933 13771 39967
rect 13771 39933 13780 39967
rect 13728 39924 13780 39933
rect 13912 39967 13964 39976
rect 13912 39933 13946 39967
rect 13946 39933 13964 39967
rect 13912 39924 13964 39933
rect 12532 39856 12584 39908
rect 12624 39856 12676 39908
rect 14280 39899 14332 39908
rect 5908 39788 5960 39840
rect 7932 39788 7984 39840
rect 11980 39788 12032 39840
rect 12716 39788 12768 39840
rect 14280 39865 14289 39899
rect 14289 39865 14323 39899
rect 14323 39865 14332 39899
rect 14280 39856 14332 39865
rect 13912 39788 13964 39840
rect 15200 39967 15252 39976
rect 15200 39933 15209 39967
rect 15209 39933 15243 39967
rect 15243 39933 15252 39967
rect 15200 39924 15252 39933
rect 19340 39924 19392 39976
rect 21456 39992 21508 40044
rect 21180 39924 21232 39976
rect 25412 39967 25464 39976
rect 25412 39933 25421 39967
rect 25421 39933 25455 39967
rect 25455 39933 25464 39967
rect 25412 39924 25464 39933
rect 25780 39924 25832 39976
rect 25964 39967 26016 39976
rect 25964 39933 25973 39967
rect 25973 39933 26007 39967
rect 26007 39933 26016 39967
rect 25964 39924 26016 39933
rect 26148 39967 26200 39976
rect 26148 39933 26157 39967
rect 26157 39933 26191 39967
rect 26191 39933 26200 39967
rect 26148 39924 26200 39933
rect 27344 39924 27396 39976
rect 27896 39924 27948 39976
rect 28080 39924 28132 39976
rect 29000 39924 29052 39976
rect 32036 40060 32088 40112
rect 33876 40060 33928 40112
rect 37372 40060 37424 40112
rect 38936 40103 38988 40112
rect 38936 40069 38945 40103
rect 38945 40069 38979 40103
rect 38979 40069 38988 40103
rect 38936 40060 38988 40069
rect 40500 40060 40552 40112
rect 48228 40128 48280 40180
rect 64880 40128 64932 40180
rect 64972 40128 65024 40180
rect 32404 39967 32456 39976
rect 32404 39933 32413 39967
rect 32413 39933 32447 39967
rect 32447 39933 32456 39967
rect 32404 39924 32456 39933
rect 34428 39992 34480 40044
rect 33692 39924 33744 39976
rect 20996 39856 21048 39908
rect 31576 39899 31628 39908
rect 16028 39788 16080 39840
rect 21364 39788 21416 39840
rect 21548 39831 21600 39840
rect 21548 39797 21557 39831
rect 21557 39797 21591 39831
rect 21591 39797 21600 39831
rect 21548 39788 21600 39797
rect 30288 39788 30340 39840
rect 31576 39865 31585 39899
rect 31585 39865 31619 39899
rect 31619 39865 31628 39899
rect 31576 39856 31628 39865
rect 32312 39788 32364 39840
rect 34336 39856 34388 39908
rect 37372 39924 37424 39976
rect 37556 39924 37608 39976
rect 38660 39992 38712 40044
rect 40592 39992 40644 40044
rect 37924 39967 37976 39976
rect 37924 39933 37933 39967
rect 37933 39933 37967 39967
rect 37967 39933 37976 39967
rect 37924 39924 37976 39933
rect 38108 39924 38160 39976
rect 40408 39924 40460 39976
rect 40960 39924 41012 39976
rect 49148 40060 49200 40112
rect 43536 40035 43588 40044
rect 43536 40001 43545 40035
rect 43545 40001 43579 40035
rect 43579 40001 43588 40035
rect 43536 39992 43588 40001
rect 48320 39992 48372 40044
rect 49332 39992 49384 40044
rect 49792 40060 49844 40112
rect 77208 40128 77260 40180
rect 79876 40128 79928 40180
rect 67548 40103 67600 40112
rect 67548 40069 67557 40103
rect 67557 40069 67591 40103
rect 67591 40069 67600 40103
rect 67548 40060 67600 40069
rect 37740 39788 37792 39840
rect 38936 39788 38988 39840
rect 40316 39788 40368 39840
rect 40960 39788 41012 39840
rect 41144 39831 41196 39840
rect 41144 39797 41153 39831
rect 41153 39797 41187 39831
rect 41187 39797 41196 39831
rect 41144 39788 41196 39797
rect 43904 39924 43956 39976
rect 44180 39967 44232 39976
rect 44180 39933 44189 39967
rect 44189 39933 44223 39967
rect 44223 39933 44232 39967
rect 44180 39924 44232 39933
rect 45100 39967 45152 39976
rect 45100 39933 45109 39967
rect 45109 39933 45143 39967
rect 45143 39933 45152 39967
rect 45100 39924 45152 39933
rect 42800 39856 42852 39908
rect 49240 39924 49292 39976
rect 49332 39899 49384 39908
rect 49332 39865 49341 39899
rect 49341 39865 49375 39899
rect 49375 39865 49384 39899
rect 49332 39856 49384 39865
rect 44272 39788 44324 39840
rect 45100 39788 45152 39840
rect 49608 39788 49660 39840
rect 53104 39992 53156 40044
rect 70768 40060 70820 40112
rect 72148 40103 72200 40112
rect 72148 40069 72157 40103
rect 72157 40069 72191 40103
rect 72191 40069 72200 40103
rect 72148 40060 72200 40069
rect 80152 40060 80204 40112
rect 51816 39924 51868 39976
rect 52000 39967 52052 39976
rect 52000 39933 52009 39967
rect 52009 39933 52043 39967
rect 52043 39933 52052 39967
rect 52000 39924 52052 39933
rect 52368 39924 52420 39976
rect 53288 39924 53340 39976
rect 54576 39924 54628 39976
rect 50068 39788 50120 39840
rect 52644 39856 52696 39908
rect 52092 39788 52144 39840
rect 53380 39831 53432 39840
rect 53380 39797 53389 39831
rect 53389 39797 53423 39831
rect 53423 39797 53432 39831
rect 53380 39788 53432 39797
rect 53564 39831 53616 39840
rect 53564 39797 53573 39831
rect 53573 39797 53607 39831
rect 53607 39797 53616 39831
rect 53564 39788 53616 39797
rect 54668 39788 54720 39840
rect 58072 39924 58124 39976
rect 58624 39924 58676 39976
rect 62948 39924 63000 39976
rect 64144 39924 64196 39976
rect 58808 39856 58860 39908
rect 61200 39856 61252 39908
rect 63500 39856 63552 39908
rect 64604 39924 64656 39976
rect 66996 39967 67048 39976
rect 66996 39933 67005 39967
rect 67005 39933 67039 39967
rect 67039 39933 67048 39967
rect 66996 39924 67048 39933
rect 67916 39924 67968 39976
rect 67456 39899 67508 39908
rect 67456 39865 67465 39899
rect 67465 39865 67499 39899
rect 67499 39865 67508 39899
rect 67456 39856 67508 39865
rect 73344 39992 73396 40044
rect 74172 40035 74224 40044
rect 74172 40001 74181 40035
rect 74181 40001 74215 40035
rect 74215 40001 74224 40035
rect 74172 39992 74224 40001
rect 79416 40035 79468 40044
rect 79416 40001 79425 40035
rect 79425 40001 79459 40035
rect 79459 40001 79468 40035
rect 79416 39992 79468 40001
rect 79508 39992 79560 40044
rect 82360 40035 82412 40044
rect 71044 39967 71096 39976
rect 56784 39831 56836 39840
rect 56784 39797 56793 39831
rect 56793 39797 56827 39831
rect 56827 39797 56836 39831
rect 56784 39788 56836 39797
rect 57888 39788 57940 39840
rect 61660 39788 61712 39840
rect 64144 39831 64196 39840
rect 64144 39797 64153 39831
rect 64153 39797 64187 39831
rect 64187 39797 64196 39831
rect 64144 39788 64196 39797
rect 64236 39788 64288 39840
rect 65708 39788 65760 39840
rect 67640 39788 67692 39840
rect 71044 39933 71053 39967
rect 71053 39933 71087 39967
rect 71087 39933 71096 39967
rect 71044 39924 71096 39933
rect 73988 39967 74040 39976
rect 73988 39933 73997 39967
rect 73997 39933 74031 39967
rect 74031 39933 74040 39967
rect 73988 39924 74040 39933
rect 74448 39967 74500 39976
rect 74448 39933 74457 39967
rect 74457 39933 74491 39967
rect 74491 39933 74500 39967
rect 74448 39924 74500 39933
rect 77484 39967 77536 39976
rect 77484 39933 77493 39967
rect 77493 39933 77527 39967
rect 77527 39933 77536 39967
rect 77484 39924 77536 39933
rect 80336 39924 80388 39976
rect 74356 39899 74408 39908
rect 70768 39788 70820 39840
rect 73896 39788 73948 39840
rect 74356 39865 74365 39899
rect 74365 39865 74399 39899
rect 74399 39865 74408 39899
rect 74356 39856 74408 39865
rect 74908 39899 74960 39908
rect 74908 39865 74917 39899
rect 74917 39865 74951 39899
rect 74951 39865 74960 39899
rect 74908 39856 74960 39865
rect 79876 39856 79928 39908
rect 80520 39967 80572 39976
rect 80520 39933 80529 39967
rect 80529 39933 80563 39967
rect 80563 39933 80572 39967
rect 80796 39967 80848 39976
rect 80520 39924 80572 39933
rect 80796 39933 80805 39967
rect 80805 39933 80839 39967
rect 80839 39933 80848 39967
rect 80796 39924 80848 39933
rect 80888 39967 80940 39976
rect 80888 39933 80897 39967
rect 80897 39933 80931 39967
rect 80931 39933 80940 39967
rect 82360 40001 82369 40035
rect 82369 40001 82403 40035
rect 82403 40001 82412 40035
rect 82360 39992 82412 40001
rect 80888 39924 80940 39933
rect 82728 39924 82780 39976
rect 84108 39924 84160 39976
rect 84936 39992 84988 40044
rect 85212 40035 85264 40044
rect 85212 40001 85221 40035
rect 85221 40001 85255 40035
rect 85255 40001 85264 40035
rect 85212 39992 85264 40001
rect 81440 39856 81492 39908
rect 86224 40060 86276 40112
rect 85764 39992 85816 40044
rect 88432 39992 88484 40044
rect 88984 39992 89036 40044
rect 85948 39967 86000 39976
rect 85948 39933 85957 39967
rect 85957 39933 85991 39967
rect 85991 39933 86000 39967
rect 85948 39924 86000 39933
rect 86500 39924 86552 39976
rect 88524 39967 88576 39976
rect 88524 39933 88533 39967
rect 88533 39933 88567 39967
rect 88567 39933 88576 39967
rect 88524 39924 88576 39933
rect 91100 39924 91152 39976
rect 77392 39788 77444 39840
rect 77576 39831 77628 39840
rect 77576 39797 77585 39831
rect 77585 39797 77619 39831
rect 77619 39797 77628 39831
rect 77576 39788 77628 39797
rect 80796 39788 80848 39840
rect 80888 39788 80940 39840
rect 84200 39788 84252 39840
rect 84568 39788 84620 39840
rect 85948 39788 86000 39840
rect 86684 39788 86736 39840
rect 86868 39788 86920 39840
rect 19606 39686 19658 39738
rect 19670 39686 19722 39738
rect 19734 39686 19786 39738
rect 19798 39686 19850 39738
rect 50326 39686 50378 39738
rect 50390 39686 50442 39738
rect 50454 39686 50506 39738
rect 50518 39686 50570 39738
rect 81046 39686 81098 39738
rect 81110 39686 81162 39738
rect 81174 39686 81226 39738
rect 81238 39686 81290 39738
rect 2780 39584 2832 39636
rect 3700 39516 3752 39568
rect 3976 39516 4028 39568
rect 4804 39516 4856 39568
rect 4988 39559 5040 39568
rect 4988 39525 4997 39559
rect 4997 39525 5031 39559
rect 5031 39525 5040 39559
rect 4988 39516 5040 39525
rect 8208 39516 8260 39568
rect 8300 39516 8352 39568
rect 16488 39584 16540 39636
rect 21548 39584 21600 39636
rect 24124 39584 24176 39636
rect 32220 39584 32272 39636
rect 33968 39584 34020 39636
rect 7472 39448 7524 39500
rect 7840 39491 7892 39500
rect 7840 39457 7849 39491
rect 7849 39457 7883 39491
rect 7883 39457 7892 39491
rect 9680 39491 9732 39500
rect 7840 39448 7892 39457
rect 9680 39457 9689 39491
rect 9689 39457 9723 39491
rect 9723 39457 9732 39491
rect 9680 39448 9732 39457
rect 11796 39491 11848 39500
rect 4620 39380 4672 39432
rect 5724 39380 5776 39432
rect 7380 39423 7432 39432
rect 7380 39389 7389 39423
rect 7389 39389 7423 39423
rect 7423 39389 7432 39423
rect 7380 39380 7432 39389
rect 11796 39457 11805 39491
rect 11805 39457 11839 39491
rect 11839 39457 11848 39491
rect 11796 39448 11848 39457
rect 13084 39491 13136 39500
rect 13084 39457 13093 39491
rect 13093 39457 13127 39491
rect 13127 39457 13136 39491
rect 13084 39448 13136 39457
rect 13544 39448 13596 39500
rect 13820 39491 13872 39500
rect 13820 39457 13829 39491
rect 13829 39457 13863 39491
rect 13863 39457 13872 39491
rect 13820 39448 13872 39457
rect 14464 39448 14516 39500
rect 12716 39380 12768 39432
rect 20996 39516 21048 39568
rect 25412 39516 25464 39568
rect 25964 39516 26016 39568
rect 15568 39448 15620 39500
rect 20720 39448 20772 39500
rect 25596 39448 25648 39500
rect 31576 39516 31628 39568
rect 31760 39516 31812 39568
rect 43628 39584 43680 39636
rect 49056 39584 49108 39636
rect 27620 39491 27672 39500
rect 27620 39457 27629 39491
rect 27629 39457 27663 39491
rect 27663 39457 27672 39491
rect 27620 39448 27672 39457
rect 32312 39491 32364 39500
rect 32312 39457 32321 39491
rect 32321 39457 32355 39491
rect 32355 39457 32364 39491
rect 32312 39448 32364 39457
rect 32772 39448 32824 39500
rect 33048 39491 33100 39500
rect 33048 39457 33057 39491
rect 33057 39457 33091 39491
rect 33091 39457 33100 39491
rect 33048 39448 33100 39457
rect 34336 39491 34388 39500
rect 34336 39457 34345 39491
rect 34345 39457 34379 39491
rect 34379 39457 34388 39491
rect 34336 39448 34388 39457
rect 27712 39380 27764 39432
rect 27804 39380 27856 39432
rect 31760 39380 31812 39432
rect 33508 39380 33560 39432
rect 34520 39380 34572 39432
rect 46112 39516 46164 39568
rect 39120 39448 39172 39500
rect 39488 39491 39540 39500
rect 39488 39457 39497 39491
rect 39497 39457 39531 39491
rect 39531 39457 39540 39491
rect 39856 39491 39908 39500
rect 39488 39448 39540 39457
rect 39856 39457 39865 39491
rect 39865 39457 39899 39491
rect 39899 39457 39908 39491
rect 39856 39448 39908 39457
rect 39948 39491 40000 39500
rect 39948 39457 39957 39491
rect 39957 39457 39991 39491
rect 39991 39457 40000 39491
rect 39948 39448 40000 39457
rect 43904 39448 43956 39500
rect 44364 39491 44416 39500
rect 39580 39380 39632 39432
rect 40868 39380 40920 39432
rect 42800 39380 42852 39432
rect 44364 39457 44373 39491
rect 44373 39457 44407 39491
rect 44407 39457 44416 39491
rect 44364 39448 44416 39457
rect 44916 39491 44968 39500
rect 44916 39457 44925 39491
rect 44925 39457 44959 39491
rect 44959 39457 44968 39491
rect 48596 39516 48648 39568
rect 48780 39516 48832 39568
rect 48872 39516 48924 39568
rect 49792 39584 49844 39636
rect 50160 39627 50212 39636
rect 50160 39593 50169 39627
rect 50169 39593 50203 39627
rect 50203 39593 50212 39627
rect 50160 39584 50212 39593
rect 50712 39627 50764 39636
rect 50712 39593 50721 39627
rect 50721 39593 50755 39627
rect 50755 39593 50764 39627
rect 50712 39584 50764 39593
rect 50804 39584 50856 39636
rect 51540 39584 51592 39636
rect 53656 39584 53708 39636
rect 49424 39516 49476 39568
rect 44916 39448 44968 39457
rect 6368 39355 6420 39364
rect 6368 39321 6377 39355
rect 6377 39321 6411 39355
rect 6411 39321 6420 39355
rect 6368 39312 6420 39321
rect 7748 39312 7800 39364
rect 45836 39380 45888 39432
rect 46756 39423 46808 39432
rect 46756 39389 46765 39423
rect 46765 39389 46799 39423
rect 46799 39389 46808 39423
rect 46756 39380 46808 39389
rect 48964 39423 49016 39432
rect 48964 39389 48973 39423
rect 48973 39389 49007 39423
rect 49007 39389 49016 39423
rect 48964 39380 49016 39389
rect 49332 39448 49384 39500
rect 50436 39516 50488 39568
rect 54668 39559 54720 39568
rect 54668 39525 54677 39559
rect 54677 39525 54711 39559
rect 54711 39525 54720 39559
rect 54668 39516 54720 39525
rect 57796 39516 57848 39568
rect 49792 39448 49844 39500
rect 50712 39448 50764 39500
rect 50436 39380 50488 39432
rect 51632 39380 51684 39432
rect 51908 39423 51960 39432
rect 51908 39389 51917 39423
rect 51917 39389 51951 39423
rect 51951 39389 51960 39423
rect 51908 39380 51960 39389
rect 52092 39491 52144 39500
rect 52092 39457 52101 39491
rect 52101 39457 52135 39491
rect 52135 39457 52144 39491
rect 52092 39448 52144 39457
rect 52644 39491 52696 39500
rect 52644 39457 52653 39491
rect 52653 39457 52687 39491
rect 52687 39457 52696 39491
rect 52644 39448 52696 39457
rect 52828 39491 52880 39500
rect 52828 39457 52837 39491
rect 52837 39457 52871 39491
rect 52871 39457 52880 39491
rect 52828 39448 52880 39457
rect 54300 39448 54352 39500
rect 58072 39491 58124 39500
rect 58072 39457 58081 39491
rect 58081 39457 58115 39491
rect 58115 39457 58124 39491
rect 58072 39448 58124 39457
rect 58164 39448 58216 39500
rect 59084 39516 59136 39568
rect 59176 39516 59228 39568
rect 52184 39380 52236 39432
rect 54668 39380 54720 39432
rect 57980 39423 58032 39432
rect 57980 39389 57989 39423
rect 57989 39389 58023 39423
rect 58023 39389 58032 39423
rect 57980 39380 58032 39389
rect 4804 39244 4856 39296
rect 6552 39287 6604 39296
rect 6552 39253 6561 39287
rect 6561 39253 6595 39287
rect 6595 39253 6604 39287
rect 6552 39244 6604 39253
rect 7840 39244 7892 39296
rect 8300 39244 8352 39296
rect 11980 39287 12032 39296
rect 11980 39253 11989 39287
rect 11989 39253 12023 39287
rect 12023 39253 12032 39287
rect 11980 39244 12032 39253
rect 12716 39287 12768 39296
rect 12716 39253 12725 39287
rect 12725 39253 12759 39287
rect 12759 39253 12768 39287
rect 12716 39244 12768 39253
rect 14096 39287 14148 39296
rect 14096 39253 14105 39287
rect 14105 39253 14139 39287
rect 14139 39253 14148 39287
rect 14096 39244 14148 39253
rect 14464 39287 14516 39296
rect 14464 39253 14473 39287
rect 14473 39253 14507 39287
rect 14507 39253 14516 39287
rect 14464 39244 14516 39253
rect 19892 39287 19944 39296
rect 19892 39253 19901 39287
rect 19901 39253 19935 39287
rect 19935 39253 19944 39287
rect 19892 39244 19944 39253
rect 20812 39244 20864 39296
rect 27804 39287 27856 39296
rect 27804 39253 27813 39287
rect 27813 39253 27847 39287
rect 27847 39253 27856 39287
rect 27804 39244 27856 39253
rect 27988 39244 28040 39296
rect 33048 39244 33100 39296
rect 33232 39244 33284 39296
rect 33876 39287 33928 39296
rect 33876 39253 33885 39287
rect 33885 39253 33919 39287
rect 33919 39253 33928 39287
rect 33876 39244 33928 39253
rect 33968 39244 34020 39296
rect 34612 39287 34664 39296
rect 34612 39253 34621 39287
rect 34621 39253 34655 39287
rect 34655 39253 34664 39287
rect 34612 39244 34664 39253
rect 34796 39244 34848 39296
rect 40316 39244 40368 39296
rect 40684 39244 40736 39296
rect 40960 39244 41012 39296
rect 42708 39244 42760 39296
rect 43444 39244 43496 39296
rect 43904 39244 43956 39296
rect 44088 39244 44140 39296
rect 44364 39244 44416 39296
rect 44916 39244 44968 39296
rect 45928 39287 45980 39296
rect 45928 39253 45937 39287
rect 45937 39253 45971 39287
rect 45971 39253 45980 39287
rect 45928 39244 45980 39253
rect 46204 39244 46256 39296
rect 47032 39287 47084 39296
rect 47032 39253 47041 39287
rect 47041 39253 47075 39287
rect 47075 39253 47084 39287
rect 47032 39244 47084 39253
rect 49884 39312 49936 39364
rect 53564 39312 53616 39364
rect 56692 39312 56744 39364
rect 60924 39448 60976 39500
rect 59084 39312 59136 39364
rect 59452 39312 59504 39364
rect 65708 39516 65760 39568
rect 71044 39584 71096 39636
rect 72608 39627 72660 39636
rect 72608 39593 72617 39627
rect 72617 39593 72651 39627
rect 72651 39593 72660 39627
rect 72608 39584 72660 39593
rect 77484 39584 77536 39636
rect 81440 39584 81492 39636
rect 61200 39491 61252 39500
rect 61200 39457 61209 39491
rect 61209 39457 61243 39491
rect 61243 39457 61252 39491
rect 61200 39448 61252 39457
rect 61844 39380 61896 39432
rect 63500 39380 63552 39432
rect 61108 39312 61160 39364
rect 53288 39244 53340 39296
rect 53380 39244 53432 39296
rect 54116 39244 54168 39296
rect 54300 39287 54352 39296
rect 54300 39253 54309 39287
rect 54309 39253 54343 39287
rect 54343 39253 54352 39287
rect 54300 39244 54352 39253
rect 54668 39244 54720 39296
rect 57980 39244 58032 39296
rect 59176 39244 59228 39296
rect 59360 39287 59412 39296
rect 59360 39253 59369 39287
rect 59369 39253 59403 39287
rect 59403 39253 59412 39287
rect 59360 39244 59412 39253
rect 59544 39244 59596 39296
rect 65340 39244 65392 39296
rect 67456 39448 67508 39500
rect 71964 39448 72016 39500
rect 72332 39448 72384 39500
rect 72424 39380 72476 39432
rect 67548 39312 67600 39364
rect 73160 39312 73212 39364
rect 66168 39244 66220 39296
rect 74908 39448 74960 39500
rect 77300 39491 77352 39500
rect 73896 39380 73948 39432
rect 77300 39457 77309 39491
rect 77309 39457 77343 39491
rect 77343 39457 77352 39491
rect 77300 39448 77352 39457
rect 78312 39448 78364 39500
rect 79876 39491 79928 39500
rect 79876 39457 79885 39491
rect 79885 39457 79919 39491
rect 79919 39457 79928 39491
rect 79876 39448 79928 39457
rect 81348 39448 81400 39500
rect 83004 39584 83056 39636
rect 85672 39584 85724 39636
rect 85948 39627 86000 39636
rect 85948 39593 85957 39627
rect 85957 39593 85991 39627
rect 85991 39593 86000 39627
rect 85948 39584 86000 39593
rect 89444 39584 89496 39636
rect 91100 39627 91152 39636
rect 91100 39593 91109 39627
rect 91109 39593 91143 39627
rect 91143 39593 91152 39627
rect 91100 39584 91152 39593
rect 83832 39448 83884 39500
rect 84568 39448 84620 39500
rect 85764 39491 85816 39500
rect 85764 39457 85773 39491
rect 85773 39457 85807 39491
rect 85807 39457 85816 39491
rect 85764 39448 85816 39457
rect 86868 39491 86920 39500
rect 86868 39457 86877 39491
rect 86877 39457 86911 39491
rect 86911 39457 86920 39491
rect 86868 39448 86920 39457
rect 89904 39491 89956 39500
rect 89904 39457 89913 39491
rect 89913 39457 89947 39491
rect 89947 39457 89956 39491
rect 89904 39448 89956 39457
rect 91008 39491 91060 39500
rect 91008 39457 91017 39491
rect 91017 39457 91051 39491
rect 91051 39457 91060 39491
rect 91008 39448 91060 39457
rect 82360 39380 82412 39432
rect 84108 39380 84160 39432
rect 84844 39423 84896 39432
rect 80520 39312 80572 39364
rect 83280 39312 83332 39364
rect 84844 39389 84853 39423
rect 84853 39389 84887 39423
rect 84887 39389 84896 39423
rect 84844 39380 84896 39389
rect 84936 39380 84988 39432
rect 88524 39380 88576 39432
rect 90088 39312 90140 39364
rect 74908 39287 74960 39296
rect 74908 39253 74917 39287
rect 74917 39253 74951 39287
rect 74951 39253 74960 39287
rect 74908 39244 74960 39253
rect 83740 39244 83792 39296
rect 84568 39244 84620 39296
rect 86224 39244 86276 39296
rect 88524 39244 88576 39296
rect 4246 39142 4298 39194
rect 4310 39142 4362 39194
rect 4374 39142 4426 39194
rect 4438 39142 4490 39194
rect 34966 39142 35018 39194
rect 35030 39142 35082 39194
rect 35094 39142 35146 39194
rect 35158 39142 35210 39194
rect 65686 39142 65738 39194
rect 65750 39142 65802 39194
rect 65814 39142 65866 39194
rect 65878 39142 65930 39194
rect 96406 39142 96458 39194
rect 96470 39142 96522 39194
rect 96534 39142 96586 39194
rect 96598 39142 96650 39194
rect 3424 39040 3476 39092
rect 7932 39040 7984 39092
rect 2780 38947 2832 38956
rect 2780 38913 2789 38947
rect 2789 38913 2823 38947
rect 2823 38913 2832 38947
rect 2780 38904 2832 38913
rect 7472 38904 7524 38956
rect 3884 38743 3936 38752
rect 3884 38709 3893 38743
rect 3893 38709 3927 38743
rect 3927 38709 3936 38743
rect 3884 38700 3936 38709
rect 8208 38879 8260 38888
rect 6276 38768 6328 38820
rect 8208 38845 8217 38879
rect 8217 38845 8251 38879
rect 8251 38845 8260 38879
rect 8208 38836 8260 38845
rect 8484 38836 8536 38888
rect 13820 39040 13872 39092
rect 20720 39083 20772 39092
rect 20720 39049 20729 39083
rect 20729 39049 20763 39083
rect 20763 39049 20772 39083
rect 20720 39040 20772 39049
rect 21364 39040 21416 39092
rect 38660 39040 38712 39092
rect 48320 39040 48372 39092
rect 12624 38972 12676 39024
rect 20812 38972 20864 39024
rect 22008 38972 22060 39024
rect 13820 38904 13872 38956
rect 10784 38879 10836 38888
rect 10784 38845 10793 38879
rect 10793 38845 10827 38879
rect 10827 38845 10836 38879
rect 10784 38836 10836 38845
rect 12072 38836 12124 38888
rect 13636 38836 13688 38888
rect 24124 38904 24176 38956
rect 26332 38904 26384 38956
rect 19248 38836 19300 38888
rect 19432 38879 19484 38888
rect 19432 38845 19441 38879
rect 19441 38845 19475 38879
rect 19475 38845 19484 38879
rect 19432 38836 19484 38845
rect 19892 38836 19944 38888
rect 20352 38836 20404 38888
rect 21640 38879 21692 38888
rect 21640 38845 21649 38879
rect 21649 38845 21683 38879
rect 21683 38845 21692 38879
rect 21640 38836 21692 38845
rect 26424 38879 26476 38888
rect 26424 38845 26433 38879
rect 26433 38845 26467 38879
rect 26467 38845 26476 38879
rect 26424 38836 26476 38845
rect 4712 38700 4764 38752
rect 9956 38743 10008 38752
rect 9956 38709 9965 38743
rect 9965 38709 9999 38743
rect 9999 38709 10008 38743
rect 9956 38700 10008 38709
rect 10784 38700 10836 38752
rect 13820 38700 13872 38752
rect 20996 38700 21048 38752
rect 27160 38768 27212 38820
rect 28264 38700 28316 38752
rect 32772 38972 32824 39024
rect 34520 38972 34572 39024
rect 39028 39015 39080 39024
rect 39028 38981 39052 39015
rect 39052 38981 39080 39015
rect 39028 38972 39080 38981
rect 46204 38972 46256 39024
rect 33876 38904 33928 38956
rect 33508 38811 33560 38820
rect 33508 38777 33517 38811
rect 33517 38777 33551 38811
rect 33551 38777 33560 38811
rect 33508 38768 33560 38777
rect 32312 38700 32364 38752
rect 38752 38904 38804 38956
rect 39580 38904 39632 38956
rect 45100 38947 45152 38956
rect 38844 38879 38896 38888
rect 38844 38845 38853 38879
rect 38853 38845 38887 38879
rect 38887 38845 38896 38879
rect 38844 38836 38896 38845
rect 40960 38836 41012 38888
rect 40224 38768 40276 38820
rect 43812 38879 43864 38888
rect 43812 38845 43821 38879
rect 43821 38845 43855 38879
rect 43855 38845 43864 38879
rect 43812 38836 43864 38845
rect 44088 38836 44140 38888
rect 45100 38913 45109 38947
rect 45109 38913 45143 38947
rect 45143 38913 45152 38947
rect 45100 38904 45152 38913
rect 44916 38836 44968 38888
rect 45928 38904 45980 38956
rect 47032 38904 47084 38956
rect 46112 38879 46164 38888
rect 46112 38845 46121 38879
rect 46121 38845 46155 38879
rect 46155 38845 46164 38879
rect 46112 38836 46164 38845
rect 46572 38836 46624 38888
rect 46664 38836 46716 38888
rect 48964 38904 49016 38956
rect 49884 39015 49936 39024
rect 49884 38981 49893 39015
rect 49893 38981 49927 39015
rect 49927 38981 49936 39015
rect 50436 39015 50488 39024
rect 49884 38972 49936 38981
rect 50436 38981 50445 39015
rect 50445 38981 50479 39015
rect 50479 38981 50488 39015
rect 50436 38972 50488 38981
rect 50712 38972 50764 39024
rect 51448 39040 51500 39092
rect 52184 39040 52236 39092
rect 61108 39040 61160 39092
rect 51080 38904 51132 38956
rect 48872 38879 48924 38888
rect 48872 38845 48881 38879
rect 48881 38845 48915 38879
rect 48915 38845 48924 38879
rect 48872 38836 48924 38845
rect 49424 38879 49476 38888
rect 49424 38845 49433 38879
rect 49433 38845 49467 38879
rect 49467 38845 49476 38879
rect 49424 38836 49476 38845
rect 49516 38836 49568 38888
rect 52552 38972 52604 39024
rect 54208 38972 54260 39024
rect 60648 38972 60700 39024
rect 60740 39015 60792 39024
rect 60740 38981 60749 39015
rect 60749 38981 60783 39015
rect 60783 38981 60792 39015
rect 60740 38972 60792 38981
rect 61016 38972 61068 39024
rect 83740 39040 83792 39092
rect 64144 38972 64196 39024
rect 65524 38972 65576 39024
rect 67640 38972 67692 39024
rect 80888 38972 80940 39024
rect 52092 38947 52144 38956
rect 52092 38913 52101 38947
rect 52101 38913 52135 38947
rect 52135 38913 52144 38947
rect 52092 38904 52144 38913
rect 52460 38947 52512 38956
rect 52460 38913 52469 38947
rect 52469 38913 52503 38947
rect 52503 38913 52512 38947
rect 52460 38904 52512 38913
rect 54208 38836 54260 38888
rect 54668 38904 54720 38956
rect 42892 38700 42944 38752
rect 43260 38700 43312 38752
rect 43812 38700 43864 38752
rect 43904 38700 43956 38752
rect 46664 38700 46716 38752
rect 48412 38700 48464 38752
rect 49516 38700 49568 38752
rect 51448 38743 51500 38752
rect 51448 38709 51457 38743
rect 51457 38709 51491 38743
rect 51491 38709 51500 38743
rect 51448 38700 51500 38709
rect 54208 38700 54260 38752
rect 57980 38836 58032 38888
rect 58256 38879 58308 38888
rect 58256 38845 58265 38879
rect 58265 38845 58299 38879
rect 58299 38845 58308 38879
rect 58256 38836 58308 38845
rect 58624 38879 58676 38888
rect 58624 38845 58633 38879
rect 58633 38845 58667 38879
rect 58667 38845 58676 38879
rect 58624 38836 58676 38845
rect 67548 38904 67600 38956
rect 70216 38904 70268 38956
rect 59084 38879 59136 38888
rect 54484 38768 54536 38820
rect 59084 38845 59093 38879
rect 59093 38845 59127 38879
rect 59127 38845 59136 38879
rect 59084 38836 59136 38845
rect 59360 38836 59412 38888
rect 61016 38836 61068 38888
rect 61200 38879 61252 38888
rect 61200 38845 61223 38879
rect 61223 38845 61252 38879
rect 61200 38836 61252 38845
rect 61660 38879 61712 38888
rect 54576 38700 54628 38752
rect 56600 38700 56652 38752
rect 58164 38700 58216 38752
rect 59452 38768 59504 38820
rect 61660 38845 61669 38879
rect 61669 38845 61703 38879
rect 61703 38845 61712 38879
rect 61660 38836 61712 38845
rect 61844 38879 61896 38888
rect 61844 38845 61853 38879
rect 61853 38845 61887 38879
rect 61887 38845 61896 38879
rect 61844 38836 61896 38845
rect 65524 38879 65576 38888
rect 65524 38845 65533 38879
rect 65533 38845 65567 38879
rect 65567 38845 65576 38879
rect 65524 38836 65576 38845
rect 66168 38836 66220 38888
rect 69664 38879 69716 38888
rect 69664 38845 69673 38879
rect 69673 38845 69707 38879
rect 69707 38845 69716 38879
rect 69664 38836 69716 38845
rect 70308 38836 70360 38888
rect 71504 38836 71556 38888
rect 72424 38904 72476 38956
rect 72332 38836 72384 38888
rect 74448 38904 74500 38956
rect 74724 38904 74776 38956
rect 82360 38904 82412 38956
rect 82728 38904 82780 38956
rect 73068 38836 73120 38888
rect 74908 38836 74960 38888
rect 65432 38700 65484 38752
rect 67732 38700 67784 38752
rect 70308 38700 70360 38752
rect 72424 38700 72476 38752
rect 73988 38700 74040 38752
rect 79508 38836 79560 38888
rect 83188 38972 83240 39024
rect 84568 39083 84620 39092
rect 84568 39049 84577 39083
rect 84577 39049 84611 39083
rect 84611 39049 84620 39083
rect 84568 39040 84620 39049
rect 85672 39083 85724 39092
rect 85672 39049 85681 39083
rect 85681 39049 85715 39083
rect 85715 39049 85724 39083
rect 85672 39040 85724 39049
rect 84200 39015 84252 39024
rect 83372 38904 83424 38956
rect 84200 38981 84209 39015
rect 84209 38981 84243 39015
rect 84243 38981 84252 39015
rect 84200 38972 84252 38981
rect 83740 38904 83792 38956
rect 84108 38947 84160 38956
rect 84108 38913 84117 38947
rect 84117 38913 84151 38947
rect 84151 38913 84160 38947
rect 84108 38904 84160 38913
rect 82820 38768 82872 38820
rect 83372 38811 83424 38820
rect 77300 38700 77352 38752
rect 77392 38700 77444 38752
rect 81532 38700 81584 38752
rect 83372 38777 83381 38811
rect 83381 38777 83415 38811
rect 83415 38777 83424 38811
rect 83372 38768 83424 38777
rect 84568 38836 84620 38888
rect 86868 38879 86920 38888
rect 86868 38845 86877 38879
rect 86877 38845 86911 38879
rect 86911 38845 86920 38879
rect 86868 38836 86920 38845
rect 86960 38879 87012 38888
rect 86960 38845 86969 38879
rect 86969 38845 87003 38879
rect 87003 38845 87012 38879
rect 86960 38836 87012 38845
rect 89076 38836 89128 38888
rect 91560 38879 91612 38888
rect 91560 38845 91569 38879
rect 91569 38845 91603 38879
rect 91603 38845 91612 38879
rect 91560 38836 91612 38845
rect 84844 38768 84896 38820
rect 89904 38768 89956 38820
rect 91100 38768 91152 38820
rect 93492 38768 93544 38820
rect 93400 38743 93452 38752
rect 93400 38709 93409 38743
rect 93409 38709 93443 38743
rect 93443 38709 93452 38743
rect 93400 38700 93452 38709
rect 19606 38598 19658 38650
rect 19670 38598 19722 38650
rect 19734 38598 19786 38650
rect 19798 38598 19850 38650
rect 50326 38598 50378 38650
rect 50390 38598 50442 38650
rect 50454 38598 50506 38650
rect 50518 38598 50570 38650
rect 81046 38598 81098 38650
rect 81110 38598 81162 38650
rect 81174 38598 81226 38650
rect 81238 38598 81290 38650
rect 2780 38496 2832 38548
rect 4804 38428 4856 38480
rect 5080 38496 5132 38548
rect 8484 38496 8536 38548
rect 11980 38496 12032 38548
rect 13544 38496 13596 38548
rect 20536 38496 20588 38548
rect 21180 38496 21232 38548
rect 22192 38496 22244 38548
rect 31484 38496 31536 38548
rect 42892 38496 42944 38548
rect 48320 38496 48372 38548
rect 61108 38496 61160 38548
rect 61292 38496 61344 38548
rect 70768 38496 70820 38548
rect 4068 38292 4120 38344
rect 18696 38428 18748 38480
rect 8576 38360 8628 38412
rect 9588 38292 9640 38344
rect 3792 38224 3844 38276
rect 8208 38156 8260 38208
rect 9956 38156 10008 38208
rect 11980 38403 12032 38412
rect 11980 38369 11989 38403
rect 11989 38369 12023 38403
rect 12023 38369 12032 38403
rect 11980 38360 12032 38369
rect 12164 38403 12216 38412
rect 12164 38369 12173 38403
rect 12173 38369 12207 38403
rect 12207 38369 12216 38403
rect 12164 38360 12216 38369
rect 14096 38360 14148 38412
rect 18788 38403 18840 38412
rect 18788 38369 18797 38403
rect 18797 38369 18831 38403
rect 18831 38369 18840 38403
rect 18788 38360 18840 38369
rect 19340 38360 19392 38412
rect 19524 38403 19576 38412
rect 19524 38369 19533 38403
rect 19533 38369 19567 38403
rect 19567 38369 19576 38403
rect 19984 38428 20036 38480
rect 20996 38428 21048 38480
rect 21088 38403 21140 38412
rect 19524 38360 19576 38369
rect 21088 38369 21097 38403
rect 21097 38369 21131 38403
rect 21131 38369 21140 38403
rect 21088 38360 21140 38369
rect 25412 38428 25464 38480
rect 27804 38428 27856 38480
rect 28816 38428 28868 38480
rect 42984 38428 43036 38480
rect 21732 38360 21784 38412
rect 22008 38360 22060 38412
rect 24308 38360 24360 38412
rect 25596 38360 25648 38412
rect 27896 38403 27948 38412
rect 27896 38369 27905 38403
rect 27905 38369 27939 38403
rect 27939 38369 27948 38403
rect 27896 38360 27948 38369
rect 28632 38403 28684 38412
rect 28632 38369 28641 38403
rect 28641 38369 28675 38403
rect 28675 38369 28684 38403
rect 28632 38360 28684 38369
rect 32864 38403 32916 38412
rect 32864 38369 32873 38403
rect 32873 38369 32907 38403
rect 32907 38369 32916 38403
rect 32864 38360 32916 38369
rect 39120 38360 39172 38412
rect 39212 38360 39264 38412
rect 39948 38360 40000 38412
rect 27344 38292 27396 38344
rect 33232 38335 33284 38344
rect 33232 38301 33241 38335
rect 33241 38301 33275 38335
rect 33275 38301 33284 38335
rect 33232 38292 33284 38301
rect 38936 38335 38988 38344
rect 38936 38301 38945 38335
rect 38945 38301 38979 38335
rect 38979 38301 38988 38335
rect 38936 38292 38988 38301
rect 40592 38360 40644 38412
rect 40500 38292 40552 38344
rect 24492 38224 24544 38276
rect 24860 38224 24912 38276
rect 32772 38224 32824 38276
rect 33324 38224 33376 38276
rect 51448 38428 51500 38480
rect 52460 38428 52512 38480
rect 44916 38403 44968 38412
rect 44916 38369 44925 38403
rect 44925 38369 44959 38403
rect 44959 38369 44968 38403
rect 44916 38360 44968 38369
rect 45376 38360 45428 38412
rect 50068 38360 50120 38412
rect 50344 38403 50396 38412
rect 50344 38369 50353 38403
rect 50353 38369 50387 38403
rect 50387 38369 50396 38403
rect 50344 38360 50396 38369
rect 46756 38292 46808 38344
rect 12716 38156 12768 38208
rect 14096 38156 14148 38208
rect 16028 38156 16080 38208
rect 19524 38156 19576 38208
rect 20352 38156 20404 38208
rect 20536 38156 20588 38208
rect 24032 38156 24084 38208
rect 26240 38156 26292 38208
rect 27160 38156 27212 38208
rect 27344 38156 27396 38208
rect 28908 38199 28960 38208
rect 28908 38165 28917 38199
rect 28917 38165 28951 38199
rect 28951 38165 28960 38199
rect 28908 38156 28960 38165
rect 33140 38199 33192 38208
rect 33140 38165 33149 38199
rect 33149 38165 33183 38199
rect 33183 38165 33192 38199
rect 33140 38156 33192 38165
rect 39120 38156 39172 38208
rect 40868 38156 40920 38208
rect 44088 38156 44140 38208
rect 45560 38156 45612 38208
rect 49884 38292 49936 38344
rect 50252 38335 50304 38344
rect 50252 38301 50261 38335
rect 50261 38301 50295 38335
rect 50295 38301 50304 38335
rect 50252 38292 50304 38301
rect 49792 38267 49844 38276
rect 49792 38233 49801 38267
rect 49801 38233 49835 38267
rect 49835 38233 49844 38267
rect 56692 38428 56744 38480
rect 56600 38403 56652 38412
rect 56600 38369 56609 38403
rect 56609 38369 56643 38403
rect 56643 38369 56652 38403
rect 56600 38360 56652 38369
rect 52460 38292 52512 38344
rect 56232 38292 56284 38344
rect 57428 38292 57480 38344
rect 57980 38292 58032 38344
rect 58164 38360 58216 38412
rect 58992 38360 59044 38412
rect 59728 38360 59780 38412
rect 62856 38403 62908 38412
rect 62856 38369 62865 38403
rect 62865 38369 62899 38403
rect 62899 38369 62908 38403
rect 62856 38360 62908 38369
rect 63500 38360 63552 38412
rect 63776 38428 63828 38480
rect 67732 38428 67784 38480
rect 69664 38428 69716 38480
rect 70124 38471 70176 38480
rect 70124 38437 70133 38471
rect 70133 38437 70167 38471
rect 70167 38437 70176 38471
rect 70124 38428 70176 38437
rect 59084 38335 59136 38344
rect 59084 38301 59093 38335
rect 59093 38301 59127 38335
rect 59127 38301 59136 38335
rect 59084 38292 59136 38301
rect 49792 38224 49844 38233
rect 48320 38156 48372 38208
rect 50252 38156 50304 38208
rect 51448 38156 51500 38208
rect 53196 38199 53248 38208
rect 53196 38165 53205 38199
rect 53205 38165 53239 38199
rect 53239 38165 53248 38199
rect 53196 38156 53248 38165
rect 53288 38156 53340 38208
rect 56692 38199 56744 38208
rect 56692 38165 56701 38199
rect 56701 38165 56735 38199
rect 56735 38165 56744 38199
rect 56692 38156 56744 38165
rect 57428 38199 57480 38208
rect 57428 38165 57437 38199
rect 57437 38165 57471 38199
rect 57471 38165 57480 38199
rect 57428 38156 57480 38165
rect 61936 38156 61988 38208
rect 62120 38199 62172 38208
rect 62120 38165 62129 38199
rect 62129 38165 62163 38199
rect 62163 38165 62172 38199
rect 62120 38156 62172 38165
rect 62580 38199 62632 38208
rect 62580 38165 62589 38199
rect 62589 38165 62623 38199
rect 62623 38165 62632 38199
rect 62580 38156 62632 38165
rect 64696 38156 64748 38208
rect 65340 38156 65392 38208
rect 67824 38292 67876 38344
rect 67364 38224 67416 38276
rect 71228 38496 71280 38548
rect 77576 38496 77628 38548
rect 84016 38496 84068 38548
rect 68928 38292 68980 38344
rect 71780 38292 71832 38344
rect 72332 38360 72384 38412
rect 73988 38360 74040 38412
rect 77392 38403 77444 38412
rect 77392 38369 77401 38403
rect 77401 38369 77435 38403
rect 77435 38369 77444 38403
rect 77392 38360 77444 38369
rect 81440 38360 81492 38412
rect 82820 38403 82872 38412
rect 82820 38369 82829 38403
rect 82829 38369 82863 38403
rect 82863 38369 82872 38403
rect 82820 38360 82872 38369
rect 82912 38403 82964 38412
rect 82912 38369 82921 38403
rect 82921 38369 82955 38403
rect 82955 38369 82964 38403
rect 89076 38539 89128 38548
rect 86960 38428 87012 38480
rect 88432 38471 88484 38480
rect 88432 38437 88441 38471
rect 88441 38437 88475 38471
rect 88475 38437 88484 38471
rect 88432 38428 88484 38437
rect 89076 38505 89085 38539
rect 89085 38505 89119 38539
rect 89119 38505 89128 38539
rect 89076 38496 89128 38505
rect 90088 38539 90140 38548
rect 90088 38505 90097 38539
rect 90097 38505 90131 38539
rect 90131 38505 90140 38539
rect 90088 38496 90140 38505
rect 93400 38496 93452 38548
rect 89444 38428 89496 38480
rect 91008 38428 91060 38480
rect 82912 38360 82964 38369
rect 72608 38292 72660 38344
rect 72792 38292 72844 38344
rect 85672 38360 85724 38412
rect 86224 38360 86276 38412
rect 91100 38403 91152 38412
rect 91100 38369 91109 38403
rect 91109 38369 91143 38403
rect 91143 38369 91152 38403
rect 91100 38360 91152 38369
rect 67456 38199 67508 38208
rect 67456 38165 67465 38199
rect 67465 38165 67499 38199
rect 67499 38165 67508 38199
rect 67456 38156 67508 38165
rect 71596 38224 71648 38276
rect 83188 38224 83240 38276
rect 72700 38156 72752 38208
rect 74172 38199 74224 38208
rect 74172 38165 74181 38199
rect 74181 38165 74215 38199
rect 74215 38165 74224 38199
rect 74172 38156 74224 38165
rect 77484 38199 77536 38208
rect 77484 38165 77493 38199
rect 77493 38165 77527 38199
rect 77527 38165 77536 38199
rect 77484 38156 77536 38165
rect 81532 38156 81584 38208
rect 81716 38156 81768 38208
rect 83096 38199 83148 38208
rect 83096 38165 83105 38199
rect 83105 38165 83139 38199
rect 83139 38165 83148 38199
rect 83096 38156 83148 38165
rect 88524 38292 88576 38344
rect 90088 38292 90140 38344
rect 90916 38292 90968 38344
rect 94596 38335 94648 38344
rect 88708 38199 88760 38208
rect 88708 38165 88717 38199
rect 88717 38165 88751 38199
rect 88751 38165 88760 38199
rect 88708 38156 88760 38165
rect 89628 38199 89680 38208
rect 89628 38165 89637 38199
rect 89637 38165 89671 38199
rect 89671 38165 89680 38199
rect 89628 38156 89680 38165
rect 89720 38156 89772 38208
rect 91008 38156 91060 38208
rect 94596 38301 94605 38335
rect 94605 38301 94639 38335
rect 94639 38301 94648 38335
rect 94596 38292 94648 38301
rect 94504 38156 94556 38208
rect 4246 38054 4298 38106
rect 4310 38054 4362 38106
rect 4374 38054 4426 38106
rect 4438 38054 4490 38106
rect 34966 38054 35018 38106
rect 35030 38054 35082 38106
rect 35094 38054 35146 38106
rect 35158 38054 35210 38106
rect 65686 38054 65738 38106
rect 65750 38054 65802 38106
rect 65814 38054 65866 38106
rect 65878 38054 65930 38106
rect 96406 38054 96458 38106
rect 96470 38054 96522 38106
rect 96534 38054 96586 38106
rect 96598 38054 96650 38106
rect 4804 37952 4856 38004
rect 10600 37952 10652 38004
rect 49792 37952 49844 38004
rect 49884 37952 49936 38004
rect 51172 37952 51224 38004
rect 51264 37952 51316 38004
rect 58992 37995 59044 38004
rect 2780 37859 2832 37868
rect 2780 37825 2789 37859
rect 2789 37825 2823 37859
rect 2823 37825 2832 37859
rect 2780 37816 2832 37825
rect 10784 37816 10836 37868
rect 12716 37859 12768 37868
rect 12716 37825 12725 37859
rect 12725 37825 12759 37859
rect 12759 37825 12768 37859
rect 12716 37816 12768 37825
rect 21180 37816 21232 37868
rect 26332 37884 26384 37936
rect 26424 37884 26476 37936
rect 27160 37884 27212 37936
rect 31484 37927 31536 37936
rect 31484 37893 31493 37927
rect 31493 37893 31527 37927
rect 31527 37893 31536 37927
rect 31484 37884 31536 37893
rect 31944 37884 31996 37936
rect 39028 37884 39080 37936
rect 45376 37927 45428 37936
rect 45376 37893 45385 37927
rect 45385 37893 45419 37927
rect 45419 37893 45428 37927
rect 45376 37884 45428 37893
rect 56324 37927 56376 37936
rect 5448 37748 5500 37800
rect 8208 37791 8260 37800
rect 8208 37757 8217 37791
rect 8217 37757 8251 37791
rect 8251 37757 8260 37791
rect 8208 37748 8260 37757
rect 8484 37748 8536 37800
rect 12164 37748 12216 37800
rect 18144 37791 18196 37800
rect 6552 37680 6604 37732
rect 18144 37757 18153 37791
rect 18153 37757 18187 37791
rect 18187 37757 18196 37791
rect 18144 37748 18196 37757
rect 18328 37748 18380 37800
rect 19156 37748 19208 37800
rect 20812 37748 20864 37800
rect 14096 37723 14148 37732
rect 14096 37689 14105 37723
rect 14105 37689 14139 37723
rect 14139 37689 14148 37723
rect 23388 37748 23440 37800
rect 25780 37791 25832 37800
rect 25780 37757 25789 37791
rect 25789 37757 25823 37791
rect 25823 37757 25832 37791
rect 25780 37748 25832 37757
rect 14096 37680 14148 37689
rect 3424 37612 3476 37664
rect 4252 37655 4304 37664
rect 4252 37621 4261 37655
rect 4261 37621 4295 37655
rect 4295 37621 4304 37655
rect 4252 37612 4304 37621
rect 13728 37612 13780 37664
rect 18328 37655 18380 37664
rect 18328 37621 18337 37655
rect 18337 37621 18371 37655
rect 18371 37621 18380 37655
rect 18328 37612 18380 37621
rect 28908 37816 28960 37868
rect 37004 37816 37056 37868
rect 39304 37816 39356 37868
rect 39948 37816 40000 37868
rect 40132 37816 40184 37868
rect 40868 37859 40920 37868
rect 40868 37825 40877 37859
rect 40877 37825 40911 37859
rect 40911 37825 40920 37859
rect 40868 37816 40920 37825
rect 41236 37859 41288 37868
rect 41236 37825 41245 37859
rect 41245 37825 41279 37859
rect 41279 37825 41288 37859
rect 41236 37816 41288 37825
rect 26148 37791 26200 37800
rect 26148 37757 26157 37791
rect 26157 37757 26191 37791
rect 26191 37757 26200 37791
rect 26148 37748 26200 37757
rect 27896 37748 27948 37800
rect 31852 37791 31904 37800
rect 31852 37757 31861 37791
rect 31861 37757 31895 37791
rect 31895 37757 31904 37791
rect 31852 37748 31904 37757
rect 31944 37791 31996 37800
rect 31944 37757 31953 37791
rect 31953 37757 31987 37791
rect 31987 37757 31996 37791
rect 33600 37791 33652 37800
rect 31944 37748 31996 37757
rect 33600 37757 33609 37791
rect 33609 37757 33643 37791
rect 33643 37757 33652 37791
rect 33600 37748 33652 37757
rect 37556 37748 37608 37800
rect 35992 37680 36044 37732
rect 40408 37748 40460 37800
rect 41144 37748 41196 37800
rect 39396 37680 39448 37732
rect 44088 37748 44140 37800
rect 44456 37791 44508 37800
rect 44456 37757 44465 37791
rect 44465 37757 44499 37791
rect 44499 37757 44508 37791
rect 44456 37748 44508 37757
rect 42892 37680 42944 37732
rect 45560 37859 45612 37868
rect 45560 37825 45569 37859
rect 45569 37825 45603 37859
rect 45603 37825 45612 37859
rect 45560 37816 45612 37825
rect 46664 37816 46716 37868
rect 49608 37816 49660 37868
rect 51356 37816 51408 37868
rect 46204 37748 46256 37800
rect 50712 37748 50764 37800
rect 51540 37748 51592 37800
rect 51816 37748 51868 37800
rect 52368 37791 52420 37800
rect 52368 37757 52377 37791
rect 52377 37757 52411 37791
rect 52411 37757 52420 37791
rect 52368 37748 52420 37757
rect 52460 37791 52512 37800
rect 52460 37757 52469 37791
rect 52469 37757 52503 37791
rect 52503 37757 52512 37791
rect 53380 37816 53432 37868
rect 56324 37893 56333 37927
rect 56333 37893 56367 37927
rect 56367 37893 56376 37927
rect 56324 37884 56376 37893
rect 58992 37961 59001 37995
rect 59001 37961 59035 37995
rect 59035 37961 59044 37995
rect 58992 37952 59044 37961
rect 60648 37952 60700 38004
rect 62120 37952 62172 38004
rect 62856 37952 62908 38004
rect 65432 37884 65484 37936
rect 59728 37816 59780 37868
rect 59912 37859 59964 37868
rect 59912 37825 59921 37859
rect 59921 37825 59955 37859
rect 59955 37825 59964 37859
rect 59912 37816 59964 37825
rect 60464 37859 60516 37868
rect 60464 37825 60473 37859
rect 60473 37825 60507 37859
rect 60507 37825 60516 37859
rect 60464 37816 60516 37825
rect 64236 37816 64288 37868
rect 64696 37859 64748 37868
rect 64696 37825 64705 37859
rect 64705 37825 64739 37859
rect 64739 37825 64748 37859
rect 64696 37816 64748 37825
rect 52460 37748 52512 37757
rect 56232 37791 56284 37800
rect 56232 37757 56241 37791
rect 56241 37757 56275 37791
rect 56275 37757 56284 37791
rect 56232 37748 56284 37757
rect 57428 37748 57480 37800
rect 58256 37748 58308 37800
rect 64328 37748 64380 37800
rect 68928 37791 68980 37800
rect 68928 37757 68937 37791
rect 68937 37757 68971 37791
rect 68971 37757 68980 37791
rect 68928 37748 68980 37757
rect 77484 37884 77536 37936
rect 82912 37952 82964 38004
rect 89444 37927 89496 37936
rect 71596 37859 71648 37868
rect 71596 37825 71605 37859
rect 71605 37825 71639 37859
rect 71639 37825 71648 37859
rect 71596 37816 71648 37825
rect 72700 37859 72752 37868
rect 72700 37825 72709 37859
rect 72709 37825 72743 37859
rect 72743 37825 72752 37859
rect 72700 37816 72752 37825
rect 76748 37859 76800 37868
rect 76748 37825 76757 37859
rect 76757 37825 76791 37859
rect 76791 37825 76800 37859
rect 76748 37816 76800 37825
rect 70492 37748 70544 37800
rect 70768 37748 70820 37800
rect 71044 37748 71096 37800
rect 71228 37791 71280 37800
rect 71228 37757 71237 37791
rect 71237 37757 71271 37791
rect 71271 37757 71280 37791
rect 71228 37748 71280 37757
rect 71320 37791 71372 37800
rect 71320 37757 71329 37791
rect 71329 37757 71363 37791
rect 71363 37757 71372 37791
rect 72240 37791 72292 37800
rect 71320 37748 71372 37757
rect 72240 37757 72249 37791
rect 72249 37757 72283 37791
rect 72283 37757 72292 37791
rect 72240 37748 72292 37757
rect 45560 37680 45612 37732
rect 48320 37680 48372 37732
rect 48412 37680 48464 37732
rect 20352 37612 20404 37664
rect 21640 37612 21692 37664
rect 21824 37655 21876 37664
rect 21824 37621 21833 37655
rect 21833 37621 21867 37655
rect 21867 37621 21876 37655
rect 21824 37612 21876 37621
rect 32036 37612 32088 37664
rect 37556 37612 37608 37664
rect 37740 37612 37792 37664
rect 38936 37612 38988 37664
rect 40132 37612 40184 37664
rect 42800 37612 42852 37664
rect 44088 37612 44140 37664
rect 46664 37612 46716 37664
rect 47860 37612 47912 37664
rect 52460 37612 52512 37664
rect 52920 37655 52972 37664
rect 52920 37621 52929 37655
rect 52929 37621 52963 37655
rect 52963 37621 52972 37655
rect 52920 37612 52972 37621
rect 53380 37612 53432 37664
rect 54208 37612 54260 37664
rect 69296 37680 69348 37732
rect 69572 37680 69624 37732
rect 72424 37748 72476 37800
rect 83096 37816 83148 37868
rect 89444 37893 89453 37927
rect 89453 37893 89487 37927
rect 89487 37893 89496 37927
rect 89444 37884 89496 37893
rect 91284 37884 91336 37936
rect 89904 37859 89956 37868
rect 77484 37791 77536 37800
rect 77484 37757 77493 37791
rect 77493 37757 77527 37791
rect 77527 37757 77536 37791
rect 77484 37748 77536 37757
rect 77668 37791 77720 37800
rect 77668 37757 77677 37791
rect 77677 37757 77711 37791
rect 77711 37757 77720 37791
rect 77668 37748 77720 37757
rect 82544 37748 82596 37800
rect 83832 37791 83884 37800
rect 83832 37757 83841 37791
rect 83841 37757 83875 37791
rect 83875 37757 83884 37791
rect 83832 37748 83884 37757
rect 85672 37791 85724 37800
rect 64236 37655 64288 37664
rect 64236 37621 64245 37655
rect 64245 37621 64279 37655
rect 64279 37621 64288 37655
rect 64236 37612 64288 37621
rect 64420 37612 64472 37664
rect 65340 37612 65392 37664
rect 68928 37612 68980 37664
rect 69112 37655 69164 37664
rect 69112 37621 69121 37655
rect 69121 37621 69155 37655
rect 69155 37621 69164 37655
rect 69112 37612 69164 37621
rect 71228 37612 71280 37664
rect 81440 37680 81492 37732
rect 85672 37757 85681 37791
rect 85681 37757 85715 37791
rect 85715 37757 85724 37791
rect 85672 37748 85724 37757
rect 89904 37825 89913 37859
rect 89913 37825 89947 37859
rect 89947 37825 89956 37859
rect 89904 37816 89956 37825
rect 91560 37859 91612 37868
rect 91560 37825 91569 37859
rect 91569 37825 91603 37859
rect 91603 37825 91612 37859
rect 91560 37816 91612 37825
rect 94596 37816 94648 37868
rect 89720 37748 89772 37800
rect 91008 37723 91060 37732
rect 77300 37612 77352 37664
rect 91008 37689 91017 37723
rect 91017 37689 91051 37723
rect 91051 37689 91060 37723
rect 91008 37680 91060 37689
rect 90732 37612 90784 37664
rect 93492 37791 93544 37800
rect 93492 37757 93501 37791
rect 93501 37757 93535 37791
rect 93535 37757 93544 37791
rect 93492 37748 93544 37757
rect 93584 37791 93636 37800
rect 93584 37757 93593 37791
rect 93593 37757 93627 37791
rect 93627 37757 93636 37791
rect 93584 37748 93636 37757
rect 95240 37791 95292 37800
rect 95240 37757 95249 37791
rect 95249 37757 95283 37791
rect 95283 37757 95292 37791
rect 95240 37748 95292 37757
rect 97080 37748 97132 37800
rect 95332 37680 95384 37732
rect 95700 37723 95752 37732
rect 95700 37689 95709 37723
rect 95709 37689 95743 37723
rect 95743 37689 95752 37723
rect 95700 37680 95752 37689
rect 96712 37655 96764 37664
rect 96712 37621 96721 37655
rect 96721 37621 96755 37655
rect 96755 37621 96764 37655
rect 96712 37612 96764 37621
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 50326 37510 50378 37562
rect 50390 37510 50442 37562
rect 50454 37510 50506 37562
rect 50518 37510 50570 37562
rect 81046 37510 81098 37562
rect 81110 37510 81162 37562
rect 81174 37510 81226 37562
rect 81238 37510 81290 37562
rect 8576 37340 8628 37392
rect 4620 37272 4672 37324
rect 16028 37408 16080 37460
rect 19432 37451 19484 37460
rect 19432 37417 19441 37451
rect 19441 37417 19475 37451
rect 19475 37417 19484 37451
rect 19432 37408 19484 37417
rect 19984 37408 20036 37460
rect 20720 37408 20772 37460
rect 20812 37408 20864 37460
rect 23388 37451 23440 37460
rect 23388 37417 23397 37451
rect 23397 37417 23431 37451
rect 23431 37417 23440 37451
rect 23388 37408 23440 37417
rect 24492 37451 24544 37460
rect 24492 37417 24501 37451
rect 24501 37417 24535 37451
rect 24535 37417 24544 37451
rect 24492 37408 24544 37417
rect 26240 37408 26292 37460
rect 28816 37408 28868 37460
rect 31852 37408 31904 37460
rect 13268 37340 13320 37392
rect 40316 37408 40368 37460
rect 40868 37451 40920 37460
rect 40868 37417 40877 37451
rect 40877 37417 40911 37451
rect 40911 37417 40920 37451
rect 40868 37408 40920 37417
rect 41420 37408 41472 37460
rect 47952 37451 48004 37460
rect 47952 37417 47961 37451
rect 47961 37417 47995 37451
rect 47995 37417 48004 37451
rect 47952 37408 48004 37417
rect 51172 37408 51224 37460
rect 57980 37451 58032 37460
rect 12164 37272 12216 37324
rect 14556 37315 14608 37324
rect 14556 37281 14565 37315
rect 14565 37281 14599 37315
rect 14599 37281 14608 37315
rect 14556 37272 14608 37281
rect 18236 37315 18288 37324
rect 18236 37281 18245 37315
rect 18245 37281 18279 37315
rect 18279 37281 18288 37315
rect 18236 37272 18288 37281
rect 18420 37315 18472 37324
rect 18420 37281 18429 37315
rect 18429 37281 18463 37315
rect 18463 37281 18472 37315
rect 18420 37272 18472 37281
rect 18788 37272 18840 37324
rect 4252 37204 4304 37256
rect 4804 37204 4856 37256
rect 8944 37204 8996 37256
rect 10048 37136 10100 37188
rect 13636 37136 13688 37188
rect 13820 37247 13872 37256
rect 13820 37213 13829 37247
rect 13829 37213 13863 37247
rect 13863 37213 13872 37247
rect 19800 37272 19852 37324
rect 21088 37315 21140 37324
rect 21088 37281 21097 37315
rect 21097 37281 21131 37315
rect 21131 37281 21140 37315
rect 21088 37272 21140 37281
rect 21824 37315 21876 37324
rect 21824 37281 21833 37315
rect 21833 37281 21867 37315
rect 21867 37281 21876 37315
rect 21824 37272 21876 37281
rect 13820 37204 13872 37213
rect 19984 37204 20036 37256
rect 20904 37247 20956 37256
rect 20904 37213 20913 37247
rect 20913 37213 20947 37247
rect 20947 37213 20956 37247
rect 20904 37204 20956 37213
rect 24768 37272 24820 37324
rect 25044 37315 25096 37324
rect 25044 37281 25053 37315
rect 25053 37281 25087 37315
rect 25087 37281 25096 37315
rect 25044 37272 25096 37281
rect 25412 37315 25464 37324
rect 25412 37281 25421 37315
rect 25421 37281 25455 37315
rect 25455 37281 25464 37315
rect 25412 37272 25464 37281
rect 26240 37272 26292 37324
rect 27344 37315 27396 37324
rect 27344 37281 27353 37315
rect 27353 37281 27387 37315
rect 27387 37281 27396 37315
rect 27344 37272 27396 37281
rect 27804 37272 27856 37324
rect 28724 37272 28776 37324
rect 32772 37272 32824 37324
rect 34704 37272 34756 37324
rect 34796 37272 34848 37324
rect 35716 37272 35768 37324
rect 36176 37315 36228 37324
rect 36176 37281 36185 37315
rect 36185 37281 36219 37315
rect 36219 37281 36228 37315
rect 36176 37272 36228 37281
rect 37740 37340 37792 37392
rect 39396 37383 39448 37392
rect 39396 37349 39405 37383
rect 39405 37349 39439 37383
rect 39439 37349 39448 37383
rect 39396 37340 39448 37349
rect 40224 37383 40276 37392
rect 40224 37349 40233 37383
rect 40233 37349 40267 37383
rect 40267 37349 40276 37383
rect 40224 37340 40276 37349
rect 24952 37204 25004 37256
rect 26056 37204 26108 37256
rect 28816 37204 28868 37256
rect 35440 37247 35492 37256
rect 35440 37213 35449 37247
rect 35449 37213 35483 37247
rect 35483 37213 35492 37247
rect 35440 37204 35492 37213
rect 37556 37247 37608 37256
rect 37556 37213 37565 37247
rect 37565 37213 37599 37247
rect 37599 37213 37608 37247
rect 37556 37204 37608 37213
rect 37740 37247 37792 37256
rect 37740 37213 37749 37247
rect 37749 37213 37783 37247
rect 37783 37213 37792 37247
rect 44732 37272 44784 37324
rect 45836 37340 45888 37392
rect 48964 37340 49016 37392
rect 40592 37247 40644 37256
rect 37740 37204 37792 37213
rect 40592 37213 40601 37247
rect 40601 37213 40635 37247
rect 40635 37213 40644 37247
rect 40592 37204 40644 37213
rect 43996 37204 44048 37256
rect 44088 37204 44140 37256
rect 47860 37315 47912 37324
rect 47860 37281 47869 37315
rect 47869 37281 47903 37315
rect 47903 37281 47912 37315
rect 47860 37272 47912 37281
rect 47952 37272 48004 37324
rect 48596 37272 48648 37324
rect 48688 37272 48740 37324
rect 50068 37315 50120 37324
rect 50068 37281 50077 37315
rect 50077 37281 50111 37315
rect 50111 37281 50120 37315
rect 50068 37272 50120 37281
rect 50804 37272 50856 37324
rect 51540 37340 51592 37392
rect 52368 37340 52420 37392
rect 52920 37340 52972 37392
rect 52552 37272 52604 37324
rect 56324 37340 56376 37392
rect 57980 37417 57989 37451
rect 57989 37417 58023 37451
rect 58023 37417 58032 37451
rect 57980 37408 58032 37417
rect 60464 37408 60516 37460
rect 69112 37408 69164 37460
rect 69572 37451 69624 37460
rect 69572 37417 69581 37451
rect 69581 37417 69615 37451
rect 69615 37417 69624 37451
rect 69572 37408 69624 37417
rect 53840 37204 53892 37256
rect 55128 37272 55180 37324
rect 54944 37247 54996 37256
rect 54944 37213 54953 37247
rect 54953 37213 54987 37247
rect 54987 37213 54996 37247
rect 54944 37204 54996 37213
rect 56232 37247 56284 37256
rect 56232 37213 56241 37247
rect 56241 37213 56275 37247
rect 56275 37213 56284 37247
rect 57336 37272 57388 37324
rect 65432 37340 65484 37392
rect 57520 37315 57572 37324
rect 57520 37281 57529 37315
rect 57529 37281 57563 37315
rect 57563 37281 57572 37315
rect 57520 37272 57572 37281
rect 63868 37272 63920 37324
rect 70768 37408 70820 37460
rect 56232 37204 56284 37213
rect 56600 37204 56652 37256
rect 62580 37204 62632 37256
rect 71228 37408 71280 37460
rect 72240 37408 72292 37460
rect 72792 37451 72844 37460
rect 72792 37417 72801 37451
rect 72801 37417 72835 37451
rect 72835 37417 72844 37451
rect 72792 37408 72844 37417
rect 73160 37408 73212 37460
rect 82820 37408 82872 37460
rect 88708 37408 88760 37460
rect 71780 37340 71832 37392
rect 71504 37272 71556 37324
rect 83004 37340 83056 37392
rect 72976 37272 73028 37324
rect 75920 37272 75972 37324
rect 83188 37272 83240 37324
rect 85580 37340 85632 37392
rect 86224 37272 86276 37324
rect 86868 37272 86920 37324
rect 69756 37247 69808 37256
rect 20812 37136 20864 37188
rect 22284 37136 22336 37188
rect 4068 37068 4120 37120
rect 7656 37068 7708 37120
rect 12532 37068 12584 37120
rect 12900 37068 12952 37120
rect 18236 37068 18288 37120
rect 20904 37068 20956 37120
rect 20996 37068 21048 37120
rect 31760 37068 31812 37120
rect 31944 37068 31996 37120
rect 32680 37068 32732 37120
rect 35992 37068 36044 37120
rect 40316 37068 40368 37120
rect 40500 37111 40552 37120
rect 40500 37077 40509 37111
rect 40509 37077 40543 37111
rect 40543 37077 40552 37111
rect 40500 37068 40552 37077
rect 67456 37136 67508 37188
rect 48504 37068 48556 37120
rect 49148 37111 49200 37120
rect 49148 37077 49157 37111
rect 49157 37077 49191 37111
rect 49191 37077 49200 37111
rect 49148 37068 49200 37077
rect 49240 37068 49292 37120
rect 50804 37068 50856 37120
rect 51632 37068 51684 37120
rect 54852 37111 54904 37120
rect 54852 37077 54861 37111
rect 54861 37077 54895 37111
rect 54895 37077 54904 37111
rect 54852 37068 54904 37077
rect 56600 37111 56652 37120
rect 56600 37077 56609 37111
rect 56609 37077 56643 37111
rect 56643 37077 56652 37111
rect 56600 37068 56652 37077
rect 62580 37111 62632 37120
rect 62580 37077 62589 37111
rect 62589 37077 62623 37111
rect 62623 37077 62632 37111
rect 62580 37068 62632 37077
rect 64788 37068 64840 37120
rect 69756 37213 69765 37247
rect 69765 37213 69799 37247
rect 69799 37213 69808 37247
rect 69756 37204 69808 37213
rect 72332 37247 72384 37256
rect 69296 37136 69348 37188
rect 72332 37213 72341 37247
rect 72341 37213 72375 37247
rect 72375 37213 72384 37247
rect 72332 37204 72384 37213
rect 77392 37204 77444 37256
rect 84476 37247 84528 37256
rect 84476 37213 84485 37247
rect 84485 37213 84519 37247
rect 84519 37213 84528 37247
rect 84476 37204 84528 37213
rect 91008 37340 91060 37392
rect 91284 37383 91336 37392
rect 91284 37349 91293 37383
rect 91293 37349 91327 37383
rect 91327 37349 91336 37383
rect 91284 37340 91336 37349
rect 91560 37340 91612 37392
rect 89720 37315 89772 37324
rect 89720 37281 89729 37315
rect 89729 37281 89763 37315
rect 89763 37281 89772 37315
rect 96712 37408 96764 37460
rect 94596 37340 94648 37392
rect 89720 37272 89772 37281
rect 93584 37204 93636 37256
rect 95700 37315 95752 37324
rect 95700 37281 95709 37315
rect 95709 37281 95743 37315
rect 95743 37281 95752 37315
rect 95700 37272 95752 37281
rect 95240 37204 95292 37256
rect 70492 37068 70544 37120
rect 72976 37111 73028 37120
rect 72976 37077 72985 37111
rect 72985 37077 73019 37111
rect 73019 37077 73028 37111
rect 72976 37068 73028 37077
rect 76748 37111 76800 37120
rect 76748 37077 76757 37111
rect 76757 37077 76791 37111
rect 76791 37077 76800 37111
rect 76748 37068 76800 37077
rect 78404 37111 78456 37120
rect 78404 37077 78413 37111
rect 78413 37077 78447 37111
rect 78447 37077 78456 37111
rect 78404 37068 78456 37077
rect 84292 37111 84344 37120
rect 84292 37077 84301 37111
rect 84301 37077 84335 37111
rect 84335 37077 84344 37111
rect 84292 37068 84344 37077
rect 85488 37068 85540 37120
rect 87420 37068 87472 37120
rect 89720 37068 89772 37120
rect 93676 37068 93728 37120
rect 95148 37136 95200 37188
rect 95056 37068 95108 37120
rect 97080 37068 97132 37120
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 65686 36966 65738 37018
rect 65750 36966 65802 37018
rect 65814 36966 65866 37018
rect 65878 36966 65930 37018
rect 96406 36966 96458 37018
rect 96470 36966 96522 37018
rect 96534 36966 96586 37018
rect 96598 36966 96650 37018
rect 3240 36864 3292 36916
rect 3700 36796 3752 36848
rect 2504 36771 2556 36780
rect 2504 36737 2513 36771
rect 2513 36737 2547 36771
rect 2547 36737 2556 36771
rect 2504 36728 2556 36737
rect 4620 36728 4672 36780
rect 9772 36796 9824 36848
rect 10048 36839 10100 36848
rect 8760 36728 8812 36780
rect 10048 36805 10057 36839
rect 10057 36805 10091 36839
rect 10091 36805 10100 36839
rect 10048 36796 10100 36805
rect 12716 36907 12768 36916
rect 12716 36873 12725 36907
rect 12725 36873 12759 36907
rect 12759 36873 12768 36907
rect 12716 36864 12768 36873
rect 28816 36864 28868 36916
rect 13544 36796 13596 36848
rect 18420 36796 18472 36848
rect 34796 36864 34848 36916
rect 35440 36864 35492 36916
rect 37004 36907 37056 36916
rect 32036 36839 32088 36848
rect 5448 36660 5500 36712
rect 7104 36660 7156 36712
rect 7656 36703 7708 36712
rect 7656 36669 7665 36703
rect 7665 36669 7699 36703
rect 7699 36669 7708 36703
rect 7656 36660 7708 36669
rect 9588 36660 9640 36712
rect 10232 36728 10284 36780
rect 13268 36728 13320 36780
rect 24952 36771 25004 36780
rect 24952 36737 24961 36771
rect 24961 36737 24995 36771
rect 24995 36737 25004 36771
rect 24952 36728 25004 36737
rect 26792 36728 26844 36780
rect 11428 36660 11480 36712
rect 12348 36660 12400 36712
rect 12900 36660 12952 36712
rect 14004 36703 14056 36712
rect 14004 36669 14013 36703
rect 14013 36669 14047 36703
rect 14047 36669 14056 36703
rect 14004 36660 14056 36669
rect 14096 36660 14148 36712
rect 18880 36660 18932 36712
rect 19064 36703 19116 36712
rect 19064 36669 19073 36703
rect 19073 36669 19107 36703
rect 19107 36669 19116 36703
rect 19064 36660 19116 36669
rect 19340 36703 19392 36712
rect 19340 36669 19349 36703
rect 19349 36669 19383 36703
rect 19383 36669 19392 36703
rect 19340 36660 19392 36669
rect 3976 36592 4028 36644
rect 12256 36592 12308 36644
rect 12808 36592 12860 36644
rect 13636 36592 13688 36644
rect 18972 36592 19024 36644
rect 4620 36524 4672 36576
rect 4896 36524 4948 36576
rect 8576 36524 8628 36576
rect 14188 36524 14240 36576
rect 14280 36524 14332 36576
rect 22284 36660 22336 36712
rect 24308 36703 24360 36712
rect 20076 36592 20128 36644
rect 24308 36669 24317 36703
rect 24317 36669 24351 36703
rect 24351 36669 24360 36703
rect 24308 36660 24360 36669
rect 25044 36703 25096 36712
rect 25044 36669 25053 36703
rect 25053 36669 25087 36703
rect 25087 36669 25096 36703
rect 25044 36660 25096 36669
rect 25412 36703 25464 36712
rect 25412 36669 25421 36703
rect 25421 36669 25455 36703
rect 25455 36669 25464 36703
rect 25412 36660 25464 36669
rect 26424 36635 26476 36644
rect 26424 36601 26433 36635
rect 26433 36601 26467 36635
rect 26467 36601 26476 36635
rect 26424 36592 26476 36601
rect 27160 36660 27212 36712
rect 28632 36728 28684 36780
rect 32036 36805 32045 36839
rect 32045 36805 32079 36839
rect 32079 36805 32088 36839
rect 32036 36796 32088 36805
rect 32128 36728 32180 36780
rect 37004 36873 37013 36907
rect 37013 36873 37047 36907
rect 37047 36873 37056 36907
rect 37004 36864 37056 36873
rect 39488 36864 39540 36916
rect 49792 36864 49844 36916
rect 35716 36796 35768 36848
rect 43168 36796 43220 36848
rect 44180 36839 44232 36848
rect 44180 36805 44189 36839
rect 44189 36805 44223 36839
rect 44223 36805 44232 36839
rect 44180 36796 44232 36805
rect 48044 36796 48096 36848
rect 50436 36796 50488 36848
rect 50712 36839 50764 36848
rect 50712 36805 50721 36839
rect 50721 36805 50755 36839
rect 50755 36805 50764 36839
rect 50712 36796 50764 36805
rect 54944 36864 54996 36916
rect 60740 36864 60792 36916
rect 38108 36728 38160 36780
rect 48504 36728 48556 36780
rect 48688 36771 48740 36780
rect 48688 36737 48697 36771
rect 48697 36737 48731 36771
rect 48731 36737 48740 36771
rect 48688 36728 48740 36737
rect 50804 36771 50856 36780
rect 50804 36737 50813 36771
rect 50813 36737 50847 36771
rect 50847 36737 50856 36771
rect 50804 36728 50856 36737
rect 51172 36771 51224 36780
rect 51172 36737 51181 36771
rect 51181 36737 51215 36771
rect 51215 36737 51224 36771
rect 51172 36728 51224 36737
rect 52460 36728 52512 36780
rect 28724 36660 28776 36712
rect 30380 36660 30432 36712
rect 31852 36660 31904 36712
rect 35992 36703 36044 36712
rect 35992 36669 36001 36703
rect 36001 36669 36035 36703
rect 36035 36669 36044 36703
rect 35992 36660 36044 36669
rect 36452 36660 36504 36712
rect 36728 36703 36780 36712
rect 36728 36669 36737 36703
rect 36737 36669 36771 36703
rect 36771 36669 36780 36703
rect 36728 36660 36780 36669
rect 39304 36703 39356 36712
rect 39304 36669 39313 36703
rect 39313 36669 39347 36703
rect 39347 36669 39356 36703
rect 39304 36660 39356 36669
rect 44456 36660 44508 36712
rect 47308 36703 47360 36712
rect 20628 36567 20680 36576
rect 20628 36533 20637 36567
rect 20637 36533 20671 36567
rect 20671 36533 20680 36567
rect 20628 36524 20680 36533
rect 24492 36567 24544 36576
rect 24492 36533 24501 36567
rect 24501 36533 24535 36567
rect 24535 36533 24544 36567
rect 24492 36524 24544 36533
rect 25136 36524 25188 36576
rect 38568 36592 38620 36644
rect 43352 36592 43404 36644
rect 47308 36669 47317 36703
rect 47317 36669 47351 36703
rect 47351 36669 47360 36703
rect 47308 36660 47360 36669
rect 32772 36567 32824 36576
rect 32772 36533 32781 36567
rect 32781 36533 32815 36567
rect 32815 36533 32824 36567
rect 32772 36524 32824 36533
rect 37832 36524 37884 36576
rect 38660 36524 38712 36576
rect 43260 36524 43312 36576
rect 48320 36524 48372 36576
rect 49240 36660 49292 36712
rect 51448 36660 51500 36712
rect 52736 36703 52788 36712
rect 52736 36669 52745 36703
rect 52745 36669 52779 36703
rect 52779 36669 52788 36703
rect 52736 36660 52788 36669
rect 50896 36592 50948 36644
rect 52460 36635 52512 36644
rect 52460 36601 52469 36635
rect 52469 36601 52503 36635
rect 52503 36601 52512 36635
rect 53840 36660 53892 36712
rect 55036 36728 55088 36780
rect 55312 36771 55364 36780
rect 55312 36737 55321 36771
rect 55321 36737 55355 36771
rect 55355 36737 55364 36771
rect 55312 36728 55364 36737
rect 56048 36796 56100 36848
rect 56600 36839 56652 36848
rect 56600 36805 56609 36839
rect 56609 36805 56643 36839
rect 56643 36805 56652 36839
rect 56600 36796 56652 36805
rect 58256 36796 58308 36848
rect 58532 36796 58584 36848
rect 91008 36864 91060 36916
rect 91284 36864 91336 36916
rect 64420 36839 64472 36848
rect 64420 36805 64429 36839
rect 64429 36805 64463 36839
rect 64463 36805 64472 36839
rect 64420 36796 64472 36805
rect 56692 36728 56744 36780
rect 52460 36592 52512 36601
rect 53748 36592 53800 36644
rect 49148 36524 49200 36576
rect 51724 36524 51776 36576
rect 51908 36524 51960 36576
rect 54116 36567 54168 36576
rect 54116 36533 54125 36567
rect 54125 36533 54159 36567
rect 54159 36533 54168 36567
rect 54116 36524 54168 36533
rect 56324 36703 56376 36712
rect 56324 36669 56333 36703
rect 56333 36669 56367 36703
rect 56367 36669 56376 36703
rect 56784 36703 56836 36712
rect 56324 36660 56376 36669
rect 56784 36669 56793 36703
rect 56793 36669 56827 36703
rect 56827 36669 56836 36703
rect 56784 36660 56836 36669
rect 64788 36771 64840 36780
rect 64788 36737 64797 36771
rect 64797 36737 64831 36771
rect 64831 36737 64840 36771
rect 64788 36728 64840 36737
rect 69020 36728 69072 36780
rect 71044 36771 71096 36780
rect 71044 36737 71053 36771
rect 71053 36737 71087 36771
rect 71087 36737 71096 36771
rect 71044 36728 71096 36737
rect 69296 36703 69348 36712
rect 57888 36592 57940 36644
rect 62120 36592 62172 36644
rect 63132 36592 63184 36644
rect 69296 36669 69305 36703
rect 69305 36669 69339 36703
rect 69339 36669 69348 36703
rect 69296 36660 69348 36669
rect 71780 36796 71832 36848
rect 72976 36796 73028 36848
rect 77300 36771 77352 36780
rect 77300 36737 77309 36771
rect 77309 36737 77343 36771
rect 77343 36737 77352 36771
rect 77300 36728 77352 36737
rect 77484 36728 77536 36780
rect 79232 36728 79284 36780
rect 71412 36703 71464 36712
rect 71412 36669 71421 36703
rect 71421 36669 71455 36703
rect 71455 36669 71464 36703
rect 71412 36660 71464 36669
rect 77392 36660 77444 36712
rect 77668 36660 77720 36712
rect 78404 36660 78456 36712
rect 78772 36660 78824 36712
rect 69756 36592 69808 36644
rect 58624 36524 58676 36576
rect 66076 36567 66128 36576
rect 66076 36533 66085 36567
rect 66085 36533 66119 36567
rect 66119 36533 66128 36567
rect 66076 36524 66128 36533
rect 77300 36524 77352 36576
rect 79784 36635 79836 36644
rect 79784 36601 79793 36635
rect 79793 36601 79827 36635
rect 79827 36601 79836 36635
rect 79784 36592 79836 36601
rect 80060 36567 80112 36576
rect 80060 36533 80069 36567
rect 80069 36533 80103 36567
rect 80103 36533 80112 36567
rect 81716 36567 81768 36576
rect 80060 36524 80112 36533
rect 81716 36533 81725 36567
rect 81725 36533 81759 36567
rect 81759 36533 81768 36567
rect 81716 36524 81768 36533
rect 84292 36524 84344 36576
rect 85212 36796 85264 36848
rect 85580 36839 85632 36848
rect 85580 36805 85589 36839
rect 85589 36805 85623 36839
rect 85623 36805 85632 36839
rect 85580 36796 85632 36805
rect 86224 36771 86276 36780
rect 86224 36737 86233 36771
rect 86233 36737 86267 36771
rect 86267 36737 86276 36771
rect 86224 36728 86276 36737
rect 88432 36728 88484 36780
rect 91284 36728 91336 36780
rect 85488 36660 85540 36712
rect 89168 36592 89220 36644
rect 90180 36635 90232 36644
rect 90180 36601 90189 36635
rect 90189 36601 90223 36635
rect 90223 36601 90232 36635
rect 90180 36592 90232 36601
rect 93400 36864 93452 36916
rect 94044 36864 94096 36916
rect 95332 36864 95384 36916
rect 95240 36728 95292 36780
rect 92756 36592 92808 36644
rect 94688 36703 94740 36712
rect 94688 36669 94697 36703
rect 94697 36669 94731 36703
rect 94731 36669 94740 36703
rect 94964 36703 95016 36712
rect 94688 36660 94740 36669
rect 94964 36669 94973 36703
rect 94973 36669 95007 36703
rect 95007 36669 95016 36703
rect 94964 36660 95016 36669
rect 95056 36703 95108 36712
rect 95056 36669 95065 36703
rect 95065 36669 95099 36703
rect 95099 36669 95108 36703
rect 95056 36660 95108 36669
rect 95332 36660 95384 36712
rect 97264 36703 97316 36712
rect 97264 36669 97273 36703
rect 97273 36669 97307 36703
rect 97307 36669 97316 36703
rect 97264 36660 97316 36669
rect 90916 36524 90968 36576
rect 94688 36524 94740 36576
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 50326 36422 50378 36474
rect 50390 36422 50442 36474
rect 50454 36422 50506 36474
rect 50518 36422 50570 36474
rect 81046 36422 81098 36474
rect 81110 36422 81162 36474
rect 81174 36422 81226 36474
rect 81238 36422 81290 36474
rect 8944 36363 8996 36372
rect 8944 36329 8953 36363
rect 8953 36329 8987 36363
rect 8987 36329 8996 36363
rect 8944 36320 8996 36329
rect 11796 36363 11848 36372
rect 11796 36329 11805 36363
rect 11805 36329 11839 36363
rect 11839 36329 11848 36363
rect 11796 36320 11848 36329
rect 5080 36252 5132 36304
rect 24492 36320 24544 36372
rect 24768 36320 24820 36372
rect 26240 36320 26292 36372
rect 26976 36320 27028 36372
rect 12900 36252 12952 36304
rect 8576 36227 8628 36236
rect 8576 36193 8585 36227
rect 8585 36193 8619 36227
rect 8619 36193 8628 36227
rect 8576 36184 8628 36193
rect 8944 36184 8996 36236
rect 11796 36184 11848 36236
rect 12992 36184 13044 36236
rect 7748 36159 7800 36168
rect 7748 36125 7757 36159
rect 7757 36125 7791 36159
rect 7791 36125 7800 36159
rect 7748 36116 7800 36125
rect 8668 36116 8720 36168
rect 13176 36159 13228 36168
rect 13176 36125 13185 36159
rect 13185 36125 13219 36159
rect 13219 36125 13228 36159
rect 13176 36116 13228 36125
rect 6000 36048 6052 36100
rect 8760 35980 8812 36032
rect 12348 36048 12400 36100
rect 12532 36048 12584 36100
rect 12716 36091 12768 36100
rect 12716 36057 12725 36091
rect 12725 36057 12759 36091
rect 12759 36057 12768 36091
rect 12716 36048 12768 36057
rect 24400 36252 24452 36304
rect 13912 36184 13964 36236
rect 18420 36227 18472 36236
rect 18420 36193 18429 36227
rect 18429 36193 18463 36227
rect 18463 36193 18472 36227
rect 18420 36184 18472 36193
rect 20904 36227 20956 36236
rect 14188 36091 14240 36100
rect 14188 36057 14197 36091
rect 14197 36057 14231 36091
rect 14231 36057 14240 36091
rect 14188 36048 14240 36057
rect 15568 36048 15620 36100
rect 13912 36023 13964 36032
rect 13912 35989 13921 36023
rect 13921 35989 13955 36023
rect 13955 35989 13964 36023
rect 13912 35980 13964 35989
rect 17316 35980 17368 36032
rect 20904 36193 20913 36227
rect 20913 36193 20947 36227
rect 20947 36193 20956 36227
rect 20904 36184 20956 36193
rect 24124 36227 24176 36236
rect 24124 36193 24133 36227
rect 24133 36193 24167 36227
rect 24167 36193 24176 36227
rect 24124 36184 24176 36193
rect 25044 36184 25096 36236
rect 25412 36184 25464 36236
rect 26976 36227 27028 36236
rect 26976 36193 26985 36227
rect 26985 36193 27019 36227
rect 27019 36193 27028 36227
rect 26976 36184 27028 36193
rect 18788 36091 18840 36100
rect 18788 36057 18797 36091
rect 18797 36057 18831 36091
rect 18831 36057 18840 36091
rect 18788 36048 18840 36057
rect 18880 36048 18932 36100
rect 20168 36048 20220 36100
rect 18144 35980 18196 36032
rect 19248 35980 19300 36032
rect 20076 35980 20128 36032
rect 20720 36116 20772 36168
rect 25136 36116 25188 36168
rect 23848 36048 23900 36100
rect 25412 36048 25464 36100
rect 27160 36048 27212 36100
rect 28448 35980 28500 36032
rect 29092 36320 29144 36372
rect 29644 36320 29696 36372
rect 29368 36184 29420 36236
rect 29552 36227 29604 36236
rect 29552 36193 29561 36227
rect 29561 36193 29595 36227
rect 29595 36193 29604 36227
rect 29552 36184 29604 36193
rect 31944 36184 31996 36236
rect 32128 36227 32180 36236
rect 32128 36193 32137 36227
rect 32137 36193 32171 36227
rect 32171 36193 32180 36227
rect 32128 36184 32180 36193
rect 35624 36227 35676 36236
rect 35624 36193 35633 36227
rect 35633 36193 35667 36227
rect 35667 36193 35676 36227
rect 36452 36252 36504 36304
rect 47308 36320 47360 36372
rect 43444 36252 43496 36304
rect 44916 36252 44968 36304
rect 51816 36320 51868 36372
rect 54852 36320 54904 36372
rect 60740 36320 60792 36372
rect 60832 36320 60884 36372
rect 63316 36320 63368 36372
rect 71504 36363 71556 36372
rect 71504 36329 71513 36363
rect 71513 36329 71547 36363
rect 71547 36329 71556 36363
rect 71504 36320 71556 36329
rect 83740 36320 83792 36372
rect 50712 36295 50764 36304
rect 50712 36261 50721 36295
rect 50721 36261 50755 36295
rect 50755 36261 50764 36295
rect 50712 36252 50764 36261
rect 51080 36252 51132 36304
rect 53380 36252 53432 36304
rect 35624 36184 35676 36193
rect 31760 36116 31812 36168
rect 29644 36048 29696 36100
rect 30104 36048 30156 36100
rect 35348 36116 35400 36168
rect 38108 36184 38160 36236
rect 39396 36184 39448 36236
rect 42800 36184 42852 36236
rect 43352 36227 43404 36236
rect 43352 36193 43361 36227
rect 43361 36193 43395 36227
rect 43395 36193 43404 36227
rect 43352 36184 43404 36193
rect 49976 36184 50028 36236
rect 50160 36227 50212 36236
rect 50160 36193 50169 36227
rect 50169 36193 50203 36227
rect 50203 36193 50212 36227
rect 50160 36184 50212 36193
rect 50344 36227 50396 36236
rect 50344 36193 50353 36227
rect 50353 36193 50387 36227
rect 50387 36193 50396 36227
rect 50344 36184 50396 36193
rect 51632 36184 51684 36236
rect 52736 36184 52788 36236
rect 54116 36184 54168 36236
rect 38936 36116 38988 36168
rect 43628 36159 43680 36168
rect 43628 36125 43637 36159
rect 43637 36125 43671 36159
rect 43671 36125 43680 36159
rect 43628 36116 43680 36125
rect 30564 35980 30616 36032
rect 35348 36023 35400 36032
rect 35348 35989 35357 36023
rect 35357 35989 35391 36023
rect 35391 35989 35400 36023
rect 35348 35980 35400 35989
rect 48780 35980 48832 36032
rect 49516 35980 49568 36032
rect 50344 35980 50396 36032
rect 51172 36023 51224 36032
rect 51172 35989 51181 36023
rect 51181 35989 51215 36023
rect 51215 35989 51224 36023
rect 51172 35980 51224 35989
rect 55956 36023 56008 36032
rect 55956 35989 55965 36023
rect 55965 35989 55999 36023
rect 55999 35989 56008 36023
rect 55956 35980 56008 35989
rect 56232 36023 56284 36032
rect 56232 35989 56241 36023
rect 56241 35989 56275 36023
rect 56275 35989 56284 36023
rect 56232 35980 56284 35989
rect 56600 36184 56652 36236
rect 58532 36227 58584 36236
rect 58532 36193 58541 36227
rect 58541 36193 58575 36227
rect 58575 36193 58584 36227
rect 58532 36184 58584 36193
rect 58624 36184 58676 36236
rect 57796 36159 57848 36168
rect 57796 36125 57805 36159
rect 57805 36125 57839 36159
rect 57839 36125 57848 36159
rect 57796 36116 57848 36125
rect 59820 36116 59872 36168
rect 62672 36159 62724 36168
rect 62672 36125 62681 36159
rect 62681 36125 62715 36159
rect 62715 36125 62724 36159
rect 62672 36116 62724 36125
rect 63132 36159 63184 36168
rect 63132 36125 63141 36159
rect 63141 36125 63175 36159
rect 63175 36125 63184 36159
rect 63132 36116 63184 36125
rect 63316 36227 63368 36236
rect 63316 36193 63325 36227
rect 63325 36193 63359 36227
rect 63359 36193 63368 36227
rect 63316 36184 63368 36193
rect 63868 36227 63920 36236
rect 63500 36116 63552 36168
rect 63868 36193 63877 36227
rect 63877 36193 63911 36227
rect 63911 36193 63920 36227
rect 63868 36184 63920 36193
rect 66076 36184 66128 36236
rect 71320 36184 71372 36236
rect 71780 36184 71832 36236
rect 72332 36184 72384 36236
rect 73068 36227 73120 36236
rect 73068 36193 73077 36227
rect 73077 36193 73111 36227
rect 73111 36193 73120 36227
rect 73068 36184 73120 36193
rect 64420 36116 64472 36168
rect 70492 36116 70544 36168
rect 73160 36116 73212 36168
rect 58440 35980 58492 36032
rect 58624 35980 58676 36032
rect 58808 36023 58860 36032
rect 58808 35989 58817 36023
rect 58817 35989 58851 36023
rect 58851 35989 58860 36023
rect 58808 35980 58860 35989
rect 70216 35980 70268 36032
rect 71504 35980 71556 36032
rect 73252 36023 73304 36032
rect 73252 35989 73261 36023
rect 73261 35989 73295 36023
rect 73295 35989 73304 36023
rect 73252 35980 73304 35989
rect 77668 36252 77720 36304
rect 80060 36252 80112 36304
rect 81716 36252 81768 36304
rect 77576 36227 77628 36236
rect 77576 36193 77585 36227
rect 77585 36193 77619 36227
rect 77619 36193 77628 36227
rect 77576 36184 77628 36193
rect 75920 36116 75972 36168
rect 77852 36116 77904 36168
rect 78036 36116 78088 36168
rect 77944 35980 77996 36032
rect 78772 36184 78824 36236
rect 79232 36227 79284 36236
rect 79232 36193 79241 36227
rect 79241 36193 79275 36227
rect 79275 36193 79284 36227
rect 79232 36184 79284 36193
rect 84476 36227 84528 36236
rect 78312 36116 78364 36168
rect 84476 36193 84485 36227
rect 84485 36193 84519 36227
rect 84519 36193 84528 36227
rect 84476 36184 84528 36193
rect 97264 36363 97316 36372
rect 97264 36329 97273 36363
rect 97273 36329 97307 36363
rect 97307 36329 97316 36363
rect 97264 36320 97316 36329
rect 88432 36252 88484 36304
rect 79600 36023 79652 36032
rect 79600 35989 79609 36023
rect 79609 35989 79643 36023
rect 79643 35989 79652 36023
rect 79600 35980 79652 35989
rect 82544 35980 82596 36032
rect 86224 36116 86276 36168
rect 89720 36184 89772 36236
rect 91744 36184 91796 36236
rect 92756 36227 92808 36236
rect 92756 36193 92765 36227
rect 92765 36193 92799 36227
rect 92799 36193 92808 36227
rect 92756 36184 92808 36193
rect 97080 36227 97132 36236
rect 97080 36193 97089 36227
rect 97089 36193 97123 36227
rect 97123 36193 97132 36227
rect 97080 36184 97132 36193
rect 90732 36116 90784 36168
rect 94596 36159 94648 36168
rect 86776 36023 86828 36032
rect 86776 35989 86785 36023
rect 86785 35989 86819 36023
rect 86819 35989 86828 36023
rect 86776 35980 86828 35989
rect 89536 35980 89588 36032
rect 90640 36023 90692 36032
rect 90640 35989 90649 36023
rect 90649 35989 90683 36023
rect 90683 35989 90692 36023
rect 90640 35980 90692 35989
rect 93952 35980 94004 36032
rect 94596 36125 94605 36159
rect 94605 36125 94639 36159
rect 94639 36125 94648 36159
rect 94596 36116 94648 36125
rect 96712 35980 96764 36032
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 65686 35878 65738 35930
rect 65750 35878 65802 35930
rect 65814 35878 65866 35930
rect 65878 35878 65930 35930
rect 96406 35878 96458 35930
rect 96470 35878 96522 35930
rect 96534 35878 96586 35930
rect 96598 35878 96650 35930
rect 5172 35708 5224 35760
rect 2872 35640 2924 35692
rect 7748 35640 7800 35692
rect 4160 35572 4212 35624
rect 5540 35572 5592 35624
rect 5724 35615 5776 35624
rect 5724 35581 5733 35615
rect 5733 35581 5767 35615
rect 5767 35581 5776 35615
rect 5724 35572 5776 35581
rect 7104 35615 7156 35624
rect 7104 35581 7113 35615
rect 7113 35581 7147 35615
rect 7147 35581 7156 35615
rect 7104 35572 7156 35581
rect 10876 35572 10928 35624
rect 3976 35504 4028 35556
rect 3240 35436 3292 35488
rect 4160 35436 4212 35488
rect 4712 35436 4764 35488
rect 9588 35504 9640 35556
rect 15200 35708 15252 35760
rect 12808 35683 12860 35692
rect 12808 35649 12817 35683
rect 12817 35649 12851 35683
rect 12851 35649 12860 35683
rect 12808 35640 12860 35649
rect 11428 35572 11480 35624
rect 14004 35640 14056 35692
rect 17960 35640 18012 35692
rect 18788 35640 18840 35692
rect 20904 35776 20956 35828
rect 25412 35776 25464 35828
rect 25504 35776 25556 35828
rect 57888 35776 57940 35828
rect 70492 35776 70544 35828
rect 71044 35776 71096 35828
rect 73068 35776 73120 35828
rect 77668 35776 77720 35828
rect 77944 35819 77996 35828
rect 77944 35785 77968 35819
rect 77968 35785 77996 35819
rect 77944 35776 77996 35785
rect 79784 35776 79836 35828
rect 86868 35776 86920 35828
rect 20720 35751 20772 35760
rect 20720 35717 20729 35751
rect 20729 35717 20763 35751
rect 20763 35717 20772 35751
rect 20720 35708 20772 35717
rect 25136 35708 25188 35760
rect 30288 35708 30340 35760
rect 32128 35751 32180 35760
rect 32128 35717 32137 35751
rect 32137 35717 32171 35751
rect 32171 35717 32180 35751
rect 32128 35708 32180 35717
rect 32772 35708 32824 35760
rect 42800 35751 42852 35760
rect 42800 35717 42809 35751
rect 42809 35717 42843 35751
rect 42843 35717 42852 35751
rect 42800 35708 42852 35717
rect 42892 35708 42944 35760
rect 44456 35751 44508 35760
rect 44456 35717 44465 35751
rect 44465 35717 44499 35751
rect 44499 35717 44508 35751
rect 44456 35708 44508 35717
rect 24124 35640 24176 35692
rect 10876 35479 10928 35488
rect 10876 35445 10885 35479
rect 10885 35445 10919 35479
rect 10919 35445 10928 35479
rect 10876 35436 10928 35445
rect 13636 35615 13688 35624
rect 13636 35581 13645 35615
rect 13645 35581 13679 35615
rect 13679 35581 13688 35615
rect 15200 35615 15252 35624
rect 13636 35572 13688 35581
rect 15200 35581 15209 35615
rect 15209 35581 15243 35615
rect 15243 35581 15252 35615
rect 15200 35572 15252 35581
rect 15568 35615 15620 35624
rect 15568 35581 15577 35615
rect 15577 35581 15611 35615
rect 15611 35581 15620 35615
rect 15568 35572 15620 35581
rect 13452 35504 13504 35556
rect 13820 35479 13872 35488
rect 13820 35445 13829 35479
rect 13829 35445 13863 35479
rect 13863 35445 13872 35479
rect 13820 35436 13872 35445
rect 14004 35479 14056 35488
rect 14004 35445 14013 35479
rect 14013 35445 14047 35479
rect 14047 35445 14056 35479
rect 14004 35436 14056 35445
rect 19064 35572 19116 35624
rect 19984 35572 20036 35624
rect 20628 35615 20680 35624
rect 20628 35581 20637 35615
rect 20637 35581 20671 35615
rect 20671 35581 20680 35615
rect 20628 35572 20680 35581
rect 19156 35504 19208 35556
rect 25136 35572 25188 35624
rect 26792 35615 26844 35624
rect 19432 35436 19484 35488
rect 19984 35436 20036 35488
rect 21824 35436 21876 35488
rect 25044 35436 25096 35488
rect 26792 35581 26801 35615
rect 26801 35581 26835 35615
rect 26835 35581 26844 35615
rect 26792 35572 26844 35581
rect 26976 35640 27028 35692
rect 30564 35683 30616 35692
rect 27160 35615 27212 35624
rect 27160 35581 27169 35615
rect 27169 35581 27203 35615
rect 27203 35581 27212 35615
rect 27160 35572 27212 35581
rect 28908 35572 28960 35624
rect 29092 35572 29144 35624
rect 30564 35649 30573 35683
rect 30573 35649 30607 35683
rect 30607 35649 30616 35683
rect 30564 35640 30616 35649
rect 35348 35683 35400 35692
rect 35348 35649 35357 35683
rect 35357 35649 35391 35683
rect 35391 35649 35400 35683
rect 35348 35640 35400 35649
rect 30104 35504 30156 35556
rect 26516 35436 26568 35488
rect 26608 35436 26660 35488
rect 30196 35436 30248 35488
rect 31300 35572 31352 35624
rect 42616 35640 42668 35692
rect 44088 35640 44140 35692
rect 49792 35708 49844 35760
rect 51356 35708 51408 35760
rect 54576 35708 54628 35760
rect 48780 35640 48832 35692
rect 36176 35572 36228 35624
rect 36452 35572 36504 35624
rect 39672 35572 39724 35624
rect 42800 35572 42852 35624
rect 41236 35504 41288 35556
rect 42064 35504 42116 35556
rect 48872 35504 48924 35556
rect 49240 35572 49292 35624
rect 54944 35640 54996 35692
rect 55128 35708 55180 35760
rect 56600 35640 56652 35692
rect 57520 35708 57572 35760
rect 56968 35683 57020 35692
rect 56968 35649 56977 35683
rect 56977 35649 57011 35683
rect 57011 35649 57020 35683
rect 58624 35683 58676 35692
rect 56968 35640 57020 35649
rect 49976 35572 50028 35624
rect 50712 35572 50764 35624
rect 55220 35615 55272 35624
rect 55220 35581 55229 35615
rect 55229 35581 55263 35615
rect 55263 35581 55272 35615
rect 55220 35572 55272 35581
rect 50896 35547 50948 35556
rect 50896 35513 50905 35547
rect 50905 35513 50939 35547
rect 50939 35513 50948 35547
rect 50896 35504 50948 35513
rect 51724 35547 51776 35556
rect 51724 35513 51732 35547
rect 51732 35513 51766 35547
rect 51766 35513 51776 35547
rect 51724 35504 51776 35513
rect 54484 35504 54536 35556
rect 55772 35615 55824 35624
rect 55772 35581 55781 35615
rect 55781 35581 55815 35615
rect 55815 35581 55824 35615
rect 55772 35572 55824 35581
rect 31760 35436 31812 35488
rect 31944 35436 31996 35488
rect 34612 35436 34664 35488
rect 35348 35436 35400 35488
rect 36268 35436 36320 35488
rect 42984 35436 43036 35488
rect 48780 35479 48832 35488
rect 48780 35445 48789 35479
rect 48789 35445 48823 35479
rect 48823 35445 48832 35479
rect 48780 35436 48832 35445
rect 48964 35479 49016 35488
rect 48964 35445 48973 35479
rect 48973 35445 49007 35479
rect 49007 35445 49016 35479
rect 48964 35436 49016 35445
rect 50712 35479 50764 35488
rect 50712 35445 50721 35479
rect 50721 35445 50755 35479
rect 50755 35445 50764 35479
rect 50712 35436 50764 35445
rect 51172 35436 51224 35488
rect 52000 35436 52052 35488
rect 52368 35479 52420 35488
rect 52368 35445 52377 35479
rect 52377 35445 52411 35479
rect 52411 35445 52420 35479
rect 52368 35436 52420 35445
rect 54576 35436 54628 35488
rect 57520 35615 57572 35624
rect 57520 35581 57529 35615
rect 57529 35581 57563 35615
rect 57563 35581 57572 35615
rect 57520 35572 57572 35581
rect 58624 35649 58633 35683
rect 58633 35649 58667 35683
rect 58667 35649 58676 35683
rect 58624 35640 58676 35649
rect 63500 35708 63552 35760
rect 63684 35751 63736 35760
rect 63684 35717 63693 35751
rect 63693 35717 63727 35751
rect 63727 35717 63736 35751
rect 63684 35708 63736 35717
rect 66260 35683 66312 35692
rect 66260 35649 66269 35683
rect 66269 35649 66303 35683
rect 66303 35649 66312 35683
rect 68744 35708 68796 35760
rect 77576 35708 77628 35760
rect 84476 35708 84528 35760
rect 66260 35640 66312 35649
rect 59084 35615 59136 35624
rect 56140 35504 56192 35556
rect 59084 35581 59093 35615
rect 59093 35581 59127 35615
rect 59127 35581 59136 35615
rect 59084 35572 59136 35581
rect 63316 35572 63368 35624
rect 64420 35615 64472 35624
rect 64420 35581 64429 35615
rect 64429 35581 64463 35615
rect 64463 35581 64472 35615
rect 64420 35572 64472 35581
rect 64604 35615 64656 35624
rect 64604 35581 64613 35615
rect 64613 35581 64647 35615
rect 64647 35581 64656 35615
rect 64604 35572 64656 35581
rect 58900 35479 58952 35488
rect 58900 35445 58909 35479
rect 58909 35445 58943 35479
rect 58943 35445 58952 35479
rect 58900 35436 58952 35445
rect 62028 35436 62080 35488
rect 70216 35640 70268 35692
rect 77484 35640 77536 35692
rect 68560 35572 68612 35624
rect 69112 35615 69164 35624
rect 69112 35581 69115 35615
rect 69115 35581 69149 35615
rect 69149 35581 69164 35615
rect 69112 35572 69164 35581
rect 71412 35572 71464 35624
rect 74264 35572 74316 35624
rect 75920 35572 75972 35624
rect 76288 35572 76340 35624
rect 76656 35572 76708 35624
rect 77392 35572 77444 35624
rect 77944 35572 77996 35624
rect 83740 35615 83792 35624
rect 83740 35581 83749 35615
rect 83749 35581 83783 35615
rect 83783 35581 83792 35615
rect 83740 35572 83792 35581
rect 65984 35504 66036 35556
rect 68652 35504 68704 35556
rect 66076 35479 66128 35488
rect 66076 35445 66085 35479
rect 66085 35445 66119 35479
rect 66119 35445 66128 35479
rect 66076 35436 66128 35445
rect 66168 35436 66220 35488
rect 69848 35436 69900 35488
rect 70492 35436 70544 35488
rect 70584 35479 70636 35488
rect 70584 35445 70593 35479
rect 70593 35445 70627 35479
rect 70627 35445 70636 35479
rect 76564 35504 76616 35556
rect 77668 35547 77720 35556
rect 77668 35513 77677 35547
rect 77677 35513 77711 35547
rect 77711 35513 77720 35547
rect 77668 35504 77720 35513
rect 78772 35504 78824 35556
rect 79784 35547 79836 35556
rect 79784 35513 79793 35547
rect 79793 35513 79827 35547
rect 79827 35513 79836 35547
rect 79784 35504 79836 35513
rect 85396 35547 85448 35556
rect 85396 35513 85405 35547
rect 85405 35513 85439 35547
rect 85439 35513 85448 35547
rect 85396 35504 85448 35513
rect 85856 35708 85908 35760
rect 94044 35708 94096 35760
rect 85764 35683 85816 35692
rect 85764 35649 85773 35683
rect 85773 35649 85807 35683
rect 85807 35649 85816 35683
rect 85764 35640 85816 35649
rect 88432 35683 88484 35692
rect 88432 35649 88441 35683
rect 88441 35649 88475 35683
rect 88475 35649 88484 35683
rect 88432 35640 88484 35649
rect 86776 35572 86828 35624
rect 88156 35615 88208 35624
rect 88156 35581 88165 35615
rect 88165 35581 88199 35615
rect 88199 35581 88208 35615
rect 88156 35572 88208 35581
rect 88248 35572 88300 35624
rect 70584 35436 70636 35445
rect 79508 35436 79560 35488
rect 80152 35436 80204 35488
rect 84292 35436 84344 35488
rect 88984 35436 89036 35488
rect 89720 35683 89772 35692
rect 89720 35649 89729 35683
rect 89729 35649 89763 35683
rect 89763 35649 89772 35683
rect 90732 35683 90784 35692
rect 89720 35640 89772 35649
rect 90732 35649 90741 35683
rect 90741 35649 90775 35683
rect 90775 35649 90784 35683
rect 90732 35640 90784 35649
rect 91284 35615 91336 35624
rect 91284 35581 91293 35615
rect 91293 35581 91327 35615
rect 91327 35581 91336 35615
rect 91284 35572 91336 35581
rect 93676 35615 93728 35624
rect 93676 35581 93685 35615
rect 93685 35581 93719 35615
rect 93719 35581 93728 35615
rect 95240 35683 95292 35692
rect 95240 35649 95249 35683
rect 95249 35649 95283 35683
rect 95283 35649 95292 35683
rect 95240 35640 95292 35649
rect 94964 35615 95016 35624
rect 93676 35572 93728 35581
rect 94136 35504 94188 35556
rect 91284 35436 91336 35488
rect 94044 35436 94096 35488
rect 94964 35581 94973 35615
rect 94973 35581 95007 35615
rect 95007 35581 95016 35615
rect 94964 35572 95016 35581
rect 96712 35572 96764 35624
rect 95056 35504 95108 35556
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 50326 35334 50378 35386
rect 50390 35334 50442 35386
rect 50454 35334 50506 35386
rect 50518 35334 50570 35386
rect 81046 35334 81098 35386
rect 81110 35334 81162 35386
rect 81174 35334 81226 35386
rect 81238 35334 81290 35386
rect 5816 35275 5868 35284
rect 5816 35241 5825 35275
rect 5825 35241 5859 35275
rect 5859 35241 5868 35275
rect 5816 35232 5868 35241
rect 7380 35275 7432 35284
rect 7380 35241 7389 35275
rect 7389 35241 7423 35275
rect 7423 35241 7432 35275
rect 7380 35232 7432 35241
rect 13912 35232 13964 35284
rect 15016 35232 15068 35284
rect 19156 35232 19208 35284
rect 19340 35232 19392 35284
rect 3884 35164 3936 35216
rect 9956 35164 10008 35216
rect 12900 35207 12952 35216
rect 12900 35173 12909 35207
rect 12909 35173 12943 35207
rect 12943 35173 12952 35207
rect 12900 35164 12952 35173
rect 5540 35096 5592 35148
rect 6276 35139 6328 35148
rect 6276 35105 6285 35139
rect 6285 35105 6319 35139
rect 6319 35105 6328 35139
rect 6276 35096 6328 35105
rect 7104 35096 7156 35148
rect 13452 35096 13504 35148
rect 13820 35164 13872 35216
rect 19708 35164 19760 35216
rect 14004 35096 14056 35148
rect 14464 35096 14516 35148
rect 18328 35096 18380 35148
rect 20720 35232 20772 35284
rect 22192 35232 22244 35284
rect 25320 35232 25372 35284
rect 30380 35275 30432 35284
rect 21824 35139 21876 35148
rect 21824 35105 21833 35139
rect 21833 35105 21867 35139
rect 21867 35105 21876 35139
rect 21824 35096 21876 35105
rect 3608 35028 3660 35080
rect 9404 35028 9456 35080
rect 14648 35071 14700 35080
rect 14648 35037 14657 35071
rect 14657 35037 14691 35071
rect 14691 35037 14700 35071
rect 14648 35028 14700 35037
rect 3424 34960 3476 35012
rect 3792 34960 3844 35012
rect 13912 34960 13964 35012
rect 4068 34892 4120 34944
rect 15660 34892 15712 34944
rect 17316 34892 17368 34944
rect 22376 35096 22428 35148
rect 24308 35139 24360 35148
rect 24308 35105 24317 35139
rect 24317 35105 24351 35139
rect 24351 35105 24360 35139
rect 24308 35096 24360 35105
rect 25320 35139 25372 35148
rect 25320 35105 25329 35139
rect 25329 35105 25363 35139
rect 25363 35105 25372 35139
rect 25320 35096 25372 35105
rect 28080 35139 28132 35148
rect 28080 35105 28089 35139
rect 28089 35105 28123 35139
rect 28123 35105 28132 35139
rect 28080 35096 28132 35105
rect 28448 35096 28500 35148
rect 18144 34960 18196 35012
rect 22100 35071 22152 35080
rect 22100 35037 22109 35071
rect 22109 35037 22143 35071
rect 22143 35037 22152 35071
rect 22100 35028 22152 35037
rect 22284 35028 22336 35080
rect 22836 35028 22888 35080
rect 22928 35028 22980 35080
rect 25044 34960 25096 35012
rect 18788 34892 18840 34944
rect 22284 34892 22336 34944
rect 23388 34935 23440 34944
rect 23388 34901 23397 34935
rect 23397 34901 23431 34935
rect 23431 34901 23440 34935
rect 23388 34892 23440 34901
rect 23664 34935 23716 34944
rect 23664 34901 23673 34935
rect 23673 34901 23707 34935
rect 23707 34901 23716 34935
rect 29092 34960 29144 35012
rect 23664 34892 23716 34901
rect 26056 34892 26108 34944
rect 27620 34892 27672 34944
rect 28080 34892 28132 34944
rect 28448 34892 28500 34944
rect 30380 35241 30389 35275
rect 30389 35241 30423 35275
rect 30423 35241 30432 35275
rect 30380 35232 30432 35241
rect 30472 35232 30524 35284
rect 31300 35164 31352 35216
rect 30104 35139 30156 35148
rect 30104 35105 30113 35139
rect 30113 35105 30147 35139
rect 30147 35105 30156 35139
rect 30104 35096 30156 35105
rect 30288 35096 30340 35148
rect 32312 35139 32364 35148
rect 31668 35028 31720 35080
rect 31760 35071 31812 35080
rect 31760 35037 31769 35071
rect 31769 35037 31803 35071
rect 31803 35037 31812 35071
rect 31760 35028 31812 35037
rect 32312 35105 32340 35139
rect 32340 35105 32364 35139
rect 32312 35096 32364 35105
rect 32864 35139 32916 35148
rect 32864 35105 32873 35139
rect 32873 35105 32907 35139
rect 32907 35105 32916 35139
rect 32864 35096 32916 35105
rect 33324 35096 33376 35148
rect 36268 35139 36320 35148
rect 36268 35105 36277 35139
rect 36277 35105 36311 35139
rect 36311 35105 36320 35139
rect 36268 35096 36320 35105
rect 33876 35071 33928 35080
rect 33876 35037 33885 35071
rect 33885 35037 33919 35071
rect 33919 35037 33928 35071
rect 33876 35028 33928 35037
rect 35624 35071 35676 35080
rect 35624 35037 35633 35071
rect 35633 35037 35667 35071
rect 35667 35037 35676 35071
rect 35624 35028 35676 35037
rect 38936 35232 38988 35284
rect 40500 35232 40552 35284
rect 42892 35232 42944 35284
rect 43996 35232 44048 35284
rect 36820 35164 36872 35216
rect 41696 35164 41748 35216
rect 42984 35164 43036 35216
rect 36636 35139 36688 35148
rect 36636 35105 36650 35139
rect 36650 35105 36688 35139
rect 36636 35096 36688 35105
rect 36728 35139 36780 35148
rect 36728 35105 36737 35139
rect 36737 35105 36771 35139
rect 36771 35105 36780 35139
rect 36728 35096 36780 35105
rect 37280 35096 37332 35148
rect 38016 35139 38068 35148
rect 37004 35071 37056 35080
rect 37004 35037 37013 35071
rect 37013 35037 37047 35071
rect 37047 35037 37056 35071
rect 37004 35028 37056 35037
rect 38016 35105 38025 35139
rect 38025 35105 38059 35139
rect 38059 35105 38068 35139
rect 38016 35096 38068 35105
rect 38660 35096 38712 35148
rect 39580 35139 39632 35148
rect 39580 35105 39589 35139
rect 39589 35105 39623 35139
rect 39623 35105 39632 35139
rect 39580 35096 39632 35105
rect 40592 35139 40644 35148
rect 40592 35105 40601 35139
rect 40601 35105 40635 35139
rect 40635 35105 40644 35139
rect 40592 35096 40644 35105
rect 41788 35139 41840 35148
rect 41788 35105 41797 35139
rect 41797 35105 41831 35139
rect 41831 35105 41840 35139
rect 41788 35096 41840 35105
rect 44088 35164 44140 35216
rect 38752 34960 38804 35012
rect 31668 34892 31720 34944
rect 33508 34892 33560 34944
rect 33600 34892 33652 34944
rect 37096 34892 37148 34944
rect 37280 34935 37332 34944
rect 37280 34901 37289 34935
rect 37289 34901 37323 34935
rect 37323 34901 37332 34935
rect 37280 34892 37332 34901
rect 40960 35071 41012 35080
rect 40960 35037 40969 35071
rect 40969 35037 41003 35071
rect 41003 35037 41012 35071
rect 40960 35028 41012 35037
rect 43444 35071 43496 35080
rect 43444 35037 43453 35071
rect 43453 35037 43487 35071
rect 43487 35037 43496 35071
rect 43444 35028 43496 35037
rect 44364 35139 44416 35148
rect 44364 35105 44373 35139
rect 44373 35105 44407 35139
rect 44407 35105 44416 35139
rect 44364 35096 44416 35105
rect 46572 35164 46624 35216
rect 48044 35232 48096 35284
rect 49884 35232 49936 35284
rect 49976 35232 50028 35284
rect 51632 35275 51684 35284
rect 47768 35164 47820 35216
rect 44180 35028 44232 35080
rect 46756 35028 46808 35080
rect 44272 34960 44324 35012
rect 49148 35096 49200 35148
rect 49608 35096 49660 35148
rect 48872 35028 48924 35080
rect 49976 35028 50028 35080
rect 50252 35139 50304 35148
rect 50252 35105 50261 35139
rect 50261 35105 50295 35139
rect 50295 35105 50304 35139
rect 51632 35241 51641 35275
rect 51641 35241 51675 35275
rect 51675 35241 51684 35275
rect 51632 35232 51684 35241
rect 52000 35232 52052 35284
rect 56140 35232 56192 35284
rect 56324 35275 56376 35284
rect 56324 35241 56333 35275
rect 56333 35241 56367 35275
rect 56367 35241 56376 35275
rect 56324 35232 56376 35241
rect 56508 35232 56560 35284
rect 52368 35164 52420 35216
rect 57980 35164 58032 35216
rect 58808 35164 58860 35216
rect 59820 35232 59872 35284
rect 64604 35164 64656 35216
rect 50252 35096 50304 35105
rect 53288 35139 53340 35148
rect 53288 35105 53297 35139
rect 53297 35105 53331 35139
rect 53331 35105 53340 35139
rect 53288 35096 53340 35105
rect 53840 35096 53892 35148
rect 55772 35096 55824 35148
rect 51356 35071 51408 35080
rect 51356 35037 51365 35071
rect 51365 35037 51399 35071
rect 51399 35037 51408 35071
rect 51356 35028 51408 35037
rect 51816 35071 51868 35080
rect 51816 35037 51825 35071
rect 51825 35037 51859 35071
rect 51859 35037 51868 35071
rect 51816 35028 51868 35037
rect 52000 35028 52052 35080
rect 56140 35028 56192 35080
rect 56416 35028 56468 35080
rect 56968 35139 57020 35148
rect 56968 35105 56977 35139
rect 56977 35105 57011 35139
rect 57011 35105 57020 35139
rect 56968 35096 57020 35105
rect 58440 35096 58492 35148
rect 58624 35096 58676 35148
rect 62764 35139 62816 35148
rect 57980 35028 58032 35080
rect 61200 35028 61252 35080
rect 46572 34935 46624 34944
rect 46572 34901 46581 34935
rect 46581 34901 46615 34935
rect 46615 34901 46624 34935
rect 46572 34892 46624 34901
rect 46756 34935 46808 34944
rect 46756 34901 46765 34935
rect 46765 34901 46799 34935
rect 46799 34901 46808 34935
rect 46756 34892 46808 34901
rect 46848 34892 46900 34944
rect 49424 34892 49476 34944
rect 49608 34892 49660 34944
rect 62028 34960 62080 35012
rect 52000 34892 52052 34944
rect 53012 34892 53064 34944
rect 54024 34935 54076 34944
rect 54024 34901 54033 34935
rect 54033 34901 54067 34935
rect 54067 34901 54076 34935
rect 54024 34892 54076 34901
rect 54208 34935 54260 34944
rect 54208 34901 54217 34935
rect 54217 34901 54251 34935
rect 54251 34901 54260 34935
rect 54208 34892 54260 34901
rect 54760 34935 54812 34944
rect 54760 34901 54769 34935
rect 54769 34901 54803 34935
rect 54803 34901 54812 34935
rect 54760 34892 54812 34901
rect 54852 34892 54904 34944
rect 56416 34935 56468 34944
rect 56416 34901 56425 34935
rect 56425 34901 56459 34935
rect 56459 34901 56468 34935
rect 56416 34892 56468 34901
rect 56968 34892 57020 34944
rect 57796 34892 57848 34944
rect 58624 34892 58676 34944
rect 61752 34935 61804 34944
rect 61752 34901 61761 34935
rect 61761 34901 61795 34935
rect 61795 34901 61804 34935
rect 61752 34892 61804 34901
rect 62764 35105 62773 35139
rect 62773 35105 62807 35139
rect 62807 35105 62816 35139
rect 62764 35096 62816 35105
rect 63040 35096 63092 35148
rect 64328 35096 64380 35148
rect 66720 35139 66772 35148
rect 66720 35105 66729 35139
rect 66729 35105 66763 35139
rect 66763 35105 66772 35139
rect 67088 35139 67140 35148
rect 66720 35096 66772 35105
rect 67088 35105 67097 35139
rect 67097 35105 67131 35139
rect 67131 35105 67140 35139
rect 67088 35096 67140 35105
rect 69204 35232 69256 35284
rect 87420 35232 87472 35284
rect 88432 35232 88484 35284
rect 67272 35164 67324 35216
rect 68928 35164 68980 35216
rect 71780 35164 71832 35216
rect 68744 35096 68796 35148
rect 73252 35096 73304 35148
rect 66352 35028 66404 35080
rect 68560 35028 68612 35080
rect 70584 35071 70636 35080
rect 70584 35037 70593 35071
rect 70593 35037 70627 35071
rect 70627 35037 70636 35071
rect 70584 35028 70636 35037
rect 74172 35096 74224 35148
rect 74632 35139 74684 35148
rect 74632 35105 74641 35139
rect 74641 35105 74675 35139
rect 74675 35105 74684 35139
rect 74632 35096 74684 35105
rect 74264 35071 74316 35080
rect 74264 35037 74273 35071
rect 74273 35037 74307 35071
rect 74307 35037 74316 35071
rect 75368 35139 75420 35148
rect 75368 35105 75377 35139
rect 75377 35105 75411 35139
rect 75411 35105 75420 35139
rect 75368 35096 75420 35105
rect 76288 35164 76340 35216
rect 75644 35096 75696 35148
rect 78312 35164 78364 35216
rect 84476 35164 84528 35216
rect 77116 35096 77168 35148
rect 79600 35096 79652 35148
rect 81348 35096 81400 35148
rect 83280 35139 83332 35148
rect 74264 35028 74316 35037
rect 67272 34960 67324 35012
rect 68744 34960 68796 35012
rect 62764 34892 62816 34944
rect 63132 34892 63184 34944
rect 63868 34935 63920 34944
rect 63868 34901 63877 34935
rect 63877 34901 63911 34935
rect 63911 34901 63920 34935
rect 63868 34892 63920 34901
rect 64512 34892 64564 34944
rect 66168 34892 66220 34944
rect 66720 34892 66772 34944
rect 67088 34892 67140 34944
rect 69848 34892 69900 34944
rect 69940 34892 69992 34944
rect 77024 34960 77076 35012
rect 82268 35028 82320 35080
rect 82544 34960 82596 35012
rect 75092 34892 75144 34944
rect 77300 34892 77352 34944
rect 78036 34935 78088 34944
rect 78036 34901 78045 34935
rect 78045 34901 78079 34935
rect 78079 34901 78088 34935
rect 78036 34892 78088 34901
rect 78956 34892 79008 34944
rect 81808 34935 81860 34944
rect 81808 34901 81817 34935
rect 81817 34901 81851 34935
rect 81851 34901 81860 34935
rect 81808 34892 81860 34901
rect 82084 34892 82136 34944
rect 83280 35105 83289 35139
rect 83289 35105 83323 35139
rect 83323 35105 83332 35139
rect 83280 35096 83332 35105
rect 84384 35139 84436 35148
rect 84384 35105 84393 35139
rect 84393 35105 84427 35139
rect 84427 35105 84436 35139
rect 84752 35207 84804 35216
rect 84752 35173 84761 35207
rect 84761 35173 84795 35207
rect 84795 35173 84804 35207
rect 84752 35164 84804 35173
rect 86040 35207 86092 35216
rect 86040 35173 86049 35207
rect 86049 35173 86083 35207
rect 86083 35173 86092 35207
rect 86040 35164 86092 35173
rect 86224 35164 86276 35216
rect 84384 35096 84436 35105
rect 85396 35139 85448 35148
rect 85396 35105 85405 35139
rect 85405 35105 85439 35139
rect 85439 35105 85448 35139
rect 85396 35096 85448 35105
rect 85580 35139 85632 35148
rect 85580 35105 85589 35139
rect 85589 35105 85623 35139
rect 85623 35105 85632 35139
rect 85580 35096 85632 35105
rect 88248 35139 88300 35148
rect 88248 35105 88257 35139
rect 88257 35105 88291 35139
rect 88291 35105 88300 35139
rect 88248 35096 88300 35105
rect 89536 35139 89588 35148
rect 89168 35028 89220 35080
rect 89536 35105 89545 35139
rect 89545 35105 89579 35139
rect 89579 35105 89588 35139
rect 89536 35096 89588 35105
rect 91744 35139 91796 35148
rect 91744 35105 91753 35139
rect 91753 35105 91787 35139
rect 91787 35105 91796 35139
rect 94136 35139 94188 35148
rect 91744 35096 91796 35105
rect 93860 35071 93912 35080
rect 93860 35037 93869 35071
rect 93869 35037 93903 35071
rect 93903 35037 93912 35071
rect 93860 35028 93912 35037
rect 94136 35105 94145 35139
rect 94145 35105 94179 35139
rect 94179 35105 94188 35139
rect 94136 35096 94188 35105
rect 83464 35003 83516 35012
rect 83464 34969 83473 35003
rect 83473 34969 83507 35003
rect 83507 34969 83516 35003
rect 83464 34960 83516 34969
rect 83556 34960 83608 35012
rect 88340 34892 88392 34944
rect 90180 34892 90232 34944
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 65686 34790 65738 34842
rect 65750 34790 65802 34842
rect 65814 34790 65866 34842
rect 65878 34790 65930 34842
rect 96406 34790 96458 34842
rect 96470 34790 96522 34842
rect 96534 34790 96586 34842
rect 96598 34790 96650 34842
rect 4620 34688 4672 34740
rect 11428 34731 11480 34740
rect 11428 34697 11437 34731
rect 11437 34697 11471 34731
rect 11471 34697 11480 34731
rect 11428 34688 11480 34697
rect 13084 34688 13136 34740
rect 13728 34688 13780 34740
rect 14464 34731 14516 34740
rect 14464 34697 14473 34731
rect 14473 34697 14507 34731
rect 14507 34697 14516 34731
rect 14464 34688 14516 34697
rect 15292 34688 15344 34740
rect 18788 34731 18840 34740
rect 18788 34697 18797 34731
rect 18797 34697 18831 34731
rect 18831 34697 18840 34731
rect 18788 34688 18840 34697
rect 19432 34688 19484 34740
rect 21180 34688 21232 34740
rect 22100 34688 22152 34740
rect 22284 34731 22336 34740
rect 22284 34697 22293 34731
rect 22293 34697 22327 34731
rect 22327 34697 22336 34731
rect 22284 34688 22336 34697
rect 14372 34620 14424 34672
rect 2504 34595 2556 34604
rect 2504 34561 2513 34595
rect 2513 34561 2547 34595
rect 2547 34561 2556 34595
rect 2504 34552 2556 34561
rect 3148 34552 3200 34604
rect 10876 34552 10928 34604
rect 22192 34620 22244 34672
rect 25320 34620 25372 34672
rect 30472 34620 30524 34672
rect 17776 34552 17828 34604
rect 20076 34552 20128 34604
rect 4068 34416 4120 34468
rect 5908 34484 5960 34536
rect 6276 34484 6328 34536
rect 7288 34527 7340 34536
rect 7288 34493 7297 34527
rect 7297 34493 7331 34527
rect 7331 34493 7340 34527
rect 7288 34484 7340 34493
rect 3884 34391 3936 34400
rect 3884 34357 3893 34391
rect 3893 34357 3927 34391
rect 3927 34357 3936 34391
rect 3884 34348 3936 34357
rect 5264 34391 5316 34400
rect 5264 34357 5273 34391
rect 5273 34357 5307 34391
rect 5307 34357 5316 34391
rect 5264 34348 5316 34357
rect 5540 34416 5592 34468
rect 12624 34416 12676 34468
rect 6920 34391 6972 34400
rect 6920 34357 6929 34391
rect 6929 34357 6963 34391
rect 6963 34357 6972 34391
rect 6920 34348 6972 34357
rect 13084 34527 13136 34536
rect 13084 34493 13093 34527
rect 13093 34493 13127 34527
rect 13127 34493 13136 34527
rect 13084 34484 13136 34493
rect 13728 34484 13780 34536
rect 14372 34484 14424 34536
rect 16580 34484 16632 34536
rect 17960 34484 18012 34536
rect 19984 34484 20036 34536
rect 20352 34484 20404 34536
rect 23388 34552 23440 34604
rect 21180 34527 21232 34536
rect 21180 34493 21189 34527
rect 21189 34493 21223 34527
rect 21223 34493 21232 34527
rect 21180 34484 21232 34493
rect 21272 34527 21324 34536
rect 21272 34493 21281 34527
rect 21281 34493 21315 34527
rect 21315 34493 21324 34527
rect 21272 34484 21324 34493
rect 32220 34595 32272 34604
rect 26056 34416 26108 34468
rect 26240 34459 26292 34468
rect 26240 34425 26249 34459
rect 26249 34425 26283 34459
rect 26283 34425 26292 34459
rect 26700 34484 26752 34536
rect 30564 34484 30616 34536
rect 30748 34527 30800 34536
rect 30748 34493 30757 34527
rect 30757 34493 30791 34527
rect 30791 34493 30800 34527
rect 30748 34484 30800 34493
rect 30932 34527 30984 34536
rect 30932 34493 30941 34527
rect 30941 34493 30975 34527
rect 30975 34493 30984 34527
rect 30932 34484 30984 34493
rect 32220 34561 32229 34595
rect 32229 34561 32263 34595
rect 32263 34561 32272 34595
rect 32220 34552 32272 34561
rect 32864 34552 32916 34604
rect 33508 34620 33560 34672
rect 36636 34688 36688 34740
rect 37004 34688 37056 34740
rect 38844 34688 38896 34740
rect 39028 34731 39080 34740
rect 39028 34697 39037 34731
rect 39037 34697 39071 34731
rect 39071 34697 39080 34731
rect 39028 34688 39080 34697
rect 39580 34731 39632 34740
rect 39580 34697 39589 34731
rect 39589 34697 39623 34731
rect 39623 34697 39632 34731
rect 39580 34688 39632 34697
rect 39672 34688 39724 34740
rect 41512 34688 41564 34740
rect 41696 34688 41748 34740
rect 42892 34688 42944 34740
rect 43628 34688 43680 34740
rect 26240 34416 26292 34425
rect 13636 34348 13688 34400
rect 19984 34348 20036 34400
rect 20352 34391 20404 34400
rect 20352 34357 20361 34391
rect 20361 34357 20395 34391
rect 20395 34357 20404 34391
rect 20352 34348 20404 34357
rect 21180 34348 21232 34400
rect 23848 34391 23900 34400
rect 23848 34357 23857 34391
rect 23857 34357 23891 34391
rect 23891 34357 23900 34391
rect 23848 34348 23900 34357
rect 26608 34391 26660 34400
rect 26608 34357 26617 34391
rect 26617 34357 26651 34391
rect 26651 34357 26660 34391
rect 26608 34348 26660 34357
rect 32312 34348 32364 34400
rect 33324 34484 33376 34536
rect 42064 34620 42116 34672
rect 81348 34688 81400 34740
rect 81440 34688 81492 34740
rect 37464 34527 37516 34536
rect 37464 34493 37473 34527
rect 37473 34493 37507 34527
rect 37507 34493 37516 34527
rect 37464 34484 37516 34493
rect 38016 34527 38068 34536
rect 38016 34493 38025 34527
rect 38025 34493 38059 34527
rect 38059 34493 38068 34527
rect 38016 34484 38068 34493
rect 38660 34484 38712 34536
rect 42984 34552 43036 34604
rect 44548 34552 44600 34604
rect 51908 34552 51960 34604
rect 37096 34348 37148 34400
rect 40040 34484 40092 34536
rect 40960 34484 41012 34536
rect 41512 34459 41564 34468
rect 41512 34425 41521 34459
rect 41521 34425 41555 34459
rect 41555 34425 41564 34459
rect 43996 34484 44048 34536
rect 51816 34484 51868 34536
rect 52644 34620 52696 34672
rect 53012 34595 53064 34604
rect 53012 34561 53021 34595
rect 53021 34561 53055 34595
rect 53055 34561 53064 34595
rect 53012 34552 53064 34561
rect 53932 34552 53984 34604
rect 59084 34620 59136 34672
rect 41512 34416 41564 34425
rect 52552 34416 52604 34468
rect 49976 34348 50028 34400
rect 52368 34348 52420 34400
rect 54116 34484 54168 34536
rect 54300 34484 54352 34536
rect 54392 34459 54444 34468
rect 54392 34425 54401 34459
rect 54401 34425 54435 34459
rect 54435 34425 54444 34459
rect 54852 34527 54904 34536
rect 54852 34493 54861 34527
rect 54861 34493 54895 34527
rect 54895 34493 54904 34527
rect 54852 34484 54904 34493
rect 54944 34484 54996 34536
rect 56140 34552 56192 34604
rect 58992 34595 59044 34604
rect 55404 34527 55456 34536
rect 55404 34493 55413 34527
rect 55413 34493 55447 34527
rect 55447 34493 55456 34527
rect 55404 34484 55456 34493
rect 55220 34459 55272 34468
rect 54392 34416 54444 34425
rect 55220 34425 55229 34459
rect 55229 34425 55263 34459
rect 55263 34425 55272 34459
rect 55220 34416 55272 34425
rect 54576 34348 54628 34400
rect 57520 34527 57572 34536
rect 56784 34459 56836 34468
rect 56784 34425 56793 34459
rect 56793 34425 56827 34459
rect 56827 34425 56836 34459
rect 57520 34493 57529 34527
rect 57529 34493 57563 34527
rect 57563 34493 57572 34527
rect 57520 34484 57572 34493
rect 58992 34561 59001 34595
rect 59001 34561 59035 34595
rect 59035 34561 59044 34595
rect 58992 34552 59044 34561
rect 57888 34484 57940 34536
rect 57980 34527 58032 34536
rect 57980 34493 57989 34527
rect 57989 34493 58023 34527
rect 58023 34493 58032 34527
rect 57980 34484 58032 34493
rect 58900 34527 58952 34536
rect 56784 34416 56836 34425
rect 57520 34348 57572 34400
rect 58900 34493 58909 34527
rect 58909 34493 58943 34527
rect 58943 34493 58952 34527
rect 58900 34484 58952 34493
rect 59084 34484 59136 34536
rect 58164 34348 58216 34400
rect 58532 34391 58584 34400
rect 58532 34357 58541 34391
rect 58541 34357 58575 34391
rect 58575 34357 58584 34391
rect 58532 34348 58584 34357
rect 62488 34459 62540 34468
rect 62488 34425 62497 34459
rect 62497 34425 62531 34459
rect 62531 34425 62540 34459
rect 63132 34527 63184 34536
rect 62488 34416 62540 34425
rect 63132 34493 63141 34527
rect 63141 34493 63175 34527
rect 63175 34493 63184 34527
rect 63132 34484 63184 34493
rect 63868 34484 63920 34536
rect 65340 34620 65392 34672
rect 66996 34620 67048 34672
rect 75644 34620 75696 34672
rect 77760 34663 77812 34672
rect 77760 34629 77769 34663
rect 77769 34629 77803 34663
rect 77803 34629 77812 34663
rect 77760 34620 77812 34629
rect 78772 34620 78824 34672
rect 79784 34620 79836 34672
rect 81532 34620 81584 34672
rect 82544 34663 82596 34672
rect 82544 34629 82553 34663
rect 82553 34629 82587 34663
rect 82587 34629 82596 34663
rect 82544 34620 82596 34629
rect 85488 34620 85540 34672
rect 88156 34688 88208 34740
rect 91284 34731 91336 34740
rect 91284 34697 91293 34731
rect 91293 34697 91327 34731
rect 91327 34697 91336 34731
rect 91284 34688 91336 34697
rect 66260 34595 66312 34604
rect 66260 34561 66269 34595
rect 66269 34561 66303 34595
rect 66303 34561 66312 34595
rect 66260 34552 66312 34561
rect 66352 34552 66404 34604
rect 75092 34552 75144 34604
rect 76472 34595 76524 34604
rect 76196 34527 76248 34536
rect 76196 34493 76205 34527
rect 76205 34493 76239 34527
rect 76239 34493 76248 34527
rect 76196 34484 76248 34493
rect 76472 34561 76481 34595
rect 76481 34561 76515 34595
rect 76515 34561 76524 34595
rect 76472 34552 76524 34561
rect 78496 34552 78548 34604
rect 78956 34595 79008 34604
rect 78956 34561 78965 34595
rect 78965 34561 78999 34595
rect 78999 34561 79008 34595
rect 78956 34552 79008 34561
rect 81348 34552 81400 34604
rect 81624 34595 81676 34604
rect 81624 34561 81633 34595
rect 81633 34561 81667 34595
rect 81667 34561 81676 34595
rect 81624 34552 81676 34561
rect 77116 34484 77168 34536
rect 77760 34484 77812 34536
rect 78588 34484 78640 34536
rect 78864 34484 78916 34536
rect 80888 34484 80940 34536
rect 81440 34527 81492 34536
rect 81440 34493 81449 34527
rect 81449 34493 81483 34527
rect 81483 34493 81492 34527
rect 81440 34484 81492 34493
rect 82360 34527 82412 34536
rect 74632 34416 74684 34468
rect 64512 34391 64564 34400
rect 64512 34357 64521 34391
rect 64521 34357 64555 34391
rect 64555 34357 64564 34391
rect 64512 34348 64564 34357
rect 65984 34348 66036 34400
rect 67364 34391 67416 34400
rect 67364 34357 67373 34391
rect 67373 34357 67407 34391
rect 67407 34357 67416 34391
rect 78496 34416 78548 34468
rect 78772 34459 78824 34468
rect 78772 34425 78781 34459
rect 78781 34425 78815 34459
rect 78815 34425 78824 34459
rect 81992 34459 82044 34468
rect 78772 34416 78824 34425
rect 81992 34425 82001 34459
rect 82001 34425 82035 34459
rect 82035 34425 82044 34459
rect 81992 34416 82044 34425
rect 82360 34493 82369 34527
rect 82369 34493 82403 34527
rect 82403 34493 82412 34527
rect 82360 34484 82412 34493
rect 82544 34484 82596 34536
rect 83464 34484 83516 34536
rect 85488 34484 85540 34536
rect 88432 34620 88484 34672
rect 88340 34552 88392 34604
rect 88248 34484 88300 34536
rect 88984 34527 89036 34536
rect 88984 34493 88993 34527
rect 88993 34493 89027 34527
rect 89027 34493 89036 34527
rect 88984 34484 89036 34493
rect 90640 34484 90692 34536
rect 85580 34391 85632 34400
rect 67364 34348 67416 34357
rect 85580 34357 85589 34391
rect 85589 34357 85623 34391
rect 85623 34357 85632 34391
rect 85580 34348 85632 34357
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 50326 34246 50378 34298
rect 50390 34246 50442 34298
rect 50454 34246 50506 34298
rect 50518 34246 50570 34298
rect 81046 34246 81098 34298
rect 81110 34246 81162 34298
rect 81174 34246 81226 34298
rect 81238 34246 81290 34298
rect 5540 34144 5592 34196
rect 6092 34187 6144 34196
rect 6092 34153 6101 34187
rect 6101 34153 6135 34187
rect 6135 34153 6144 34187
rect 6092 34144 6144 34153
rect 9772 34144 9824 34196
rect 10232 34144 10284 34196
rect 11520 34187 11572 34196
rect 11520 34153 11529 34187
rect 11529 34153 11563 34187
rect 11563 34153 11572 34187
rect 11520 34144 11572 34153
rect 3792 34076 3844 34128
rect 18052 34144 18104 34196
rect 27528 34144 27580 34196
rect 56048 34144 56100 34196
rect 13728 34119 13780 34128
rect 13728 34085 13737 34119
rect 13737 34085 13771 34119
rect 13771 34085 13780 34119
rect 13728 34076 13780 34085
rect 15660 34076 15712 34128
rect 21180 34076 21232 34128
rect 24308 34076 24360 34128
rect 24400 34076 24452 34128
rect 48780 34076 48832 34128
rect 52368 34076 52420 34128
rect 67364 34076 67416 34128
rect 4804 34008 4856 34060
rect 5448 34008 5500 34060
rect 6276 34051 6328 34060
rect 6276 34017 6285 34051
rect 6285 34017 6319 34051
rect 6319 34017 6328 34051
rect 6276 34008 6328 34017
rect 6552 34051 6604 34060
rect 6552 34017 6561 34051
rect 6561 34017 6595 34051
rect 6595 34017 6604 34051
rect 6552 34008 6604 34017
rect 9772 34008 9824 34060
rect 10140 34008 10192 34060
rect 11980 34008 12032 34060
rect 13176 34051 13228 34060
rect 13176 34017 13185 34051
rect 13185 34017 13219 34051
rect 13219 34017 13228 34051
rect 13176 34008 13228 34017
rect 13912 34008 13964 34060
rect 15292 34051 15344 34060
rect 15292 34017 15301 34051
rect 15301 34017 15335 34051
rect 15335 34017 15344 34051
rect 15292 34008 15344 34017
rect 20168 34008 20220 34060
rect 21456 34008 21508 34060
rect 23112 34008 23164 34060
rect 56416 34008 56468 34060
rect 12348 33983 12400 33992
rect 12348 33949 12357 33983
rect 12357 33949 12391 33983
rect 12391 33949 12400 33983
rect 12348 33940 12400 33949
rect 15844 33940 15896 33992
rect 11888 33872 11940 33924
rect 20444 33872 20496 33924
rect 11244 33804 11296 33856
rect 12716 33804 12768 33856
rect 13912 33847 13964 33856
rect 13912 33813 13921 33847
rect 13921 33813 13955 33847
rect 13955 33813 13964 33847
rect 13912 33804 13964 33813
rect 19984 33804 20036 33856
rect 21272 33940 21324 33992
rect 21364 33983 21416 33992
rect 21364 33949 21373 33983
rect 21373 33949 21407 33983
rect 21407 33949 21416 33983
rect 21364 33940 21416 33949
rect 22008 33940 22060 33992
rect 23664 33940 23716 33992
rect 22468 33872 22520 33924
rect 24400 33872 24452 33924
rect 61752 33940 61804 33992
rect 21732 33804 21784 33856
rect 23204 33804 23256 33856
rect 62488 33872 62540 33924
rect 24584 33804 24636 33856
rect 49976 33804 50028 33856
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 24768 33736 24820 33788
rect 46572 33736 46624 33788
rect 4804 33643 4856 33652
rect 4804 33609 4813 33643
rect 4813 33609 4847 33643
rect 4847 33609 4856 33643
rect 4804 33600 4856 33609
rect 9312 33600 9364 33652
rect 21640 33600 21692 33652
rect 22192 33643 22244 33652
rect 22192 33609 22201 33643
rect 22201 33609 22235 33643
rect 22235 33609 22244 33643
rect 22192 33600 22244 33609
rect 23848 33600 23900 33652
rect 24400 33600 24452 33652
rect 24584 33600 24636 33652
rect 24860 33600 24912 33652
rect 55956 33600 56008 33652
rect 11244 33575 11296 33584
rect 11244 33541 11253 33575
rect 11253 33541 11287 33575
rect 11287 33541 11296 33575
rect 11244 33532 11296 33541
rect 4068 33396 4120 33448
rect 5632 33396 5684 33448
rect 12440 33439 12492 33448
rect 12440 33405 12449 33439
rect 12449 33405 12483 33439
rect 12483 33405 12492 33439
rect 12716 33439 12768 33448
rect 12440 33396 12492 33405
rect 12716 33405 12725 33439
rect 12725 33405 12759 33439
rect 12759 33405 12768 33439
rect 12716 33396 12768 33405
rect 11704 33260 11756 33312
rect 13728 33260 13780 33312
rect 20352 33464 20404 33516
rect 15200 33396 15252 33448
rect 54484 33532 54536 33584
rect 21640 33464 21692 33516
rect 30748 33464 30800 33516
rect 20352 33371 20404 33380
rect 20352 33337 20361 33371
rect 20361 33337 20395 33371
rect 20395 33337 20404 33371
rect 20352 33328 20404 33337
rect 20996 33396 21048 33448
rect 21272 33439 21324 33448
rect 21272 33405 21277 33439
rect 21277 33405 21311 33439
rect 21311 33405 21324 33439
rect 21272 33396 21324 33405
rect 21548 33396 21600 33448
rect 52092 33396 52144 33448
rect 20812 33328 20864 33380
rect 21732 33328 21784 33380
rect 54576 33328 54628 33380
rect 21272 33260 21324 33312
rect 21364 33260 21416 33312
rect 22376 33260 22428 33312
rect 22652 33260 22704 33312
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 3424 33056 3476 33108
rect 7012 33056 7064 33108
rect 40040 33056 40092 33108
rect 52092 33056 52144 33108
rect 54392 33056 54444 33108
rect 11428 32988 11480 33040
rect 3516 32920 3568 32972
rect 4620 32920 4672 32972
rect 6092 32920 6144 32972
rect 11796 32963 11848 32972
rect 11796 32929 11805 32963
rect 11805 32929 11839 32963
rect 11839 32929 11848 32963
rect 11796 32920 11848 32929
rect 12716 32988 12768 33040
rect 13176 32988 13228 33040
rect 12532 32920 12584 32972
rect 15292 32963 15344 32972
rect 3516 32784 3568 32836
rect 3700 32784 3752 32836
rect 2412 32716 2464 32768
rect 4068 32716 4120 32768
rect 4804 32716 4856 32768
rect 8484 32716 8536 32768
rect 11980 32784 12032 32836
rect 15292 32929 15301 32963
rect 15301 32929 15335 32963
rect 15335 32929 15344 32963
rect 15292 32920 15344 32929
rect 17500 32988 17552 33040
rect 17960 32963 18012 32972
rect 17960 32929 17969 32963
rect 17969 32929 18003 32963
rect 18003 32929 18012 32963
rect 17960 32920 18012 32929
rect 18328 32988 18380 33040
rect 19616 32963 19668 32972
rect 19616 32929 19625 32963
rect 19625 32929 19659 32963
rect 19659 32929 19668 32963
rect 19616 32920 19668 32929
rect 30932 32988 30984 33040
rect 37280 32920 37332 32972
rect 14280 32784 14332 32836
rect 14464 32784 14516 32836
rect 21732 32852 21784 32904
rect 22192 32895 22244 32904
rect 22192 32861 22201 32895
rect 22201 32861 22235 32895
rect 22235 32861 22244 32895
rect 22192 32852 22244 32861
rect 31760 32852 31812 32904
rect 12348 32716 12400 32768
rect 13820 32716 13872 32768
rect 15476 32759 15528 32768
rect 15476 32725 15485 32759
rect 15485 32725 15519 32759
rect 15519 32725 15528 32759
rect 15476 32716 15528 32725
rect 17132 32759 17184 32768
rect 17132 32725 17141 32759
rect 17141 32725 17175 32759
rect 17175 32725 17184 32759
rect 17132 32716 17184 32725
rect 18052 32716 18104 32768
rect 19248 32716 19300 32768
rect 19892 32716 19944 32768
rect 21732 32759 21784 32768
rect 21732 32725 21741 32759
rect 21741 32725 21775 32759
rect 21775 32725 21784 32759
rect 21732 32716 21784 32725
rect 34612 32784 34664 32836
rect 37464 32716 37516 32768
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 28356 32580 28408 32632
rect 48964 32580 49016 32632
rect 3700 32444 3752 32496
rect 66168 32512 66220 32564
rect 4620 32444 4672 32496
rect 5356 32444 5408 32496
rect 2872 32376 2924 32428
rect 5816 32376 5868 32428
rect 5908 32376 5960 32428
rect 10324 32376 10376 32428
rect 11796 32376 11848 32428
rect 12532 32376 12584 32428
rect 19892 32444 19944 32496
rect 20812 32487 20864 32496
rect 19616 32419 19668 32428
rect 3700 32308 3752 32360
rect 4068 32308 4120 32360
rect 5448 32308 5500 32360
rect 4804 32240 4856 32292
rect 9680 32351 9732 32360
rect 9680 32317 9689 32351
rect 9689 32317 9723 32351
rect 9723 32317 9732 32351
rect 9680 32308 9732 32317
rect 11244 32308 11296 32360
rect 11980 32308 12032 32360
rect 14464 32351 14516 32360
rect 14464 32317 14473 32351
rect 14473 32317 14507 32351
rect 14507 32317 14516 32351
rect 14464 32308 14516 32317
rect 14740 32240 14792 32292
rect 16948 32308 17000 32360
rect 18144 32351 18196 32360
rect 18144 32317 18153 32351
rect 18153 32317 18187 32351
rect 18187 32317 18196 32351
rect 18144 32308 18196 32317
rect 16396 32240 16448 32292
rect 18052 32240 18104 32292
rect 19616 32385 19625 32419
rect 19625 32385 19659 32419
rect 19659 32385 19668 32419
rect 19616 32376 19668 32385
rect 20812 32453 20821 32487
rect 20821 32453 20855 32487
rect 20855 32453 20864 32487
rect 20812 32444 20864 32453
rect 20904 32444 20956 32496
rect 21548 32376 21600 32428
rect 24860 32376 24912 32428
rect 49608 32444 49660 32496
rect 62580 32376 62632 32428
rect 3884 32172 3936 32224
rect 5540 32172 5592 32224
rect 8576 32172 8628 32224
rect 13176 32172 13228 32224
rect 15476 32172 15528 32224
rect 15568 32172 15620 32224
rect 20260 32172 20312 32224
rect 21824 32240 21876 32292
rect 46756 32240 46808 32292
rect 63684 32172 63736 32224
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 5448 31968 5500 32020
rect 10876 32011 10928 32020
rect 10876 31977 10885 32011
rect 10885 31977 10919 32011
rect 10919 31977 10928 32011
rect 10876 31968 10928 31977
rect 13176 31968 13228 32020
rect 14280 31968 14332 32020
rect 14740 31968 14792 32020
rect 15568 31968 15620 32020
rect 16580 31968 16632 32020
rect 16856 31968 16908 32020
rect 17776 32011 17828 32020
rect 17776 31977 17785 32011
rect 17785 31977 17819 32011
rect 17819 31977 17828 32011
rect 17776 31968 17828 31977
rect 18144 31968 18196 32020
rect 20260 31968 20312 32020
rect 21732 32011 21784 32020
rect 21732 31977 21741 32011
rect 21741 31977 21775 32011
rect 21775 31977 21784 32011
rect 21732 31968 21784 31977
rect 21824 31968 21876 32020
rect 52092 31968 52144 32020
rect 4068 31875 4120 31884
rect 3148 31807 3200 31816
rect 3148 31773 3157 31807
rect 3157 31773 3191 31807
rect 3191 31773 3200 31807
rect 3148 31764 3200 31773
rect 3792 31696 3844 31748
rect 4068 31841 4077 31875
rect 4077 31841 4111 31875
rect 4111 31841 4120 31875
rect 4068 31832 4120 31841
rect 4988 31832 5040 31884
rect 5632 31875 5684 31884
rect 5632 31841 5641 31875
rect 5641 31841 5675 31875
rect 5675 31841 5684 31875
rect 5632 31832 5684 31841
rect 8576 31875 8628 31884
rect 8576 31841 8585 31875
rect 8585 31841 8619 31875
rect 8619 31841 8628 31875
rect 8576 31832 8628 31841
rect 9680 31943 9732 31952
rect 9680 31909 9689 31943
rect 9689 31909 9723 31943
rect 9723 31909 9732 31943
rect 9680 31900 9732 31909
rect 9956 31900 10008 31952
rect 21640 31900 21692 31952
rect 10232 31875 10284 31884
rect 8392 31764 8444 31816
rect 4620 31696 4672 31748
rect 10232 31841 10241 31875
rect 10241 31841 10275 31875
rect 10275 31841 10284 31875
rect 10232 31832 10284 31841
rect 10876 31832 10928 31884
rect 14280 31832 14332 31884
rect 15292 31832 15344 31884
rect 15476 31875 15528 31884
rect 15476 31841 15485 31875
rect 15485 31841 15519 31875
rect 15519 31841 15528 31875
rect 15476 31832 15528 31841
rect 16580 31875 16632 31884
rect 16580 31841 16589 31875
rect 16589 31841 16623 31875
rect 16623 31841 16632 31875
rect 17684 31875 17736 31884
rect 16580 31832 16632 31841
rect 17684 31841 17693 31875
rect 17693 31841 17727 31875
rect 17727 31841 17736 31875
rect 17684 31832 17736 31841
rect 10324 31764 10376 31816
rect 17040 31764 17092 31816
rect 17868 31764 17920 31816
rect 20904 31764 20956 31816
rect 22008 31832 22060 31884
rect 22284 31832 22336 31884
rect 35624 31900 35676 31952
rect 23020 31832 23072 31884
rect 51540 31832 51592 31884
rect 55312 31764 55364 31816
rect 8668 31671 8720 31680
rect 8668 31637 8677 31671
rect 8677 31637 8711 31671
rect 8711 31637 8720 31671
rect 8668 31628 8720 31637
rect 16396 31628 16448 31680
rect 17040 31628 17092 31680
rect 62672 31696 62724 31748
rect 81440 31696 81492 31748
rect 81716 31696 81768 31748
rect 23296 31628 23348 31680
rect 51080 31628 51132 31680
rect 54852 31628 54904 31680
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 4620 31424 4672 31476
rect 11704 31467 11756 31476
rect 2412 31263 2464 31272
rect 2412 31229 2421 31263
rect 2421 31229 2455 31263
rect 2455 31229 2464 31263
rect 2412 31220 2464 31229
rect 3792 31263 3844 31272
rect 3792 31229 3801 31263
rect 3801 31229 3835 31263
rect 3835 31229 3844 31263
rect 3792 31220 3844 31229
rect 4620 31220 4672 31272
rect 8668 31288 8720 31340
rect 11704 31433 11713 31467
rect 11713 31433 11747 31467
rect 11747 31433 11756 31467
rect 11704 31424 11756 31433
rect 11796 31424 11848 31476
rect 26976 31492 27028 31544
rect 52000 31560 52052 31612
rect 55220 31560 55272 31612
rect 16948 31399 17000 31408
rect 16948 31365 16957 31399
rect 16957 31365 16991 31399
rect 16991 31365 17000 31399
rect 16948 31356 17000 31365
rect 18328 31356 18380 31408
rect 21548 31399 21600 31408
rect 8484 31263 8536 31272
rect 8484 31229 8493 31263
rect 8493 31229 8527 31263
rect 8527 31229 8536 31263
rect 8484 31220 8536 31229
rect 9864 31220 9916 31272
rect 11704 31220 11756 31272
rect 14372 31263 14424 31272
rect 14372 31229 14381 31263
rect 14381 31229 14415 31263
rect 14415 31229 14424 31263
rect 14372 31220 14424 31229
rect 15384 31288 15436 31340
rect 20076 31288 20128 31340
rect 21548 31365 21557 31399
rect 21557 31365 21591 31399
rect 21591 31365 21600 31399
rect 21548 31356 21600 31365
rect 22744 31356 22796 31408
rect 23296 31356 23348 31408
rect 23388 31356 23440 31408
rect 54300 31492 54352 31544
rect 53840 31424 53892 31476
rect 54116 31424 54168 31476
rect 52368 31356 52420 31408
rect 55404 31356 55456 31408
rect 2688 31084 2740 31136
rect 3792 31127 3844 31136
rect 3792 31093 3801 31127
rect 3801 31093 3835 31127
rect 3835 31093 3844 31127
rect 3792 31084 3844 31093
rect 4804 31084 4856 31136
rect 10140 31195 10192 31204
rect 10140 31161 10149 31195
rect 10149 31161 10183 31195
rect 10183 31161 10192 31195
rect 10140 31152 10192 31161
rect 10968 31195 11020 31204
rect 10968 31161 10977 31195
rect 10977 31161 11011 31195
rect 11011 31161 11020 31195
rect 10968 31152 11020 31161
rect 11796 31152 11848 31204
rect 16028 31220 16080 31272
rect 20168 31263 20220 31272
rect 20168 31229 20177 31263
rect 20177 31229 20211 31263
rect 20211 31229 20220 31263
rect 20168 31220 20220 31229
rect 53840 31288 53892 31340
rect 54024 31288 54076 31340
rect 20720 31263 20772 31272
rect 20720 31229 20729 31263
rect 20729 31229 20763 31263
rect 20763 31229 20772 31263
rect 22560 31263 22612 31272
rect 20720 31220 20772 31229
rect 22560 31229 22569 31263
rect 22569 31229 22603 31263
rect 22603 31229 22612 31263
rect 22560 31220 22612 31229
rect 43444 31220 43496 31272
rect 56784 31220 56836 31272
rect 9864 31084 9916 31136
rect 15292 31084 15344 31136
rect 16028 31084 16080 31136
rect 16212 31127 16264 31136
rect 16212 31093 16221 31127
rect 16221 31093 16255 31127
rect 16255 31093 16264 31127
rect 16212 31084 16264 31093
rect 20996 31084 21048 31136
rect 22192 31084 22244 31136
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 3424 30880 3476 30932
rect 4068 30787 4120 30796
rect 4068 30753 4077 30787
rect 4077 30753 4111 30787
rect 4111 30753 4120 30787
rect 4068 30744 4120 30753
rect 5080 30880 5132 30932
rect 15476 30880 15528 30932
rect 20168 30880 20220 30932
rect 20720 30880 20772 30932
rect 22100 30880 22152 30932
rect 7564 30744 7616 30796
rect 3056 30676 3108 30728
rect 7012 30676 7064 30728
rect 10324 30744 10376 30796
rect 10968 30744 11020 30796
rect 14004 30812 14056 30864
rect 17960 30812 18012 30864
rect 22560 30812 22612 30864
rect 11060 30676 11112 30728
rect 11428 30719 11480 30728
rect 11428 30685 11437 30719
rect 11437 30685 11471 30719
rect 11471 30685 11480 30719
rect 11428 30676 11480 30685
rect 14188 30787 14240 30796
rect 14188 30753 14197 30787
rect 14197 30753 14231 30787
rect 14231 30753 14240 30787
rect 14188 30744 14240 30753
rect 20812 30744 20864 30796
rect 22744 30880 22796 30932
rect 26792 31016 26844 31068
rect 53932 31016 53984 31068
rect 27068 30948 27120 31000
rect 81808 30948 81860 31000
rect 26884 30880 26936 30932
rect 81532 30880 81584 30932
rect 16212 30719 16264 30728
rect 16212 30685 16221 30719
rect 16221 30685 16255 30719
rect 16255 30685 16264 30719
rect 16212 30676 16264 30685
rect 16488 30719 16540 30728
rect 16488 30685 16497 30719
rect 16497 30685 16531 30719
rect 16531 30685 16540 30719
rect 16488 30676 16540 30685
rect 14372 30540 14424 30592
rect 22836 30676 22888 30728
rect 17592 30583 17644 30592
rect 17592 30549 17601 30583
rect 17601 30549 17635 30583
rect 17635 30549 17644 30583
rect 17592 30540 17644 30549
rect 17776 30540 17828 30592
rect 20996 30583 21048 30592
rect 20996 30549 21005 30583
rect 21005 30549 21039 30583
rect 21039 30549 21048 30583
rect 20996 30540 21048 30549
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 54024 30472 54076 30524
rect 54852 30472 54904 30524
rect 4068 30268 4120 30320
rect 6000 30311 6052 30320
rect 6000 30277 6009 30311
rect 6009 30277 6043 30311
rect 6043 30277 6052 30311
rect 6000 30268 6052 30277
rect 9312 30311 9364 30320
rect 9312 30277 9321 30311
rect 9321 30277 9355 30311
rect 9355 30277 9364 30311
rect 9312 30268 9364 30277
rect 11060 30268 11112 30320
rect 11428 30336 11480 30388
rect 12992 30336 13044 30388
rect 16488 30379 16540 30388
rect 16488 30345 16497 30379
rect 16497 30345 16531 30379
rect 16531 30345 16540 30379
rect 16488 30336 16540 30345
rect 11888 30268 11940 30320
rect 2688 30132 2740 30184
rect 4712 30132 4764 30184
rect 9404 30132 9456 30184
rect 10600 30132 10652 30184
rect 16488 30200 16540 30252
rect 16856 30311 16908 30320
rect 16856 30277 16865 30311
rect 16865 30277 16899 30311
rect 16899 30277 16908 30311
rect 16856 30268 16908 30277
rect 11060 30175 11112 30184
rect 11060 30141 11069 30175
rect 11069 30141 11103 30175
rect 11103 30141 11112 30175
rect 11060 30132 11112 30141
rect 11244 30132 11296 30184
rect 11428 30132 11480 30184
rect 10876 30064 10928 30116
rect 3608 30039 3660 30048
rect 3608 30005 3617 30039
rect 3617 30005 3651 30039
rect 3651 30005 3660 30039
rect 3608 29996 3660 30005
rect 4712 29996 4764 30048
rect 9404 29996 9456 30048
rect 10692 29996 10744 30048
rect 14648 29996 14700 30048
rect 15476 30175 15528 30184
rect 15476 30141 15485 30175
rect 15485 30141 15519 30175
rect 15519 30141 15528 30175
rect 15476 30132 15528 30141
rect 18144 30200 18196 30252
rect 22744 30336 22796 30388
rect 23388 30336 23440 30388
rect 22652 30268 22704 30320
rect 16396 30064 16448 30116
rect 16304 29996 16356 30048
rect 22100 30132 22152 30184
rect 24492 30200 24544 30252
rect 26700 30200 26752 30252
rect 20260 29996 20312 30048
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 3332 29835 3384 29844
rect 3332 29801 3341 29835
rect 3341 29801 3375 29835
rect 3375 29801 3384 29835
rect 3332 29792 3384 29801
rect 2688 29699 2740 29708
rect 2688 29665 2697 29699
rect 2697 29665 2731 29699
rect 2731 29665 2740 29699
rect 2688 29656 2740 29665
rect 2964 29631 3016 29640
rect 2964 29597 2973 29631
rect 2973 29597 3007 29631
rect 3007 29597 3016 29631
rect 2964 29588 3016 29597
rect 2504 29520 2556 29572
rect 7656 29656 7708 29708
rect 9312 29792 9364 29844
rect 14556 29792 14608 29844
rect 22100 29835 22152 29844
rect 22100 29801 22109 29835
rect 22109 29801 22143 29835
rect 22143 29801 22152 29835
rect 22100 29792 22152 29801
rect 22652 29792 22704 29844
rect 10876 29724 10928 29776
rect 26424 29724 26476 29776
rect 14372 29656 14424 29708
rect 5264 29588 5316 29640
rect 9864 29631 9916 29640
rect 4068 29452 4120 29504
rect 7288 29495 7340 29504
rect 7288 29461 7297 29495
rect 7297 29461 7331 29495
rect 7331 29461 7340 29495
rect 9864 29597 9873 29631
rect 9873 29597 9907 29631
rect 9907 29597 9916 29631
rect 9864 29588 9916 29597
rect 10784 29588 10836 29640
rect 8484 29563 8536 29572
rect 8484 29529 8493 29563
rect 8493 29529 8527 29563
rect 8527 29529 8536 29563
rect 8484 29520 8536 29529
rect 14648 29520 14700 29572
rect 7288 29452 7340 29461
rect 11336 29452 11388 29504
rect 15292 29699 15344 29708
rect 15292 29665 15301 29699
rect 15301 29665 15335 29699
rect 15335 29665 15344 29699
rect 15292 29656 15344 29665
rect 15384 29656 15436 29708
rect 15016 29588 15068 29640
rect 17500 29656 17552 29708
rect 20812 29656 20864 29708
rect 22652 29656 22704 29708
rect 16396 29520 16448 29572
rect 14924 29452 14976 29504
rect 15016 29495 15068 29504
rect 15016 29461 15025 29495
rect 15025 29461 15059 29495
rect 15059 29461 15068 29495
rect 15016 29452 15068 29461
rect 20812 29452 20864 29504
rect 53840 29452 53892 29504
rect 54208 29452 54260 29504
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 10784 29291 10836 29300
rect 10784 29257 10793 29291
rect 10793 29257 10827 29291
rect 10827 29257 10836 29291
rect 10784 29248 10836 29257
rect 14004 29248 14056 29300
rect 15016 29248 15068 29300
rect 15200 29248 15252 29300
rect 8484 29155 8536 29164
rect 6920 29044 6972 29096
rect 8484 29121 8493 29155
rect 8493 29121 8527 29155
rect 8527 29121 8536 29155
rect 8484 29112 8536 29121
rect 9404 29112 9456 29164
rect 9864 29044 9916 29096
rect 10692 29087 10744 29096
rect 10692 29053 10701 29087
rect 10701 29053 10735 29087
rect 10735 29053 10744 29087
rect 10692 29044 10744 29053
rect 12440 29044 12492 29096
rect 15476 29180 15528 29232
rect 15200 29044 15252 29096
rect 17132 29044 17184 29096
rect 19340 29044 19392 29096
rect 2596 28908 2648 28960
rect 3976 28976 4028 29028
rect 21824 29044 21876 29096
rect 24768 29112 24820 29164
rect 22560 29087 22612 29096
rect 22560 29053 22569 29087
rect 22569 29053 22603 29087
rect 22603 29053 22612 29087
rect 22560 29044 22612 29053
rect 23480 29044 23532 29096
rect 3884 28951 3936 28960
rect 3884 28917 3893 28951
rect 3893 28917 3927 28951
rect 3927 28917 3936 28951
rect 3884 28908 3936 28917
rect 4068 28908 4120 28960
rect 14740 28951 14792 28960
rect 14740 28917 14749 28951
rect 14749 28917 14783 28951
rect 14783 28917 14792 28951
rect 14740 28908 14792 28917
rect 20720 28976 20772 29028
rect 22652 28951 22704 28960
rect 22652 28917 22661 28951
rect 22661 28917 22695 28951
rect 22695 28917 22704 28951
rect 22652 28908 22704 28917
rect 27344 28908 27396 28960
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 3976 28704 4028 28756
rect 4528 28568 4580 28620
rect 13728 28500 13780 28552
rect 10968 28432 11020 28484
rect 11796 28364 11848 28416
rect 15200 28704 15252 28756
rect 19892 28636 19944 28688
rect 20168 28636 20220 28688
rect 20352 28636 20404 28688
rect 20536 28636 20588 28688
rect 15292 28611 15344 28620
rect 15292 28577 15301 28611
rect 15301 28577 15335 28611
rect 15335 28577 15344 28611
rect 15292 28568 15344 28577
rect 16580 28611 16632 28620
rect 16580 28577 16589 28611
rect 16589 28577 16623 28611
rect 16623 28577 16632 28611
rect 16580 28568 16632 28577
rect 19340 28611 19392 28620
rect 19340 28577 19349 28611
rect 19349 28577 19383 28611
rect 19383 28577 19392 28611
rect 19340 28568 19392 28577
rect 19524 28611 19576 28620
rect 19524 28577 19533 28611
rect 19533 28577 19567 28611
rect 19567 28577 19576 28611
rect 19524 28568 19576 28577
rect 18420 28500 18472 28552
rect 20352 28500 20404 28552
rect 22560 28543 22612 28552
rect 22560 28509 22569 28543
rect 22569 28509 22603 28543
rect 22603 28509 22612 28543
rect 22560 28500 22612 28509
rect 15384 28364 15436 28416
rect 15660 28364 15712 28416
rect 16396 28407 16448 28416
rect 16396 28373 16405 28407
rect 16405 28373 16439 28407
rect 16439 28373 16448 28407
rect 16396 28364 16448 28373
rect 18420 28407 18472 28416
rect 18420 28373 18429 28407
rect 18429 28373 18463 28407
rect 18463 28373 18472 28407
rect 18420 28364 18472 28373
rect 20352 28364 20404 28416
rect 26516 28364 26568 28416
rect 54300 28364 54352 28416
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 13820 28160 13872 28212
rect 18420 28160 18472 28212
rect 21824 28203 21876 28212
rect 21824 28169 21833 28203
rect 21833 28169 21867 28203
rect 21867 28169 21876 28203
rect 21824 28160 21876 28169
rect 2504 28067 2556 28076
rect 2504 28033 2513 28067
rect 2513 28033 2547 28067
rect 2547 28033 2556 28067
rect 2504 28024 2556 28033
rect 7840 28024 7892 28076
rect 14740 28024 14792 28076
rect 20720 28067 20772 28076
rect 20720 28033 20729 28067
rect 20729 28033 20763 28067
rect 20763 28033 20772 28067
rect 20720 28024 20772 28033
rect 2596 27956 2648 28008
rect 7932 27999 7984 28008
rect 7932 27965 7941 27999
rect 7941 27965 7975 27999
rect 7975 27965 7984 27999
rect 7932 27956 7984 27965
rect 8300 27999 8352 28008
rect 6920 27888 6972 27940
rect 8300 27965 8309 27999
rect 8309 27965 8343 27999
rect 8343 27965 8352 27999
rect 8300 27956 8352 27965
rect 11980 27956 12032 28008
rect 14924 27956 14976 28008
rect 16396 27956 16448 28008
rect 20352 27956 20404 28008
rect 11060 27888 11112 27940
rect 3884 27863 3936 27872
rect 3884 27829 3893 27863
rect 3893 27829 3927 27863
rect 3927 27829 3936 27863
rect 3884 27820 3936 27829
rect 4620 27820 4672 27872
rect 11428 27863 11480 27872
rect 11428 27829 11437 27863
rect 11437 27829 11471 27863
rect 11471 27829 11480 27863
rect 11428 27820 11480 27829
rect 14280 27820 14332 27872
rect 15292 27820 15344 27872
rect 20812 27820 20864 27872
rect 21364 27820 21416 27872
rect 24400 27820 24452 27872
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 9588 27616 9640 27668
rect 7656 27523 7708 27532
rect 7656 27489 7665 27523
rect 7665 27489 7699 27523
rect 7699 27489 7708 27523
rect 7656 27480 7708 27489
rect 9496 27548 9548 27600
rect 12532 27591 12584 27600
rect 8484 27523 8536 27532
rect 8484 27489 8493 27523
rect 8493 27489 8527 27523
rect 8527 27489 8536 27523
rect 8484 27480 8536 27489
rect 12532 27557 12541 27591
rect 12541 27557 12575 27591
rect 12575 27557 12584 27591
rect 12532 27548 12584 27557
rect 9772 27523 9824 27532
rect 9772 27489 9781 27523
rect 9781 27489 9815 27523
rect 9815 27489 9824 27523
rect 9772 27480 9824 27489
rect 6644 27276 6696 27328
rect 8392 27412 8444 27464
rect 9496 27412 9548 27464
rect 12532 27412 12584 27464
rect 12992 27455 13044 27464
rect 12992 27421 13001 27455
rect 13001 27421 13035 27455
rect 13035 27421 13044 27455
rect 12992 27412 13044 27421
rect 7104 27344 7156 27396
rect 16304 27523 16356 27532
rect 16304 27489 16313 27523
rect 16313 27489 16347 27523
rect 16347 27489 16356 27523
rect 16304 27480 16356 27489
rect 17224 27523 17276 27532
rect 17224 27489 17233 27523
rect 17233 27489 17267 27523
rect 17267 27489 17276 27523
rect 17224 27480 17276 27489
rect 18328 27480 18380 27532
rect 53840 27548 53892 27600
rect 54116 27548 54168 27600
rect 21364 27480 21416 27532
rect 21456 27412 21508 27464
rect 21916 27455 21968 27464
rect 21916 27421 21925 27455
rect 21925 27421 21959 27455
rect 21959 27421 21968 27455
rect 21916 27412 21968 27421
rect 22928 27412 22980 27464
rect 23204 27412 23256 27464
rect 7656 27276 7708 27328
rect 11428 27276 11480 27328
rect 13084 27276 13136 27328
rect 17868 27276 17920 27328
rect 20812 27276 20864 27328
rect 21456 27319 21508 27328
rect 21456 27285 21465 27319
rect 21465 27285 21499 27319
rect 21499 27285 21508 27319
rect 21456 27276 21508 27285
rect 28356 27344 28408 27396
rect 23204 27319 23256 27328
rect 23204 27285 23213 27319
rect 23213 27285 23247 27319
rect 23247 27285 23256 27319
rect 23204 27276 23256 27285
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 2780 27072 2832 27124
rect 3424 27072 3476 27124
rect 4068 27072 4120 27124
rect 25688 27072 25740 27124
rect 4620 27004 4672 27056
rect 6828 27004 6880 27056
rect 2504 26979 2556 26988
rect 2504 26945 2513 26979
rect 2513 26945 2547 26979
rect 2547 26945 2556 26979
rect 2504 26936 2556 26945
rect 3608 26936 3660 26988
rect 4068 26936 4120 26988
rect 7104 26979 7156 26988
rect 6828 26911 6880 26920
rect 6828 26877 6837 26911
rect 6837 26877 6871 26911
rect 6871 26877 6880 26911
rect 6828 26868 6880 26877
rect 7104 26945 7113 26979
rect 7113 26945 7147 26979
rect 7147 26945 7156 26979
rect 7104 26936 7156 26945
rect 11428 26868 11480 26920
rect 6920 26800 6972 26852
rect 12716 26800 12768 26852
rect 12992 27004 13044 27056
rect 18328 27047 18380 27056
rect 18328 27013 18337 27047
rect 18337 27013 18371 27047
rect 18371 27013 18380 27047
rect 18328 27004 18380 27013
rect 19892 27004 19944 27056
rect 20628 27004 20680 27056
rect 12992 26868 13044 26920
rect 13176 26911 13228 26920
rect 13176 26877 13185 26911
rect 13185 26877 13219 26911
rect 13219 26877 13228 26911
rect 13176 26868 13228 26877
rect 19248 26868 19300 26920
rect 21916 26936 21968 26988
rect 18696 26800 18748 26852
rect 3424 26732 3476 26784
rect 3608 26732 3660 26784
rect 3884 26775 3936 26784
rect 3884 26741 3893 26775
rect 3893 26741 3927 26775
rect 3927 26741 3936 26775
rect 3884 26732 3936 26741
rect 6736 26732 6788 26784
rect 8392 26775 8444 26784
rect 8392 26741 8401 26775
rect 8401 26741 8435 26775
rect 8435 26741 8444 26775
rect 8392 26732 8444 26741
rect 8576 26775 8628 26784
rect 8576 26741 8585 26775
rect 8585 26741 8619 26775
rect 8619 26741 8628 26775
rect 8576 26732 8628 26741
rect 13728 26732 13780 26784
rect 17224 26732 17276 26784
rect 20628 26911 20680 26920
rect 20628 26877 20637 26911
rect 20637 26877 20671 26911
rect 20671 26877 20680 26911
rect 20628 26868 20680 26877
rect 20168 26800 20220 26852
rect 20720 26732 20772 26784
rect 23296 26732 23348 26784
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 3332 26528 3384 26580
rect 3516 26528 3568 26580
rect 10968 26528 11020 26580
rect 6736 26435 6788 26444
rect 6736 26401 6745 26435
rect 6745 26401 6779 26435
rect 6779 26401 6788 26435
rect 6736 26392 6788 26401
rect 6828 26324 6880 26376
rect 8576 26460 8628 26512
rect 12532 26528 12584 26580
rect 12440 26460 12492 26512
rect 10232 26256 10284 26308
rect 12348 26392 12400 26444
rect 13728 26435 13780 26444
rect 13728 26401 13737 26435
rect 13737 26401 13771 26435
rect 13771 26401 13780 26435
rect 13728 26392 13780 26401
rect 15292 26435 15344 26444
rect 15292 26401 15301 26435
rect 15301 26401 15335 26435
rect 15335 26401 15344 26435
rect 24308 26528 24360 26580
rect 19248 26503 19300 26512
rect 19248 26469 19257 26503
rect 19257 26469 19291 26503
rect 19291 26469 19300 26503
rect 19248 26460 19300 26469
rect 23388 26460 23440 26512
rect 17868 26435 17920 26444
rect 15292 26392 15344 26401
rect 17868 26401 17877 26435
rect 17877 26401 17911 26435
rect 17911 26401 17920 26435
rect 17868 26392 17920 26401
rect 19340 26392 19392 26444
rect 20536 26392 20588 26444
rect 23204 26435 23256 26444
rect 23204 26401 23213 26435
rect 23213 26401 23247 26435
rect 23247 26401 23256 26435
rect 23204 26392 23256 26401
rect 23296 26435 23348 26444
rect 23296 26401 23305 26435
rect 23305 26401 23339 26435
rect 23339 26401 23348 26435
rect 23296 26392 23348 26401
rect 24860 26392 24912 26444
rect 19432 26367 19484 26376
rect 19432 26333 19441 26367
rect 19441 26333 19475 26367
rect 19475 26333 19484 26367
rect 19432 26324 19484 26333
rect 13820 26256 13872 26308
rect 8024 26231 8076 26240
rect 8024 26197 8033 26231
rect 8033 26197 8067 26231
rect 8067 26197 8076 26231
rect 8024 26188 8076 26197
rect 12440 26188 12492 26240
rect 18236 26188 18288 26240
rect 21088 26231 21140 26240
rect 21088 26197 21097 26231
rect 21097 26197 21131 26231
rect 21131 26197 21140 26231
rect 21088 26188 21140 26197
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 4068 25984 4120 26036
rect 12440 25984 12492 26036
rect 12532 25984 12584 26036
rect 2964 25848 3016 25900
rect 2504 25823 2556 25832
rect 2504 25789 2513 25823
rect 2513 25789 2547 25823
rect 2547 25789 2556 25823
rect 4620 25916 4672 25968
rect 7840 25848 7892 25900
rect 2504 25780 2556 25789
rect 12440 25823 12492 25832
rect 12440 25789 12449 25823
rect 12449 25789 12483 25823
rect 12483 25789 12492 25823
rect 15292 25984 15344 26036
rect 13820 25891 13872 25900
rect 13820 25857 13829 25891
rect 13829 25857 13863 25891
rect 13863 25857 13872 25891
rect 13820 25848 13872 25857
rect 14004 25848 14056 25900
rect 12440 25780 12492 25789
rect 19432 25780 19484 25832
rect 19892 25823 19944 25832
rect 8024 25712 8076 25764
rect 3884 25687 3936 25696
rect 3884 25653 3893 25687
rect 3893 25653 3927 25687
rect 3927 25653 3936 25687
rect 3884 25644 3936 25653
rect 7932 25687 7984 25696
rect 7932 25653 7941 25687
rect 7941 25653 7975 25687
rect 7975 25653 7984 25687
rect 7932 25644 7984 25653
rect 8576 25687 8628 25696
rect 8576 25653 8585 25687
rect 8585 25653 8619 25687
rect 8619 25653 8628 25687
rect 8576 25644 8628 25653
rect 19892 25789 19901 25823
rect 19901 25789 19935 25823
rect 19935 25789 19944 25823
rect 19892 25780 19944 25789
rect 20812 25644 20864 25696
rect 20904 25644 20956 25696
rect 24768 25644 24820 25696
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 8576 25440 8628 25492
rect 7472 25372 7524 25424
rect 10232 25372 10284 25424
rect 3516 25304 3568 25356
rect 3976 25304 4028 25356
rect 11888 25347 11940 25356
rect 6000 25279 6052 25288
rect 6000 25245 6009 25279
rect 6009 25245 6043 25279
rect 6043 25245 6052 25279
rect 6000 25236 6052 25245
rect 11888 25313 11897 25347
rect 11897 25313 11931 25347
rect 11931 25313 11940 25347
rect 14188 25372 14240 25424
rect 11888 25304 11940 25313
rect 16580 25304 16632 25356
rect 17224 25304 17276 25356
rect 11980 25279 12032 25288
rect 11980 25245 11989 25279
rect 11989 25245 12023 25279
rect 12023 25245 12032 25279
rect 11980 25236 12032 25245
rect 12716 25236 12768 25288
rect 7932 25100 7984 25152
rect 12348 25168 12400 25220
rect 21088 25440 21140 25492
rect 19892 25372 19944 25424
rect 20628 25304 20680 25356
rect 21088 25347 21140 25356
rect 21088 25313 21097 25347
rect 21097 25313 21131 25347
rect 21131 25313 21140 25347
rect 21088 25304 21140 25313
rect 21548 25304 21600 25356
rect 21824 25347 21876 25356
rect 21824 25313 21833 25347
rect 21833 25313 21867 25347
rect 21867 25313 21876 25347
rect 21824 25304 21876 25313
rect 20720 25236 20772 25288
rect 22008 25168 22060 25220
rect 12716 25100 12768 25152
rect 20720 25143 20772 25152
rect 20720 25109 20729 25143
rect 20729 25109 20763 25143
rect 20763 25109 20772 25143
rect 20720 25100 20772 25109
rect 22100 25143 22152 25152
rect 22100 25109 22109 25143
rect 22109 25109 22143 25143
rect 22143 25109 22152 25143
rect 22100 25100 22152 25109
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 4896 24760 4948 24812
rect 2504 24735 2556 24744
rect 2504 24701 2513 24735
rect 2513 24701 2547 24735
rect 2547 24701 2556 24735
rect 2504 24692 2556 24701
rect 7932 24760 7984 24812
rect 8484 24803 8536 24812
rect 8484 24769 8493 24803
rect 8493 24769 8527 24803
rect 8527 24769 8536 24803
rect 8484 24760 8536 24769
rect 7104 24735 7156 24744
rect 7104 24701 7113 24735
rect 7113 24701 7147 24735
rect 7147 24701 7156 24735
rect 7104 24692 7156 24701
rect 12348 24692 12400 24744
rect 12624 24692 12676 24744
rect 4068 24624 4120 24676
rect 13452 24667 13504 24676
rect 3240 24556 3292 24608
rect 7932 24556 7984 24608
rect 9036 24556 9088 24608
rect 11428 24556 11480 24608
rect 12532 24599 12584 24608
rect 12532 24565 12541 24599
rect 12541 24565 12575 24599
rect 12575 24565 12584 24599
rect 12532 24556 12584 24565
rect 12624 24556 12676 24608
rect 13452 24633 13461 24667
rect 13461 24633 13495 24667
rect 13495 24633 13504 24667
rect 16488 24692 16540 24744
rect 13452 24624 13504 24633
rect 13544 24556 13596 24608
rect 13728 24599 13780 24608
rect 13728 24565 13737 24599
rect 13737 24565 13771 24599
rect 13771 24565 13780 24599
rect 13728 24556 13780 24565
rect 14648 24556 14700 24608
rect 19340 24556 19392 24608
rect 20536 24556 20588 24608
rect 20812 24556 20864 24608
rect 22100 24760 22152 24812
rect 26792 24692 26844 24744
rect 23572 24624 23624 24676
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 6000 24352 6052 24404
rect 7472 24352 7524 24404
rect 12348 24352 12400 24404
rect 13452 24352 13504 24404
rect 13544 24352 13596 24404
rect 17316 24352 17368 24404
rect 6092 24216 6144 24268
rect 7012 24284 7064 24336
rect 12716 24284 12768 24336
rect 7472 24259 7524 24268
rect 7472 24225 7481 24259
rect 7481 24225 7515 24259
rect 7515 24225 7524 24259
rect 7472 24216 7524 24225
rect 11428 24216 11480 24268
rect 18328 24284 18380 24336
rect 11244 24148 11296 24200
rect 6644 24080 6696 24132
rect 6828 24080 6880 24132
rect 12624 24012 12676 24064
rect 18420 24216 18472 24268
rect 20168 24352 20220 24404
rect 20628 24352 20680 24404
rect 21824 24352 21876 24404
rect 20904 24259 20956 24268
rect 20904 24225 20913 24259
rect 20913 24225 20947 24259
rect 20947 24225 20956 24259
rect 20904 24216 20956 24225
rect 23572 24284 23624 24336
rect 12900 24012 12952 24064
rect 15568 24191 15620 24200
rect 15568 24157 15577 24191
rect 15577 24157 15611 24191
rect 15611 24157 15620 24191
rect 15568 24148 15620 24157
rect 16488 24148 16540 24200
rect 17040 24148 17092 24200
rect 18880 24191 18932 24200
rect 18880 24157 18889 24191
rect 18889 24157 18923 24191
rect 18923 24157 18932 24191
rect 18880 24148 18932 24157
rect 23480 24216 23532 24268
rect 53840 24216 53892 24268
rect 54760 24216 54812 24268
rect 24124 24148 24176 24200
rect 16580 24080 16632 24132
rect 22284 24012 22336 24064
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 2780 23715 2832 23724
rect 2780 23681 2789 23715
rect 2789 23681 2823 23715
rect 2823 23681 2832 23715
rect 2780 23672 2832 23681
rect 2504 23647 2556 23656
rect 2504 23613 2513 23647
rect 2513 23613 2547 23647
rect 2547 23613 2556 23647
rect 2504 23604 2556 23613
rect 8484 23808 8536 23860
rect 8024 23740 8076 23792
rect 12256 23808 12308 23860
rect 12716 23808 12768 23860
rect 15568 23808 15620 23860
rect 18788 23808 18840 23860
rect 20996 23808 21048 23860
rect 12808 23740 12860 23792
rect 12256 23672 12308 23724
rect 13636 23672 13688 23724
rect 17776 23672 17828 23724
rect 20720 23740 20772 23792
rect 9864 23604 9916 23656
rect 10876 23647 10928 23656
rect 10876 23613 10885 23647
rect 10885 23613 10919 23647
rect 10919 23613 10928 23647
rect 10876 23604 10928 23613
rect 11244 23604 11296 23656
rect 12440 23647 12492 23656
rect 12440 23613 12449 23647
rect 12449 23613 12483 23647
rect 12483 23613 12492 23647
rect 12440 23604 12492 23613
rect 12808 23604 12860 23656
rect 12532 23536 12584 23588
rect 14464 23647 14516 23656
rect 14464 23613 14473 23647
rect 14473 23613 14507 23647
rect 14507 23613 14516 23647
rect 14648 23647 14700 23656
rect 14464 23604 14516 23613
rect 14648 23613 14657 23647
rect 14657 23613 14691 23647
rect 14691 23613 14700 23647
rect 14648 23604 14700 23613
rect 3884 23511 3936 23520
rect 3884 23477 3893 23511
rect 3893 23477 3927 23511
rect 3927 23477 3936 23511
rect 3884 23468 3936 23477
rect 4620 23468 4672 23520
rect 6920 23468 6972 23520
rect 10876 23468 10928 23520
rect 18604 23536 18656 23588
rect 18880 23604 18932 23656
rect 20168 23604 20220 23656
rect 21548 23647 21600 23656
rect 21548 23613 21557 23647
rect 21557 23613 21591 23647
rect 21591 23613 21600 23647
rect 21548 23604 21600 23613
rect 22284 23647 22336 23656
rect 22284 23613 22293 23647
rect 22293 23613 22327 23647
rect 22327 23613 22336 23647
rect 22284 23604 22336 23613
rect 17776 23511 17828 23520
rect 17776 23477 17785 23511
rect 17785 23477 17819 23511
rect 17819 23477 17828 23511
rect 17776 23468 17828 23477
rect 19248 23511 19300 23520
rect 19248 23477 19257 23511
rect 19257 23477 19291 23511
rect 19291 23477 19300 23511
rect 19248 23468 19300 23477
rect 20168 23511 20220 23520
rect 20168 23477 20177 23511
rect 20177 23477 20211 23511
rect 20211 23477 20220 23511
rect 20168 23468 20220 23477
rect 22560 23511 22612 23520
rect 22560 23477 22569 23511
rect 22569 23477 22603 23511
rect 22603 23477 22612 23511
rect 22560 23468 22612 23477
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 4068 23264 4120 23316
rect 23020 23264 23072 23316
rect 7104 23196 7156 23248
rect 6184 23171 6236 23180
rect 6184 23137 6193 23171
rect 6193 23137 6227 23171
rect 6227 23137 6236 23171
rect 6184 23128 6236 23137
rect 6920 23128 6972 23180
rect 7748 23128 7800 23180
rect 11888 23128 11940 23180
rect 12624 23196 12676 23248
rect 20168 23196 20220 23248
rect 12808 23171 12860 23180
rect 12808 23137 12817 23171
rect 12817 23137 12851 23171
rect 12851 23137 12860 23171
rect 12808 23128 12860 23137
rect 12992 23171 13044 23180
rect 12992 23137 13001 23171
rect 13001 23137 13035 23171
rect 13035 23137 13044 23171
rect 12992 23128 13044 23137
rect 19248 23128 19300 23180
rect 22560 23128 22612 23180
rect 5264 23060 5316 23112
rect 12532 23103 12584 23112
rect 12532 23069 12541 23103
rect 12541 23069 12575 23103
rect 12575 23069 12584 23103
rect 12532 23060 12584 23069
rect 19616 23060 19668 23112
rect 20812 23060 20864 23112
rect 21640 23060 21692 23112
rect 7288 22992 7340 23044
rect 6184 22924 6236 22976
rect 7472 22924 7524 22976
rect 9772 22967 9824 22976
rect 9772 22933 9781 22967
rect 9781 22933 9815 22967
rect 9815 22933 9824 22967
rect 9772 22924 9824 22933
rect 12072 22967 12124 22976
rect 12072 22933 12081 22967
rect 12081 22933 12115 22967
rect 12115 22933 12124 22967
rect 12072 22924 12124 22933
rect 23480 22967 23532 22976
rect 23480 22933 23489 22967
rect 23489 22933 23523 22967
rect 23523 22933 23532 22967
rect 23480 22924 23532 22933
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 81624 22856 81676 22908
rect 82268 22856 82320 22908
rect 3148 22720 3200 22772
rect 4620 22720 4672 22772
rect 9036 22763 9088 22772
rect 9036 22729 9045 22763
rect 9045 22729 9079 22763
rect 9079 22729 9088 22763
rect 9036 22720 9088 22729
rect 9680 22763 9732 22772
rect 9680 22729 9689 22763
rect 9689 22729 9723 22763
rect 9723 22729 9732 22763
rect 9680 22720 9732 22729
rect 12532 22584 12584 22636
rect 12808 22584 12860 22636
rect 2504 22559 2556 22568
rect 2504 22525 2513 22559
rect 2513 22525 2547 22559
rect 2547 22525 2556 22559
rect 2504 22516 2556 22525
rect 7932 22516 7984 22568
rect 9680 22516 9732 22568
rect 13912 22720 13964 22772
rect 19616 22627 19668 22636
rect 19616 22593 19625 22627
rect 19625 22593 19659 22627
rect 19659 22593 19668 22627
rect 19616 22584 19668 22593
rect 5632 22448 5684 22500
rect 12440 22491 12492 22500
rect 12440 22457 12449 22491
rect 12449 22457 12483 22491
rect 12483 22457 12492 22491
rect 12440 22448 12492 22457
rect 12624 22448 12676 22500
rect 14648 22516 14700 22568
rect 19892 22559 19944 22568
rect 19892 22525 19901 22559
rect 19901 22525 19935 22559
rect 19935 22525 19944 22559
rect 19892 22516 19944 22525
rect 18420 22448 18472 22500
rect 21272 22491 21324 22500
rect 21272 22457 21281 22491
rect 21281 22457 21315 22491
rect 21315 22457 21324 22491
rect 21272 22448 21324 22457
rect 9956 22380 10008 22432
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 4620 22176 4672 22228
rect 7932 22219 7984 22228
rect 4712 22040 4764 22092
rect 7932 22185 7941 22219
rect 7941 22185 7975 22219
rect 7975 22185 7984 22219
rect 7932 22176 7984 22185
rect 12716 22176 12768 22228
rect 18328 22219 18380 22228
rect 18328 22185 18337 22219
rect 18337 22185 18371 22219
rect 18371 22185 18380 22219
rect 18328 22176 18380 22185
rect 7748 22108 7800 22160
rect 7472 22083 7524 22092
rect 7472 22049 7481 22083
rect 7481 22049 7515 22083
rect 7515 22049 7524 22083
rect 7472 22040 7524 22049
rect 4068 21836 4120 21888
rect 6644 21879 6696 21888
rect 6644 21845 6653 21879
rect 6653 21845 6687 21879
rect 6687 21845 6696 21879
rect 9128 22040 9180 22092
rect 12440 22040 12492 22092
rect 13268 22108 13320 22160
rect 18696 22108 18748 22160
rect 9496 21972 9548 22024
rect 9864 21947 9916 21956
rect 9864 21913 9873 21947
rect 9873 21913 9907 21947
rect 9907 21913 9916 21947
rect 9864 21904 9916 21913
rect 12716 21972 12768 22024
rect 12808 21972 12860 22024
rect 13820 22040 13872 22092
rect 14188 22040 14240 22092
rect 14464 22040 14516 22092
rect 18420 22040 18472 22092
rect 20076 22176 20128 22228
rect 21272 22151 21324 22160
rect 21272 22117 21281 22151
rect 21281 22117 21315 22151
rect 21315 22117 21324 22151
rect 21272 22108 21324 22117
rect 24492 22040 24544 22092
rect 14096 21972 14148 22024
rect 18052 21972 18104 22024
rect 19064 21972 19116 22024
rect 28448 21904 28500 21956
rect 6644 21836 6696 21845
rect 9956 21836 10008 21888
rect 11704 21836 11756 21888
rect 12256 21879 12308 21888
rect 12256 21845 12265 21879
rect 12265 21845 12299 21879
rect 12299 21845 12308 21879
rect 12256 21836 12308 21845
rect 14096 21836 14148 21888
rect 15844 21836 15896 21888
rect 19156 21836 19208 21888
rect 24124 21879 24176 21888
rect 24124 21845 24133 21879
rect 24133 21845 24167 21879
rect 24167 21845 24176 21879
rect 24124 21836 24176 21845
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 5172 21632 5224 21684
rect 7748 21632 7800 21684
rect 9312 21675 9364 21684
rect 9312 21641 9321 21675
rect 9321 21641 9355 21675
rect 9355 21641 9364 21675
rect 9312 21632 9364 21641
rect 2504 21471 2556 21480
rect 2504 21437 2513 21471
rect 2513 21437 2547 21471
rect 2547 21437 2556 21471
rect 4620 21564 4672 21616
rect 6644 21564 6696 21616
rect 17132 21632 17184 21684
rect 19892 21632 19944 21684
rect 14096 21564 14148 21616
rect 5632 21496 5684 21548
rect 6184 21496 6236 21548
rect 2504 21428 2556 21437
rect 5724 21428 5776 21480
rect 9772 21496 9824 21548
rect 12440 21539 12492 21548
rect 12440 21505 12449 21539
rect 12449 21505 12483 21539
rect 12483 21505 12492 21539
rect 12716 21539 12768 21548
rect 12440 21496 12492 21505
rect 12716 21505 12725 21539
rect 12725 21505 12759 21539
rect 12759 21505 12768 21539
rect 12716 21496 12768 21505
rect 22376 21496 22428 21548
rect 22928 21496 22980 21548
rect 6736 21360 6788 21412
rect 9128 21471 9180 21480
rect 9128 21437 9137 21471
rect 9137 21437 9171 21471
rect 9171 21437 9180 21471
rect 9128 21428 9180 21437
rect 9312 21428 9364 21480
rect 14464 21428 14516 21480
rect 18604 21471 18656 21480
rect 3148 21292 3200 21344
rect 12532 21360 12584 21412
rect 12256 21292 12308 21344
rect 12716 21292 12768 21344
rect 18604 21437 18613 21471
rect 18613 21437 18647 21471
rect 18647 21437 18656 21471
rect 18604 21428 18656 21437
rect 19064 21471 19116 21480
rect 19064 21437 19073 21471
rect 19073 21437 19107 21471
rect 19107 21437 19116 21471
rect 19064 21428 19116 21437
rect 19156 21471 19208 21480
rect 19156 21437 19165 21471
rect 19165 21437 19199 21471
rect 19199 21437 19208 21471
rect 19156 21428 19208 21437
rect 21180 21428 21232 21480
rect 22468 21428 22520 21480
rect 18788 21292 18840 21344
rect 22284 21335 22336 21344
rect 22284 21301 22293 21335
rect 22293 21301 22327 21335
rect 22327 21301 22336 21335
rect 22284 21292 22336 21301
rect 22560 21335 22612 21344
rect 22560 21301 22569 21335
rect 22569 21301 22603 21335
rect 22603 21301 22612 21335
rect 22560 21292 22612 21301
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 7104 21088 7156 21140
rect 7564 21020 7616 21072
rect 7840 21063 7892 21072
rect 7840 21029 7849 21063
rect 7849 21029 7883 21063
rect 7883 21029 7892 21063
rect 7840 21020 7892 21029
rect 7288 20995 7340 21004
rect 7288 20961 7297 20995
rect 7297 20961 7331 20995
rect 7331 20961 7340 20995
rect 7288 20952 7340 20961
rect 15292 20995 15344 21004
rect 15292 20961 15301 20995
rect 15301 20961 15335 20995
rect 15335 20961 15344 20995
rect 15292 20952 15344 20961
rect 15660 20952 15712 21004
rect 21640 20995 21692 21004
rect 21640 20961 21649 20995
rect 21649 20961 21683 20995
rect 21683 20961 21692 20995
rect 21640 20952 21692 20961
rect 7196 20884 7248 20936
rect 12440 20884 12492 20936
rect 12992 20927 13044 20936
rect 12992 20893 13001 20927
rect 13001 20893 13035 20927
rect 13035 20893 13044 20927
rect 12992 20884 13044 20893
rect 14556 20884 14608 20936
rect 22376 21088 22428 21140
rect 22560 21088 22612 21140
rect 21916 20927 21968 20936
rect 21916 20893 21925 20927
rect 21925 20893 21959 20927
rect 21959 20893 21968 20927
rect 21916 20884 21968 20893
rect 13820 20816 13872 20868
rect 12900 20748 12952 20800
rect 13728 20748 13780 20800
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 4620 20544 4672 20596
rect 2504 20451 2556 20460
rect 2504 20417 2513 20451
rect 2513 20417 2547 20451
rect 2547 20417 2556 20451
rect 2504 20408 2556 20417
rect 3516 20408 3568 20460
rect 6920 20383 6972 20392
rect 6920 20349 6929 20383
rect 6929 20349 6963 20383
rect 6963 20349 6972 20383
rect 6920 20340 6972 20349
rect 3884 20247 3936 20256
rect 3884 20213 3893 20247
rect 3893 20213 3927 20247
rect 3927 20213 3936 20247
rect 3884 20204 3936 20213
rect 8116 20340 8168 20392
rect 8760 20544 8812 20596
rect 15384 20587 15436 20596
rect 15384 20553 15393 20587
rect 15393 20553 15427 20587
rect 15427 20553 15436 20587
rect 15384 20544 15436 20553
rect 19984 20544 20036 20596
rect 13728 20451 13780 20460
rect 13728 20417 13737 20451
rect 13737 20417 13771 20451
rect 13771 20417 13780 20451
rect 13728 20408 13780 20417
rect 13912 20340 13964 20392
rect 8024 20315 8076 20324
rect 8024 20281 8033 20315
rect 8033 20281 8067 20315
rect 8067 20281 8076 20315
rect 8024 20272 8076 20281
rect 8484 20204 8536 20256
rect 19432 20204 19484 20256
rect 19984 20340 20036 20392
rect 20812 20383 20864 20392
rect 20812 20349 20821 20383
rect 20821 20349 20855 20383
rect 20855 20349 20864 20383
rect 20812 20340 20864 20349
rect 22560 20340 22612 20392
rect 23112 20544 23164 20596
rect 20628 20204 20680 20256
rect 20812 20204 20864 20256
rect 21272 20204 21324 20256
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 6184 20043 6236 20052
rect 6184 20009 6193 20043
rect 6193 20009 6227 20043
rect 6227 20009 6236 20043
rect 6184 20000 6236 20009
rect 8116 20043 8168 20052
rect 8116 20009 8125 20043
rect 8125 20009 8159 20043
rect 8159 20009 8168 20043
rect 8116 20000 8168 20009
rect 14556 20043 14608 20052
rect 14556 20009 14565 20043
rect 14565 20009 14599 20043
rect 14599 20009 14608 20043
rect 14556 20000 14608 20009
rect 22560 20043 22612 20052
rect 22560 20009 22569 20043
rect 22569 20009 22603 20043
rect 22603 20009 22612 20043
rect 22560 20000 22612 20009
rect 9128 19932 9180 19984
rect 12992 19932 13044 19984
rect 5356 19796 5408 19848
rect 6552 19864 6604 19916
rect 7012 19907 7064 19916
rect 7012 19873 7021 19907
rect 7021 19873 7055 19907
rect 7055 19873 7064 19907
rect 7012 19864 7064 19873
rect 7288 19796 7340 19848
rect 7472 19796 7524 19848
rect 8116 19864 8168 19916
rect 9312 19864 9364 19916
rect 7840 19839 7892 19848
rect 7840 19805 7849 19839
rect 7849 19805 7883 19839
rect 7883 19805 7892 19839
rect 7840 19796 7892 19805
rect 8484 19660 8536 19712
rect 10784 19660 10836 19712
rect 13636 19907 13688 19916
rect 13636 19873 13645 19907
rect 13645 19873 13679 19907
rect 13679 19873 13688 19907
rect 13636 19864 13688 19873
rect 13820 19907 13872 19916
rect 13820 19873 13829 19907
rect 13829 19873 13863 19907
rect 13863 19873 13872 19907
rect 13820 19864 13872 19873
rect 12716 19796 12768 19848
rect 14188 19864 14240 19916
rect 14924 19864 14976 19916
rect 15292 19907 15344 19916
rect 15292 19873 15301 19907
rect 15301 19873 15335 19907
rect 15335 19873 15344 19907
rect 15292 19864 15344 19873
rect 21272 19907 21324 19916
rect 21272 19873 21281 19907
rect 21281 19873 21315 19907
rect 21315 19873 21324 19907
rect 21272 19864 21324 19873
rect 19432 19796 19484 19848
rect 20996 19839 21048 19848
rect 20996 19805 21005 19839
rect 21005 19805 21039 19839
rect 21039 19805 21048 19839
rect 20996 19796 21048 19805
rect 12716 19703 12768 19712
rect 12716 19669 12725 19703
rect 12725 19669 12759 19703
rect 12759 19669 12768 19703
rect 12716 19660 12768 19669
rect 15384 19660 15436 19712
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 15292 19456 15344 19508
rect 19984 19499 20036 19508
rect 19984 19465 19993 19499
rect 19993 19465 20027 19499
rect 20027 19465 20036 19499
rect 19984 19456 20036 19465
rect 14556 19388 14608 19440
rect 8300 19320 8352 19372
rect 12348 19320 12400 19372
rect 13820 19320 13872 19372
rect 14924 19363 14976 19372
rect 14924 19329 14933 19363
rect 14933 19329 14967 19363
rect 14967 19329 14976 19363
rect 14924 19320 14976 19329
rect 7196 19252 7248 19304
rect 7012 19227 7064 19236
rect 7012 19193 7021 19227
rect 7021 19193 7055 19227
rect 7055 19193 7064 19227
rect 7012 19184 7064 19193
rect 7104 19184 7156 19236
rect 8392 19252 8444 19304
rect 8668 19252 8720 19304
rect 9404 19295 9456 19304
rect 9404 19261 9413 19295
rect 9413 19261 9447 19295
rect 9447 19261 9456 19295
rect 9404 19252 9456 19261
rect 9772 19252 9824 19304
rect 7656 19184 7708 19236
rect 8484 19184 8536 19236
rect 12624 19252 12676 19304
rect 13912 19252 13964 19304
rect 14096 19295 14148 19304
rect 14096 19261 14105 19295
rect 14105 19261 14139 19295
rect 14139 19261 14148 19295
rect 14096 19252 14148 19261
rect 14372 19295 14424 19304
rect 5908 19116 5960 19168
rect 8668 19116 8720 19168
rect 8852 19159 8904 19168
rect 8852 19125 8861 19159
rect 8861 19125 8895 19159
rect 8895 19125 8904 19159
rect 13636 19184 13688 19236
rect 14372 19261 14381 19295
rect 14381 19261 14415 19295
rect 14415 19261 14424 19295
rect 14372 19252 14424 19261
rect 15200 19252 15252 19304
rect 18052 19295 18104 19304
rect 18052 19261 18061 19295
rect 18061 19261 18095 19295
rect 18095 19261 18104 19295
rect 18052 19252 18104 19261
rect 16120 19184 16172 19236
rect 8852 19116 8904 19125
rect 10324 19159 10376 19168
rect 10324 19125 10333 19159
rect 10333 19125 10367 19159
rect 10367 19125 10376 19159
rect 10324 19116 10376 19125
rect 12532 19116 12584 19168
rect 13452 19159 13504 19168
rect 13452 19125 13461 19159
rect 13461 19125 13495 19159
rect 13495 19125 13504 19159
rect 13452 19116 13504 19125
rect 14096 19116 14148 19168
rect 21916 19456 21968 19508
rect 54116 19363 54168 19372
rect 54116 19329 54125 19363
rect 54125 19329 54159 19363
rect 54159 19329 54168 19363
rect 54116 19320 54168 19329
rect 22284 19252 22336 19304
rect 18144 19159 18196 19168
rect 18144 19125 18153 19159
rect 18153 19125 18187 19159
rect 18187 19125 18196 19159
rect 18144 19116 18196 19125
rect 20720 19116 20772 19168
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 3332 18912 3384 18964
rect 22836 18912 22888 18964
rect 5356 18844 5408 18896
rect 6736 18844 6788 18896
rect 5908 18819 5960 18828
rect 5908 18785 5917 18819
rect 5917 18785 5951 18819
rect 5951 18785 5960 18819
rect 5908 18776 5960 18785
rect 6000 18819 6052 18828
rect 6000 18785 6009 18819
rect 6009 18785 6043 18819
rect 6043 18785 6052 18819
rect 6000 18776 6052 18785
rect 7104 18776 7156 18828
rect 7656 18819 7708 18828
rect 7656 18785 7665 18819
rect 7665 18785 7699 18819
rect 7699 18785 7708 18819
rect 7656 18776 7708 18785
rect 7840 18819 7892 18828
rect 7840 18785 7849 18819
rect 7849 18785 7883 18819
rect 7883 18785 7892 18819
rect 7840 18776 7892 18785
rect 8116 18819 8168 18828
rect 8116 18785 8125 18819
rect 8125 18785 8159 18819
rect 8159 18785 8168 18819
rect 8116 18776 8168 18785
rect 9036 18844 9088 18896
rect 16580 18844 16632 18896
rect 13636 18819 13688 18828
rect 6460 18751 6512 18760
rect 6460 18717 6469 18751
rect 6469 18717 6503 18751
rect 6503 18717 6512 18751
rect 6460 18708 6512 18717
rect 13636 18785 13645 18819
rect 13645 18785 13679 18819
rect 13679 18785 13688 18819
rect 13636 18776 13688 18785
rect 14004 18819 14056 18828
rect 14004 18785 14013 18819
rect 14013 18785 14047 18819
rect 14047 18785 14056 18819
rect 14004 18776 14056 18785
rect 14372 18819 14424 18828
rect 14372 18785 14381 18819
rect 14381 18785 14415 18819
rect 14415 18785 14424 18819
rect 14372 18776 14424 18785
rect 15384 18819 15436 18828
rect 15384 18785 15393 18819
rect 15393 18785 15427 18819
rect 15427 18785 15436 18819
rect 15384 18776 15436 18785
rect 17960 18819 18012 18828
rect 17960 18785 17969 18819
rect 17969 18785 18003 18819
rect 18003 18785 18012 18819
rect 17960 18776 18012 18785
rect 18052 18819 18104 18828
rect 18052 18785 18061 18819
rect 18061 18785 18095 18819
rect 18095 18785 18104 18819
rect 18052 18776 18104 18785
rect 7472 18640 7524 18692
rect 10324 18640 10376 18692
rect 7748 18572 7800 18624
rect 9128 18615 9180 18624
rect 9128 18581 9137 18615
rect 9137 18581 9171 18615
rect 9171 18581 9180 18615
rect 9128 18572 9180 18581
rect 15844 18708 15896 18760
rect 21732 18708 21784 18760
rect 22192 18751 22244 18760
rect 22192 18717 22201 18751
rect 22201 18717 22235 18751
rect 22235 18717 22244 18751
rect 22192 18708 22244 18717
rect 14004 18640 14056 18692
rect 14372 18572 14424 18624
rect 15568 18615 15620 18624
rect 15568 18581 15577 18615
rect 15577 18581 15611 18615
rect 15611 18581 15620 18615
rect 15568 18572 15620 18581
rect 18236 18615 18288 18624
rect 18236 18581 18245 18615
rect 18245 18581 18279 18615
rect 18279 18581 18288 18615
rect 18236 18572 18288 18581
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 4252 18232 4304 18284
rect 4988 18368 5040 18420
rect 6000 18368 6052 18420
rect 9036 18411 9088 18420
rect 9036 18377 9045 18411
rect 9045 18377 9079 18411
rect 9079 18377 9088 18411
rect 9036 18368 9088 18377
rect 12624 18368 12676 18420
rect 15292 18368 15344 18420
rect 18696 18411 18748 18420
rect 18696 18377 18705 18411
rect 18705 18377 18739 18411
rect 18739 18377 18748 18411
rect 18696 18368 18748 18377
rect 22192 18411 22244 18420
rect 22192 18377 22201 18411
rect 22201 18377 22235 18411
rect 22235 18377 22244 18411
rect 22192 18368 22244 18377
rect 6460 18300 6512 18352
rect 9680 18300 9732 18352
rect 10784 18300 10836 18352
rect 12532 18300 12584 18352
rect 13636 18232 13688 18284
rect 5632 18207 5684 18216
rect 5632 18173 5641 18207
rect 5641 18173 5675 18207
rect 5675 18173 5684 18207
rect 5632 18164 5684 18173
rect 8024 18207 8076 18216
rect 8024 18173 8033 18207
rect 8033 18173 8067 18207
rect 8067 18173 8076 18207
rect 8024 18164 8076 18173
rect 8300 18096 8352 18148
rect 3884 18071 3936 18080
rect 3884 18037 3893 18071
rect 3893 18037 3927 18071
rect 3927 18037 3936 18071
rect 3884 18028 3936 18037
rect 4252 18028 4304 18080
rect 4988 18028 5040 18080
rect 9036 18164 9088 18216
rect 9220 18164 9272 18216
rect 13084 18164 13136 18216
rect 9404 18096 9456 18148
rect 8576 18028 8628 18080
rect 9496 18028 9548 18080
rect 14004 18164 14056 18216
rect 14096 18028 14148 18080
rect 15384 18164 15436 18216
rect 18052 18164 18104 18216
rect 20168 18300 20220 18352
rect 21180 18300 21232 18352
rect 21824 18300 21876 18352
rect 16948 18139 17000 18148
rect 16948 18105 16957 18139
rect 16957 18105 16991 18139
rect 16991 18105 17000 18139
rect 16948 18096 17000 18105
rect 18696 18096 18748 18148
rect 20720 18164 20772 18216
rect 21180 18207 21232 18216
rect 21180 18173 21189 18207
rect 21189 18173 21223 18207
rect 21223 18173 21232 18207
rect 21180 18164 21232 18173
rect 21640 18207 21692 18216
rect 21640 18173 21649 18207
rect 21649 18173 21683 18207
rect 21683 18173 21692 18207
rect 21640 18164 21692 18173
rect 21824 18164 21876 18216
rect 17592 18028 17644 18080
rect 19432 18028 19484 18080
rect 22284 18096 22336 18148
rect 19984 18028 20036 18080
rect 20720 18028 20772 18080
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 6552 17824 6604 17876
rect 12992 17824 13044 17876
rect 14004 17824 14056 17876
rect 21640 17824 21692 17876
rect 26976 17892 27028 17944
rect 4620 17688 4672 17740
rect 6552 17731 6604 17740
rect 6552 17697 6561 17731
rect 6561 17697 6595 17731
rect 6595 17697 6604 17731
rect 6552 17688 6604 17697
rect 6736 17688 6788 17740
rect 5908 17552 5960 17604
rect 12072 17688 12124 17740
rect 18052 17688 18104 17740
rect 19432 17688 19484 17740
rect 8024 17620 8076 17672
rect 18328 17620 18380 17672
rect 9128 17552 9180 17604
rect 12072 17552 12124 17604
rect 15936 17552 15988 17604
rect 16672 17552 16724 17604
rect 7012 17484 7064 17536
rect 7656 17484 7708 17536
rect 8300 17484 8352 17536
rect 13084 17484 13136 17536
rect 14188 17484 14240 17536
rect 18420 17527 18472 17536
rect 18420 17493 18429 17527
rect 18429 17493 18463 17527
rect 18463 17493 18472 17527
rect 18420 17484 18472 17493
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 6552 17280 6604 17332
rect 5816 17212 5868 17264
rect 10232 17212 10284 17264
rect 5724 17187 5776 17196
rect 5724 17153 5733 17187
rect 5733 17153 5767 17187
rect 5767 17153 5776 17187
rect 5724 17144 5776 17153
rect 3884 17119 3936 17128
rect 3884 17085 3893 17119
rect 3893 17085 3927 17119
rect 3927 17085 3936 17119
rect 3884 17076 3936 17085
rect 4620 17008 4672 17060
rect 2872 16940 2924 16992
rect 5356 17076 5408 17128
rect 7012 17076 7064 17128
rect 14188 17187 14240 17196
rect 14188 17153 14197 17187
rect 14197 17153 14231 17187
rect 14231 17153 14240 17187
rect 14188 17144 14240 17153
rect 15568 17280 15620 17332
rect 15936 17280 15988 17332
rect 19984 17323 20036 17332
rect 19984 17289 19993 17323
rect 19993 17289 20027 17323
rect 20027 17289 20036 17323
rect 19984 17280 20036 17289
rect 20168 17323 20220 17332
rect 20168 17289 20177 17323
rect 20177 17289 20211 17323
rect 20211 17289 20220 17323
rect 20168 17280 20220 17289
rect 16488 17212 16540 17264
rect 19892 17255 19944 17264
rect 7472 17119 7524 17128
rect 7472 17085 7481 17119
rect 7481 17085 7515 17119
rect 7515 17085 7524 17119
rect 7472 17076 7524 17085
rect 7656 17119 7708 17128
rect 7656 17085 7665 17119
rect 7665 17085 7699 17119
rect 7699 17085 7708 17119
rect 7656 17076 7708 17085
rect 8300 17119 8352 17128
rect 8300 17085 8309 17119
rect 8309 17085 8343 17119
rect 8343 17085 8352 17119
rect 8300 17076 8352 17085
rect 9128 17119 9180 17128
rect 9128 17085 9137 17119
rect 9137 17085 9171 17119
rect 9171 17085 9180 17119
rect 9128 17076 9180 17085
rect 10968 17119 11020 17128
rect 10968 17085 10977 17119
rect 10977 17085 11011 17119
rect 11011 17085 11020 17119
rect 10968 17076 11020 17085
rect 11152 17076 11204 17128
rect 14740 17119 14792 17128
rect 14740 17085 14749 17119
rect 14749 17085 14783 17119
rect 14783 17085 14792 17119
rect 14740 17076 14792 17085
rect 18144 17144 18196 17196
rect 15200 17119 15252 17128
rect 15200 17085 15209 17119
rect 15209 17085 15243 17119
rect 15243 17085 15252 17119
rect 15200 17076 15252 17085
rect 11520 17051 11572 17060
rect 11520 17017 11529 17051
rect 11529 17017 11563 17051
rect 11563 17017 11572 17051
rect 11520 17008 11572 17017
rect 17040 17076 17092 17128
rect 18236 17119 18288 17128
rect 18236 17085 18245 17119
rect 18245 17085 18279 17119
rect 18279 17085 18288 17119
rect 18236 17076 18288 17085
rect 18604 17119 18656 17128
rect 18604 17085 18613 17119
rect 18613 17085 18647 17119
rect 18647 17085 18656 17119
rect 18604 17076 18656 17085
rect 19156 17144 19208 17196
rect 19064 17119 19116 17128
rect 19064 17085 19073 17119
rect 19073 17085 19107 17119
rect 19107 17085 19116 17119
rect 19064 17076 19116 17085
rect 18972 17008 19024 17060
rect 19892 17221 19901 17255
rect 19901 17221 19935 17255
rect 19935 17221 19944 17255
rect 19892 17212 19944 17221
rect 20812 17187 20864 17196
rect 20812 17153 20821 17187
rect 20821 17153 20855 17187
rect 20855 17153 20864 17187
rect 20812 17144 20864 17153
rect 19432 17076 19484 17128
rect 21548 17119 21600 17128
rect 21548 17085 21557 17119
rect 21557 17085 21591 17119
rect 21591 17085 21600 17119
rect 21548 17076 21600 17085
rect 27068 17280 27120 17332
rect 21824 17212 21876 17264
rect 24124 17076 24176 17128
rect 7840 16940 7892 16992
rect 9312 16983 9364 16992
rect 9312 16949 9321 16983
rect 9321 16949 9355 16983
rect 9355 16949 9364 16983
rect 9312 16940 9364 16949
rect 10968 16940 11020 16992
rect 12440 16940 12492 16992
rect 15568 16983 15620 16992
rect 15568 16949 15577 16983
rect 15577 16949 15611 16983
rect 15611 16949 15620 16983
rect 15568 16940 15620 16949
rect 18052 16940 18104 16992
rect 19064 16940 19116 16992
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 3884 16736 3936 16788
rect 5356 16736 5408 16788
rect 7288 16736 7340 16788
rect 8024 16736 8076 16788
rect 14740 16736 14792 16788
rect 17224 16736 17276 16788
rect 21548 16736 21600 16788
rect 4620 16668 4672 16720
rect 4896 16643 4948 16652
rect 4896 16609 4905 16643
rect 4905 16609 4939 16643
rect 4939 16609 4948 16643
rect 4896 16600 4948 16609
rect 5632 16600 5684 16652
rect 9220 16668 9272 16720
rect 11336 16668 11388 16720
rect 11796 16668 11848 16720
rect 18328 16668 18380 16720
rect 21824 16668 21876 16720
rect 6736 16643 6788 16652
rect 5816 16532 5868 16584
rect 6736 16609 6745 16643
rect 6745 16609 6779 16643
rect 6779 16609 6788 16643
rect 6736 16600 6788 16609
rect 7840 16643 7892 16652
rect 7840 16609 7849 16643
rect 7849 16609 7883 16643
rect 7883 16609 7892 16643
rect 7840 16600 7892 16609
rect 9312 16600 9364 16652
rect 11060 16600 11112 16652
rect 11520 16600 11572 16652
rect 7012 16532 7064 16584
rect 13084 16643 13136 16652
rect 13084 16609 13093 16643
rect 13093 16609 13127 16643
rect 13127 16609 13136 16643
rect 13084 16600 13136 16609
rect 16672 16643 16724 16652
rect 16672 16609 16681 16643
rect 16681 16609 16715 16643
rect 16715 16609 16724 16643
rect 16672 16600 16724 16609
rect 16948 16643 17000 16652
rect 16948 16609 16957 16643
rect 16957 16609 16991 16643
rect 16991 16609 17000 16643
rect 16948 16600 17000 16609
rect 17224 16643 17276 16652
rect 17224 16609 17233 16643
rect 17233 16609 17267 16643
rect 17267 16609 17276 16643
rect 17224 16600 17276 16609
rect 17316 16600 17368 16652
rect 17592 16643 17644 16652
rect 11888 16575 11940 16584
rect 11888 16541 11897 16575
rect 11897 16541 11931 16575
rect 11931 16541 11940 16575
rect 12992 16575 13044 16584
rect 11888 16532 11940 16541
rect 12992 16541 13001 16575
rect 13001 16541 13035 16575
rect 13035 16541 13044 16575
rect 12992 16532 13044 16541
rect 13544 16575 13596 16584
rect 13544 16541 13553 16575
rect 13553 16541 13587 16575
rect 13587 16541 13596 16575
rect 13544 16532 13596 16541
rect 17592 16609 17601 16643
rect 17601 16609 17635 16643
rect 17635 16609 17644 16643
rect 17592 16600 17644 16609
rect 18512 16643 18564 16652
rect 18512 16609 18521 16643
rect 18521 16609 18555 16643
rect 18555 16609 18564 16643
rect 18512 16600 18564 16609
rect 18972 16643 19024 16652
rect 18972 16609 18981 16643
rect 18981 16609 19015 16643
rect 19015 16609 19024 16643
rect 18972 16600 19024 16609
rect 22652 16600 22704 16652
rect 23572 16600 23624 16652
rect 17960 16575 18012 16584
rect 17960 16541 17969 16575
rect 17969 16541 18003 16575
rect 18003 16541 18012 16575
rect 17960 16532 18012 16541
rect 7472 16464 7524 16516
rect 11704 16507 11756 16516
rect 11704 16473 11713 16507
rect 11713 16473 11747 16507
rect 11747 16473 11756 16507
rect 11704 16464 11756 16473
rect 12440 16464 12492 16516
rect 26884 16464 26936 16516
rect 4804 16439 4856 16448
rect 4804 16405 4813 16439
rect 4813 16405 4847 16439
rect 4847 16405 4856 16439
rect 4804 16396 4856 16405
rect 16580 16396 16632 16448
rect 17592 16396 17644 16448
rect 19064 16396 19116 16448
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 5356 16192 5408 16244
rect 20628 16192 20680 16244
rect 7472 16124 7524 16176
rect 9956 16056 10008 16108
rect 10784 16099 10836 16108
rect 2504 16031 2556 16040
rect 2504 15997 2513 16031
rect 2513 15997 2547 16031
rect 2547 15997 2556 16031
rect 2504 15988 2556 15997
rect 3056 15988 3108 16040
rect 7012 16031 7064 16040
rect 4804 15920 4856 15972
rect 7012 15997 7021 16031
rect 7021 15997 7055 16031
rect 7055 15997 7064 16031
rect 7012 15988 7064 15997
rect 7288 16031 7340 16040
rect 7288 15997 7297 16031
rect 7297 15997 7331 16031
rect 7331 15997 7340 16031
rect 7288 15988 7340 15997
rect 10784 16065 10793 16099
rect 10793 16065 10827 16099
rect 10827 16065 10836 16099
rect 10784 16056 10836 16065
rect 11152 16056 11204 16108
rect 18052 16099 18104 16108
rect 10416 16031 10468 16040
rect 10416 15997 10425 16031
rect 10425 15997 10459 16031
rect 10459 15997 10468 16031
rect 10416 15988 10468 15997
rect 18052 16065 18061 16099
rect 18061 16065 18095 16099
rect 18095 16065 18104 16099
rect 18052 16056 18104 16065
rect 5356 15920 5408 15972
rect 7932 15920 7984 15972
rect 10692 15963 10744 15972
rect 10692 15929 10701 15963
rect 10701 15929 10735 15963
rect 10735 15929 10744 15963
rect 10692 15920 10744 15929
rect 3884 15895 3936 15904
rect 3884 15861 3893 15895
rect 3893 15861 3927 15895
rect 3927 15861 3936 15895
rect 3884 15852 3936 15861
rect 4620 15852 4672 15904
rect 4988 15852 5040 15904
rect 15200 15988 15252 16040
rect 18420 16031 18472 16040
rect 18420 15997 18429 16031
rect 18429 15997 18463 16031
rect 18463 15997 18472 16031
rect 18420 15988 18472 15997
rect 18604 16031 18656 16040
rect 18604 15997 18613 16031
rect 18613 15997 18647 16031
rect 18647 15997 18656 16031
rect 18604 15988 18656 15997
rect 18972 16031 19024 16040
rect 12992 15963 13044 15972
rect 12992 15929 13001 15963
rect 13001 15929 13035 15963
rect 13035 15929 13044 15963
rect 12992 15920 13044 15929
rect 17224 15920 17276 15972
rect 18972 15997 18981 16031
rect 18981 15997 19015 16031
rect 19015 15997 19024 16031
rect 18972 15988 19024 15997
rect 21088 16031 21140 16040
rect 21088 15997 21097 16031
rect 21097 15997 21131 16031
rect 21131 15997 21140 16031
rect 21088 15988 21140 15997
rect 21548 16031 21600 16040
rect 21548 15997 21557 16031
rect 21557 15997 21591 16031
rect 21591 15997 21600 16031
rect 21548 15988 21600 15997
rect 19892 15920 19944 15972
rect 22192 15963 22244 15972
rect 22192 15929 22201 15963
rect 22201 15929 22235 15963
rect 22235 15929 22244 15963
rect 22192 15920 22244 15929
rect 13268 15852 13320 15904
rect 17868 15852 17920 15904
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 3700 15648 3752 15700
rect 3792 15623 3844 15632
rect 3792 15589 3801 15623
rect 3801 15589 3835 15623
rect 3835 15589 3844 15623
rect 3792 15580 3844 15589
rect 5448 15512 5500 15564
rect 10140 15648 10192 15700
rect 13820 15648 13872 15700
rect 14648 15648 14700 15700
rect 15108 15691 15160 15700
rect 15108 15657 15117 15691
rect 15117 15657 15151 15691
rect 15151 15657 15160 15691
rect 15108 15648 15160 15657
rect 16396 15648 16448 15700
rect 20996 15648 21048 15700
rect 7932 15623 7984 15632
rect 7932 15589 7941 15623
rect 7941 15589 7975 15623
rect 7975 15589 7984 15623
rect 7932 15580 7984 15589
rect 10416 15580 10468 15632
rect 10692 15580 10744 15632
rect 12808 15512 12860 15564
rect 2504 15444 2556 15496
rect 4528 15444 4580 15496
rect 8392 15487 8444 15496
rect 8392 15453 8401 15487
rect 8401 15453 8435 15487
rect 8435 15453 8444 15487
rect 8392 15444 8444 15453
rect 11336 15444 11388 15496
rect 12532 15444 12584 15496
rect 13544 15512 13596 15564
rect 16120 15555 16172 15564
rect 16120 15521 16129 15555
rect 16129 15521 16163 15555
rect 16163 15521 16172 15555
rect 16396 15555 16448 15564
rect 16120 15512 16172 15521
rect 16396 15521 16405 15555
rect 16405 15521 16439 15555
rect 16439 15521 16448 15555
rect 16396 15512 16448 15521
rect 16580 15555 16632 15564
rect 16580 15521 16589 15555
rect 16589 15521 16623 15555
rect 16623 15521 16632 15555
rect 16580 15512 16632 15521
rect 19432 15512 19484 15564
rect 19892 15512 19944 15564
rect 23572 15623 23624 15632
rect 23572 15589 23581 15623
rect 23581 15589 23615 15623
rect 23615 15589 23624 15623
rect 23572 15580 23624 15589
rect 22192 15555 22244 15564
rect 22192 15521 22201 15555
rect 22201 15521 22235 15555
rect 22235 15521 22244 15555
rect 22192 15512 22244 15521
rect 12992 15444 13044 15496
rect 13360 15487 13412 15496
rect 13360 15453 13369 15487
rect 13369 15453 13403 15487
rect 13403 15453 13412 15487
rect 13360 15444 13412 15453
rect 13636 15444 13688 15496
rect 11060 15419 11112 15428
rect 11060 15385 11069 15419
rect 11069 15385 11103 15419
rect 11103 15385 11112 15419
rect 11060 15376 11112 15385
rect 11152 15376 11204 15428
rect 5448 15308 5500 15360
rect 7104 15308 7156 15360
rect 13820 15308 13872 15360
rect 19432 15308 19484 15360
rect 21916 15308 21968 15360
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 7012 15104 7064 15156
rect 7564 15104 7616 15156
rect 8668 15104 8720 15156
rect 2504 15011 2556 15020
rect 2504 14977 2513 15011
rect 2513 14977 2547 15011
rect 2547 14977 2556 15011
rect 2504 14968 2556 14977
rect 5540 15036 5592 15088
rect 11244 15104 11296 15156
rect 20352 15104 20404 15156
rect 21916 15147 21968 15156
rect 21916 15113 21925 15147
rect 21925 15113 21959 15147
rect 21959 15113 21968 15147
rect 21916 15104 21968 15113
rect 13084 15036 13136 15088
rect 15752 15036 15804 15088
rect 4620 14968 4672 15020
rect 5448 14968 5500 15020
rect 4988 14900 5040 14952
rect 7932 14943 7984 14952
rect 7932 14909 7941 14943
rect 7941 14909 7975 14943
rect 7975 14909 7984 14943
rect 7932 14900 7984 14909
rect 11888 14968 11940 15020
rect 12624 14968 12676 15020
rect 13176 14968 13228 15020
rect 10416 14943 10468 14952
rect 10416 14909 10425 14943
rect 10425 14909 10459 14943
rect 10459 14909 10468 14943
rect 10416 14900 10468 14909
rect 11244 14900 11296 14952
rect 8392 14832 8444 14884
rect 13544 14943 13596 14952
rect 13544 14909 13553 14943
rect 13553 14909 13587 14943
rect 13587 14909 13596 14943
rect 13544 14900 13596 14909
rect 15200 14900 15252 14952
rect 15292 14900 15344 14952
rect 14924 14832 14976 14884
rect 15752 14900 15804 14952
rect 20996 14968 21048 15020
rect 20628 14943 20680 14952
rect 20628 14909 20637 14943
rect 20637 14909 20671 14943
rect 20671 14909 20680 14943
rect 20628 14900 20680 14909
rect 3884 14807 3936 14816
rect 3884 14773 3893 14807
rect 3893 14773 3927 14807
rect 3927 14773 3936 14807
rect 3884 14764 3936 14773
rect 4988 14807 5040 14816
rect 4988 14773 4997 14807
rect 4997 14773 5031 14807
rect 5031 14773 5040 14807
rect 4988 14764 5040 14773
rect 7104 14764 7156 14816
rect 10600 14764 10652 14816
rect 13912 14764 13964 14816
rect 14740 14764 14792 14816
rect 16120 14807 16172 14816
rect 16120 14773 16129 14807
rect 16129 14773 16163 14807
rect 16163 14773 16172 14807
rect 16120 14764 16172 14773
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 6736 14560 6788 14612
rect 7932 14560 7984 14612
rect 5356 14424 5408 14476
rect 15292 14560 15344 14612
rect 15752 14603 15804 14612
rect 15752 14569 15761 14603
rect 15761 14569 15795 14603
rect 15795 14569 15804 14603
rect 15752 14560 15804 14569
rect 10600 14535 10652 14544
rect 10600 14501 10609 14535
rect 10609 14501 10643 14535
rect 10643 14501 10652 14535
rect 10600 14492 10652 14501
rect 13360 14492 13412 14544
rect 16488 14560 16540 14612
rect 17776 14560 17828 14612
rect 5356 14263 5408 14272
rect 5356 14229 5365 14263
rect 5365 14229 5399 14263
rect 5399 14229 5408 14263
rect 5356 14220 5408 14229
rect 8668 14263 8720 14272
rect 8668 14229 8677 14263
rect 8677 14229 8711 14263
rect 8711 14229 8720 14263
rect 8668 14220 8720 14229
rect 11152 14424 11204 14476
rect 12532 14467 12584 14476
rect 12532 14433 12541 14467
rect 12541 14433 12575 14467
rect 12575 14433 12584 14467
rect 12532 14424 12584 14433
rect 20628 14492 20680 14544
rect 15200 14424 15252 14476
rect 16120 14467 16172 14476
rect 13636 14356 13688 14408
rect 15752 14356 15804 14408
rect 16120 14433 16129 14467
rect 16129 14433 16163 14467
rect 16163 14433 16172 14467
rect 16120 14424 16172 14433
rect 19432 14424 19484 14476
rect 23480 14424 23532 14476
rect 10324 14288 10376 14340
rect 9588 14220 9640 14272
rect 15476 14220 15528 14272
rect 18788 14220 18840 14272
rect 21824 14220 21876 14272
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 4712 14016 4764 14068
rect 5448 14016 5500 14068
rect 9588 14059 9640 14068
rect 9588 14025 9597 14059
rect 9597 14025 9631 14059
rect 9631 14025 9640 14059
rect 9588 14016 9640 14025
rect 10876 14016 10928 14068
rect 10968 14016 11020 14068
rect 13084 14016 13136 14068
rect 14924 14016 14976 14068
rect 10600 13948 10652 14000
rect 15200 13948 15252 14000
rect 6092 13923 6144 13932
rect 4528 13812 4580 13864
rect 6092 13889 6101 13923
rect 6101 13889 6135 13923
rect 6135 13889 6144 13923
rect 6092 13880 6144 13889
rect 13268 13880 13320 13932
rect 15476 13923 15528 13932
rect 8300 13855 8352 13864
rect 8300 13821 8309 13855
rect 8309 13821 8343 13855
rect 8343 13821 8352 13855
rect 8300 13812 8352 13821
rect 9680 13812 9732 13864
rect 12164 13812 12216 13864
rect 15476 13889 15485 13923
rect 15485 13889 15519 13923
rect 15519 13889 15528 13923
rect 15476 13880 15528 13889
rect 5540 13744 5592 13796
rect 6644 13744 6696 13796
rect 18328 13948 18380 14000
rect 15752 13812 15804 13864
rect 18236 13812 18288 13864
rect 19156 14016 19208 14068
rect 19340 14016 19392 14068
rect 20720 14059 20772 14068
rect 20720 14025 20729 14059
rect 20729 14025 20763 14059
rect 20763 14025 20772 14059
rect 20720 14016 20772 14025
rect 20812 13812 20864 13864
rect 21824 13855 21876 13864
rect 16672 13787 16724 13796
rect 16672 13753 16681 13787
rect 16681 13753 16715 13787
rect 16715 13753 16724 13787
rect 16672 13744 16724 13753
rect 21824 13821 21833 13855
rect 21833 13821 21867 13855
rect 21867 13821 21876 13855
rect 21824 13812 21876 13821
rect 22192 13787 22244 13796
rect 22192 13753 22201 13787
rect 22201 13753 22235 13787
rect 22235 13753 22244 13787
rect 22192 13744 22244 13753
rect 3884 13719 3936 13728
rect 3884 13685 3893 13719
rect 3893 13685 3927 13719
rect 3927 13685 3936 13719
rect 3884 13676 3936 13685
rect 5816 13719 5868 13728
rect 5816 13685 5825 13719
rect 5825 13685 5859 13719
rect 5859 13685 5868 13719
rect 5816 13676 5868 13685
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 6092 13515 6144 13524
rect 6092 13481 6101 13515
rect 6101 13481 6135 13515
rect 6135 13481 6144 13515
rect 6092 13472 6144 13481
rect 7288 13515 7340 13524
rect 7288 13481 7297 13515
rect 7297 13481 7331 13515
rect 7331 13481 7340 13515
rect 7288 13472 7340 13481
rect 7840 13472 7892 13524
rect 8300 13472 8352 13524
rect 4068 13336 4120 13388
rect 12716 13472 12768 13524
rect 4528 13311 4580 13320
rect 4528 13277 4537 13311
rect 4537 13277 4571 13311
rect 4571 13277 4580 13311
rect 4528 13268 4580 13277
rect 5724 13268 5776 13320
rect 7288 13268 7340 13320
rect 7472 13268 7524 13320
rect 8668 13336 8720 13388
rect 9680 13379 9732 13388
rect 9680 13345 9689 13379
rect 9689 13345 9723 13379
rect 9723 13345 9732 13379
rect 9680 13336 9732 13345
rect 11704 13379 11756 13388
rect 11704 13345 11713 13379
rect 11713 13345 11747 13379
rect 11747 13345 11756 13379
rect 11704 13336 11756 13345
rect 14004 13336 14056 13388
rect 15108 13472 15160 13524
rect 21732 13515 21784 13524
rect 21732 13481 21741 13515
rect 21741 13481 21775 13515
rect 21775 13481 21784 13515
rect 21732 13472 21784 13481
rect 23480 13515 23532 13524
rect 23480 13481 23489 13515
rect 23489 13481 23523 13515
rect 23523 13481 23532 13515
rect 23480 13472 23532 13481
rect 18236 13447 18288 13456
rect 18236 13413 18245 13447
rect 18245 13413 18279 13447
rect 18279 13413 18288 13447
rect 18236 13404 18288 13413
rect 14924 13379 14976 13388
rect 14924 13345 14933 13379
rect 14933 13345 14967 13379
rect 14967 13345 14976 13379
rect 14924 13336 14976 13345
rect 16672 13336 16724 13388
rect 22008 13336 22060 13388
rect 22192 13379 22244 13388
rect 22192 13345 22201 13379
rect 22201 13345 22235 13379
rect 22235 13345 22244 13379
rect 22192 13336 22244 13345
rect 9864 13243 9916 13252
rect 9864 13209 9873 13243
rect 9873 13209 9907 13243
rect 9907 13209 9916 13243
rect 9864 13200 9916 13209
rect 12716 13175 12768 13184
rect 12716 13141 12725 13175
rect 12725 13141 12759 13175
rect 12759 13141 12768 13175
rect 12716 13132 12768 13141
rect 15384 13132 15436 13184
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 5540 12928 5592 12980
rect 5724 12971 5776 12980
rect 5724 12937 5733 12971
rect 5733 12937 5767 12971
rect 5767 12937 5776 12971
rect 5724 12928 5776 12937
rect 5264 12767 5316 12776
rect 5264 12733 5273 12767
rect 5273 12733 5307 12767
rect 5307 12733 5316 12767
rect 5264 12724 5316 12733
rect 5816 12724 5868 12776
rect 8392 12928 8444 12980
rect 8576 12928 8628 12980
rect 11704 12928 11756 12980
rect 20536 12971 20588 12980
rect 14004 12903 14056 12912
rect 14004 12869 14013 12903
rect 14013 12869 14047 12903
rect 14047 12869 14056 12903
rect 14004 12860 14056 12869
rect 12716 12835 12768 12844
rect 12716 12801 12725 12835
rect 12725 12801 12759 12835
rect 12759 12801 12768 12835
rect 12716 12792 12768 12801
rect 13084 12792 13136 12844
rect 20536 12937 20545 12971
rect 20545 12937 20579 12971
rect 20579 12937 20588 12971
rect 20536 12928 20588 12937
rect 9864 12724 9916 12776
rect 4896 12656 4948 12708
rect 7472 12656 7524 12708
rect 6920 12588 6972 12640
rect 12348 12588 12400 12640
rect 13452 12588 13504 12640
rect 15752 12767 15804 12776
rect 15752 12733 15761 12767
rect 15761 12733 15795 12767
rect 15795 12733 15804 12767
rect 15752 12724 15804 12733
rect 16580 12724 16632 12776
rect 20812 12767 20864 12776
rect 20812 12733 20821 12767
rect 20821 12733 20855 12767
rect 20855 12733 20864 12767
rect 20812 12724 20864 12733
rect 22284 12724 22336 12776
rect 16212 12631 16264 12640
rect 16212 12597 16221 12631
rect 16221 12597 16255 12631
rect 16255 12597 16264 12631
rect 16212 12588 16264 12597
rect 21824 12631 21876 12640
rect 21824 12597 21833 12631
rect 21833 12597 21867 12631
rect 21867 12597 21876 12631
rect 21824 12588 21876 12597
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 5264 12384 5316 12436
rect 8484 12427 8536 12436
rect 8484 12393 8493 12427
rect 8493 12393 8527 12427
rect 8527 12393 8536 12427
rect 8484 12384 8536 12393
rect 11980 12384 12032 12436
rect 17960 12384 18012 12436
rect 4896 12291 4948 12300
rect 4896 12257 4905 12291
rect 4905 12257 4939 12291
rect 4939 12257 4948 12291
rect 4896 12248 4948 12257
rect 5264 12248 5316 12300
rect 6736 12291 6788 12300
rect 6736 12257 6745 12291
rect 6745 12257 6779 12291
rect 6779 12257 6788 12291
rect 6736 12248 6788 12257
rect 6920 12291 6972 12300
rect 6920 12257 6929 12291
rect 6929 12257 6963 12291
rect 6963 12257 6972 12291
rect 6920 12248 6972 12257
rect 17316 12359 17368 12368
rect 17316 12325 17325 12359
rect 17325 12325 17359 12359
rect 17359 12325 17368 12359
rect 17316 12316 17368 12325
rect 16212 12248 16264 12300
rect 18328 12291 18380 12300
rect 18328 12257 18337 12291
rect 18337 12257 18371 12291
rect 18371 12257 18380 12291
rect 18328 12248 18380 12257
rect 21364 12248 21416 12300
rect 22008 12384 22060 12436
rect 23388 12316 23440 12368
rect 21824 12248 21876 12300
rect 5172 12180 5224 12232
rect 7472 12180 7524 12232
rect 12348 12180 12400 12232
rect 16120 12180 16172 12232
rect 5172 12044 5224 12096
rect 7288 12044 7340 12096
rect 8300 12087 8352 12096
rect 8300 12053 8309 12087
rect 8309 12053 8343 12087
rect 8343 12053 8352 12087
rect 8300 12044 8352 12053
rect 16396 12044 16448 12096
rect 19340 12044 19392 12096
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 7380 11840 7432 11892
rect 8392 11883 8444 11892
rect 8392 11849 8401 11883
rect 8401 11849 8435 11883
rect 8435 11849 8444 11883
rect 8392 11840 8444 11849
rect 16580 11883 16632 11892
rect 16580 11849 16589 11883
rect 16589 11849 16623 11883
rect 16623 11849 16632 11883
rect 16580 11840 16632 11849
rect 4620 11772 4672 11824
rect 2504 11679 2556 11688
rect 2504 11645 2513 11679
rect 2513 11645 2547 11679
rect 2547 11645 2556 11679
rect 7288 11747 7340 11756
rect 7288 11713 7297 11747
rect 7297 11713 7331 11747
rect 7331 11713 7340 11747
rect 7288 11704 7340 11713
rect 2504 11636 2556 11645
rect 7104 11636 7156 11688
rect 8852 11636 8904 11688
rect 17316 11840 17368 11892
rect 19892 11840 19944 11892
rect 21364 11883 21416 11892
rect 21364 11849 21373 11883
rect 21373 11849 21407 11883
rect 21407 11849 21416 11883
rect 21364 11840 21416 11849
rect 22284 11883 22336 11892
rect 22284 11849 22293 11883
rect 22293 11849 22327 11883
rect 22327 11849 22336 11883
rect 22284 11840 22336 11849
rect 20812 11704 20864 11756
rect 23388 11636 23440 11688
rect 3884 11543 3936 11552
rect 3884 11509 3893 11543
rect 3893 11509 3927 11543
rect 3927 11509 3936 11543
rect 3884 11500 3936 11509
rect 20904 11543 20956 11552
rect 20904 11509 20913 11543
rect 20913 11509 20947 11543
rect 20947 11509 20956 11543
rect 20904 11500 20956 11509
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 8484 11339 8536 11348
rect 8484 11305 8493 11339
rect 8493 11305 8527 11339
rect 8527 11305 8536 11339
rect 8484 11296 8536 11305
rect 8852 11339 8904 11348
rect 8852 11305 8861 11339
rect 8861 11305 8895 11339
rect 8895 11305 8904 11339
rect 8852 11296 8904 11305
rect 7104 11203 7156 11212
rect 7104 11169 7113 11203
rect 7113 11169 7147 11203
rect 7147 11169 7156 11203
rect 7104 11160 7156 11169
rect 12900 11160 12952 11212
rect 14004 11160 14056 11212
rect 16396 11203 16448 11212
rect 16396 11169 16405 11203
rect 16405 11169 16439 11203
rect 16439 11169 16448 11203
rect 16396 11160 16448 11169
rect 7380 11135 7432 11144
rect 7380 11101 7389 11135
rect 7389 11101 7423 11135
rect 7423 11101 7432 11135
rect 7380 11092 7432 11101
rect 12716 11135 12768 11144
rect 12716 11101 12725 11135
rect 12725 11101 12759 11135
rect 12759 11101 12768 11135
rect 12716 11092 12768 11101
rect 13820 11092 13872 11144
rect 19432 11296 19484 11348
rect 24216 11296 24268 11348
rect 19340 11160 19392 11212
rect 13728 11024 13780 11076
rect 16212 11067 16264 11076
rect 16212 11033 16221 11067
rect 16221 11033 16255 11067
rect 16255 11033 16264 11067
rect 16212 11024 16264 11033
rect 12808 10956 12860 11008
rect 16580 10956 16632 11008
rect 19892 11024 19944 11076
rect 18328 10956 18380 11008
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 4620 10752 4672 10804
rect 7380 10752 7432 10804
rect 8116 10752 8168 10804
rect 12808 10752 12860 10804
rect 12900 10752 12952 10804
rect 14004 10752 14056 10804
rect 19892 10752 19944 10804
rect 2504 10659 2556 10668
rect 2504 10625 2513 10659
rect 2513 10625 2547 10659
rect 2547 10625 2556 10659
rect 2504 10616 2556 10625
rect 6736 10616 6788 10668
rect 2780 10591 2832 10600
rect 2780 10557 2789 10591
rect 2789 10557 2823 10591
rect 2823 10557 2832 10591
rect 2780 10548 2832 10557
rect 6552 10548 6604 10600
rect 6828 10591 6880 10600
rect 6828 10557 6837 10591
rect 6837 10557 6871 10591
rect 6871 10557 6880 10591
rect 6828 10548 6880 10557
rect 8024 10616 8076 10668
rect 12164 10616 12216 10668
rect 12716 10659 12768 10668
rect 12716 10625 12725 10659
rect 12725 10625 12759 10659
rect 12759 10625 12768 10659
rect 12716 10616 12768 10625
rect 15384 10684 15436 10736
rect 16580 10684 16632 10736
rect 17776 10684 17828 10736
rect 18328 10659 18380 10668
rect 8300 10548 8352 10600
rect 18328 10625 18337 10659
rect 18337 10625 18371 10659
rect 18371 10625 18380 10659
rect 18328 10616 18380 10625
rect 20536 10659 20588 10668
rect 20536 10625 20545 10659
rect 20545 10625 20579 10659
rect 20579 10625 20588 10659
rect 20536 10616 20588 10625
rect 20904 10616 20956 10668
rect 3884 10455 3936 10464
rect 3884 10421 3893 10455
rect 3893 10421 3927 10455
rect 3927 10421 3936 10455
rect 3884 10412 3936 10421
rect 6552 10455 6604 10464
rect 6552 10421 6561 10455
rect 6561 10421 6595 10455
rect 6595 10421 6604 10455
rect 6552 10412 6604 10421
rect 16212 10412 16264 10464
rect 21456 10412 21508 10464
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 13636 10208 13688 10260
rect 20536 10208 20588 10260
rect 2780 10140 2832 10192
rect 7012 10072 7064 10124
rect 13544 10072 13596 10124
rect 13912 10072 13964 10124
rect 21456 10072 21508 10124
rect 12256 10047 12308 10056
rect 12256 10013 12265 10047
rect 12265 10013 12299 10047
rect 12299 10013 12308 10047
rect 12256 10004 12308 10013
rect 12532 10047 12584 10056
rect 12532 10013 12541 10047
rect 12541 10013 12575 10047
rect 12575 10013 12584 10047
rect 12532 10004 12584 10013
rect 7748 9936 7800 9988
rect 13912 9936 13964 9988
rect 7012 9911 7064 9920
rect 7012 9877 7021 9911
rect 7021 9877 7055 9911
rect 7055 9877 7064 9911
rect 7012 9868 7064 9877
rect 14004 9911 14056 9920
rect 14004 9877 14013 9911
rect 14013 9877 14047 9911
rect 14047 9877 14056 9911
rect 14004 9868 14056 9877
rect 16212 9868 16264 9920
rect 22468 9911 22520 9920
rect 22468 9877 22477 9911
rect 22477 9877 22511 9911
rect 22511 9877 22520 9911
rect 22468 9868 22520 9877
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 20536 9664 20588 9716
rect 7748 9639 7800 9648
rect 7748 9605 7757 9639
rect 7757 9605 7791 9639
rect 7791 9605 7800 9639
rect 7748 9596 7800 9605
rect 2780 9571 2832 9580
rect 2780 9537 2789 9571
rect 2789 9537 2823 9571
rect 2823 9537 2832 9571
rect 12348 9596 12400 9648
rect 14004 9596 14056 9648
rect 2780 9528 2832 9537
rect 2504 9503 2556 9512
rect 2504 9469 2513 9503
rect 2513 9469 2547 9503
rect 2547 9469 2556 9503
rect 12532 9528 12584 9580
rect 13820 9571 13872 9580
rect 13820 9537 13829 9571
rect 13829 9537 13863 9571
rect 13863 9537 13872 9571
rect 13820 9528 13872 9537
rect 2504 9460 2556 9469
rect 2780 9324 2832 9376
rect 9404 9503 9456 9512
rect 7932 9435 7984 9444
rect 7932 9401 7941 9435
rect 7941 9401 7975 9435
rect 7975 9401 7984 9435
rect 7932 9392 7984 9401
rect 3884 9367 3936 9376
rect 3884 9333 3893 9367
rect 3893 9333 3927 9367
rect 3927 9333 3936 9367
rect 3884 9324 3936 9333
rect 9404 9469 9413 9503
rect 9413 9469 9447 9503
rect 9447 9469 9456 9503
rect 9404 9460 9456 9469
rect 10140 9460 10192 9512
rect 8116 9392 8168 9444
rect 11980 9324 12032 9376
rect 13636 9460 13688 9512
rect 13728 9324 13780 9376
rect 15292 9324 15344 9376
rect 20076 9460 20128 9512
rect 20536 9324 20588 9376
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 7932 9120 7984 9172
rect 14096 9163 14148 9172
rect 14096 9129 14105 9163
rect 14105 9129 14139 9163
rect 14139 9129 14148 9163
rect 14096 9120 14148 9129
rect 19432 9163 19484 9172
rect 19432 9129 19441 9163
rect 19441 9129 19475 9163
rect 19475 9129 19484 9163
rect 19432 9120 19484 9129
rect 20536 9120 20588 9172
rect 7840 9052 7892 9104
rect 7748 9027 7800 9036
rect 7748 8993 7757 9027
rect 7757 8993 7791 9027
rect 7791 8993 7800 9027
rect 7748 8984 7800 8993
rect 12072 9052 12124 9104
rect 13820 9052 13872 9104
rect 9680 9027 9732 9036
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 8300 8916 8352 8968
rect 8392 8916 8444 8968
rect 14004 8984 14056 9036
rect 15292 9027 15344 9036
rect 15292 8993 15301 9027
rect 15301 8993 15335 9027
rect 15335 8993 15344 9027
rect 15292 8984 15344 8993
rect 10968 8916 11020 8968
rect 12348 8916 12400 8968
rect 12992 8959 13044 8968
rect 12992 8925 13001 8959
rect 13001 8925 13035 8959
rect 13035 8925 13044 8959
rect 12992 8916 13044 8925
rect 4068 8848 4120 8900
rect 12624 8848 12676 8900
rect 22468 8984 22520 9036
rect 2780 8780 2832 8832
rect 8208 8823 8260 8832
rect 8208 8789 8217 8823
rect 8217 8789 8251 8823
rect 8251 8789 8260 8823
rect 8208 8780 8260 8789
rect 19340 8780 19392 8832
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 8392 8619 8444 8628
rect 8392 8585 8401 8619
rect 8401 8585 8435 8619
rect 8435 8585 8444 8619
rect 8392 8576 8444 8585
rect 10140 8619 10192 8628
rect 10140 8585 10149 8619
rect 10149 8585 10183 8619
rect 10183 8585 10192 8619
rect 10140 8576 10192 8585
rect 20076 8619 20128 8628
rect 16212 8508 16264 8560
rect 20076 8585 20085 8619
rect 20085 8585 20119 8619
rect 20119 8585 20128 8619
rect 20076 8576 20128 8585
rect 20536 8619 20588 8628
rect 20536 8585 20545 8619
rect 20545 8585 20579 8619
rect 20579 8585 20588 8619
rect 20536 8576 20588 8585
rect 20720 8508 20772 8560
rect 8208 8440 8260 8492
rect 12992 8440 13044 8492
rect 13820 8440 13872 8492
rect 6828 8415 6880 8424
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 7104 8415 7156 8424
rect 7104 8381 7113 8415
rect 7113 8381 7147 8415
rect 7147 8381 7156 8415
rect 7104 8372 7156 8381
rect 9772 8372 9824 8424
rect 10140 8372 10192 8424
rect 14004 8415 14056 8424
rect 14004 8381 14013 8415
rect 14013 8381 14047 8415
rect 14047 8381 14056 8415
rect 14004 8372 14056 8381
rect 14096 8372 14148 8424
rect 4620 8304 4672 8356
rect 5448 8304 5500 8356
rect 22284 8440 22336 8492
rect 19340 8372 19392 8424
rect 3884 8279 3936 8288
rect 3884 8245 3893 8279
rect 3893 8245 3927 8279
rect 3927 8245 3936 8279
rect 3884 8236 3936 8245
rect 4068 8236 4120 8288
rect 6552 8236 6604 8288
rect 6828 8236 6880 8288
rect 8208 8236 8260 8288
rect 9864 8279 9916 8288
rect 9864 8245 9873 8279
rect 9873 8245 9907 8279
rect 9907 8245 9916 8279
rect 9864 8236 9916 8245
rect 12900 8236 12952 8288
rect 13912 8236 13964 8288
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 8300 8032 8352 8084
rect 7104 7964 7156 8016
rect 9680 8007 9732 8016
rect 7104 7828 7156 7880
rect 8484 7939 8536 7948
rect 8484 7905 8493 7939
rect 8493 7905 8527 7939
rect 8527 7905 8536 7939
rect 9680 7973 9689 8007
rect 9689 7973 9723 8007
rect 9723 7973 9732 8007
rect 9680 7964 9732 7973
rect 8484 7896 8536 7905
rect 9772 7896 9824 7948
rect 8576 7828 8628 7880
rect 12164 7896 12216 7948
rect 17868 8032 17920 8084
rect 15476 7939 15528 7948
rect 15476 7905 15485 7939
rect 15485 7905 15519 7939
rect 15519 7905 15528 7939
rect 15476 7896 15528 7905
rect 15568 7939 15620 7948
rect 15568 7905 15577 7939
rect 15577 7905 15611 7939
rect 15611 7905 15620 7939
rect 15568 7896 15620 7905
rect 12900 7828 12952 7880
rect 9036 7760 9088 7812
rect 9680 7760 9732 7812
rect 7012 7692 7064 7744
rect 13636 7735 13688 7744
rect 13636 7701 13645 7735
rect 13645 7701 13679 7735
rect 13679 7701 13688 7735
rect 13636 7692 13688 7701
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 8576 7531 8628 7540
rect 8576 7497 8585 7531
rect 8585 7497 8619 7531
rect 8619 7497 8628 7531
rect 8576 7488 8628 7497
rect 14372 7488 14424 7540
rect 15108 7488 15160 7540
rect 15384 7488 15436 7540
rect 20720 7531 20772 7540
rect 20720 7497 20729 7531
rect 20729 7497 20763 7531
rect 20763 7497 20772 7531
rect 20720 7488 20772 7497
rect 22284 7531 22336 7540
rect 22284 7497 22293 7531
rect 22293 7497 22327 7531
rect 22327 7497 22336 7531
rect 22284 7488 22336 7497
rect 9772 7352 9824 7404
rect 12808 7352 12860 7404
rect 19340 7395 19392 7404
rect 19340 7361 19349 7395
rect 19349 7361 19383 7395
rect 19383 7361 19392 7395
rect 19340 7352 19392 7361
rect 2504 7327 2556 7336
rect 2504 7293 2513 7327
rect 2513 7293 2547 7327
rect 2547 7293 2556 7327
rect 2504 7284 2556 7293
rect 6828 7284 6880 7336
rect 7288 7327 7340 7336
rect 7288 7293 7297 7327
rect 7297 7293 7331 7327
rect 7331 7293 7340 7327
rect 7288 7284 7340 7293
rect 15292 7284 15344 7336
rect 22284 7284 22336 7336
rect 3884 7191 3936 7200
rect 3884 7157 3893 7191
rect 3893 7157 3927 7191
rect 3927 7157 3936 7191
rect 3884 7148 3936 7157
rect 4620 7148 4672 7200
rect 8208 7148 8260 7200
rect 10968 7148 11020 7200
rect 19984 7191 20036 7200
rect 19984 7157 19993 7191
rect 19993 7157 20027 7191
rect 20027 7157 20036 7191
rect 19984 7148 20036 7157
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 15108 6987 15160 6996
rect 15108 6953 15117 6987
rect 15117 6953 15151 6987
rect 15151 6953 15160 6987
rect 20720 6987 20772 6996
rect 15108 6944 15160 6953
rect 7104 6919 7156 6928
rect 7104 6885 7113 6919
rect 7113 6885 7147 6919
rect 7147 6885 7156 6919
rect 7104 6876 7156 6885
rect 15292 6919 15344 6928
rect 15292 6885 15301 6919
rect 15301 6885 15335 6919
rect 15335 6885 15344 6919
rect 15292 6876 15344 6885
rect 4068 6808 4120 6860
rect 5172 6808 5224 6860
rect 10968 6808 11020 6860
rect 12992 6808 13044 6860
rect 13912 6808 13964 6860
rect 5448 6783 5500 6792
rect 5448 6749 5457 6783
rect 5457 6749 5491 6783
rect 5491 6749 5500 6783
rect 5448 6740 5500 6749
rect 5724 6783 5776 6792
rect 5724 6749 5733 6783
rect 5733 6749 5767 6783
rect 5767 6749 5776 6783
rect 5724 6740 5776 6749
rect 11428 6783 11480 6792
rect 11428 6749 11437 6783
rect 11437 6749 11471 6783
rect 11471 6749 11480 6783
rect 11428 6740 11480 6749
rect 12164 6740 12216 6792
rect 15476 6808 15528 6860
rect 20720 6953 20729 6987
rect 20729 6953 20763 6987
rect 20763 6953 20772 6987
rect 20720 6944 20772 6953
rect 22284 6987 22336 6996
rect 22284 6953 22293 6987
rect 22293 6953 22327 6987
rect 22327 6953 22336 6987
rect 22284 6944 22336 6953
rect 16304 6851 16356 6860
rect 16304 6817 16313 6851
rect 16313 6817 16347 6851
rect 16347 6817 16356 6851
rect 16304 6808 16356 6817
rect 19984 6808 20036 6860
rect 15660 6740 15712 6792
rect 16212 6783 16264 6792
rect 15108 6672 15160 6724
rect 16212 6749 16221 6783
rect 16221 6749 16255 6783
rect 16255 6749 16264 6783
rect 16212 6740 16264 6749
rect 20720 6740 20772 6792
rect 11336 6604 11388 6656
rect 12808 6604 12860 6656
rect 12992 6647 13044 6656
rect 12992 6613 13001 6647
rect 13001 6613 13035 6647
rect 13035 6613 13044 6647
rect 12992 6604 13044 6613
rect 19892 6647 19944 6656
rect 19892 6613 19901 6647
rect 19901 6613 19935 6647
rect 19935 6613 19944 6647
rect 19892 6604 19944 6613
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 2504 6239 2556 6248
rect 2504 6205 2513 6239
rect 2513 6205 2547 6239
rect 2547 6205 2556 6239
rect 2504 6196 2556 6205
rect 9680 6400 9732 6452
rect 16304 6400 16356 6452
rect 7288 6264 7340 6316
rect 9864 6264 9916 6316
rect 20720 6264 20772 6316
rect 8576 6196 8628 6248
rect 8852 6239 8904 6248
rect 8852 6205 8861 6239
rect 8861 6205 8895 6239
rect 8895 6205 8904 6239
rect 8852 6196 8904 6205
rect 9036 6239 9088 6248
rect 9036 6205 9045 6239
rect 9045 6205 9079 6239
rect 9079 6205 9088 6239
rect 9036 6196 9088 6205
rect 15108 6196 15160 6248
rect 15660 6196 15712 6248
rect 16212 6196 16264 6248
rect 20904 6196 20956 6248
rect 16856 6128 16908 6180
rect 3884 6103 3936 6112
rect 3884 6069 3893 6103
rect 3893 6069 3927 6103
rect 3927 6069 3936 6103
rect 3884 6060 3936 6069
rect 4068 6060 4120 6112
rect 4620 6060 4672 6112
rect 5908 6060 5960 6112
rect 15568 6060 15620 6112
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 5908 5899 5960 5908
rect 5908 5865 5917 5899
rect 5917 5865 5951 5899
rect 5951 5865 5960 5899
rect 5908 5856 5960 5865
rect 6828 5856 6880 5908
rect 15200 5856 15252 5908
rect 15384 5856 15436 5908
rect 15660 5856 15712 5908
rect 20720 5856 20772 5908
rect 21732 5899 21784 5908
rect 5724 5831 5776 5840
rect 5724 5797 5733 5831
rect 5733 5797 5767 5831
rect 5767 5797 5776 5831
rect 5724 5788 5776 5797
rect 11428 5788 11480 5840
rect 9864 5720 9916 5772
rect 14004 5788 14056 5840
rect 15108 5788 15160 5840
rect 12164 5763 12216 5772
rect 12164 5729 12173 5763
rect 12173 5729 12207 5763
rect 12207 5729 12216 5763
rect 12164 5720 12216 5729
rect 12532 5763 12584 5772
rect 12532 5729 12541 5763
rect 12541 5729 12575 5763
rect 12575 5729 12584 5763
rect 12532 5720 12584 5729
rect 15568 5763 15620 5772
rect 4068 5695 4120 5704
rect 4068 5661 4077 5695
rect 4077 5661 4111 5695
rect 4111 5661 4120 5695
rect 4068 5652 4120 5661
rect 5632 5652 5684 5704
rect 9036 5652 9088 5704
rect 15200 5652 15252 5704
rect 15568 5729 15577 5763
rect 15577 5729 15611 5763
rect 15611 5729 15620 5763
rect 15568 5720 15620 5729
rect 19892 5720 19944 5772
rect 16212 5652 16264 5704
rect 21364 5652 21416 5704
rect 21732 5865 21741 5899
rect 21741 5865 21775 5899
rect 21775 5865 21784 5899
rect 21732 5856 21784 5865
rect 19340 5516 19392 5568
rect 23480 5559 23532 5568
rect 23480 5525 23489 5559
rect 23489 5525 23523 5559
rect 23523 5525 23532 5559
rect 23480 5516 23532 5525
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 4068 5312 4120 5364
rect 5632 5355 5684 5364
rect 5632 5321 5641 5355
rect 5641 5321 5675 5355
rect 5675 5321 5684 5355
rect 5632 5312 5684 5321
rect 8852 5312 8904 5364
rect 15200 5312 15252 5364
rect 16856 5355 16908 5364
rect 2780 5219 2832 5228
rect 2780 5185 2789 5219
rect 2789 5185 2823 5219
rect 2823 5185 2832 5219
rect 2780 5176 2832 5185
rect 4068 5176 4120 5228
rect 5540 5176 5592 5228
rect 16856 5321 16865 5355
rect 16865 5321 16899 5355
rect 16899 5321 16908 5355
rect 16856 5312 16908 5321
rect 20904 5355 20956 5364
rect 20904 5321 20913 5355
rect 20913 5321 20947 5355
rect 20947 5321 20956 5355
rect 20904 5312 20956 5321
rect 21364 5355 21416 5364
rect 21364 5321 21373 5355
rect 21373 5321 21407 5355
rect 21407 5321 21416 5355
rect 21364 5312 21416 5321
rect 19892 5176 19944 5228
rect 2504 5151 2556 5160
rect 2504 5117 2513 5151
rect 2513 5117 2547 5151
rect 2547 5117 2556 5151
rect 2504 5108 2556 5117
rect 5816 5108 5868 5160
rect 6920 5151 6972 5160
rect 6920 5117 6929 5151
rect 6929 5117 6963 5151
rect 6963 5117 6972 5151
rect 6920 5108 6972 5117
rect 7196 5151 7248 5160
rect 7196 5117 7205 5151
rect 7205 5117 7239 5151
rect 7239 5117 7248 5151
rect 7196 5108 7248 5117
rect 16672 5108 16724 5160
rect 20720 5108 20772 5160
rect 3884 5015 3936 5024
rect 3884 4981 3893 5015
rect 3893 4981 3927 5015
rect 3927 4981 3936 5015
rect 3884 4972 3936 4981
rect 8760 5015 8812 5024
rect 8760 4981 8769 5015
rect 8769 4981 8803 5015
rect 8803 4981 8812 5015
rect 8760 4972 8812 4981
rect 10508 4972 10560 5024
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 6920 4768 6972 4820
rect 8760 4768 8812 4820
rect 16672 4811 16724 4820
rect 16672 4777 16681 4811
rect 16681 4777 16715 4811
rect 16715 4777 16724 4811
rect 16672 4768 16724 4777
rect 7196 4743 7248 4752
rect 7196 4709 7205 4743
rect 7205 4709 7239 4743
rect 7239 4709 7248 4743
rect 7196 4700 7248 4709
rect 12532 4700 12584 4752
rect 5264 4632 5316 4684
rect 5908 4632 5960 4684
rect 10508 4632 10560 4684
rect 5816 4607 5868 4616
rect 5816 4573 5825 4607
rect 5825 4573 5859 4607
rect 5859 4573 5868 4607
rect 5816 4564 5868 4573
rect 11060 4607 11112 4616
rect 11060 4573 11069 4607
rect 11069 4573 11103 4607
rect 11103 4573 11112 4607
rect 11060 4564 11112 4573
rect 19340 4632 19392 4684
rect 12992 4496 13044 4548
rect 13176 4428 13228 4480
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 3976 4224 4028 4276
rect 11060 4224 11112 4276
rect 2504 4131 2556 4140
rect 2504 4097 2513 4131
rect 2513 4097 2547 4131
rect 2547 4097 2556 4131
rect 2504 4088 2556 4097
rect 3976 4088 4028 4140
rect 13176 4088 13228 4140
rect 5816 4020 5868 4072
rect 11336 4063 11388 4072
rect 11336 4029 11345 4063
rect 11345 4029 11379 4063
rect 11379 4029 11388 4063
rect 11336 4020 11388 4029
rect 8116 3952 8168 4004
rect 3884 3927 3936 3936
rect 3884 3893 3893 3927
rect 3893 3893 3927 3927
rect 3927 3893 3936 3927
rect 3884 3884 3936 3893
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 4068 3680 4120 3732
rect 7104 3680 7156 3732
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 5264 3179 5316 3188
rect 5264 3145 5273 3179
rect 5273 3145 5307 3179
rect 5307 3145 5316 3179
rect 5264 3136 5316 3145
rect 10508 3179 10560 3188
rect 3976 3000 4028 3052
rect 10508 3145 10517 3179
rect 10517 3145 10551 3179
rect 10551 3145 10560 3179
rect 10508 3136 10560 3145
rect 10324 3000 10376 3052
rect 7564 2932 7616 2984
rect 2780 2796 2832 2848
rect 10048 2839 10100 2848
rect 10048 2805 10057 2839
rect 10057 2805 10091 2839
rect 10091 2805 10100 2839
rect 10048 2796 10100 2805
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 3516 2592 3568 2644
rect 10048 2592 10100 2644
rect 2872 2524 2924 2576
rect 4988 2524 5040 2576
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 52552 892 52604 944
rect 53380 892 53432 944
rect 2780 416 2832 468
rect 5356 416 5408 468
<< metal2 >>
rect 3606 45928 3662 45937
rect 3606 45863 3662 45872
rect 2778 44704 2834 44713
rect 2778 44639 2834 44648
rect 2792 43314 2820 44639
rect 3514 44160 3570 44169
rect 3514 44095 3570 44104
rect 2780 43308 2832 43314
rect 2780 43250 2832 43256
rect 3148 43308 3200 43314
rect 3148 43250 3200 43256
rect 2688 42764 2740 42770
rect 2688 42706 2740 42712
rect 2700 42634 2728 42706
rect 2688 42628 2740 42634
rect 2688 42570 2740 42576
rect 2780 42560 2832 42566
rect 2780 42502 2832 42508
rect 3056 42560 3108 42566
rect 3056 42502 3108 42508
rect 1490 40624 1546 40633
rect 1490 40559 1546 40568
rect 1504 40186 1532 40559
rect 1492 40180 1544 40186
rect 1492 40122 1544 40128
rect 2792 40050 2820 42502
rect 3068 42226 3096 42502
rect 3056 42220 3108 42226
rect 3056 42162 3108 42168
rect 3160 42106 3188 43250
rect 3528 42906 3556 44095
rect 3516 42900 3568 42906
rect 3516 42842 3568 42848
rect 3068 42078 3188 42106
rect 2964 41472 3016 41478
rect 2964 41414 3016 41420
rect 2872 40724 2924 40730
rect 2872 40666 2924 40672
rect 2780 40044 2832 40050
rect 2780 39986 2832 39992
rect 2780 39636 2832 39642
rect 2780 39578 2832 39584
rect 2792 38962 2820 39578
rect 2780 38956 2832 38962
rect 2780 38898 2832 38904
rect 2780 38548 2832 38554
rect 2780 38490 2832 38496
rect 2792 37874 2820 38490
rect 2780 37868 2832 37874
rect 2780 37810 2832 37816
rect 2504 36780 2556 36786
rect 2504 36722 2556 36728
rect 2516 34610 2544 36722
rect 2884 35698 2912 40666
rect 2976 40100 3004 41414
rect 3068 40168 3096 42078
rect 3068 40140 3556 40168
rect 2976 40072 3096 40100
rect 2964 39976 3016 39982
rect 2964 39918 3016 39924
rect 2872 35692 2924 35698
rect 2872 35634 2924 35640
rect 2504 34604 2556 34610
rect 2504 34546 2556 34552
rect 2412 32768 2464 32774
rect 2412 32710 2464 32716
rect 2424 31278 2452 32710
rect 2412 31272 2464 31278
rect 2412 31214 2464 31220
rect 2516 29578 2544 34546
rect 2872 32428 2924 32434
rect 2872 32370 2924 32376
rect 2688 31136 2740 31142
rect 2688 31078 2740 31084
rect 2700 30190 2728 31078
rect 2688 30184 2740 30190
rect 2688 30126 2740 30132
rect 2700 29714 2728 30126
rect 2688 29708 2740 29714
rect 2688 29650 2740 29656
rect 2504 29572 2556 29578
rect 2504 29514 2556 29520
rect 2516 28082 2544 29514
rect 2596 28960 2648 28966
rect 2596 28902 2648 28908
rect 2504 28076 2556 28082
rect 2504 28018 2556 28024
rect 2516 26994 2544 28018
rect 2608 28014 2636 28902
rect 2596 28008 2648 28014
rect 2596 27950 2648 27956
rect 2780 27124 2832 27130
rect 2780 27066 2832 27072
rect 2504 26988 2556 26994
rect 2504 26930 2556 26936
rect 2516 25838 2544 26930
rect 2504 25832 2556 25838
rect 2504 25774 2556 25780
rect 2504 24744 2556 24750
rect 2504 24686 2556 24692
rect 2516 23662 2544 24686
rect 2792 23730 2820 27066
rect 2884 24154 2912 32370
rect 2976 29889 3004 39918
rect 3068 31113 3096 40072
rect 3330 40080 3386 40089
rect 3330 40015 3386 40024
rect 3240 39908 3292 39914
rect 3240 39850 3292 39856
rect 3252 38978 3280 39850
rect 3160 38950 3280 38978
rect 3160 34610 3188 38950
rect 3238 38856 3294 38865
rect 3238 38791 3294 38800
rect 3252 36922 3280 38791
rect 3240 36916 3292 36922
rect 3240 36858 3292 36864
rect 3240 35488 3292 35494
rect 3240 35430 3292 35436
rect 3148 34604 3200 34610
rect 3148 34546 3200 34552
rect 3252 34105 3280 35430
rect 3238 34096 3294 34105
rect 3238 34031 3294 34040
rect 3344 33946 3372 40015
rect 3424 39976 3476 39982
rect 3424 39918 3476 39924
rect 3436 39098 3464 39918
rect 3424 39092 3476 39098
rect 3424 39034 3476 39040
rect 3424 37664 3476 37670
rect 3424 37606 3476 37612
rect 3436 35329 3464 37606
rect 3422 35320 3478 35329
rect 3422 35255 3478 35264
rect 3424 35012 3476 35018
rect 3424 34954 3476 34960
rect 3252 33918 3372 33946
rect 3148 31816 3200 31822
rect 3148 31758 3200 31764
rect 3054 31104 3110 31113
rect 3054 31039 3110 31048
rect 3056 30728 3108 30734
rect 3056 30670 3108 30676
rect 2962 29880 3018 29889
rect 2962 29815 3018 29824
rect 2964 29640 3016 29646
rect 2964 29582 3016 29588
rect 2976 25906 3004 29582
rect 3068 28937 3096 30670
rect 3054 28928 3110 28937
rect 3054 28863 3110 28872
rect 3160 28744 3188 31758
rect 3068 28716 3188 28744
rect 2964 25900 3016 25906
rect 2964 25842 3016 25848
rect 2884 24126 3004 24154
rect 2780 23724 2832 23730
rect 2780 23666 2832 23672
rect 2504 23656 2556 23662
rect 2504 23598 2556 23604
rect 2516 22574 2544 23598
rect 2504 22568 2556 22574
rect 2504 22510 2556 22516
rect 2516 21486 2544 22510
rect 2504 21480 2556 21486
rect 2504 21422 2556 21428
rect 2516 20466 2544 21422
rect 2504 20460 2556 20466
rect 2504 20402 2556 20408
rect 2872 16992 2924 16998
rect 2976 16969 3004 24126
rect 2872 16934 2924 16940
rect 2962 16960 3018 16969
rect 2884 16538 2912 16934
rect 2962 16895 3018 16904
rect 2884 16510 3004 16538
rect 2504 16040 2556 16046
rect 2504 15982 2556 15988
rect 2516 15502 2544 15982
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 2516 15026 2544 15438
rect 2504 15020 2556 15026
rect 2504 14962 2556 14968
rect 2504 11688 2556 11694
rect 2504 11630 2556 11636
rect 2516 10674 2544 11630
rect 2504 10668 2556 10674
rect 2504 10610 2556 10616
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2792 10198 2820 10542
rect 2780 10192 2832 10198
rect 2780 10134 2832 10140
rect 2780 9580 2832 9586
rect 2780 9522 2832 9528
rect 2504 9512 2556 9518
rect 2504 9454 2556 9460
rect 2516 7342 2544 9454
rect 2792 9382 2820 9522
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2504 7336 2556 7342
rect 2504 7278 2556 7284
rect 2516 6254 2544 7278
rect 2504 6248 2556 6254
rect 2504 6190 2556 6196
rect 2516 5166 2544 6190
rect 2792 5234 2820 8774
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 2504 5160 2556 5166
rect 2504 5102 2556 5108
rect 2516 4146 2544 5102
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2792 921 2820 2790
rect 2870 2680 2926 2689
rect 2870 2615 2926 2624
rect 2884 2582 2912 2615
rect 2872 2576 2924 2582
rect 2872 2518 2924 2524
rect 2976 1465 3004 16510
rect 3068 16046 3096 28716
rect 3252 25684 3280 33918
rect 3436 33810 3464 34954
rect 3344 33782 3464 33810
rect 3344 29850 3372 33782
rect 3424 33108 3476 33114
rect 3424 33050 3476 33056
rect 3436 31793 3464 33050
rect 3528 32978 3556 40140
rect 3620 35086 3648 45863
rect 53378 45440 53434 46240
rect 4066 45384 4122 45393
rect 4066 45319 4122 45328
rect 4080 44198 4108 45319
rect 4068 44192 4120 44198
rect 4068 44134 4120 44140
rect 19580 44092 19876 44112
rect 19636 44090 19660 44092
rect 19716 44090 19740 44092
rect 19796 44090 19820 44092
rect 19658 44038 19660 44090
rect 19722 44038 19734 44090
rect 19796 44038 19798 44090
rect 19636 44036 19660 44038
rect 19716 44036 19740 44038
rect 19796 44036 19820 44038
rect 19580 44016 19876 44036
rect 50300 44092 50596 44112
rect 50356 44090 50380 44092
rect 50436 44090 50460 44092
rect 50516 44090 50540 44092
rect 50378 44038 50380 44090
rect 50442 44038 50454 44090
rect 50516 44038 50518 44090
rect 50356 44036 50380 44038
rect 50436 44036 50460 44038
rect 50516 44036 50540 44038
rect 50300 44016 50596 44036
rect 17868 43920 17920 43926
rect 17868 43862 17920 43868
rect 45928 43920 45980 43926
rect 45928 43862 45980 43868
rect 15660 43784 15712 43790
rect 15660 43726 15712 43732
rect 4220 43548 4516 43568
rect 4276 43546 4300 43548
rect 4356 43546 4380 43548
rect 4436 43546 4460 43548
rect 4298 43494 4300 43546
rect 4362 43494 4374 43546
rect 4436 43494 4438 43546
rect 4276 43492 4300 43494
rect 4356 43492 4380 43494
rect 4436 43492 4460 43494
rect 4220 43472 4516 43492
rect 8576 43308 8628 43314
rect 8576 43250 8628 43256
rect 7840 43240 7892 43246
rect 7840 43182 7892 43188
rect 3884 43104 3936 43110
rect 3884 43046 3936 43052
rect 4804 43104 4856 43110
rect 4804 43046 4856 43052
rect 3700 42220 3752 42226
rect 3700 42162 3752 42168
rect 3712 39574 3740 42162
rect 3896 41177 3924 43046
rect 4068 42764 4120 42770
rect 4068 42706 4120 42712
rect 4080 42362 4108 42706
rect 4220 42460 4516 42480
rect 4276 42458 4300 42460
rect 4356 42458 4380 42460
rect 4436 42458 4460 42460
rect 4298 42406 4300 42458
rect 4362 42406 4374 42458
rect 4436 42406 4438 42458
rect 4276 42404 4300 42406
rect 4356 42404 4380 42406
rect 4436 42404 4460 42406
rect 4220 42384 4516 42404
rect 4068 42356 4120 42362
rect 4068 42298 4120 42304
rect 4816 42022 4844 43046
rect 7564 42900 7616 42906
rect 7564 42842 7616 42848
rect 6552 42560 6604 42566
rect 6552 42502 6604 42508
rect 6920 42560 6972 42566
rect 6920 42502 6972 42508
rect 4804 42016 4856 42022
rect 4804 41958 4856 41964
rect 4220 41372 4516 41392
rect 4276 41370 4300 41372
rect 4356 41370 4380 41372
rect 4436 41370 4460 41372
rect 4298 41318 4300 41370
rect 4362 41318 4374 41370
rect 4436 41318 4438 41370
rect 4276 41316 4300 41318
rect 4356 41316 4380 41318
rect 4436 41316 4460 41318
rect 4220 41296 4516 41316
rect 4816 41274 4844 41958
rect 5080 41540 5132 41546
rect 5080 41482 5132 41488
rect 4804 41268 4856 41274
rect 4804 41210 4856 41216
rect 3882 41168 3938 41177
rect 3882 41103 3938 41112
rect 3792 41064 3844 41070
rect 3792 41006 3844 41012
rect 3804 40118 3832 41006
rect 4816 40610 4844 41210
rect 4988 40724 5040 40730
rect 4988 40666 5040 40672
rect 4816 40582 4936 40610
rect 4804 40520 4856 40526
rect 4804 40462 4856 40468
rect 4220 40284 4516 40304
rect 4276 40282 4300 40284
rect 4356 40282 4380 40284
rect 4436 40282 4460 40284
rect 4298 40230 4300 40282
rect 4362 40230 4374 40282
rect 4436 40230 4438 40282
rect 4276 40228 4300 40230
rect 4356 40228 4380 40230
rect 4436 40228 4460 40230
rect 4220 40208 4516 40228
rect 3792 40112 3844 40118
rect 3792 40054 3844 40060
rect 4816 39982 4844 40462
rect 4804 39976 4856 39982
rect 4804 39918 4856 39924
rect 4816 39574 4844 39918
rect 3700 39568 3752 39574
rect 3700 39510 3752 39516
rect 3976 39568 4028 39574
rect 3976 39510 4028 39516
rect 4804 39568 4856 39574
rect 4804 39510 4856 39516
rect 3988 39409 4016 39510
rect 4620 39432 4672 39438
rect 3974 39400 4030 39409
rect 4620 39374 4672 39380
rect 3974 39335 4030 39344
rect 4220 39196 4516 39216
rect 4276 39194 4300 39196
rect 4356 39194 4380 39196
rect 4436 39194 4460 39196
rect 4298 39142 4300 39194
rect 4362 39142 4374 39194
rect 4436 39142 4438 39194
rect 4276 39140 4300 39142
rect 4356 39140 4380 39142
rect 4436 39140 4460 39142
rect 4220 39120 4516 39140
rect 3884 38752 3936 38758
rect 3884 38694 3936 38700
rect 3792 38276 3844 38282
rect 3792 38218 3844 38224
rect 3700 36848 3752 36854
rect 3700 36790 3752 36796
rect 3608 35080 3660 35086
rect 3608 35022 3660 35028
rect 3516 32972 3568 32978
rect 3516 32914 3568 32920
rect 3712 32842 3740 36790
rect 3804 35018 3832 38218
rect 3896 37641 3924 38694
rect 4068 38344 4120 38350
rect 4068 38286 4120 38292
rect 4080 38185 4108 38286
rect 4066 38176 4122 38185
rect 4066 38111 4122 38120
rect 4220 38108 4516 38128
rect 4276 38106 4300 38108
rect 4356 38106 4380 38108
rect 4436 38106 4460 38108
rect 4298 38054 4300 38106
rect 4362 38054 4374 38106
rect 4436 38054 4438 38106
rect 4276 38052 4300 38054
rect 4356 38052 4380 38054
rect 4436 38052 4460 38054
rect 4220 38032 4516 38052
rect 4252 37664 4304 37670
rect 3882 37632 3938 37641
rect 4252 37606 4304 37612
rect 3882 37567 3938 37576
rect 4264 37262 4292 37606
rect 4632 37330 4660 39374
rect 4816 39302 4844 39510
rect 4804 39296 4856 39302
rect 4804 39238 4856 39244
rect 4712 38752 4764 38758
rect 4712 38694 4764 38700
rect 4620 37324 4672 37330
rect 4620 37266 4672 37272
rect 4252 37256 4304 37262
rect 4252 37198 4304 37204
rect 4068 37120 4120 37126
rect 3974 37088 4030 37097
rect 4068 37062 4120 37068
rect 3974 37023 4030 37032
rect 3988 36650 4016 37023
rect 3976 36644 4028 36650
rect 3976 36586 4028 36592
rect 4080 36417 4108 37062
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 4620 36780 4672 36786
rect 4724 36768 4752 38694
rect 4816 38486 4844 39238
rect 4804 38480 4856 38486
rect 4804 38422 4856 38428
rect 4816 38010 4844 38422
rect 4804 38004 4856 38010
rect 4804 37946 4856 37952
rect 4804 37256 4856 37262
rect 4908 37244 4936 40582
rect 5000 39574 5028 40666
rect 4988 39568 5040 39574
rect 4988 39510 5040 39516
rect 5092 38554 5120 41482
rect 5632 40996 5684 41002
rect 5632 40938 5684 40944
rect 5644 40594 5672 40938
rect 5632 40588 5684 40594
rect 5632 40530 5684 40536
rect 5724 40384 5776 40390
rect 5724 40326 5776 40332
rect 6368 40384 6420 40390
rect 6368 40326 6420 40332
rect 5736 40118 5764 40326
rect 5724 40112 5776 40118
rect 5724 40054 5776 40060
rect 5908 39840 5960 39846
rect 5908 39782 5960 39788
rect 5724 39432 5776 39438
rect 5724 39374 5776 39380
rect 5080 38548 5132 38554
rect 5080 38490 5132 38496
rect 5448 37800 5500 37806
rect 5448 37742 5500 37748
rect 4856 37216 4936 37244
rect 4804 37198 4856 37204
rect 4672 36740 4752 36768
rect 4620 36722 4672 36728
rect 4632 36582 4660 36722
rect 4620 36576 4672 36582
rect 4620 36518 4672 36524
rect 4066 36408 4122 36417
rect 4066 36343 4122 36352
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4066 35864 4122 35873
rect 4220 35856 4516 35876
rect 4066 35799 4122 35808
rect 3976 35556 4028 35562
rect 3976 35498 4028 35504
rect 3884 35216 3936 35222
rect 3884 35158 3936 35164
rect 3792 35012 3844 35018
rect 3792 34954 3844 34960
rect 3896 34649 3924 35158
rect 3882 34640 3938 34649
rect 3882 34575 3938 34584
rect 3884 34400 3936 34406
rect 3884 34342 3936 34348
rect 3792 34128 3844 34134
rect 3792 34070 3844 34076
rect 3516 32836 3568 32842
rect 3516 32778 3568 32784
rect 3700 32836 3752 32842
rect 3700 32778 3752 32784
rect 3422 31784 3478 31793
rect 3422 31719 3478 31728
rect 3424 30932 3476 30938
rect 3424 30874 3476 30880
rect 3332 29844 3384 29850
rect 3332 29786 3384 29792
rect 3330 28928 3386 28937
rect 3330 28863 3386 28872
rect 3344 26772 3372 28863
rect 3436 27130 3464 30874
rect 3424 27124 3476 27130
rect 3424 27066 3476 27072
rect 3424 26784 3476 26790
rect 3344 26744 3424 26772
rect 3424 26726 3476 26732
rect 3528 26586 3556 32778
rect 3700 32496 3752 32502
rect 3700 32438 3752 32444
rect 3712 32366 3740 32438
rect 3700 32360 3752 32366
rect 3700 32302 3752 32308
rect 3804 31872 3832 34070
rect 3896 32881 3924 34342
rect 3882 32872 3938 32881
rect 3882 32807 3938 32816
rect 3884 32224 3936 32230
rect 3884 32166 3936 32172
rect 3712 31844 3832 31872
rect 3608 30048 3660 30054
rect 3608 29990 3660 29996
rect 3620 26994 3648 29990
rect 3608 26988 3660 26994
rect 3608 26930 3660 26936
rect 3608 26784 3660 26790
rect 3608 26726 3660 26732
rect 3332 26580 3384 26586
rect 3332 26522 3384 26528
rect 3516 26580 3568 26586
rect 3516 26522 3568 26528
rect 3160 25656 3280 25684
rect 3160 22778 3188 25656
rect 3240 24608 3292 24614
rect 3240 24550 3292 24556
rect 3252 23497 3280 24550
rect 3238 23488 3294 23497
rect 3238 23423 3294 23432
rect 3148 22772 3200 22778
rect 3148 22714 3200 22720
rect 3148 21344 3200 21350
rect 3148 21286 3200 21292
rect 3160 19825 3188 21286
rect 3344 20505 3372 26522
rect 3516 25356 3568 25362
rect 3516 25298 3568 25304
rect 3330 20496 3386 20505
rect 3528 20466 3556 25298
rect 3330 20431 3386 20440
rect 3516 20460 3568 20466
rect 3516 20402 3568 20408
rect 3146 19816 3202 19825
rect 3146 19751 3202 19760
rect 3330 19272 3386 19281
rect 3330 19207 3386 19216
rect 3344 18970 3372 19207
rect 3332 18964 3384 18970
rect 3332 18906 3384 18912
rect 3056 16040 3108 16046
rect 3056 15982 3108 15988
rect 3620 15745 3648 26726
rect 3712 18057 3740 31844
rect 3792 31748 3844 31754
rect 3792 31690 3844 31696
rect 3804 31278 3832 31690
rect 3792 31272 3844 31278
rect 3792 31214 3844 31220
rect 3792 31136 3844 31142
rect 3792 31078 3844 31084
rect 3698 18048 3754 18057
rect 3698 17983 3754 17992
rect 3698 16280 3754 16289
rect 3698 16215 3754 16224
rect 3606 15736 3662 15745
rect 3712 15706 3740 16215
rect 3606 15671 3662 15680
rect 3700 15700 3752 15706
rect 3700 15642 3752 15648
rect 3804 15638 3832 31078
rect 3896 30569 3924 32166
rect 3882 30560 3938 30569
rect 3882 30495 3938 30504
rect 3988 29034 4016 35498
rect 4080 34950 4108 35799
rect 4160 35624 4212 35630
rect 4160 35566 4212 35572
rect 4172 35494 4200 35566
rect 4160 35488 4212 35494
rect 4160 35430 4212 35436
rect 4068 34944 4120 34950
rect 4068 34886 4120 34892
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 4220 34768 4516 34788
rect 4632 34746 4660 36518
rect 4712 35488 4764 35494
rect 4816 35476 4844 37198
rect 5460 36718 5488 37742
rect 5448 36712 5500 36718
rect 5448 36654 5500 36660
rect 4896 36576 4948 36582
rect 4896 36518 4948 36524
rect 4764 35448 4844 35476
rect 4712 35430 4764 35436
rect 4620 34740 4672 34746
rect 4620 34682 4672 34688
rect 4068 34468 4120 34474
rect 4068 34410 4120 34416
rect 4080 33561 4108 34410
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 4066 33552 4122 33561
rect 4724 33538 4752 35430
rect 4804 34060 4856 34066
rect 4804 34002 4856 34008
rect 4816 33658 4844 34002
rect 4804 33652 4856 33658
rect 4804 33594 4856 33600
rect 4724 33510 4844 33538
rect 4066 33487 4122 33496
rect 4068 33448 4120 33454
rect 4068 33390 4120 33396
rect 4080 32774 4108 33390
rect 4620 32972 4672 32978
rect 4620 32914 4672 32920
rect 4068 32768 4120 32774
rect 4068 32710 4120 32716
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 4632 32502 4660 32914
rect 4816 32774 4844 33510
rect 4804 32768 4856 32774
rect 4804 32710 4856 32716
rect 4620 32496 4672 32502
rect 4620 32438 4672 32444
rect 4068 32360 4120 32366
rect 4068 32302 4120 32308
rect 4080 31890 4108 32302
rect 4816 32298 4844 32710
rect 4804 32292 4856 32298
rect 4804 32234 4856 32240
rect 4068 31884 4120 31890
rect 4068 31826 4120 31832
rect 4620 31748 4672 31754
rect 4620 31690 4672 31696
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 4632 31482 4660 31690
rect 4620 31476 4672 31482
rect 4620 31418 4672 31424
rect 4632 31278 4660 31418
rect 4620 31272 4672 31278
rect 4620 31214 4672 31220
rect 4804 31136 4856 31142
rect 4804 31078 4856 31084
rect 4068 30796 4120 30802
rect 4068 30738 4120 30744
rect 4080 30326 4108 30738
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 4068 30320 4120 30326
rect 4068 30262 4120 30268
rect 4712 30184 4764 30190
rect 4632 30132 4712 30138
rect 4632 30126 4764 30132
rect 4632 30110 4752 30126
rect 4068 29504 4120 29510
rect 4068 29446 4120 29452
rect 4080 29345 4108 29446
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4066 29336 4122 29345
rect 4220 29328 4516 29348
rect 4066 29271 4122 29280
rect 4632 29186 4660 30110
rect 4712 30048 4764 30054
rect 4712 29990 4764 29996
rect 4540 29158 4660 29186
rect 3976 29028 4028 29034
rect 3976 28970 4028 28976
rect 3884 28960 3936 28966
rect 3884 28902 3936 28908
rect 4068 28960 4120 28966
rect 4068 28902 4120 28908
rect 3896 28121 3924 28902
rect 4080 28801 4108 28902
rect 4066 28792 4122 28801
rect 3976 28756 4028 28762
rect 4066 28727 4122 28736
rect 3976 28698 4028 28704
rect 3882 28112 3938 28121
rect 3882 28047 3938 28056
rect 3884 27872 3936 27878
rect 3884 27814 3936 27820
rect 3896 27033 3924 27814
rect 3882 27024 3938 27033
rect 3882 26959 3938 26968
rect 3884 26784 3936 26790
rect 3884 26726 3936 26732
rect 3896 25809 3924 26726
rect 3882 25800 3938 25809
rect 3882 25735 3938 25744
rect 3884 25696 3936 25702
rect 3884 25638 3936 25644
rect 3896 24585 3924 25638
rect 3988 25362 4016 28698
rect 4540 28626 4568 29158
rect 4528 28620 4580 28626
rect 4528 28562 4580 28568
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 4620 27872 4672 27878
rect 4620 27814 4672 27820
rect 4066 27568 4122 27577
rect 4066 27503 4122 27512
rect 4080 27130 4108 27503
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 4068 27124 4120 27130
rect 4068 27066 4120 27072
rect 4632 27062 4660 27814
rect 4620 27056 4672 27062
rect 4620 26998 4672 27004
rect 4068 26988 4120 26994
rect 4068 26930 4120 26936
rect 4080 26353 4108 26930
rect 4066 26344 4122 26353
rect 4066 26279 4122 26288
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 4068 26036 4120 26042
rect 4068 25978 4120 25984
rect 3976 25356 4028 25362
rect 3976 25298 4028 25304
rect 4080 25265 4108 25978
rect 4632 25974 4660 26998
rect 4620 25968 4672 25974
rect 4620 25910 4672 25916
rect 4066 25256 4122 25265
rect 4066 25191 4122 25200
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 4068 24676 4120 24682
rect 4068 24618 4120 24624
rect 3882 24576 3938 24585
rect 3882 24511 3938 24520
rect 4080 24041 4108 24618
rect 4066 24032 4122 24041
rect 4066 23967 4122 23976
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4220 23888 4516 23908
rect 3884 23520 3936 23526
rect 3884 23462 3936 23468
rect 4620 23520 4672 23526
rect 4620 23462 4672 23468
rect 3896 22273 3924 23462
rect 4068 23316 4120 23322
rect 4068 23258 4120 23264
rect 4080 22817 4108 23258
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4066 22808 4122 22817
rect 4220 22800 4516 22820
rect 4632 22778 4660 23462
rect 4066 22743 4122 22752
rect 4620 22772 4672 22778
rect 4620 22714 4672 22720
rect 3882 22264 3938 22273
rect 4632 22234 4660 22714
rect 3882 22199 3938 22208
rect 4620 22228 4672 22234
rect 4620 22170 4672 22176
rect 4068 21888 4120 21894
rect 4068 21830 4120 21836
rect 4080 21049 4108 21830
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 4632 21622 4660 22170
rect 4724 22098 4752 29990
rect 4712 22092 4764 22098
rect 4712 22034 4764 22040
rect 4620 21616 4672 21622
rect 4620 21558 4672 21564
rect 4066 21040 4122 21049
rect 4066 20975 4122 20984
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 4632 20602 4660 21558
rect 4620 20596 4672 20602
rect 4620 20538 4672 20544
rect 3884 20256 3936 20262
rect 3884 20198 3936 20204
rect 3896 18737 3924 20198
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 3882 18728 3938 18737
rect 3882 18663 3938 18672
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 4252 18284 4304 18290
rect 4252 18226 4304 18232
rect 4264 18086 4292 18226
rect 3884 18080 3936 18086
rect 3884 18022 3936 18028
rect 4252 18080 4304 18086
rect 4252 18022 4304 18028
rect 3896 17513 3924 18022
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 3882 17504 3938 17513
rect 3882 17439 3938 17448
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 3884 17128 3936 17134
rect 3884 17070 3936 17076
rect 3896 16794 3924 17070
rect 4632 17066 4660 17682
rect 4620 17060 4672 17066
rect 4620 17002 4672 17008
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 4632 16726 4660 17002
rect 4620 16720 4672 16726
rect 4620 16662 4672 16668
rect 4816 16538 4844 31078
rect 4908 24818 4936 36518
rect 5080 36304 5132 36310
rect 5080 36246 5132 36252
rect 4988 31884 5040 31890
rect 4988 31826 5040 31832
rect 4896 24812 4948 24818
rect 4896 24754 4948 24760
rect 5000 18426 5028 31826
rect 5092 30938 5120 36246
rect 5172 35760 5224 35766
rect 5172 35702 5224 35708
rect 5080 30932 5132 30938
rect 5080 30874 5132 30880
rect 5184 21690 5212 35702
rect 5264 34400 5316 34406
rect 5264 34342 5316 34348
rect 5276 29646 5304 34342
rect 5460 34066 5488 36654
rect 5736 35630 5764 39374
rect 5540 35624 5592 35630
rect 5540 35566 5592 35572
rect 5724 35624 5776 35630
rect 5724 35566 5776 35572
rect 5552 35154 5580 35566
rect 5816 35284 5868 35290
rect 5816 35226 5868 35232
rect 5540 35148 5592 35154
rect 5540 35090 5592 35096
rect 5552 34474 5580 35090
rect 5540 34468 5592 34474
rect 5540 34410 5592 34416
rect 5552 34202 5580 34410
rect 5540 34196 5592 34202
rect 5540 34138 5592 34144
rect 5448 34060 5500 34066
rect 5448 34002 5500 34008
rect 5632 33448 5684 33454
rect 5632 33390 5684 33396
rect 5356 32496 5408 32502
rect 5356 32438 5408 32444
rect 5264 29640 5316 29646
rect 5264 29582 5316 29588
rect 5368 24154 5396 32438
rect 5448 32360 5500 32366
rect 5448 32302 5500 32308
rect 5460 32026 5488 32302
rect 5540 32224 5592 32230
rect 5540 32166 5592 32172
rect 5448 32020 5500 32026
rect 5448 31962 5500 31968
rect 5368 24126 5488 24154
rect 5264 23112 5316 23118
rect 5264 23054 5316 23060
rect 5172 21684 5224 21690
rect 5172 21626 5224 21632
rect 4988 18420 5040 18426
rect 4988 18362 5040 18368
rect 4988 18080 5040 18086
rect 4988 18022 5040 18028
rect 4896 16652 4948 16658
rect 4896 16594 4948 16600
rect 4724 16510 4844 16538
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 4620 15904 4672 15910
rect 4620 15846 4672 15852
rect 3792 15632 3844 15638
rect 3792 15574 3844 15580
rect 3896 15065 3924 15846
rect 4528 15496 4580 15502
rect 4632 15484 4660 15846
rect 4580 15456 4660 15484
rect 4528 15438 4580 15444
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 3882 15056 3938 15065
rect 4632 15026 4660 15456
rect 3882 14991 3938 15000
rect 4620 15020 4672 15026
rect 4620 14962 4672 14968
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 3896 13977 3924 14758
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 4724 14074 4752 16510
rect 4804 16448 4856 16454
rect 4804 16390 4856 16396
rect 4816 15978 4844 16390
rect 4804 15972 4856 15978
rect 4804 15914 4856 15920
rect 4908 15484 4936 16594
rect 5000 15910 5028 18022
rect 5276 17218 5304 23054
rect 5356 19848 5408 19854
rect 5356 19790 5408 19796
rect 5368 18902 5396 19790
rect 5356 18896 5408 18902
rect 5356 18838 5408 18844
rect 5184 17190 5304 17218
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 4908 15456 5028 15484
rect 5000 14958 5028 15456
rect 4988 14952 5040 14958
rect 4988 14894 5040 14900
rect 5000 14822 5028 14894
rect 4988 14816 5040 14822
rect 4988 14758 5040 14764
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 3882 13968 3938 13977
rect 3882 13903 3938 13912
rect 4528 13864 4580 13870
rect 4528 13806 4580 13812
rect 3884 13728 3936 13734
rect 3884 13670 3936 13676
rect 3896 12753 3924 13670
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 4080 13297 4108 13330
rect 4540 13326 4568 13806
rect 4528 13320 4580 13326
rect 4066 13288 4122 13297
rect 4580 13280 4660 13308
rect 4528 13262 4580 13268
rect 4066 13223 4122 13232
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 3882 12744 3938 12753
rect 3882 12679 3938 12688
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4632 11830 4660 13280
rect 4896 12708 4948 12714
rect 4896 12650 4948 12656
rect 4908 12306 4936 12650
rect 4896 12300 4948 12306
rect 4896 12242 4948 12248
rect 4620 11824 4672 11830
rect 4620 11766 4672 11772
rect 3884 11552 3936 11558
rect 3882 11520 3884 11529
rect 3936 11520 3938 11529
rect 3882 11455 3938 11464
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 4632 10810 4660 11766
rect 4620 10804 4672 10810
rect 4620 10746 4672 10752
rect 3884 10464 3936 10470
rect 3882 10432 3884 10441
rect 3936 10432 3938 10441
rect 3882 10367 3938 10376
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 3884 9376 3936 9382
rect 3884 9318 3936 9324
rect 3896 9217 3924 9318
rect 3882 9208 3938 9217
rect 3882 9143 3938 9152
rect 4068 8900 4120 8906
rect 4068 8842 4120 8848
rect 4080 8673 4108 8842
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4066 8664 4122 8673
rect 4220 8656 4516 8676
rect 4066 8599 4122 8608
rect 4632 8362 4660 10746
rect 4620 8356 4672 8362
rect 4620 8298 4672 8304
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 3896 7993 3924 8230
rect 3882 7984 3938 7993
rect 3882 7919 3938 7928
rect 4080 7449 4108 8230
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 4066 7440 4122 7449
rect 4066 7375 4122 7384
rect 3884 7200 3936 7206
rect 3884 7142 3936 7148
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 3896 6769 3924 7142
rect 4068 6860 4120 6866
rect 4068 6802 4120 6808
rect 3882 6760 3938 6769
rect 3882 6695 3938 6704
rect 4080 6225 4108 6802
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 4066 6216 4122 6225
rect 4066 6151 4122 6160
rect 4632 6118 4660 7142
rect 3884 6112 3936 6118
rect 3884 6054 3936 6060
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 3896 5681 3924 6054
rect 4080 5710 4108 6054
rect 4068 5704 4120 5710
rect 3882 5672 3938 5681
rect 4068 5646 4120 5652
rect 3882 5607 3938 5616
rect 4080 5370 4108 5646
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4068 5364 4120 5370
rect 3988 5324 4068 5352
rect 3884 5024 3936 5030
rect 3884 4966 3936 4972
rect 3896 4457 3924 4966
rect 3882 4448 3938 4457
rect 3882 4383 3938 4392
rect 3988 4282 4016 5324
rect 4068 5306 4120 5312
rect 4068 5228 4120 5234
rect 4068 5170 4120 5176
rect 4080 5001 4108 5170
rect 4066 4992 4122 5001
rect 4066 4927 4122 4936
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 3976 4276 4028 4282
rect 3976 4218 4028 4224
rect 3988 4146 4016 4218
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3896 3233 3924 3878
rect 3882 3224 3938 3233
rect 3882 3159 3938 3168
rect 3988 3058 4016 4082
rect 4066 3904 4122 3913
rect 4066 3839 4122 3848
rect 4080 3738 4108 3839
rect 4068 3732 4120 3738
rect 4068 3674 4120 3680
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3528 2145 3556 2586
rect 5000 2582 5028 14758
rect 5184 12238 5212 17190
rect 5368 17134 5396 18838
rect 5356 17128 5408 17134
rect 5356 17070 5408 17076
rect 5368 16794 5396 17070
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5368 16250 5396 16730
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 5356 15972 5408 15978
rect 5356 15914 5408 15920
rect 5368 14482 5396 15914
rect 5460 15570 5488 24126
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5460 15026 5488 15302
rect 5552 15094 5580 32166
rect 5644 31890 5672 33390
rect 5828 32434 5856 35226
rect 5920 34542 5948 39782
rect 6380 39370 6408 40326
rect 6368 39364 6420 39370
rect 6368 39306 6420 39312
rect 6564 39302 6592 42502
rect 6932 41614 6960 42502
rect 7472 41676 7524 41682
rect 7472 41618 7524 41624
rect 6920 41608 6972 41614
rect 6920 41550 6972 41556
rect 6932 41478 6960 41550
rect 6920 41472 6972 41478
rect 6920 41414 6972 41420
rect 7484 40934 7512 41618
rect 7472 40928 7524 40934
rect 7472 40870 7524 40876
rect 7484 40594 7512 40870
rect 7472 40588 7524 40594
rect 7472 40530 7524 40536
rect 7288 40384 7340 40390
rect 7288 40326 7340 40332
rect 6552 39296 6604 39302
rect 6552 39238 6604 39244
rect 6276 38820 6328 38826
rect 6276 38762 6328 38768
rect 6000 36100 6052 36106
rect 6000 36042 6052 36048
rect 5908 34536 5960 34542
rect 5908 34478 5960 34484
rect 5816 32428 5868 32434
rect 5816 32370 5868 32376
rect 5908 32428 5960 32434
rect 5908 32370 5960 32376
rect 5920 32337 5948 32370
rect 5906 32328 5962 32337
rect 5906 32263 5962 32272
rect 5632 31884 5684 31890
rect 5632 31826 5684 31832
rect 6012 30326 6040 36042
rect 6288 35154 6316 38762
rect 6552 37732 6604 37738
rect 6552 37674 6604 37680
rect 6276 35148 6328 35154
rect 6276 35090 6328 35096
rect 6276 34536 6328 34542
rect 6276 34478 6328 34484
rect 6092 34196 6144 34202
rect 6092 34138 6144 34144
rect 6104 32978 6132 34138
rect 6288 34066 6316 34478
rect 6564 34066 6592 37674
rect 7104 36712 7156 36718
rect 7104 36654 7156 36660
rect 7116 35630 7144 36654
rect 7104 35624 7156 35630
rect 7104 35566 7156 35572
rect 7116 35154 7144 35566
rect 7104 35148 7156 35154
rect 7104 35090 7156 35096
rect 7300 34542 7328 40326
rect 7472 39500 7524 39506
rect 7472 39442 7524 39448
rect 7380 39432 7432 39438
rect 7378 39400 7380 39409
rect 7432 39400 7434 39409
rect 7378 39335 7434 39344
rect 7484 38962 7512 39442
rect 7472 38956 7524 38962
rect 7472 38898 7524 38904
rect 7380 35284 7432 35290
rect 7380 35226 7432 35232
rect 7288 34536 7340 34542
rect 7288 34478 7340 34484
rect 6920 34400 6972 34406
rect 6920 34342 6972 34348
rect 6276 34060 6328 34066
rect 6276 34002 6328 34008
rect 6552 34060 6604 34066
rect 6552 34002 6604 34008
rect 6092 32972 6144 32978
rect 6092 32914 6144 32920
rect 6000 30320 6052 30326
rect 6000 30262 6052 30268
rect 6932 29102 6960 34342
rect 7012 33108 7064 33114
rect 7012 33050 7064 33056
rect 7024 30734 7052 33050
rect 7012 30728 7064 30734
rect 7012 30670 7064 30676
rect 7288 29504 7340 29510
rect 7288 29446 7340 29452
rect 6920 29096 6972 29102
rect 6920 29038 6972 29044
rect 6920 27940 6972 27946
rect 6920 27882 6972 27888
rect 6644 27328 6696 27334
rect 6644 27270 6696 27276
rect 6000 25288 6052 25294
rect 6000 25230 6052 25236
rect 6012 24410 6040 25230
rect 6000 24404 6052 24410
rect 6000 24346 6052 24352
rect 6092 24268 6144 24274
rect 6092 24210 6144 24216
rect 6104 24154 6132 24210
rect 6104 24126 6224 24154
rect 6656 24138 6684 27270
rect 6828 27056 6880 27062
rect 6828 26998 6880 27004
rect 6840 26926 6868 26998
rect 6828 26920 6880 26926
rect 6828 26862 6880 26868
rect 6736 26784 6788 26790
rect 6736 26726 6788 26732
rect 6748 26450 6776 26726
rect 6736 26444 6788 26450
rect 6736 26386 6788 26392
rect 6840 26382 6868 26862
rect 6932 26858 6960 27882
rect 7104 27396 7156 27402
rect 7104 27338 7156 27344
rect 7116 26994 7144 27338
rect 7104 26988 7156 26994
rect 7104 26930 7156 26936
rect 6920 26852 6972 26858
rect 6920 26794 6972 26800
rect 6828 26376 6880 26382
rect 6828 26318 6880 26324
rect 7104 24744 7156 24750
rect 7104 24686 7156 24692
rect 7012 24336 7064 24342
rect 7012 24278 7064 24284
rect 6196 23186 6224 24126
rect 6644 24132 6696 24138
rect 6644 24074 6696 24080
rect 6828 24132 6880 24138
rect 6828 24074 6880 24080
rect 6184 23180 6236 23186
rect 6184 23122 6236 23128
rect 6196 22982 6224 23122
rect 6184 22976 6236 22982
rect 6184 22918 6236 22924
rect 5632 22500 5684 22506
rect 5632 22442 5684 22448
rect 5644 21554 5672 22442
rect 6644 21888 6696 21894
rect 6644 21830 6696 21836
rect 6656 21622 6684 21830
rect 6644 21616 6696 21622
rect 6644 21558 6696 21564
rect 5632 21548 5684 21554
rect 5632 21490 5684 21496
rect 6184 21548 6236 21554
rect 6184 21490 6236 21496
rect 5724 21480 5776 21486
rect 5724 21422 5776 21428
rect 5632 18216 5684 18222
rect 5632 18158 5684 18164
rect 5644 16658 5672 18158
rect 5736 17202 5764 21422
rect 6196 20058 6224 21490
rect 6184 20052 6236 20058
rect 6184 19994 6236 20000
rect 6552 19916 6604 19922
rect 6552 19858 6604 19864
rect 5908 19168 5960 19174
rect 5908 19110 5960 19116
rect 5920 18834 5948 19110
rect 5908 18828 5960 18834
rect 5908 18770 5960 18776
rect 6000 18828 6052 18834
rect 6000 18770 6052 18776
rect 5920 17610 5948 18770
rect 6012 18426 6040 18770
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 6472 18358 6500 18702
rect 6460 18352 6512 18358
rect 6460 18294 6512 18300
rect 6564 17882 6592 19858
rect 6552 17876 6604 17882
rect 6552 17818 6604 17824
rect 6564 17746 6592 17818
rect 6552 17740 6604 17746
rect 6552 17682 6604 17688
rect 5908 17604 5960 17610
rect 5908 17546 5960 17552
rect 6564 17338 6592 17682
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 5816 17264 5868 17270
rect 5816 17206 5868 17212
rect 5724 17196 5776 17202
rect 5724 17138 5776 17144
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 5828 16590 5856 17206
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 5540 15088 5592 15094
rect 5540 15030 5592 15036
rect 5448 15020 5500 15026
rect 5448 14962 5500 14968
rect 5356 14476 5408 14482
rect 5356 14418 5408 14424
rect 5368 14278 5396 14418
rect 5356 14272 5408 14278
rect 5356 14214 5408 14220
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 5276 12442 5304 12718
rect 5264 12436 5316 12442
rect 5264 12378 5316 12384
rect 5276 12306 5304 12378
rect 5264 12300 5316 12306
rect 5264 12242 5316 12248
rect 5172 12232 5224 12238
rect 5172 12174 5224 12180
rect 5184 12102 5212 12174
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 5184 6866 5212 12038
rect 5172 6860 5224 6866
rect 5172 6802 5224 6808
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 5276 3194 5304 4626
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 4988 2576 5040 2582
rect 4988 2518 5040 2524
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 3514 2136 3570 2145
rect 4220 2128 4516 2148
rect 3514 2071 3570 2080
rect 2962 1456 3018 1465
rect 2962 1391 3018 1400
rect 2778 912 2834 921
rect 2778 847 2834 856
rect 5368 474 5396 14214
rect 5460 14074 5488 14962
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 6092 13932 6144 13938
rect 6092 13874 6144 13880
rect 5540 13796 5592 13802
rect 5540 13738 5592 13744
rect 5552 12986 5580 13738
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5736 12986 5764 13262
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5724 12980 5776 12986
rect 5724 12922 5776 12928
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5460 6798 5488 8298
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5552 5234 5580 12922
rect 5828 12782 5856 13670
rect 6104 13530 6132 13874
rect 6656 13802 6684 21558
rect 6736 21412 6788 21418
rect 6736 21354 6788 21360
rect 6748 18902 6776 21354
rect 6736 18896 6788 18902
rect 6736 18838 6788 18844
rect 6736 17740 6788 17746
rect 6736 17682 6788 17688
rect 6748 16658 6776 17682
rect 6736 16652 6788 16658
rect 6736 16594 6788 16600
rect 6748 14618 6776 16594
rect 6736 14612 6788 14618
rect 6736 14554 6788 14560
rect 6644 13796 6696 13802
rect 6644 13738 6696 13744
rect 6092 13524 6144 13530
rect 6092 13466 6144 13472
rect 5816 12776 5868 12782
rect 5816 12718 5868 12724
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6748 10674 6776 12242
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6840 10606 6868 24074
rect 6920 23520 6972 23526
rect 6920 23462 6972 23468
rect 6932 23186 6960 23462
rect 6920 23180 6972 23186
rect 6920 23122 6972 23128
rect 6932 20398 6960 23122
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 7024 19922 7052 24278
rect 7116 23254 7144 24686
rect 7104 23248 7156 23254
rect 7104 23190 7156 23196
rect 7300 23050 7328 29446
rect 7288 23044 7340 23050
rect 7288 22986 7340 22992
rect 7104 21140 7156 21146
rect 7104 21082 7156 21088
rect 7012 19916 7064 19922
rect 7012 19858 7064 19864
rect 7116 19281 7144 21082
rect 7288 21004 7340 21010
rect 7288 20946 7340 20952
rect 7196 20936 7248 20942
rect 7196 20878 7248 20884
rect 7208 19310 7236 20878
rect 7300 19854 7328 20946
rect 7288 19848 7340 19854
rect 7288 19790 7340 19796
rect 7196 19304 7248 19310
rect 7102 19272 7158 19281
rect 7012 19236 7064 19242
rect 7196 19246 7248 19252
rect 7102 19207 7104 19216
rect 7012 19178 7064 19184
rect 7156 19207 7158 19216
rect 7104 19178 7156 19184
rect 7024 17542 7052 19178
rect 7116 18834 7144 19178
rect 7208 19145 7236 19246
rect 7194 19136 7250 19145
rect 7194 19071 7250 19080
rect 7104 18828 7156 18834
rect 7104 18770 7156 18776
rect 7012 17536 7064 17542
rect 7012 17478 7064 17484
rect 7012 17128 7064 17134
rect 7012 17070 7064 17076
rect 7024 16590 7052 17070
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7012 16584 7064 16590
rect 7012 16526 7064 16532
rect 7024 16046 7052 16526
rect 7300 16046 7328 16730
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 7024 15162 7052 15982
rect 7104 15360 7156 15366
rect 7104 15302 7156 15308
rect 7012 15156 7064 15162
rect 7012 15098 7064 15104
rect 7116 14822 7144 15302
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 6920 12640 6972 12646
rect 6920 12582 6972 12588
rect 6932 12306 6960 12582
rect 6920 12300 6972 12306
rect 6920 12242 6972 12248
rect 7116 11778 7144 14758
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7300 13326 7328 13466
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7300 12186 7328 13262
rect 7024 11750 7144 11778
rect 7208 12158 7328 12186
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6564 10470 6592 10542
rect 6552 10464 6604 10470
rect 6552 10406 6604 10412
rect 6564 8294 6592 10406
rect 7024 10130 7052 11750
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7116 11218 7144 11630
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 7024 9926 7052 10066
rect 7012 9920 7064 9926
rect 7012 9862 7064 9868
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6840 8294 6868 8366
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6840 7342 6868 8230
rect 7024 7750 7052 9862
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 7116 8022 7144 8366
rect 7104 8016 7156 8022
rect 7104 7958 7156 7964
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5736 5846 5764 6734
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 5920 5914 5948 6054
rect 6840 5914 6868 7278
rect 7116 6934 7144 7822
rect 7104 6928 7156 6934
rect 7104 6870 7156 6876
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 5724 5840 5776 5846
rect 5724 5782 5776 5788
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5644 5370 5672 5646
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5816 5160 5868 5166
rect 5816 5102 5868 5108
rect 5828 4622 5856 5102
rect 5920 4690 5948 5850
rect 7208 5250 7236 12158
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7300 11762 7328 12038
rect 7392 11898 7420 35226
rect 7576 30802 7604 42842
rect 7852 41818 7880 43182
rect 8116 42764 8168 42770
rect 8116 42706 8168 42712
rect 8024 42628 8076 42634
rect 8024 42570 8076 42576
rect 7840 41812 7892 41818
rect 7840 41754 7892 41760
rect 7932 41676 7984 41682
rect 7932 41618 7984 41624
rect 7944 39846 7972 41618
rect 8036 40526 8064 42570
rect 8128 41682 8156 42706
rect 8588 42226 8616 43250
rect 12348 43240 12400 43246
rect 12348 43182 12400 43188
rect 15476 43240 15528 43246
rect 15476 43182 15528 43188
rect 8944 43104 8996 43110
rect 8944 43046 8996 43052
rect 8852 42560 8904 42566
rect 8852 42502 8904 42508
rect 8864 42226 8892 42502
rect 8576 42220 8628 42226
rect 8576 42162 8628 42168
rect 8852 42220 8904 42226
rect 8852 42162 8904 42168
rect 8116 41676 8168 41682
rect 8116 41618 8168 41624
rect 8956 41274 8984 43046
rect 12360 42906 12388 43182
rect 12532 43104 12584 43110
rect 12532 43046 12584 43052
rect 12348 42900 12400 42906
rect 12348 42842 12400 42848
rect 10784 42696 10836 42702
rect 10784 42638 10836 42644
rect 11520 42696 11572 42702
rect 11520 42638 11572 42644
rect 10048 42560 10100 42566
rect 10048 42502 10100 42508
rect 10060 42226 10088 42502
rect 10048 42220 10100 42226
rect 10048 42162 10100 42168
rect 10796 42158 10824 42638
rect 10784 42152 10836 42158
rect 10784 42094 10836 42100
rect 10508 42016 10560 42022
rect 10508 41958 10560 41964
rect 11428 42016 11480 42022
rect 11428 41958 11480 41964
rect 9128 41744 9180 41750
rect 9128 41686 9180 41692
rect 8392 41268 8444 41274
rect 8392 41210 8444 41216
rect 8944 41268 8996 41274
rect 8944 41210 8996 41216
rect 8404 41070 8432 41210
rect 8392 41064 8444 41070
rect 8392 41006 8444 41012
rect 8208 40656 8260 40662
rect 8208 40598 8260 40604
rect 8024 40520 8076 40526
rect 8024 40462 8076 40468
rect 8220 39982 8248 40598
rect 8484 40588 8536 40594
rect 8484 40530 8536 40536
rect 8496 39982 8524 40530
rect 9140 40118 9168 41686
rect 10520 41682 10548 41958
rect 10508 41676 10560 41682
rect 10508 41618 10560 41624
rect 11060 41676 11112 41682
rect 11060 41618 11112 41624
rect 10324 41608 10376 41614
rect 10324 41550 10376 41556
rect 9680 41132 9732 41138
rect 9680 41074 9732 41080
rect 9692 40186 9720 41074
rect 10336 40390 10364 41550
rect 11072 41478 11100 41618
rect 11060 41472 11112 41478
rect 11060 41414 11112 41420
rect 10968 40520 11020 40526
rect 10968 40462 11020 40468
rect 10980 40390 11008 40462
rect 10324 40384 10376 40390
rect 10324 40326 10376 40332
rect 10968 40384 11020 40390
rect 10968 40326 11020 40332
rect 9680 40180 9732 40186
rect 9680 40122 9732 40128
rect 9128 40112 9180 40118
rect 9128 40054 9180 40060
rect 8576 40044 8628 40050
rect 8944 40044 8996 40050
rect 8628 40004 8944 40032
rect 8576 39986 8628 39992
rect 8944 39986 8996 39992
rect 8208 39976 8260 39982
rect 8208 39918 8260 39924
rect 8484 39976 8536 39982
rect 8484 39918 8536 39924
rect 7932 39840 7984 39846
rect 7932 39782 7984 39788
rect 7838 39536 7894 39545
rect 7838 39471 7840 39480
rect 7892 39471 7894 39480
rect 7840 39442 7892 39448
rect 7746 39400 7802 39409
rect 7746 39335 7748 39344
rect 7800 39335 7802 39344
rect 7748 39306 7800 39312
rect 7852 39302 7880 39442
rect 7840 39296 7892 39302
rect 7840 39238 7892 39244
rect 7944 39098 7972 39782
rect 8220 39574 8248 39918
rect 8208 39568 8260 39574
rect 8300 39568 8352 39574
rect 8208 39510 8260 39516
rect 8298 39536 8300 39545
rect 8352 39536 8354 39545
rect 7932 39092 7984 39098
rect 7932 39034 7984 39040
rect 8220 38894 8248 39510
rect 8298 39471 8354 39480
rect 8300 39296 8352 39302
rect 8300 39238 8352 39244
rect 8208 38888 8260 38894
rect 8208 38830 8260 38836
rect 8220 38214 8248 38830
rect 8208 38208 8260 38214
rect 8208 38150 8260 38156
rect 8220 37806 8248 38150
rect 8208 37800 8260 37806
rect 8208 37742 8260 37748
rect 7656 37120 7708 37126
rect 7656 37062 7708 37068
rect 7668 36718 7696 37062
rect 7656 36712 7708 36718
rect 7656 36654 7708 36660
rect 7748 36168 7800 36174
rect 7748 36110 7800 36116
rect 7760 35698 7788 36110
rect 7748 35692 7800 35698
rect 7748 35634 7800 35640
rect 7564 30796 7616 30802
rect 7564 30738 7616 30744
rect 7470 26208 7526 26217
rect 7470 26143 7526 26152
rect 7484 25430 7512 26143
rect 7472 25424 7524 25430
rect 7472 25366 7524 25372
rect 7484 24410 7512 25366
rect 7472 24404 7524 24410
rect 7472 24346 7524 24352
rect 7484 24274 7512 24346
rect 7472 24268 7524 24274
rect 7472 24210 7524 24216
rect 7472 22976 7524 22982
rect 7472 22918 7524 22924
rect 7484 22098 7512 22918
rect 7472 22092 7524 22098
rect 7472 22034 7524 22040
rect 7576 21078 7604 30738
rect 7656 29708 7708 29714
rect 7656 29650 7708 29656
rect 7668 27538 7696 29650
rect 7840 28076 7892 28082
rect 7840 28018 7892 28024
rect 7656 27532 7708 27538
rect 7656 27474 7708 27480
rect 7668 27334 7696 27474
rect 7656 27328 7708 27334
rect 7656 27270 7708 27276
rect 7852 25906 7880 28018
rect 8312 28014 8340 39238
rect 8496 38894 8524 39918
rect 9692 39506 9720 40122
rect 9680 39500 9732 39506
rect 9680 39442 9732 39448
rect 8484 38888 8536 38894
rect 8484 38830 8536 38836
rect 8496 38554 8524 38830
rect 9956 38752 10008 38758
rect 9956 38694 10008 38700
rect 8484 38548 8536 38554
rect 8484 38490 8536 38496
rect 8496 37806 8524 38490
rect 8576 38412 8628 38418
rect 8576 38354 8628 38360
rect 8484 37800 8536 37806
rect 8484 37742 8536 37748
rect 8588 37398 8616 38354
rect 9588 38344 9640 38350
rect 9588 38286 9640 38292
rect 8576 37392 8628 37398
rect 8576 37334 8628 37340
rect 8588 36582 8616 37334
rect 8944 37256 8996 37262
rect 8944 37198 8996 37204
rect 8760 36780 8812 36786
rect 8760 36722 8812 36728
rect 8576 36576 8628 36582
rect 8576 36518 8628 36524
rect 8588 36242 8616 36518
rect 8576 36236 8628 36242
rect 8576 36178 8628 36184
rect 8668 36168 8720 36174
rect 8772 36122 8800 36722
rect 8956 36378 8984 37198
rect 9600 36718 9628 38286
rect 9968 38214 9996 38694
rect 9956 38208 10008 38214
rect 9956 38150 10008 38156
rect 9772 36848 9824 36854
rect 9772 36790 9824 36796
rect 9588 36712 9640 36718
rect 9588 36654 9640 36660
rect 8944 36372 8996 36378
rect 8944 36314 8996 36320
rect 8956 36242 8984 36314
rect 8944 36236 8996 36242
rect 8944 36178 8996 36184
rect 8720 36116 8800 36122
rect 8668 36110 8800 36116
rect 8680 36094 8800 36110
rect 8772 36038 8800 36094
rect 8760 36032 8812 36038
rect 8760 35974 8812 35980
rect 8484 32768 8536 32774
rect 8484 32710 8536 32716
rect 8390 31920 8446 31929
rect 8390 31855 8446 31864
rect 8404 31822 8432 31855
rect 8392 31816 8444 31822
rect 8392 31758 8444 31764
rect 8496 31278 8524 32710
rect 8576 32224 8628 32230
rect 8576 32166 8628 32172
rect 8588 31890 8616 32166
rect 8576 31884 8628 31890
rect 8576 31826 8628 31832
rect 8668 31680 8720 31686
rect 8668 31622 8720 31628
rect 8680 31346 8708 31622
rect 8668 31340 8720 31346
rect 8668 31282 8720 31288
rect 8484 31272 8536 31278
rect 8484 31214 8536 31220
rect 8484 29572 8536 29578
rect 8484 29514 8536 29520
rect 8496 29170 8524 29514
rect 8484 29164 8536 29170
rect 8484 29106 8536 29112
rect 7932 28008 7984 28014
rect 7932 27950 7984 27956
rect 8300 28008 8352 28014
rect 8300 27950 8352 27956
rect 7840 25900 7892 25906
rect 7840 25842 7892 25848
rect 7748 23180 7800 23186
rect 7748 23122 7800 23128
rect 7760 22166 7788 23122
rect 7748 22160 7800 22166
rect 7748 22102 7800 22108
rect 7760 21690 7788 22102
rect 7748 21684 7800 21690
rect 7748 21626 7800 21632
rect 7852 21078 7880 25842
rect 7944 25702 7972 27950
rect 8484 27532 8536 27538
rect 8484 27474 8536 27480
rect 8392 27464 8444 27470
rect 8496 27441 8524 27474
rect 8392 27406 8444 27412
rect 8482 27432 8538 27441
rect 8404 26790 8432 27406
rect 8482 27367 8538 27376
rect 8392 26784 8444 26790
rect 8392 26726 8444 26732
rect 8576 26784 8628 26790
rect 8576 26726 8628 26732
rect 8024 26240 8076 26246
rect 8024 26182 8076 26188
rect 8036 25770 8064 26182
rect 8024 25764 8076 25770
rect 8024 25706 8076 25712
rect 7932 25696 7984 25702
rect 7932 25638 7984 25644
rect 7932 25152 7984 25158
rect 7932 25094 7984 25100
rect 7944 24818 7972 25094
rect 7932 24812 7984 24818
rect 7932 24754 7984 24760
rect 7944 24614 7972 24754
rect 7932 24608 7984 24614
rect 7932 24550 7984 24556
rect 8024 23792 8076 23798
rect 8024 23734 8076 23740
rect 7932 22568 7984 22574
rect 7932 22510 7984 22516
rect 7944 22234 7972 22510
rect 7932 22228 7984 22234
rect 7932 22170 7984 22176
rect 8036 21604 8064 23734
rect 7944 21576 8064 21604
rect 7564 21072 7616 21078
rect 7564 21014 7616 21020
rect 7840 21072 7892 21078
rect 7840 21014 7892 21020
rect 7472 19848 7524 19854
rect 7472 19790 7524 19796
rect 7840 19848 7892 19854
rect 7840 19790 7892 19796
rect 7484 18698 7512 19790
rect 7656 19236 7708 19242
rect 7656 19178 7708 19184
rect 7668 18834 7696 19178
rect 7852 18834 7880 19790
rect 7656 18828 7708 18834
rect 7656 18770 7708 18776
rect 7840 18828 7892 18834
rect 7840 18770 7892 18776
rect 7472 18692 7524 18698
rect 7472 18634 7524 18640
rect 7484 17134 7512 18634
rect 7748 18624 7800 18630
rect 7748 18566 7800 18572
rect 7656 17536 7708 17542
rect 7656 17478 7708 17484
rect 7668 17134 7696 17478
rect 7472 17128 7524 17134
rect 7472 17070 7524 17076
rect 7656 17128 7708 17134
rect 7656 17070 7708 17076
rect 7484 16522 7512 17070
rect 7472 16516 7524 16522
rect 7472 16458 7524 16464
rect 7484 16182 7512 16458
rect 7472 16176 7524 16182
rect 7472 16118 7524 16124
rect 7564 15156 7616 15162
rect 7564 15098 7616 15104
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7484 12714 7512 13262
rect 7472 12708 7524 12714
rect 7472 12650 7524 12656
rect 7472 12232 7524 12238
rect 7470 12200 7472 12209
rect 7524 12200 7526 12209
rect 7470 12135 7526 12144
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7288 11756 7340 11762
rect 7288 11698 7340 11704
rect 7380 11144 7432 11150
rect 7380 11086 7432 11092
rect 7392 10810 7420 11086
rect 7380 10804 7432 10810
rect 7380 10746 7432 10752
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 7300 6322 7328 7278
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7116 5222 7236 5250
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6932 4826 6960 5102
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 5816 4616 5868 4622
rect 5816 4558 5868 4564
rect 5828 4078 5856 4558
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 7116 3738 7144 5222
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 7208 4758 7236 5102
rect 7196 4752 7248 4758
rect 7196 4694 7248 4700
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 7576 2990 7604 15098
rect 7760 12322 7788 18566
rect 7840 16992 7892 16998
rect 7840 16934 7892 16940
rect 7852 16658 7880 16934
rect 7840 16652 7892 16658
rect 7840 16594 7892 16600
rect 7944 16130 7972 21576
rect 8116 20392 8168 20398
rect 8116 20334 8168 20340
rect 8024 20324 8076 20330
rect 8024 20266 8076 20272
rect 8036 18222 8064 20266
rect 8128 20058 8156 20334
rect 8116 20052 8168 20058
rect 8116 19994 8168 20000
rect 8128 19922 8156 19994
rect 8116 19916 8168 19922
rect 8116 19858 8168 19864
rect 8300 19372 8352 19378
rect 8300 19314 8352 19320
rect 8116 18828 8168 18834
rect 8116 18770 8168 18776
rect 8128 18737 8156 18770
rect 8114 18728 8170 18737
rect 8114 18663 8170 18672
rect 8024 18216 8076 18222
rect 8024 18158 8076 18164
rect 8312 18154 8340 19314
rect 8404 19310 8432 26726
rect 8588 26518 8616 26726
rect 8576 26512 8628 26518
rect 8576 26454 8628 26460
rect 8576 25696 8628 25702
rect 8576 25638 8628 25644
rect 8588 25498 8616 25638
rect 8576 25492 8628 25498
rect 8576 25434 8628 25440
rect 8484 24812 8536 24818
rect 8484 24754 8536 24760
rect 8496 23866 8524 24754
rect 8484 23860 8536 23866
rect 8484 23802 8536 23808
rect 8772 20602 8800 35974
rect 9600 35562 9628 36654
rect 9588 35556 9640 35562
rect 9588 35498 9640 35504
rect 9404 35080 9456 35086
rect 9404 35022 9456 35028
rect 9312 33652 9364 33658
rect 9312 33594 9364 33600
rect 9324 30326 9352 33594
rect 9416 31396 9444 35022
rect 9784 34202 9812 36790
rect 9968 35222 9996 38150
rect 10048 37188 10100 37194
rect 10048 37130 10100 37136
rect 10060 36854 10088 37130
rect 10048 36848 10100 36854
rect 10048 36790 10100 36796
rect 10232 36780 10284 36786
rect 10232 36722 10284 36728
rect 9956 35216 10008 35222
rect 9956 35158 10008 35164
rect 10244 34202 10272 36722
rect 9772 34196 9824 34202
rect 9772 34138 9824 34144
rect 10232 34196 10284 34202
rect 10232 34138 10284 34144
rect 9784 34066 9812 34138
rect 9772 34060 9824 34066
rect 9772 34002 9824 34008
rect 10140 34060 10192 34066
rect 10140 34002 10192 34008
rect 9680 32360 9732 32366
rect 9680 32302 9732 32308
rect 9692 31958 9720 32302
rect 9680 31952 9732 31958
rect 9956 31952 10008 31958
rect 9680 31894 9732 31900
rect 9954 31920 9956 31929
rect 10008 31920 10010 31929
rect 9954 31855 10010 31864
rect 9678 31512 9734 31521
rect 9678 31447 9734 31456
rect 9692 31396 9720 31447
rect 9416 31368 9720 31396
rect 9864 31272 9916 31278
rect 9864 31214 9916 31220
rect 9876 31142 9904 31214
rect 10152 31210 10180 34002
rect 10244 31890 10272 34138
rect 10336 32434 10364 40326
rect 10784 38888 10836 38894
rect 10784 38830 10836 38836
rect 10796 38758 10824 38830
rect 10784 38752 10836 38758
rect 10784 38694 10836 38700
rect 10600 38004 10652 38010
rect 10600 37946 10652 37952
rect 10324 32428 10376 32434
rect 10324 32370 10376 32376
rect 10232 31884 10284 31890
rect 10232 31826 10284 31832
rect 10324 31816 10376 31822
rect 10324 31758 10376 31764
rect 10140 31204 10192 31210
rect 10140 31146 10192 31152
rect 9864 31136 9916 31142
rect 9864 31078 9916 31084
rect 9312 30320 9364 30326
rect 9312 30262 9364 30268
rect 9324 29850 9352 30262
rect 9404 30184 9456 30190
rect 9404 30126 9456 30132
rect 9416 30054 9444 30126
rect 9404 30048 9456 30054
rect 9404 29990 9456 29996
rect 9312 29844 9364 29850
rect 9312 29786 9364 29792
rect 9416 29170 9444 29990
rect 9876 29646 9904 31078
rect 9864 29640 9916 29646
rect 9864 29582 9916 29588
rect 9404 29164 9456 29170
rect 9404 29106 9456 29112
rect 9036 24608 9088 24614
rect 9036 24550 9088 24556
rect 9048 22778 9076 24550
rect 9036 22772 9088 22778
rect 9036 22714 9088 22720
rect 9128 22092 9180 22098
rect 9128 22034 9180 22040
rect 9140 21486 9168 22034
rect 9312 21684 9364 21690
rect 9312 21626 9364 21632
rect 9324 21486 9352 21626
rect 9128 21480 9180 21486
rect 9128 21422 9180 21428
rect 9312 21480 9364 21486
rect 9312 21422 9364 21428
rect 8760 20596 8812 20602
rect 8760 20538 8812 20544
rect 8484 20256 8536 20262
rect 8484 20198 8536 20204
rect 8496 19718 8524 20198
rect 9140 19990 9168 21422
rect 9128 19984 9180 19990
rect 9128 19926 9180 19932
rect 9312 19916 9364 19922
rect 9312 19858 9364 19864
rect 8484 19712 8536 19718
rect 8484 19654 8536 19660
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 8668 19304 8720 19310
rect 8668 19246 8720 19252
rect 8850 19272 8906 19281
rect 8484 19236 8536 19242
rect 8484 19178 8536 19184
rect 8496 19145 8524 19178
rect 8680 19174 8708 19246
rect 8850 19207 8906 19216
rect 8864 19174 8892 19207
rect 8668 19168 8720 19174
rect 8482 19136 8538 19145
rect 8668 19110 8720 19116
rect 8852 19168 8904 19174
rect 8852 19110 8904 19116
rect 8482 19071 8538 19080
rect 9036 18896 9088 18902
rect 9036 18838 9088 18844
rect 8482 18728 8538 18737
rect 8482 18663 8538 18672
rect 8300 18148 8352 18154
rect 8300 18090 8352 18096
rect 8024 17672 8076 17678
rect 8024 17614 8076 17620
rect 8036 16794 8064 17614
rect 8300 17536 8352 17542
rect 8300 17478 8352 17484
rect 8312 17134 8340 17478
rect 8300 17128 8352 17134
rect 8300 17070 8352 17076
rect 8024 16788 8076 16794
rect 8024 16730 8076 16736
rect 7852 16102 7972 16130
rect 7852 13530 7880 16102
rect 7932 15972 7984 15978
rect 7932 15914 7984 15920
rect 7944 15638 7972 15914
rect 7932 15632 7984 15638
rect 7932 15574 7984 15580
rect 8392 15496 8444 15502
rect 8392 15438 8444 15444
rect 7932 14952 7984 14958
rect 7932 14894 7984 14900
rect 7944 14618 7972 14894
rect 8404 14890 8432 15438
rect 8392 14884 8444 14890
rect 8392 14826 8444 14832
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8312 13530 8340 13806
rect 7840 13524 7892 13530
rect 7840 13466 7892 13472
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8392 12980 8444 12986
rect 8392 12922 8444 12928
rect 7760 12294 7880 12322
rect 7748 9988 7800 9994
rect 7748 9930 7800 9936
rect 7760 9654 7788 9930
rect 7748 9648 7800 9654
rect 7748 9590 7800 9596
rect 7760 9042 7788 9590
rect 7852 9110 7880 12294
rect 8300 12096 8352 12102
rect 8300 12038 8352 12044
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8022 10704 8078 10713
rect 8022 10639 8024 10648
rect 8076 10639 8078 10648
rect 8024 10610 8076 10616
rect 8128 10033 8156 10746
rect 8312 10606 8340 12038
rect 8404 11898 8432 12922
rect 8496 12442 8524 18663
rect 9048 18426 9076 18838
rect 9126 18728 9182 18737
rect 9126 18663 9182 18672
rect 9140 18630 9168 18663
rect 9128 18624 9180 18630
rect 9128 18566 9180 18572
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 9048 18222 9076 18362
rect 9036 18216 9088 18222
rect 9036 18158 9088 18164
rect 9220 18216 9272 18222
rect 9220 18158 9272 18164
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 8588 12986 8616 18022
rect 9128 17604 9180 17610
rect 9128 17546 9180 17552
rect 9140 17134 9168 17546
rect 9128 17128 9180 17134
rect 9128 17070 9180 17076
rect 9232 16726 9260 18158
rect 9324 16998 9352 19858
rect 9416 19310 9444 29106
rect 9876 29102 9904 29582
rect 9864 29096 9916 29102
rect 9864 29038 9916 29044
rect 9588 27668 9640 27674
rect 9588 27610 9640 27616
rect 9496 27600 9548 27606
rect 9600 27577 9628 27610
rect 9496 27542 9548 27548
rect 9586 27568 9642 27577
rect 9508 27470 9536 27542
rect 9586 27503 9642 27512
rect 9772 27532 9824 27538
rect 9772 27474 9824 27480
rect 9496 27464 9548 27470
rect 9784 27441 9812 27474
rect 9496 27406 9548 27412
rect 9770 27432 9826 27441
rect 9770 27367 9826 27376
rect 9864 23656 9916 23662
rect 9864 23598 9916 23604
rect 9772 22976 9824 22982
rect 9772 22918 9824 22924
rect 9678 22808 9734 22817
rect 9678 22743 9680 22752
rect 9732 22743 9734 22752
rect 9680 22714 9732 22720
rect 9692 22574 9720 22714
rect 9680 22568 9732 22574
rect 9680 22510 9732 22516
rect 9496 22024 9548 22030
rect 9496 21966 9548 21972
rect 9508 21593 9536 21966
rect 9494 21584 9550 21593
rect 9784 21554 9812 22918
rect 9876 21962 9904 23598
rect 9956 22432 10008 22438
rect 9956 22374 10008 22380
rect 9864 21956 9916 21962
rect 9864 21898 9916 21904
rect 9968 21894 9996 22374
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 9494 21519 9550 21528
rect 9772 21548 9824 21554
rect 9772 21490 9824 21496
rect 9784 19310 9812 21490
rect 9404 19304 9456 19310
rect 9404 19246 9456 19252
rect 9772 19304 9824 19310
rect 9772 19246 9824 19252
rect 9680 18352 9732 18358
rect 9680 18294 9732 18300
rect 9404 18148 9456 18154
rect 9404 18090 9456 18096
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 9220 16720 9272 16726
rect 9220 16662 9272 16668
rect 9324 16658 9352 16934
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 8668 15156 8720 15162
rect 8668 15098 8720 15104
rect 8680 14521 8708 15098
rect 8666 14512 8722 14521
rect 8666 14447 8722 14456
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8680 13394 8708 14214
rect 8668 13388 8720 13394
rect 8668 13330 8720 13336
rect 8576 12980 8628 12986
rect 8576 12922 8628 12928
rect 8484 12436 8536 12442
rect 8484 12378 8536 12384
rect 8392 11892 8444 11898
rect 8392 11834 8444 11840
rect 8496 11354 8524 12378
rect 8852 11688 8904 11694
rect 8852 11630 8904 11636
rect 8864 11354 8892 11630
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8114 10024 8170 10033
rect 8114 9959 8170 9968
rect 9416 9518 9444 18090
rect 9496 18080 9548 18086
rect 9494 18048 9496 18057
rect 9548 18048 9550 18057
rect 9494 17983 9550 17992
rect 9588 14272 9640 14278
rect 9588 14214 9640 14220
rect 9600 14074 9628 14214
rect 9588 14068 9640 14074
rect 9588 14010 9640 14016
rect 9692 13870 9720 18294
rect 9968 16114 9996 21830
rect 9956 16108 10008 16114
rect 9956 16050 10008 16056
rect 10152 15706 10180 31146
rect 10336 30802 10364 31758
rect 10324 30796 10376 30802
rect 10324 30738 10376 30744
rect 10612 30190 10640 37946
rect 10796 37874 10824 38694
rect 10784 37868 10836 37874
rect 10784 37810 10836 37816
rect 11440 36718 11468 41958
rect 11532 41818 11560 42638
rect 11796 42356 11848 42362
rect 11796 42298 11848 42304
rect 11520 41812 11572 41818
rect 11520 41754 11572 41760
rect 11808 41750 11836 42298
rect 12544 41818 12572 43046
rect 15488 42770 15516 43182
rect 15476 42764 15528 42770
rect 15476 42706 15528 42712
rect 13728 42560 13780 42566
rect 13728 42502 13780 42508
rect 13740 41818 13768 42502
rect 15672 42226 15700 43726
rect 17040 43648 17092 43654
rect 17040 43590 17092 43596
rect 16672 43240 16724 43246
rect 16672 43182 16724 43188
rect 16488 43104 16540 43110
rect 16488 43046 16540 43052
rect 16500 42770 16528 43046
rect 16488 42764 16540 42770
rect 16488 42706 16540 42712
rect 16684 42294 16712 43182
rect 17052 42770 17080 43590
rect 17040 42764 17092 42770
rect 17040 42706 17092 42712
rect 16672 42288 16724 42294
rect 16672 42230 16724 42236
rect 15660 42220 15712 42226
rect 15660 42162 15712 42168
rect 16764 42220 16816 42226
rect 16764 42162 16816 42168
rect 12532 41812 12584 41818
rect 12532 41754 12584 41760
rect 13728 41812 13780 41818
rect 13728 41754 13780 41760
rect 11796 41744 11848 41750
rect 11796 41686 11848 41692
rect 14188 41676 14240 41682
rect 14188 41618 14240 41624
rect 12532 41608 12584 41614
rect 12532 41550 12584 41556
rect 11980 40588 12032 40594
rect 11980 40530 12032 40536
rect 12072 40588 12124 40594
rect 12072 40530 12124 40536
rect 11992 39846 12020 40530
rect 12084 39982 12112 40530
rect 12440 40180 12492 40186
rect 12440 40122 12492 40128
rect 12072 39976 12124 39982
rect 12072 39918 12124 39924
rect 11980 39840 12032 39846
rect 11980 39782 12032 39788
rect 11796 39500 11848 39506
rect 11796 39442 11848 39448
rect 11808 37777 11836 39442
rect 11992 39302 12020 39782
rect 11980 39296 12032 39302
rect 11980 39238 12032 39244
rect 12084 38894 12112 39918
rect 12072 38888 12124 38894
rect 12072 38830 12124 38836
rect 11980 38548 12032 38554
rect 11980 38490 12032 38496
rect 11992 38418 12020 38490
rect 11980 38412 12032 38418
rect 11980 38354 12032 38360
rect 12164 38412 12216 38418
rect 12164 38354 12216 38360
rect 12176 37806 12204 38354
rect 12164 37800 12216 37806
rect 11794 37768 11850 37777
rect 12164 37742 12216 37748
rect 11794 37703 11850 37712
rect 11428 36712 11480 36718
rect 11428 36654 11480 36660
rect 11440 35986 11468 36654
rect 11808 36378 11836 37703
rect 12176 37330 12204 37742
rect 12164 37324 12216 37330
rect 12164 37266 12216 37272
rect 12254 36816 12310 36825
rect 12254 36751 12310 36760
rect 12268 36650 12296 36751
rect 12348 36712 12400 36718
rect 12346 36680 12348 36689
rect 12400 36680 12402 36689
rect 12256 36644 12308 36650
rect 12346 36615 12402 36624
rect 12256 36586 12308 36592
rect 11796 36372 11848 36378
rect 11796 36314 11848 36320
rect 11808 36242 11836 36314
rect 11796 36236 11848 36242
rect 11796 36178 11848 36184
rect 12348 36100 12400 36106
rect 12348 36042 12400 36048
rect 12360 35986 12388 36042
rect 12452 35986 12480 40122
rect 12544 39914 12572 41550
rect 13084 41472 13136 41478
rect 13084 41414 13136 41420
rect 12992 41064 13044 41070
rect 12992 41006 13044 41012
rect 13004 40730 13032 41006
rect 12992 40724 13044 40730
rect 12992 40666 13044 40672
rect 12716 40588 12768 40594
rect 12716 40530 12768 40536
rect 12728 40118 12756 40530
rect 12716 40112 12768 40118
rect 12716 40054 12768 40060
rect 12808 40044 12860 40050
rect 12808 39986 12860 39992
rect 12820 39930 12848 39986
rect 12532 39908 12584 39914
rect 12532 39850 12584 39856
rect 12624 39908 12676 39914
rect 12624 39850 12676 39856
rect 12728 39902 12848 39930
rect 12636 39030 12664 39850
rect 12728 39846 12756 39902
rect 12716 39840 12768 39846
rect 12716 39782 12768 39788
rect 12728 39438 12756 39782
rect 13096 39506 13124 41414
rect 14200 41206 14228 41618
rect 14280 41472 14332 41478
rect 14280 41414 14332 41420
rect 14188 41200 14240 41206
rect 14188 41142 14240 41148
rect 13728 41064 13780 41070
rect 13728 41006 13780 41012
rect 13636 40928 13688 40934
rect 13636 40870 13688 40876
rect 13544 40588 13596 40594
rect 13544 40530 13596 40536
rect 13556 40186 13584 40530
rect 13544 40180 13596 40186
rect 13544 40122 13596 40128
rect 13084 39500 13136 39506
rect 13084 39442 13136 39448
rect 13544 39500 13596 39506
rect 13544 39442 13596 39448
rect 12716 39432 12768 39438
rect 12716 39374 12768 39380
rect 12728 39302 12756 39374
rect 12716 39296 12768 39302
rect 12716 39238 12768 39244
rect 12624 39024 12676 39030
rect 12624 38966 12676 38972
rect 12728 38570 12756 39238
rect 12636 38542 12756 38570
rect 13556 38554 13584 39442
rect 13648 38894 13676 40870
rect 13740 40594 13768 41006
rect 14292 41002 14320 41414
rect 14280 40996 14332 41002
rect 14280 40938 14332 40944
rect 13728 40588 13780 40594
rect 13728 40530 13780 40536
rect 14292 40526 14320 40938
rect 15384 40928 15436 40934
rect 15384 40870 15436 40876
rect 14280 40520 14332 40526
rect 14280 40462 14332 40468
rect 13728 40384 13780 40390
rect 13728 40326 13780 40332
rect 13740 40118 13768 40326
rect 15396 40186 15424 40870
rect 15384 40180 15436 40186
rect 15384 40122 15436 40128
rect 13728 40112 13780 40118
rect 13728 40054 13780 40060
rect 13740 39982 13768 40054
rect 13728 39976 13780 39982
rect 13728 39918 13780 39924
rect 13912 39976 13964 39982
rect 13912 39918 13964 39924
rect 15200 39976 15252 39982
rect 15200 39918 15252 39924
rect 13924 39846 13952 39918
rect 14280 39908 14332 39914
rect 14280 39850 14332 39856
rect 13912 39840 13964 39846
rect 13912 39782 13964 39788
rect 14292 39545 14320 39850
rect 14278 39536 14334 39545
rect 13820 39500 13872 39506
rect 14278 39471 14334 39480
rect 14464 39500 14516 39506
rect 13820 39442 13872 39448
rect 14464 39442 14516 39448
rect 13832 39098 13860 39442
rect 14476 39302 14504 39442
rect 14096 39296 14148 39302
rect 14464 39296 14516 39302
rect 14096 39238 14148 39244
rect 14462 39264 14464 39273
rect 14516 39264 14518 39273
rect 13820 39092 13872 39098
rect 13820 39034 13872 39040
rect 14108 39001 14136 39238
rect 14462 39199 14518 39208
rect 14094 38992 14150 39001
rect 13820 38956 13872 38962
rect 14094 38927 14150 38936
rect 13820 38898 13872 38904
rect 13636 38888 13688 38894
rect 13636 38830 13688 38836
rect 13832 38758 13860 38898
rect 13820 38752 13872 38758
rect 13820 38694 13872 38700
rect 13544 38548 13596 38554
rect 12532 37120 12584 37126
rect 12532 37062 12584 37068
rect 12544 36106 12572 37062
rect 12532 36100 12584 36106
rect 12532 36042 12584 36048
rect 11440 35958 11560 35986
rect 12360 35958 12572 35986
rect 10876 35624 10928 35630
rect 10876 35566 10928 35572
rect 11428 35624 11480 35630
rect 11428 35566 11480 35572
rect 10888 35494 10916 35566
rect 10876 35488 10928 35494
rect 10876 35430 10928 35436
rect 10888 34610 10916 35430
rect 11440 34746 11468 35566
rect 11428 34740 11480 34746
rect 11428 34682 11480 34688
rect 10876 34604 10928 34610
rect 10876 34546 10928 34552
rect 10888 32026 10916 34546
rect 11244 33856 11296 33862
rect 11244 33798 11296 33804
rect 11256 33590 11284 33798
rect 11244 33584 11296 33590
rect 11244 33526 11296 33532
rect 11256 32366 11284 33526
rect 11440 33046 11468 34682
rect 11532 34202 11560 35958
rect 11520 34196 11572 34202
rect 11520 34138 11572 34144
rect 11980 34060 12032 34066
rect 11980 34002 12032 34008
rect 11888 33924 11940 33930
rect 11888 33866 11940 33872
rect 11704 33312 11756 33318
rect 11704 33254 11756 33260
rect 11428 33040 11480 33046
rect 11428 32982 11480 32988
rect 11244 32360 11296 32366
rect 11244 32302 11296 32308
rect 10876 32020 10928 32026
rect 10876 31962 10928 31968
rect 10888 31890 10916 31962
rect 10876 31884 10928 31890
rect 10876 31826 10928 31832
rect 10888 30682 10916 31826
rect 10968 31204 11020 31210
rect 10968 31146 11020 31152
rect 10980 30802 11008 31146
rect 10968 30796 11020 30802
rect 10968 30738 11020 30744
rect 11060 30728 11112 30734
rect 10888 30654 11008 30682
rect 11060 30670 11112 30676
rect 10600 30184 10652 30190
rect 10600 30126 10652 30132
rect 10876 30116 10928 30122
rect 10876 30058 10928 30064
rect 10692 30048 10744 30054
rect 10692 29990 10744 29996
rect 10704 29102 10732 29990
rect 10888 29782 10916 30058
rect 10876 29776 10928 29782
rect 10876 29718 10928 29724
rect 10784 29640 10836 29646
rect 10784 29582 10836 29588
rect 10796 29306 10824 29582
rect 10784 29300 10836 29306
rect 10784 29242 10836 29248
rect 10692 29096 10744 29102
rect 10692 29038 10744 29044
rect 10980 28490 11008 30654
rect 11072 30326 11100 30670
rect 11060 30320 11112 30326
rect 11060 30262 11112 30268
rect 11256 30190 11284 32302
rect 11716 31482 11744 33254
rect 11796 32972 11848 32978
rect 11796 32914 11848 32920
rect 11808 32434 11836 32914
rect 11796 32428 11848 32434
rect 11796 32370 11848 32376
rect 11794 31512 11850 31521
rect 11704 31476 11756 31482
rect 11794 31447 11796 31456
rect 11704 31418 11756 31424
rect 11848 31447 11850 31456
rect 11796 31418 11848 31424
rect 11716 31278 11744 31418
rect 11704 31272 11756 31278
rect 11704 31214 11756 31220
rect 11796 31204 11848 31210
rect 11796 31146 11848 31152
rect 11428 30728 11480 30734
rect 11428 30670 11480 30676
rect 11440 30394 11468 30670
rect 11428 30388 11480 30394
rect 11428 30330 11480 30336
rect 11060 30184 11112 30190
rect 11060 30126 11112 30132
rect 11244 30184 11296 30190
rect 11244 30126 11296 30132
rect 11428 30184 11480 30190
rect 11428 30126 11480 30132
rect 10968 28484 11020 28490
rect 10968 28426 11020 28432
rect 10980 26586 11008 28426
rect 11072 27946 11100 30126
rect 11440 30002 11468 30126
rect 11348 29974 11468 30002
rect 11348 29510 11376 29974
rect 11336 29504 11388 29510
rect 11336 29446 11388 29452
rect 11060 27940 11112 27946
rect 11060 27882 11112 27888
rect 10968 26580 11020 26586
rect 10968 26522 11020 26528
rect 10232 26308 10284 26314
rect 10232 26250 10284 26256
rect 10244 25430 10272 26250
rect 10232 25424 10284 25430
rect 10232 25366 10284 25372
rect 10244 17270 10272 25366
rect 11244 24200 11296 24206
rect 11244 24142 11296 24148
rect 11256 23662 11284 24142
rect 10876 23656 10928 23662
rect 10876 23598 10928 23604
rect 11244 23656 11296 23662
rect 11244 23598 11296 23604
rect 10888 23526 10916 23598
rect 10876 23520 10928 23526
rect 10876 23462 10928 23468
rect 10784 19712 10836 19718
rect 10784 19654 10836 19660
rect 10324 19168 10376 19174
rect 10324 19110 10376 19116
rect 10336 18698 10364 19110
rect 10324 18692 10376 18698
rect 10324 18634 10376 18640
rect 10796 18358 10824 19654
rect 11348 19360 11376 29446
rect 11808 28506 11836 31146
rect 11900 30326 11928 33866
rect 11992 32842 12020 34002
rect 12348 33992 12400 33998
rect 12348 33934 12400 33940
rect 11980 32836 12032 32842
rect 11980 32778 12032 32784
rect 11992 32366 12020 32778
rect 12360 32774 12388 33934
rect 12440 33448 12492 33454
rect 12440 33390 12492 33396
rect 12348 32768 12400 32774
rect 12348 32710 12400 32716
rect 11980 32360 12032 32366
rect 11980 32302 12032 32308
rect 11888 30320 11940 30326
rect 11888 30262 11940 30268
rect 11808 28478 11928 28506
rect 11796 28416 11848 28422
rect 11796 28358 11848 28364
rect 11428 27872 11480 27878
rect 11428 27814 11480 27820
rect 11440 27334 11468 27814
rect 11428 27328 11480 27334
rect 11428 27270 11480 27276
rect 11440 26926 11468 27270
rect 11428 26920 11480 26926
rect 11428 26862 11480 26868
rect 11428 24608 11480 24614
rect 11428 24550 11480 24556
rect 11440 24274 11468 24550
rect 11428 24268 11480 24274
rect 11428 24210 11480 24216
rect 11704 21888 11756 21894
rect 11704 21830 11756 21836
rect 11256 19332 11376 19360
rect 10784 18352 10836 18358
rect 10784 18294 10836 18300
rect 10232 17264 10284 17270
rect 10232 17206 10284 17212
rect 10796 16114 10824 18294
rect 10968 17128 11020 17134
rect 10968 17070 11020 17076
rect 11152 17128 11204 17134
rect 11152 17070 11204 17076
rect 10980 16998 11008 17070
rect 10968 16992 11020 16998
rect 10888 16952 10968 16980
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10416 16040 10468 16046
rect 10416 15982 10468 15988
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10428 15638 10456 15982
rect 10692 15972 10744 15978
rect 10692 15914 10744 15920
rect 10704 15638 10732 15914
rect 10416 15632 10468 15638
rect 10416 15574 10468 15580
rect 10692 15632 10744 15638
rect 10692 15574 10744 15580
rect 10428 14958 10456 15574
rect 10416 14952 10468 14958
rect 10416 14894 10468 14900
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10612 14550 10640 14758
rect 10600 14544 10652 14550
rect 10600 14486 10652 14492
rect 10324 14340 10376 14346
rect 10324 14282 10376 14288
rect 9680 13864 9732 13870
rect 9680 13806 9732 13812
rect 9692 13394 9720 13806
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9864 13252 9916 13258
rect 9864 13194 9916 13200
rect 9876 12782 9904 13194
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 9404 9512 9456 9518
rect 9404 9454 9456 9460
rect 10140 9512 10192 9518
rect 10140 9454 10192 9460
rect 7932 9444 7984 9450
rect 7932 9386 7984 9392
rect 8116 9444 8168 9450
rect 8116 9386 8168 9392
rect 7944 9178 7972 9386
rect 7932 9172 7984 9178
rect 7932 9114 7984 9120
rect 7840 9104 7892 9110
rect 7840 9046 7892 9052
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 8128 4010 8156 9386
rect 9680 9036 9732 9042
rect 9680 8978 9732 8984
rect 8300 8968 8352 8974
rect 8300 8910 8352 8916
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8208 8832 8260 8838
rect 8208 8774 8260 8780
rect 8220 8498 8248 8774
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 8220 7206 8248 8230
rect 8312 8090 8340 8910
rect 8404 8634 8432 8910
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 8404 8378 8432 8570
rect 8404 8350 8524 8378
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8496 7954 8524 8350
rect 9692 8022 9720 8978
rect 10152 8634 10180 9454
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10152 8430 10180 8570
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 10140 8424 10192 8430
rect 10140 8366 10192 8372
rect 9680 8016 9732 8022
rect 9680 7958 9732 7964
rect 9784 7954 9812 8366
rect 9864 8288 9916 8294
rect 9864 8230 9916 8236
rect 8484 7948 8536 7954
rect 8484 7890 8536 7896
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 8576 7880 8628 7886
rect 8576 7822 8628 7828
rect 8588 7546 8616 7822
rect 9036 7812 9088 7818
rect 9036 7754 9088 7760
rect 9680 7812 9732 7818
rect 9680 7754 9732 7760
rect 8576 7540 8628 7546
rect 8576 7482 8628 7488
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8588 6254 8616 7482
rect 9048 6254 9076 7754
rect 9692 6458 9720 7754
rect 9770 7440 9826 7449
rect 9770 7375 9772 7384
rect 9824 7375 9826 7384
rect 9772 7346 9824 7352
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9876 6322 9904 8230
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 9036 6248 9088 6254
rect 9036 6190 9088 6196
rect 8864 5370 8892 6190
rect 9048 5710 9076 6190
rect 9876 5778 9904 6258
rect 9864 5772 9916 5778
rect 9864 5714 9916 5720
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 8772 4826 8800 4966
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8116 4004 8168 4010
rect 8116 3946 8168 3952
rect 10336 3058 10364 14282
rect 10888 14074 10916 16952
rect 10968 16934 11020 16940
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 11072 15434 11100 16594
rect 11164 16114 11192 17070
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 11060 15428 11112 15434
rect 11060 15370 11112 15376
rect 11152 15428 11204 15434
rect 11152 15370 11204 15376
rect 11164 14482 11192 15370
rect 11256 15162 11284 19332
rect 11520 17060 11572 17066
rect 11520 17002 11572 17008
rect 11336 16720 11388 16726
rect 11336 16662 11388 16668
rect 11348 15502 11376 16662
rect 11532 16658 11560 17002
rect 11520 16652 11572 16658
rect 11520 16594 11572 16600
rect 11716 16522 11744 21830
rect 11808 16726 11836 28358
rect 11900 25362 11928 28478
rect 11992 28014 12020 32302
rect 12452 29186 12480 33390
rect 12544 32978 12572 35958
rect 12636 34474 12664 38542
rect 13544 38490 13596 38496
rect 12716 38208 12768 38214
rect 12716 38150 12768 38156
rect 12728 37874 12756 38150
rect 12716 37868 12768 37874
rect 12716 37810 12768 37816
rect 13268 37392 13320 37398
rect 13268 37334 13320 37340
rect 12900 37120 12952 37126
rect 12900 37062 12952 37068
rect 12716 36916 12768 36922
rect 12716 36858 12768 36864
rect 12728 36106 12756 36858
rect 12912 36718 12940 37062
rect 13280 36786 13308 37334
rect 13556 36854 13584 38490
rect 13728 37664 13780 37670
rect 13728 37606 13780 37612
rect 13636 37188 13688 37194
rect 13636 37130 13688 37136
rect 13544 36848 13596 36854
rect 13544 36790 13596 36796
rect 13268 36780 13320 36786
rect 13268 36722 13320 36728
rect 12900 36712 12952 36718
rect 12900 36654 12952 36660
rect 13648 36650 13676 37130
rect 12808 36644 12860 36650
rect 12808 36586 12860 36592
rect 13636 36644 13688 36650
rect 13636 36586 13688 36592
rect 12716 36100 12768 36106
rect 12716 36042 12768 36048
rect 12624 34468 12676 34474
rect 12624 34410 12676 34416
rect 12728 33862 12756 36042
rect 12820 35698 12848 36586
rect 12900 36304 12952 36310
rect 12900 36246 12952 36252
rect 12808 35692 12860 35698
rect 12808 35634 12860 35640
rect 12912 35222 12940 36246
rect 12992 36236 13044 36242
rect 12992 36178 13044 36184
rect 12900 35216 12952 35222
rect 12900 35158 12952 35164
rect 12716 33856 12768 33862
rect 12716 33798 12768 33804
rect 12716 33448 12768 33454
rect 12716 33390 12768 33396
rect 12728 33046 12756 33390
rect 12716 33040 12768 33046
rect 12716 32982 12768 32988
rect 12532 32972 12584 32978
rect 12532 32914 12584 32920
rect 12544 32434 12572 32914
rect 12532 32428 12584 32434
rect 12532 32370 12584 32376
rect 13004 30394 13032 36178
rect 13176 36168 13228 36174
rect 13174 36136 13176 36145
rect 13228 36136 13230 36145
rect 13174 36071 13230 36080
rect 13636 35624 13688 35630
rect 13636 35566 13688 35572
rect 13452 35556 13504 35562
rect 13452 35498 13504 35504
rect 13464 35154 13492 35498
rect 13452 35148 13504 35154
rect 13452 35090 13504 35096
rect 13084 34740 13136 34746
rect 13084 34682 13136 34688
rect 13096 34542 13124 34682
rect 13084 34536 13136 34542
rect 13084 34478 13136 34484
rect 13648 34406 13676 35566
rect 13740 34746 13768 37606
rect 13832 37262 13860 38694
rect 14096 38412 14148 38418
rect 14096 38354 14148 38360
rect 14108 38214 14136 38354
rect 14096 38208 14148 38214
rect 14096 38150 14148 38156
rect 14108 37738 14136 38150
rect 14096 37732 14148 37738
rect 14096 37674 14148 37680
rect 14554 37360 14610 37369
rect 14554 37295 14556 37304
rect 14608 37295 14610 37304
rect 14556 37266 14608 37272
rect 13820 37256 13872 37262
rect 13820 37198 13872 37204
rect 14016 36774 14320 36802
rect 14016 36718 14044 36774
rect 14004 36712 14056 36718
rect 14096 36712 14148 36718
rect 14004 36654 14056 36660
rect 14094 36680 14096 36689
rect 14148 36680 14150 36689
rect 14094 36615 14150 36624
rect 14292 36582 14320 36774
rect 14188 36576 14240 36582
rect 14188 36518 14240 36524
rect 14280 36576 14332 36582
rect 14280 36518 14332 36524
rect 13912 36236 13964 36242
rect 13912 36178 13964 36184
rect 13924 36038 13952 36178
rect 14200 36106 14228 36518
rect 14188 36100 14240 36106
rect 14188 36042 14240 36048
rect 13912 36032 13964 36038
rect 13912 35974 13964 35980
rect 13820 35488 13872 35494
rect 13820 35430 13872 35436
rect 13832 35222 13860 35430
rect 13924 35290 13952 35974
rect 14004 35692 14056 35698
rect 14004 35634 14056 35640
rect 14016 35494 14044 35634
rect 14004 35488 14056 35494
rect 14004 35430 14056 35436
rect 13912 35284 13964 35290
rect 13912 35226 13964 35232
rect 13820 35216 13872 35222
rect 13820 35158 13872 35164
rect 14016 35154 14044 35430
rect 14004 35148 14056 35154
rect 14004 35090 14056 35096
rect 13912 35012 13964 35018
rect 13912 34954 13964 34960
rect 13728 34740 13780 34746
rect 13728 34682 13780 34688
rect 13728 34536 13780 34542
rect 13728 34478 13780 34484
rect 13636 34400 13688 34406
rect 13636 34342 13688 34348
rect 13176 34060 13228 34066
rect 13176 34002 13228 34008
rect 13188 33046 13216 34002
rect 13648 33300 13676 34342
rect 13740 34134 13768 34478
rect 13728 34128 13780 34134
rect 13728 34070 13780 34076
rect 13924 34066 13952 34954
rect 13912 34060 13964 34066
rect 13912 34002 13964 34008
rect 13924 33862 13952 34002
rect 13912 33856 13964 33862
rect 13912 33798 13964 33804
rect 13728 33312 13780 33318
rect 13648 33272 13728 33300
rect 13728 33254 13780 33260
rect 13176 33040 13228 33046
rect 13176 32982 13228 32988
rect 13188 32230 13216 32982
rect 13176 32224 13228 32230
rect 13176 32166 13228 32172
rect 13176 32020 13228 32026
rect 13176 31962 13228 31968
rect 12992 30388 13044 30394
rect 12992 30330 13044 30336
rect 12452 29158 12572 29186
rect 12440 29096 12492 29102
rect 12440 29038 12492 29044
rect 11980 28008 12032 28014
rect 11980 27950 12032 27956
rect 11888 25356 11940 25362
rect 11888 25298 11940 25304
rect 11900 23186 11928 25298
rect 11992 25294 12020 27950
rect 12452 27577 12480 29038
rect 12544 27606 12572 29158
rect 12532 27600 12584 27606
rect 12438 27568 12494 27577
rect 12532 27542 12584 27548
rect 12438 27503 12494 27512
rect 12452 26518 12480 27503
rect 12544 27470 12572 27542
rect 12532 27464 12584 27470
rect 12532 27406 12584 27412
rect 12992 27464 13044 27470
rect 12992 27406 13044 27412
rect 12544 26586 12572 27406
rect 13004 27062 13032 27406
rect 13084 27328 13136 27334
rect 13084 27270 13136 27276
rect 12992 27056 13044 27062
rect 12992 26998 13044 27004
rect 12992 26920 13044 26926
rect 13096 26874 13124 27270
rect 13188 26926 13216 31962
rect 13740 28558 13768 33254
rect 13820 32768 13872 32774
rect 13820 32710 13872 32716
rect 13728 28552 13780 28558
rect 13728 28494 13780 28500
rect 13832 28218 13860 32710
rect 13820 28212 13872 28218
rect 13820 28154 13872 28160
rect 13044 26868 13124 26874
rect 12992 26862 13124 26868
rect 13176 26920 13228 26926
rect 13832 26874 13860 28154
rect 13176 26862 13228 26868
rect 12716 26852 12768 26858
rect 12716 26794 12768 26800
rect 13004 26846 13124 26862
rect 13648 26846 13860 26874
rect 12532 26580 12584 26586
rect 12532 26522 12584 26528
rect 12440 26512 12492 26518
rect 12440 26454 12492 26460
rect 12348 26444 12400 26450
rect 12348 26386 12400 26392
rect 11980 25288 12032 25294
rect 11980 25230 12032 25236
rect 12360 25226 12388 26386
rect 12440 26240 12492 26246
rect 12440 26182 12492 26188
rect 12452 26042 12480 26182
rect 12544 26042 12572 26522
rect 12440 26036 12492 26042
rect 12440 25978 12492 25984
rect 12532 26036 12584 26042
rect 12532 25978 12584 25984
rect 12440 25832 12492 25838
rect 12440 25774 12492 25780
rect 12348 25220 12400 25226
rect 12348 25162 12400 25168
rect 12360 24750 12388 25162
rect 12348 24744 12400 24750
rect 12348 24686 12400 24692
rect 12348 24404 12400 24410
rect 12348 24346 12400 24352
rect 12256 23860 12308 23866
rect 12256 23802 12308 23808
rect 12268 23730 12296 23802
rect 12256 23724 12308 23730
rect 12256 23666 12308 23672
rect 11888 23180 11940 23186
rect 11888 23122 11940 23128
rect 12072 22976 12124 22982
rect 12072 22918 12124 22924
rect 12084 17746 12112 22918
rect 12256 21888 12308 21894
rect 12256 21830 12308 21836
rect 12268 21350 12296 21830
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 12360 19378 12388 24346
rect 12452 23662 12480 25774
rect 12728 25294 12756 26794
rect 12716 25288 12768 25294
rect 12768 25248 12848 25276
rect 12716 25230 12768 25236
rect 12716 25152 12768 25158
rect 12716 25094 12768 25100
rect 12624 24744 12676 24750
rect 12624 24686 12676 24692
rect 12636 24614 12664 24686
rect 12532 24608 12584 24614
rect 12532 24550 12584 24556
rect 12624 24608 12676 24614
rect 12624 24550 12676 24556
rect 12440 23656 12492 23662
rect 12440 23598 12492 23604
rect 12544 23594 12572 24550
rect 12636 24070 12664 24550
rect 12728 24342 12756 25094
rect 12716 24336 12768 24342
rect 12716 24278 12768 24284
rect 12624 24064 12676 24070
rect 12624 24006 12676 24012
rect 12532 23588 12584 23594
rect 12532 23530 12584 23536
rect 12544 23118 12572 23530
rect 12636 23497 12664 24006
rect 12728 23866 12756 24278
rect 12716 23860 12768 23866
rect 12716 23802 12768 23808
rect 12820 23798 12848 25248
rect 12900 24064 12952 24070
rect 12900 24006 12952 24012
rect 12808 23792 12860 23798
rect 12728 23740 12808 23746
rect 12728 23734 12860 23740
rect 12728 23718 12848 23734
rect 12622 23488 12678 23497
rect 12622 23423 12678 23432
rect 12624 23248 12676 23254
rect 12624 23190 12676 23196
rect 12532 23112 12584 23118
rect 12532 23054 12584 23060
rect 12532 22636 12584 22642
rect 12532 22578 12584 22584
rect 12440 22500 12492 22506
rect 12440 22442 12492 22448
rect 12452 22098 12480 22442
rect 12440 22092 12492 22098
rect 12440 22034 12492 22040
rect 12440 21548 12492 21554
rect 12440 21490 12492 21496
rect 12452 20942 12480 21490
rect 12544 21418 12572 22578
rect 12636 22506 12664 23190
rect 12624 22500 12676 22506
rect 12624 22442 12676 22448
rect 12532 21412 12584 21418
rect 12532 21354 12584 21360
rect 12440 20936 12492 20942
rect 12440 20878 12492 20884
rect 12348 19372 12400 19378
rect 12348 19314 12400 19320
rect 12636 19310 12664 22442
rect 12728 22234 12756 23718
rect 12808 23656 12860 23662
rect 12808 23598 12860 23604
rect 12820 23186 12848 23598
rect 12808 23180 12860 23186
rect 12808 23122 12860 23128
rect 12820 22642 12848 23122
rect 12808 22636 12860 22642
rect 12808 22578 12860 22584
rect 12716 22228 12768 22234
rect 12716 22170 12768 22176
rect 12716 22024 12768 22030
rect 12716 21966 12768 21972
rect 12808 22024 12860 22030
rect 12808 21966 12860 21972
rect 12728 21554 12756 21966
rect 12716 21548 12768 21554
rect 12716 21490 12768 21496
rect 12716 21344 12768 21350
rect 12820 21332 12848 21966
rect 12768 21304 12848 21332
rect 12716 21286 12768 21292
rect 12728 19854 12756 21286
rect 12912 20806 12940 24006
rect 13004 23186 13032 26846
rect 13452 24676 13504 24682
rect 13452 24618 13504 24624
rect 13464 24410 13492 24618
rect 13544 24608 13596 24614
rect 13544 24550 13596 24556
rect 13556 24410 13584 24550
rect 13452 24404 13504 24410
rect 13452 24346 13504 24352
rect 13544 24404 13596 24410
rect 13544 24346 13596 24352
rect 13648 23730 13676 26846
rect 13728 26784 13780 26790
rect 13728 26726 13780 26732
rect 13740 26450 13768 26726
rect 13728 26444 13780 26450
rect 13728 26386 13780 26392
rect 13740 24614 13768 26386
rect 13820 26308 13872 26314
rect 13820 26250 13872 26256
rect 13832 25906 13860 26250
rect 13820 25900 13872 25906
rect 13820 25842 13872 25848
rect 13728 24608 13780 24614
rect 13728 24550 13780 24556
rect 13636 23724 13688 23730
rect 13636 23666 13688 23672
rect 12992 23180 13044 23186
rect 12992 23122 13044 23128
rect 13924 22778 13952 33798
rect 14292 32842 14320 36518
rect 15212 35766 15240 39918
rect 15568 39500 15620 39506
rect 15568 39442 15620 39448
rect 15474 37768 15530 37777
rect 15474 37703 15530 37712
rect 15200 35760 15252 35766
rect 15200 35702 15252 35708
rect 15212 35630 15240 35702
rect 15200 35624 15252 35630
rect 15200 35566 15252 35572
rect 15016 35284 15068 35290
rect 15016 35226 15068 35232
rect 14464 35148 14516 35154
rect 14464 35090 14516 35096
rect 14476 34746 14504 35090
rect 14648 35080 14700 35086
rect 14646 35048 14648 35057
rect 14700 35048 14702 35057
rect 14646 34983 14702 34992
rect 14464 34740 14516 34746
rect 14464 34682 14516 34688
rect 14372 34672 14424 34678
rect 14372 34614 14424 34620
rect 14384 34542 14412 34614
rect 14372 34536 14424 34542
rect 14372 34478 14424 34484
rect 14280 32836 14332 32842
rect 14280 32778 14332 32784
rect 14292 32026 14320 32778
rect 14280 32020 14332 32026
rect 14280 31962 14332 31968
rect 14292 31890 14320 31962
rect 14280 31884 14332 31890
rect 14280 31826 14332 31832
rect 14384 31278 14412 34478
rect 14464 32836 14516 32842
rect 14464 32778 14516 32784
rect 14476 32366 14504 32778
rect 14464 32360 14516 32366
rect 14464 32302 14516 32308
rect 14740 32292 14792 32298
rect 14740 32234 14792 32240
rect 14752 32026 14780 32234
rect 14740 32020 14792 32026
rect 14740 31962 14792 31968
rect 14372 31272 14424 31278
rect 14372 31214 14424 31220
rect 14004 30864 14056 30870
rect 14004 30806 14056 30812
rect 14016 29306 14044 30806
rect 14188 30796 14240 30802
rect 14188 30738 14240 30744
rect 14004 29300 14056 29306
rect 14004 29242 14056 29248
rect 14016 25906 14044 29242
rect 14004 25900 14056 25906
rect 14004 25842 14056 25848
rect 14200 25430 14228 30738
rect 14384 30598 14412 31214
rect 14372 30592 14424 30598
rect 14372 30534 14424 30540
rect 14384 29714 14412 30534
rect 14648 30048 14700 30054
rect 14648 29990 14700 29996
rect 14556 29844 14608 29850
rect 14556 29786 14608 29792
rect 14372 29708 14424 29714
rect 14372 29650 14424 29656
rect 14280 27872 14332 27878
rect 14280 27814 14332 27820
rect 14188 25424 14240 25430
rect 14188 25366 14240 25372
rect 13912 22772 13964 22778
rect 13912 22714 13964 22720
rect 13268 22160 13320 22166
rect 13268 22102 13320 22108
rect 12992 20936 13044 20942
rect 12992 20878 13044 20884
rect 12900 20800 12952 20806
rect 12900 20742 12952 20748
rect 13004 19990 13032 20878
rect 12992 19984 13044 19990
rect 12992 19926 13044 19932
rect 12716 19848 12768 19854
rect 12716 19790 12768 19796
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 12624 19304 12676 19310
rect 12624 19246 12676 19252
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12544 18358 12572 19110
rect 12636 18426 12664 19246
rect 12624 18420 12676 18426
rect 12624 18362 12676 18368
rect 12532 18352 12584 18358
rect 12532 18294 12584 18300
rect 12072 17740 12124 17746
rect 12072 17682 12124 17688
rect 12072 17604 12124 17610
rect 12072 17546 12124 17552
rect 11796 16720 11848 16726
rect 11796 16662 11848 16668
rect 11888 16584 11940 16590
rect 11888 16526 11940 16532
rect 11704 16516 11756 16522
rect 11704 16458 11756 16464
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 11256 14958 11284 15098
rect 11900 15026 11928 16526
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11244 14952 11296 14958
rect 11244 14894 11296 14900
rect 11152 14476 11204 14482
rect 11152 14418 11204 14424
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 10600 14000 10652 14006
rect 10980 13954 11008 14010
rect 10652 13948 11008 13954
rect 10600 13942 11008 13948
rect 10612 13926 11008 13942
rect 11704 13388 11756 13394
rect 11704 13330 11756 13336
rect 11716 12986 11744 13330
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11992 9382 12020 12378
rect 11980 9376 12032 9382
rect 11980 9318 12032 9324
rect 12084 9110 12112 17546
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12452 16522 12480 16934
rect 12440 16516 12492 16522
rect 12440 16458 12492 16464
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12544 14482 12572 15438
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 12176 10674 12204 13806
rect 12348 12640 12400 12646
rect 12348 12582 12400 12588
rect 12360 12238 12388 12582
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12164 10668 12216 10674
rect 12164 10610 12216 10616
rect 12256 10056 12308 10062
rect 12532 10056 12584 10062
rect 12308 10016 12388 10044
rect 12256 9998 12308 10004
rect 12360 9654 12388 10016
rect 12532 9998 12584 10004
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 12072 9104 12124 9110
rect 12072 9046 12124 9052
rect 12360 8974 12388 9590
rect 12544 9586 12572 9998
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 10980 7206 11008 8910
rect 12636 8906 12664 14962
rect 12728 13530 12756 19654
rect 13084 18216 13136 18222
rect 13084 18158 13136 18164
rect 12992 17876 13044 17882
rect 12992 17818 13044 17824
rect 13004 16590 13032 17818
rect 13096 17542 13124 18158
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 13096 16658 13124 17478
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 13280 15994 13308 22102
rect 14200 22098 14228 25366
rect 13820 22092 13872 22098
rect 13820 22034 13872 22040
rect 14188 22092 14240 22098
rect 14188 22034 14240 22040
rect 13832 20874 13860 22034
rect 14096 22024 14148 22030
rect 14096 21966 14148 21972
rect 14108 21894 14136 21966
rect 14096 21888 14148 21894
rect 14096 21830 14148 21836
rect 14108 21622 14136 21830
rect 14096 21616 14148 21622
rect 14096 21558 14148 21564
rect 13820 20868 13872 20874
rect 13820 20810 13872 20816
rect 13728 20800 13780 20806
rect 13728 20742 13780 20748
rect 13740 20466 13768 20742
rect 13728 20460 13780 20466
rect 13728 20402 13780 20408
rect 13832 19922 13860 20810
rect 13912 20392 13964 20398
rect 13912 20334 13964 20340
rect 13636 19916 13688 19922
rect 13636 19858 13688 19864
rect 13820 19916 13872 19922
rect 13820 19858 13872 19864
rect 13648 19242 13676 19858
rect 13832 19378 13860 19858
rect 13820 19372 13872 19378
rect 13820 19314 13872 19320
rect 13924 19310 13952 20334
rect 14200 19922 14228 22034
rect 14188 19916 14240 19922
rect 14188 19858 14240 19864
rect 14292 19802 14320 27814
rect 14464 23656 14516 23662
rect 14464 23598 14516 23604
rect 14476 22098 14504 23598
rect 14568 22420 14596 29786
rect 14660 29578 14688 29990
rect 15028 29646 15056 35226
rect 15292 34740 15344 34746
rect 15292 34682 15344 34688
rect 15304 34066 15332 34682
rect 15292 34060 15344 34066
rect 15292 34002 15344 34008
rect 15200 33448 15252 33454
rect 15200 33390 15252 33396
rect 15016 29640 15068 29646
rect 15016 29582 15068 29588
rect 14648 29572 14700 29578
rect 14648 29514 14700 29520
rect 15028 29510 15056 29582
rect 14924 29504 14976 29510
rect 14924 29446 14976 29452
rect 15016 29504 15068 29510
rect 15016 29446 15068 29452
rect 14740 28960 14792 28966
rect 14740 28902 14792 28908
rect 14752 28082 14780 28902
rect 14740 28076 14792 28082
rect 14740 28018 14792 28024
rect 14936 28014 14964 29446
rect 15028 29306 15056 29446
rect 15212 29306 15240 33390
rect 15292 32972 15344 32978
rect 15292 32914 15344 32920
rect 15304 31890 15332 32914
rect 15488 32774 15516 37703
rect 15580 36106 15608 39442
rect 15568 36100 15620 36106
rect 15568 36042 15620 36048
rect 15580 35630 15608 36042
rect 15568 35624 15620 35630
rect 15568 35566 15620 35572
rect 15672 34950 15700 42162
rect 16212 42152 16264 42158
rect 16212 42094 16264 42100
rect 16224 42022 16252 42094
rect 16776 42022 16804 42162
rect 16948 42084 17000 42090
rect 16948 42026 17000 42032
rect 16212 42016 16264 42022
rect 16212 41958 16264 41964
rect 16764 42016 16816 42022
rect 16764 41958 16816 41964
rect 16776 41818 16804 41958
rect 16960 41818 16988 42026
rect 17880 42022 17908 43862
rect 28264 43852 28316 43858
rect 28264 43794 28316 43800
rect 26240 43716 26292 43722
rect 26240 43658 26292 43664
rect 18420 43648 18472 43654
rect 18420 43590 18472 43596
rect 18432 43450 18460 43590
rect 18420 43444 18472 43450
rect 18420 43386 18472 43392
rect 18144 43104 18196 43110
rect 18144 43046 18196 43052
rect 18156 42242 18184 43046
rect 18328 42560 18380 42566
rect 18328 42502 18380 42508
rect 18064 42226 18184 42242
rect 18052 42220 18184 42226
rect 18104 42214 18184 42220
rect 18052 42162 18104 42168
rect 17868 42016 17920 42022
rect 17868 41958 17920 41964
rect 16764 41812 16816 41818
rect 16764 41754 16816 41760
rect 16948 41812 17000 41818
rect 16948 41754 17000 41760
rect 16776 41682 16804 41754
rect 16028 41676 16080 41682
rect 16028 41618 16080 41624
rect 16488 41676 16540 41682
rect 16488 41618 16540 41624
rect 16764 41676 16816 41682
rect 16764 41618 16816 41624
rect 16040 40526 16068 41618
rect 16500 41478 16528 41618
rect 16960 41614 16988 41754
rect 16948 41608 17000 41614
rect 16948 41550 17000 41556
rect 16488 41472 16540 41478
rect 16488 41414 16540 41420
rect 16028 40520 16080 40526
rect 16028 40462 16080 40468
rect 16040 39846 16068 40462
rect 16028 39840 16080 39846
rect 16028 39782 16080 39788
rect 16500 39642 16528 41414
rect 17880 40730 17908 41958
rect 18156 41546 18184 42214
rect 18340 42158 18368 42502
rect 18432 42226 18460 43386
rect 21180 43240 21232 43246
rect 21180 43182 21232 43188
rect 20168 43104 20220 43110
rect 20168 43046 20220 43052
rect 19580 43004 19876 43024
rect 19636 43002 19660 43004
rect 19716 43002 19740 43004
rect 19796 43002 19820 43004
rect 19658 42950 19660 43002
rect 19722 42950 19734 43002
rect 19796 42950 19798 43002
rect 19636 42948 19660 42950
rect 19716 42948 19740 42950
rect 19796 42948 19820 42950
rect 19580 42928 19876 42948
rect 18420 42220 18472 42226
rect 18420 42162 18472 42168
rect 18328 42152 18380 42158
rect 18328 42094 18380 42100
rect 20180 42022 20208 43046
rect 21192 42906 21220 43182
rect 21456 43104 21508 43110
rect 21456 43046 21508 43052
rect 22100 43104 22152 43110
rect 22100 43046 22152 43052
rect 21180 42900 21232 42906
rect 21180 42842 21232 42848
rect 20904 42696 20956 42702
rect 20904 42638 20956 42644
rect 20168 42016 20220 42022
rect 20168 41958 20220 41964
rect 19580 41916 19876 41936
rect 19636 41914 19660 41916
rect 19716 41914 19740 41916
rect 19796 41914 19820 41916
rect 19658 41862 19660 41914
rect 19722 41862 19734 41914
rect 19796 41862 19798 41914
rect 19636 41860 19660 41862
rect 19716 41860 19740 41862
rect 19796 41860 19820 41862
rect 19580 41840 19876 41860
rect 18144 41540 18196 41546
rect 18144 41482 18196 41488
rect 19340 41064 19392 41070
rect 19340 41006 19392 41012
rect 19984 41064 20036 41070
rect 19984 41006 20036 41012
rect 17868 40724 17920 40730
rect 17868 40666 17920 40672
rect 16580 40588 16632 40594
rect 16580 40530 16632 40536
rect 16488 39636 16540 39642
rect 16488 39578 16540 39584
rect 16028 38208 16080 38214
rect 16028 38150 16080 38156
rect 16040 37466 16068 38150
rect 16028 37460 16080 37466
rect 16028 37402 16080 37408
rect 15660 34944 15712 34950
rect 15660 34886 15712 34892
rect 16592 34542 16620 40530
rect 19352 39982 19380 41006
rect 19580 40828 19876 40848
rect 19636 40826 19660 40828
rect 19716 40826 19740 40828
rect 19796 40826 19820 40828
rect 19658 40774 19660 40826
rect 19722 40774 19734 40826
rect 19796 40774 19798 40826
rect 19636 40772 19660 40774
rect 19716 40772 19740 40774
rect 19796 40772 19820 40774
rect 19580 40752 19876 40772
rect 19340 39976 19392 39982
rect 19340 39918 19392 39924
rect 19062 39264 19118 39273
rect 19246 39264 19302 39273
rect 19118 39222 19246 39250
rect 19062 39199 19118 39208
rect 19246 39199 19302 39208
rect 19352 38978 19380 39918
rect 19580 39740 19876 39760
rect 19636 39738 19660 39740
rect 19716 39738 19740 39740
rect 19796 39738 19820 39740
rect 19658 39686 19660 39738
rect 19722 39686 19734 39738
rect 19796 39686 19798 39738
rect 19636 39684 19660 39686
rect 19716 39684 19740 39686
rect 19796 39684 19820 39686
rect 19580 39664 19876 39684
rect 19892 39296 19944 39302
rect 19892 39238 19944 39244
rect 19260 38950 19380 38978
rect 19260 38894 19288 38950
rect 19904 38894 19932 39238
rect 19248 38888 19300 38894
rect 19248 38830 19300 38836
rect 19432 38888 19484 38894
rect 19432 38830 19484 38836
rect 19892 38888 19944 38894
rect 19892 38830 19944 38836
rect 18696 38480 18748 38486
rect 19444 38457 19472 38830
rect 19580 38652 19876 38672
rect 19636 38650 19660 38652
rect 19716 38650 19740 38652
rect 19796 38650 19820 38652
rect 19658 38598 19660 38650
rect 19722 38598 19734 38650
rect 19796 38598 19798 38650
rect 19636 38596 19660 38598
rect 19716 38596 19740 38598
rect 19796 38596 19820 38598
rect 19580 38576 19876 38596
rect 18696 38422 18748 38428
rect 19430 38448 19486 38457
rect 18144 37800 18196 37806
rect 18142 37768 18144 37777
rect 18328 37800 18380 37806
rect 18196 37768 18198 37777
rect 18328 37742 18380 37748
rect 18142 37703 18198 37712
rect 18156 36038 18184 37703
rect 18340 37670 18368 37742
rect 18328 37664 18380 37670
rect 18328 37606 18380 37612
rect 18236 37324 18288 37330
rect 18236 37266 18288 37272
rect 18248 37126 18276 37266
rect 18236 37120 18288 37126
rect 18236 37062 18288 37068
rect 17316 36032 17368 36038
rect 17316 35974 17368 35980
rect 18144 36032 18196 36038
rect 18144 35974 18196 35980
rect 17328 34950 17356 35974
rect 17960 35692 18012 35698
rect 17960 35634 18012 35640
rect 17972 35034 18000 35634
rect 17972 35018 18184 35034
rect 17972 35012 18196 35018
rect 17972 35006 18144 35012
rect 18144 34954 18196 34960
rect 17316 34944 17368 34950
rect 17316 34886 17368 34892
rect 16580 34536 16632 34542
rect 16580 34478 16632 34484
rect 15660 34128 15712 34134
rect 15660 34070 15712 34076
rect 15476 32768 15528 32774
rect 15476 32710 15528 32716
rect 15476 32224 15528 32230
rect 15396 32184 15476 32212
rect 15292 31884 15344 31890
rect 15292 31826 15344 31832
rect 15396 31346 15424 32184
rect 15476 32166 15528 32172
rect 15568 32224 15620 32230
rect 15568 32166 15620 32172
rect 15580 32026 15608 32166
rect 15568 32020 15620 32026
rect 15568 31962 15620 31968
rect 15476 31884 15528 31890
rect 15476 31826 15528 31832
rect 15384 31340 15436 31346
rect 15384 31282 15436 31288
rect 15292 31136 15344 31142
rect 15292 31078 15344 31084
rect 15304 29714 15332 31078
rect 15488 30938 15516 31826
rect 15672 31498 15700 34070
rect 15844 33992 15896 33998
rect 15844 33934 15896 33940
rect 15580 31470 15700 31498
rect 15476 30932 15528 30938
rect 15476 30874 15528 30880
rect 15476 30184 15528 30190
rect 15476 30126 15528 30132
rect 15292 29708 15344 29714
rect 15292 29650 15344 29656
rect 15384 29708 15436 29714
rect 15384 29650 15436 29656
rect 15016 29300 15068 29306
rect 15016 29242 15068 29248
rect 15200 29300 15252 29306
rect 15200 29242 15252 29248
rect 15212 29102 15240 29242
rect 15200 29096 15252 29102
rect 15200 29038 15252 29044
rect 15212 28762 15240 29038
rect 15200 28756 15252 28762
rect 15200 28698 15252 28704
rect 15292 28620 15344 28626
rect 15292 28562 15344 28568
rect 14924 28008 14976 28014
rect 14924 27950 14976 27956
rect 15304 27878 15332 28562
rect 15396 28422 15424 29650
rect 15488 29238 15516 30126
rect 15476 29232 15528 29238
rect 15476 29174 15528 29180
rect 15384 28416 15436 28422
rect 15384 28358 15436 28364
rect 15292 27872 15344 27878
rect 15292 27814 15344 27820
rect 15292 26444 15344 26450
rect 15292 26386 15344 26392
rect 15304 26042 15332 26386
rect 15292 26036 15344 26042
rect 15292 25978 15344 25984
rect 14648 24608 14700 24614
rect 14648 24550 14700 24556
rect 14660 23662 14688 24550
rect 15580 24290 15608 31470
rect 15660 28416 15712 28422
rect 15660 28358 15712 28364
rect 15396 24262 15608 24290
rect 14648 23656 14700 23662
rect 14648 23598 14700 23604
rect 14660 22574 14688 23598
rect 14648 22568 14700 22574
rect 14648 22510 14700 22516
rect 14568 22392 14688 22420
rect 14464 22092 14516 22098
rect 14464 22034 14516 22040
rect 14476 21486 14504 22034
rect 14464 21480 14516 21486
rect 14464 21422 14516 21428
rect 14556 20936 14608 20942
rect 14556 20878 14608 20884
rect 14568 20058 14596 20878
rect 14556 20052 14608 20058
rect 14556 19994 14608 20000
rect 14016 19774 14320 19802
rect 13912 19304 13964 19310
rect 13912 19246 13964 19252
rect 13636 19236 13688 19242
rect 13636 19178 13688 19184
rect 13452 19168 13504 19174
rect 13452 19110 13504 19116
rect 12992 15972 13044 15978
rect 12992 15914 13044 15920
rect 13188 15966 13308 15994
rect 12808 15564 12860 15570
rect 12860 15524 12940 15552
rect 12808 15506 12860 15512
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12728 12850 12756 13126
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12912 11218 12940 15524
rect 13004 15502 13032 15914
rect 12992 15496 13044 15502
rect 12992 15438 13044 15444
rect 13084 15088 13136 15094
rect 13084 15030 13136 15036
rect 13096 14074 13124 15030
rect 13188 15026 13216 15966
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 13176 15020 13228 15026
rect 13176 14962 13228 14968
rect 13280 14657 13308 15846
rect 13360 15496 13412 15502
rect 13360 15438 13412 15444
rect 13266 14648 13322 14657
rect 13266 14583 13322 14592
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13096 12850 13124 14010
rect 13280 13938 13308 14583
rect 13372 14550 13400 15438
rect 13360 14544 13412 14550
rect 13360 14486 13412 14492
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 13084 12844 13136 12850
rect 13084 12786 13136 12792
rect 13464 12646 13492 19110
rect 14016 18834 14044 19774
rect 14568 19446 14596 19994
rect 14556 19440 14608 19446
rect 14556 19382 14608 19388
rect 14096 19304 14148 19310
rect 14096 19246 14148 19252
rect 14372 19304 14424 19310
rect 14372 19246 14424 19252
rect 14108 19174 14136 19246
rect 14096 19168 14148 19174
rect 14096 19110 14148 19116
rect 14384 18834 14412 19246
rect 13636 18828 13688 18834
rect 13636 18770 13688 18776
rect 14004 18828 14056 18834
rect 14004 18770 14056 18776
rect 14372 18828 14424 18834
rect 14372 18770 14424 18776
rect 13648 18290 13676 18770
rect 14004 18692 14056 18698
rect 14004 18634 14056 18640
rect 13636 18284 13688 18290
rect 13636 18226 13688 18232
rect 14016 18222 14044 18634
rect 14372 18624 14424 18630
rect 14372 18566 14424 18572
rect 14004 18216 14056 18222
rect 14004 18158 14056 18164
rect 14016 17882 14044 18158
rect 14096 18080 14148 18086
rect 14096 18022 14148 18028
rect 14004 17876 14056 17882
rect 14004 17818 14056 17824
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 13556 15570 13584 16526
rect 13820 15700 13872 15706
rect 13820 15642 13872 15648
rect 13544 15564 13596 15570
rect 13544 15506 13596 15512
rect 13556 14958 13584 15506
rect 13636 15496 13688 15502
rect 13636 15438 13688 15444
rect 13544 14952 13596 14958
rect 13544 14894 13596 14900
rect 13648 14498 13676 15438
rect 13832 15366 13860 15642
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 13912 14816 13964 14822
rect 13912 14758 13964 14764
rect 13556 14470 13676 14498
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 12716 11144 12768 11150
rect 12716 11086 12768 11092
rect 12728 10674 12756 11086
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12820 10810 12848 10950
rect 12912 10810 12940 11154
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12900 10804 12952 10810
rect 12900 10746 12952 10752
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 13556 10130 13584 14470
rect 13636 14408 13688 14414
rect 13636 14350 13688 14356
rect 13648 10266 13676 14350
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13728 11076 13780 11082
rect 13728 11018 13780 11024
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13544 10124 13596 10130
rect 13544 10066 13596 10072
rect 13648 9518 13676 10202
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13740 9382 13768 11018
rect 13832 9586 13860 11086
rect 13924 10130 13952 14758
rect 14004 13388 14056 13394
rect 14004 13330 14056 13336
rect 14016 12918 14044 13330
rect 14004 12912 14056 12918
rect 14004 12854 14056 12860
rect 14004 11212 14056 11218
rect 14004 11154 14056 11160
rect 14016 10810 14044 11154
rect 14004 10804 14056 10810
rect 14004 10746 14056 10752
rect 13912 10124 13964 10130
rect 13912 10066 13964 10072
rect 13912 9988 13964 9994
rect 13912 9930 13964 9936
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13832 9110 13860 9522
rect 13820 9104 13872 9110
rect 13820 9046 13872 9052
rect 12992 8968 13044 8974
rect 12992 8910 13044 8916
rect 12624 8900 12676 8906
rect 12624 8842 12676 8848
rect 13004 8498 13032 8910
rect 13832 8498 13860 9046
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13924 8294 13952 9930
rect 14004 9920 14056 9926
rect 14004 9862 14056 9868
rect 14016 9654 14044 9862
rect 14004 9648 14056 9654
rect 14004 9590 14056 9596
rect 14016 9042 14044 9590
rect 14108 9178 14136 18022
rect 14188 17536 14240 17542
rect 14188 17478 14240 17484
rect 14200 17202 14228 17478
rect 14188 17196 14240 17202
rect 14188 17138 14240 17144
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 14004 9036 14056 9042
rect 14004 8978 14056 8984
rect 14108 8430 14136 9114
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 10968 7200 11020 7206
rect 10968 7142 11020 7148
rect 10980 6866 11008 7142
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 12176 6798 12204 7890
rect 12912 7886 12940 8230
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 13636 7744 13688 7750
rect 13636 7686 13688 7692
rect 13648 7449 13676 7686
rect 13634 7440 13690 7449
rect 12808 7404 12860 7410
rect 13634 7375 13690 7384
rect 12808 7346 12860 7352
rect 11428 6792 11480 6798
rect 11428 6734 11480 6740
rect 12164 6792 12216 6798
rect 12164 6734 12216 6740
rect 11336 6656 11388 6662
rect 11336 6598 11388 6604
rect 10508 5024 10560 5030
rect 10508 4966 10560 4972
rect 10520 4690 10548 4966
rect 10508 4684 10560 4690
rect 10508 4626 10560 4632
rect 10520 3194 10548 4626
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11072 4282 11100 4558
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 11348 4078 11376 6598
rect 11440 5846 11468 6734
rect 11428 5840 11480 5846
rect 11428 5782 11480 5788
rect 12176 5778 12204 6734
rect 12820 6662 12848 7346
rect 13924 6866 13952 8230
rect 12992 6860 13044 6866
rect 12992 6802 13044 6808
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 13004 6662 13032 6802
rect 12808 6656 12860 6662
rect 12808 6598 12860 6604
rect 12992 6656 13044 6662
rect 12992 6598 13044 6604
rect 12164 5772 12216 5778
rect 12164 5714 12216 5720
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12544 4758 12572 5714
rect 12532 4752 12584 4758
rect 12532 4694 12584 4700
rect 13004 4554 13032 6598
rect 14016 5846 14044 8366
rect 14384 7546 14412 18566
rect 14660 15706 14688 22392
rect 15292 21004 15344 21010
rect 15292 20946 15344 20952
rect 15304 19922 15332 20946
rect 15396 20602 15424 24262
rect 15568 24200 15620 24206
rect 15568 24142 15620 24148
rect 15580 23866 15608 24142
rect 15568 23860 15620 23866
rect 15568 23802 15620 23808
rect 15672 21010 15700 28358
rect 15856 21894 15884 33934
rect 16396 32292 16448 32298
rect 16396 32234 16448 32240
rect 16408 31686 16436 32234
rect 16592 32026 16620 34478
rect 17132 32768 17184 32774
rect 17132 32710 17184 32716
rect 16948 32360 17000 32366
rect 16948 32302 17000 32308
rect 16580 32020 16632 32026
rect 16580 31962 16632 31968
rect 16856 32020 16908 32026
rect 16856 31962 16908 31968
rect 16592 31890 16620 31962
rect 16580 31884 16632 31890
rect 16580 31826 16632 31832
rect 16396 31680 16448 31686
rect 16396 31622 16448 31628
rect 16028 31272 16080 31278
rect 16028 31214 16080 31220
rect 16040 31142 16068 31214
rect 16028 31136 16080 31142
rect 16028 31078 16080 31084
rect 16212 31136 16264 31142
rect 16212 31078 16264 31084
rect 16224 30734 16252 31078
rect 16212 30728 16264 30734
rect 16212 30670 16264 30676
rect 16408 30122 16436 31622
rect 16488 30728 16540 30734
rect 16488 30670 16540 30676
rect 16500 30394 16528 30670
rect 16488 30388 16540 30394
rect 16488 30330 16540 30336
rect 16868 30326 16896 31962
rect 16960 31414 16988 32302
rect 17040 31816 17092 31822
rect 17040 31758 17092 31764
rect 17052 31686 17080 31758
rect 17040 31680 17092 31686
rect 17040 31622 17092 31628
rect 16948 31408 17000 31414
rect 16948 31350 17000 31356
rect 16856 30320 16908 30326
rect 16856 30262 16908 30268
rect 16488 30252 16540 30258
rect 16488 30194 16540 30200
rect 16396 30116 16448 30122
rect 16396 30058 16448 30064
rect 16304 30048 16356 30054
rect 16304 29990 16356 29996
rect 16316 27538 16344 29990
rect 16396 29572 16448 29578
rect 16396 29514 16448 29520
rect 16408 28422 16436 29514
rect 16396 28416 16448 28422
rect 16396 28358 16448 28364
rect 16408 28014 16436 28358
rect 16396 28008 16448 28014
rect 16396 27950 16448 27956
rect 16304 27532 16356 27538
rect 16304 27474 16356 27480
rect 16500 24750 16528 30194
rect 17144 29102 17172 32710
rect 17132 29096 17184 29102
rect 17132 29038 17184 29044
rect 16580 28620 16632 28626
rect 16580 28562 16632 28568
rect 16592 25362 16620 28562
rect 16580 25356 16632 25362
rect 16580 25298 16632 25304
rect 16488 24744 16540 24750
rect 16488 24686 16540 24692
rect 16500 24206 16528 24686
rect 16488 24200 16540 24206
rect 16488 24142 16540 24148
rect 16592 24138 16620 25298
rect 17040 24200 17092 24206
rect 17040 24142 17092 24148
rect 16580 24132 16632 24138
rect 16580 24074 16632 24080
rect 15844 21888 15896 21894
rect 15844 21830 15896 21836
rect 15660 21004 15712 21010
rect 15660 20946 15712 20952
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 14924 19916 14976 19922
rect 14924 19858 14976 19864
rect 15292 19916 15344 19922
rect 15292 19858 15344 19864
rect 14936 19378 14964 19858
rect 15396 19802 15424 20538
rect 15304 19774 15424 19802
rect 15304 19514 15332 19774
rect 15384 19712 15436 19718
rect 15384 19654 15436 19660
rect 15292 19508 15344 19514
rect 15292 19450 15344 19456
rect 14924 19372 14976 19378
rect 14924 19314 14976 19320
rect 15200 19304 15252 19310
rect 15304 19292 15332 19450
rect 15252 19264 15332 19292
rect 15200 19246 15252 19252
rect 15304 18426 15332 19264
rect 15396 18834 15424 19654
rect 15384 18828 15436 18834
rect 15384 18770 15436 18776
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15396 18222 15424 18770
rect 15856 18766 15884 21830
rect 16120 19236 16172 19242
rect 16120 19178 16172 19184
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15568 18624 15620 18630
rect 15568 18566 15620 18572
rect 15384 18216 15436 18222
rect 15384 18158 15436 18164
rect 15580 17338 15608 18566
rect 15936 17604 15988 17610
rect 15936 17546 15988 17552
rect 15948 17338 15976 17546
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15936 17332 15988 17338
rect 15936 17274 15988 17280
rect 14740 17128 14792 17134
rect 14740 17070 14792 17076
rect 15200 17128 15252 17134
rect 15200 17070 15252 17076
rect 14752 16794 14780 17070
rect 14740 16788 14792 16794
rect 14740 16730 14792 16736
rect 14648 15700 14700 15706
rect 14648 15642 14700 15648
rect 14752 14822 14780 16730
rect 15212 16046 15240 17070
rect 15568 16992 15620 16998
rect 15568 16934 15620 16940
rect 15200 16040 15252 16046
rect 15200 15982 15252 15988
rect 15108 15700 15160 15706
rect 15108 15642 15160 15648
rect 14924 14884 14976 14890
rect 14924 14826 14976 14832
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14936 14074 14964 14826
rect 14924 14068 14976 14074
rect 14924 14010 14976 14016
rect 14936 13394 14964 14010
rect 15120 13530 15148 15642
rect 15200 14952 15252 14958
rect 15200 14894 15252 14900
rect 15292 14952 15344 14958
rect 15292 14894 15344 14900
rect 15212 14482 15240 14894
rect 15304 14618 15332 14894
rect 15292 14612 15344 14618
rect 15292 14554 15344 14560
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15212 14006 15240 14418
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 15488 13938 15516 14214
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15396 10742 15424 13126
rect 15384 10736 15436 10742
rect 15384 10678 15436 10684
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15304 9042 15332 9318
rect 15292 9036 15344 9042
rect 15292 8978 15344 8984
rect 15396 7546 15424 10678
rect 15580 7954 15608 16934
rect 16132 15570 16160 19178
rect 16580 18896 16632 18902
rect 16580 18838 16632 18844
rect 16488 17264 16540 17270
rect 16488 17206 16540 17212
rect 16394 16008 16450 16017
rect 16394 15943 16450 15952
rect 16408 15706 16436 15943
rect 16396 15700 16448 15706
rect 16396 15642 16448 15648
rect 16408 15570 16436 15642
rect 16120 15564 16172 15570
rect 16120 15506 16172 15512
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 15752 15088 15804 15094
rect 15752 15030 15804 15036
rect 15764 14958 15792 15030
rect 15752 14952 15804 14958
rect 15752 14894 15804 14900
rect 15764 14618 15792 14894
rect 16120 14816 16172 14822
rect 16120 14758 16172 14764
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 15764 14414 15792 14554
rect 16132 14482 16160 14758
rect 16500 14618 16528 17206
rect 16592 16454 16620 18838
rect 16948 18148 17000 18154
rect 16948 18090 17000 18096
rect 16672 17604 16724 17610
rect 16672 17546 16724 17552
rect 16684 16658 16712 17546
rect 16960 16658 16988 18090
rect 17052 17134 17080 24142
rect 17144 21690 17172 29038
rect 17224 27532 17276 27538
rect 17224 27474 17276 27480
rect 17236 26790 17264 27474
rect 17224 26784 17276 26790
rect 17224 26726 17276 26732
rect 17236 25362 17264 26726
rect 17224 25356 17276 25362
rect 17224 25298 17276 25304
rect 17328 24410 17356 34886
rect 17776 34604 17828 34610
rect 17776 34546 17828 34552
rect 17500 33040 17552 33046
rect 17500 32982 17552 32988
rect 17512 29714 17540 32982
rect 17788 32026 17816 34546
rect 17960 34536 18012 34542
rect 17960 34478 18012 34484
rect 17972 32978 18000 34478
rect 18052 34196 18104 34202
rect 18052 34138 18104 34144
rect 18064 33833 18092 34138
rect 18050 33824 18106 33833
rect 18050 33759 18106 33768
rect 17960 32972 18012 32978
rect 17960 32914 18012 32920
rect 18052 32768 18104 32774
rect 18052 32710 18104 32716
rect 18064 32298 18092 32710
rect 18144 32360 18196 32366
rect 18144 32302 18196 32308
rect 18052 32292 18104 32298
rect 18052 32234 18104 32240
rect 18156 32026 18184 32302
rect 17776 32020 17828 32026
rect 17776 31962 17828 31968
rect 18144 32020 18196 32026
rect 18144 31962 18196 31968
rect 17696 31890 17816 31906
rect 17684 31884 17816 31890
rect 17736 31878 17816 31884
rect 17684 31826 17736 31832
rect 17788 31770 17816 31878
rect 17868 31816 17920 31822
rect 17788 31764 17868 31770
rect 17788 31758 17920 31764
rect 17788 31742 17908 31758
rect 17788 30598 17816 31742
rect 17960 30864 18012 30870
rect 17960 30806 18012 30812
rect 17592 30592 17644 30598
rect 17592 30534 17644 30540
rect 17776 30592 17828 30598
rect 17776 30534 17828 30540
rect 17500 29708 17552 29714
rect 17500 29650 17552 29656
rect 17316 24404 17368 24410
rect 17316 24346 17368 24352
rect 17132 21684 17184 21690
rect 17132 21626 17184 21632
rect 17604 18086 17632 30534
rect 17868 27328 17920 27334
rect 17868 27270 17920 27276
rect 17880 26450 17908 27270
rect 17868 26444 17920 26450
rect 17868 26386 17920 26392
rect 17776 23724 17828 23730
rect 17776 23666 17828 23672
rect 17788 23526 17816 23666
rect 17776 23520 17828 23526
rect 17776 23462 17828 23468
rect 17592 18080 17644 18086
rect 17592 18022 17644 18028
rect 17040 17128 17092 17134
rect 17040 17070 17092 17076
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 17236 16658 17264 16730
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16948 16652 17000 16658
rect 16948 16594 17000 16600
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 17592 16652 17644 16658
rect 17592 16594 17644 16600
rect 16580 16448 16632 16454
rect 16580 16390 16632 16396
rect 16592 15570 16620 16390
rect 17236 15978 17264 16594
rect 17224 15972 17276 15978
rect 17224 15914 17276 15920
rect 16580 15564 16632 15570
rect 16580 15506 16632 15512
rect 16488 14612 16540 14618
rect 16488 14554 16540 14560
rect 16120 14476 16172 14482
rect 16120 14418 16172 14424
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15764 12782 15792 13806
rect 16672 13796 16724 13802
rect 16672 13738 16724 13744
rect 16684 13394 16712 13738
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 15752 12776 15804 12782
rect 15752 12718 15804 12724
rect 16580 12776 16632 12782
rect 16580 12718 16632 12724
rect 16212 12640 16264 12646
rect 16212 12582 16264 12588
rect 16224 12306 16252 12582
rect 16212 12300 16264 12306
rect 16212 12242 16264 12248
rect 16120 12232 16172 12238
rect 16172 12180 16252 12186
rect 16120 12174 16252 12180
rect 16132 12158 16252 12174
rect 16224 11082 16252 12158
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 16408 11218 16436 12038
rect 16592 11898 16620 12718
rect 17328 12374 17356 16594
rect 17604 16454 17632 16594
rect 17592 16448 17644 16454
rect 17592 16390 17644 16396
rect 17788 14618 17816 23462
rect 17972 18834 18000 30806
rect 18144 30252 18196 30258
rect 18144 30194 18196 30200
rect 18052 22024 18104 22030
rect 18052 21966 18104 21972
rect 18064 19310 18092 21966
rect 18052 19304 18104 19310
rect 18052 19246 18104 19252
rect 18156 19258 18184 30194
rect 18248 26246 18276 37062
rect 18340 35154 18368 37606
rect 18420 37324 18472 37330
rect 18420 37266 18472 37272
rect 18432 36854 18460 37266
rect 18420 36848 18472 36854
rect 18420 36790 18472 36796
rect 18432 36242 18460 36790
rect 18420 36236 18472 36242
rect 18420 36178 18472 36184
rect 18328 35148 18380 35154
rect 18328 35090 18380 35096
rect 18328 33040 18380 33046
rect 18328 32982 18380 32988
rect 18340 31414 18368 32982
rect 18328 31408 18380 31414
rect 18328 31350 18380 31356
rect 18420 28552 18472 28558
rect 18420 28494 18472 28500
rect 18432 28422 18460 28494
rect 18420 28416 18472 28422
rect 18420 28358 18472 28364
rect 18432 28218 18460 28358
rect 18420 28212 18472 28218
rect 18420 28154 18472 28160
rect 18328 27532 18380 27538
rect 18328 27474 18380 27480
rect 18340 27062 18368 27474
rect 18328 27056 18380 27062
rect 18328 26998 18380 27004
rect 18708 26858 18736 38422
rect 18788 38412 18840 38418
rect 18788 38354 18840 38360
rect 19340 38412 19392 38418
rect 19430 38383 19486 38392
rect 19524 38412 19576 38418
rect 19340 38354 19392 38360
rect 19524 38354 19576 38360
rect 18800 37330 18828 38354
rect 19156 37800 19208 37806
rect 19352 37777 19380 38354
rect 19430 38312 19486 38321
rect 19430 38247 19486 38256
rect 19156 37742 19208 37748
rect 19338 37768 19394 37777
rect 19168 37346 19196 37742
rect 19338 37703 19394 37712
rect 19444 37466 19472 38247
rect 19536 38214 19564 38354
rect 19524 38208 19576 38214
rect 19524 38150 19576 38156
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 19432 37460 19484 37466
rect 19432 37402 19484 37408
rect 19168 37330 19840 37346
rect 18788 37324 18840 37330
rect 19168 37324 19852 37330
rect 19168 37318 19800 37324
rect 18788 37266 18840 37272
rect 19800 37266 19852 37272
rect 19338 37224 19394 37233
rect 19338 37159 19394 37168
rect 19352 36836 19380 37159
rect 19260 36825 19380 36836
rect 19246 36816 19380 36825
rect 19302 36808 19380 36816
rect 19246 36751 19302 36760
rect 18880 36712 18932 36718
rect 19064 36712 19116 36718
rect 18880 36654 18932 36660
rect 18970 36680 19026 36689
rect 18892 36106 18920 36654
rect 19064 36654 19116 36660
rect 19340 36712 19392 36718
rect 19904 36689 19932 38830
rect 19996 38486 20024 41006
rect 19984 38480 20036 38486
rect 19984 38422 20036 38428
rect 19984 37460 20036 37466
rect 19984 37402 20036 37408
rect 19996 37262 20024 37402
rect 19984 37256 20036 37262
rect 20180 37233 20208 41958
rect 20916 41614 20944 42638
rect 21192 42294 21220 42842
rect 21468 42702 21496 43046
rect 22008 42764 22060 42770
rect 22008 42706 22060 42712
rect 21456 42696 21508 42702
rect 21456 42638 21508 42644
rect 21916 42560 21968 42566
rect 21916 42502 21968 42508
rect 21928 42362 21956 42502
rect 21824 42356 21876 42362
rect 21824 42298 21876 42304
rect 21916 42356 21968 42362
rect 21916 42298 21968 42304
rect 21180 42288 21232 42294
rect 21180 42230 21232 42236
rect 21364 42288 21416 42294
rect 21836 42265 21864 42298
rect 21364 42230 21416 42236
rect 21822 42256 21878 42265
rect 21180 42016 21232 42022
rect 21180 41958 21232 41964
rect 21192 41682 21220 41958
rect 21180 41676 21232 41682
rect 21180 41618 21232 41624
rect 20904 41608 20956 41614
rect 20904 41550 20956 41556
rect 21376 41478 21404 42230
rect 21822 42191 21878 42200
rect 22020 42106 22048 42706
rect 21560 42090 22048 42106
rect 21548 42084 22048 42090
rect 21600 42078 22048 42084
rect 21548 42026 21600 42032
rect 22112 42022 22140 43046
rect 26056 42900 26108 42906
rect 26056 42842 26108 42848
rect 23848 42832 23900 42838
rect 23848 42774 23900 42780
rect 22560 42560 22612 42566
rect 22560 42502 22612 42508
rect 23112 42560 23164 42566
rect 23112 42502 23164 42508
rect 22572 42158 22600 42502
rect 22560 42152 22612 42158
rect 22560 42094 22612 42100
rect 21732 42016 21784 42022
rect 21732 41958 21784 41964
rect 22100 42016 22152 42022
rect 22100 41958 22152 41964
rect 22836 42016 22888 42022
rect 22836 41958 22888 41964
rect 20720 41472 20772 41478
rect 20720 41414 20772 41420
rect 21364 41472 21416 41478
rect 21364 41414 21416 41420
rect 20732 40730 20760 41414
rect 21640 40996 21692 41002
rect 21640 40938 21692 40944
rect 21456 40928 21508 40934
rect 21456 40870 21508 40876
rect 20720 40724 20772 40730
rect 20720 40666 20772 40672
rect 21468 40050 21496 40870
rect 21456 40044 21508 40050
rect 21456 39986 21508 39992
rect 21180 39976 21232 39982
rect 21180 39918 21232 39924
rect 20996 39908 21048 39914
rect 20996 39850 21048 39856
rect 21008 39574 21036 39850
rect 20996 39568 21048 39574
rect 20996 39510 21048 39516
rect 20720 39500 20772 39506
rect 20720 39442 20772 39448
rect 20732 39098 20760 39442
rect 20812 39296 20864 39302
rect 20812 39238 20864 39244
rect 20720 39092 20772 39098
rect 20720 39034 20772 39040
rect 20824 39030 20852 39238
rect 20812 39024 20864 39030
rect 20732 38972 20812 38978
rect 20732 38966 20864 38972
rect 20732 38950 20852 38966
rect 20352 38888 20404 38894
rect 20352 38830 20404 38836
rect 20364 38214 20392 38830
rect 20536 38548 20588 38554
rect 20536 38490 20588 38496
rect 20548 38214 20576 38490
rect 20352 38208 20404 38214
rect 20352 38150 20404 38156
rect 20536 38208 20588 38214
rect 20536 38150 20588 38156
rect 20364 37670 20392 38150
rect 20352 37664 20404 37670
rect 20352 37606 20404 37612
rect 20732 37466 20760 38950
rect 20824 38901 20852 38950
rect 20996 38752 21048 38758
rect 20996 38694 21048 38700
rect 21008 38486 21036 38694
rect 21192 38554 21220 39918
rect 21364 39840 21416 39846
rect 21364 39782 21416 39788
rect 21548 39840 21600 39846
rect 21548 39782 21600 39788
rect 21376 39098 21404 39782
rect 21560 39642 21588 39782
rect 21548 39636 21600 39642
rect 21548 39578 21600 39584
rect 21652 39273 21680 40938
rect 21744 40526 21772 41958
rect 21916 41540 21968 41546
rect 21916 41482 21968 41488
rect 21928 40730 21956 41482
rect 21916 40724 21968 40730
rect 21916 40666 21968 40672
rect 21928 40594 21956 40666
rect 22112 40594 22140 41958
rect 22284 41472 22336 41478
rect 22284 41414 22336 41420
rect 22296 41070 22324 41414
rect 22284 41064 22336 41070
rect 22284 41006 22336 41012
rect 22376 40928 22428 40934
rect 22376 40870 22428 40876
rect 22388 40594 22416 40870
rect 21916 40588 21968 40594
rect 21916 40530 21968 40536
rect 22100 40588 22152 40594
rect 22100 40530 22152 40536
rect 22376 40588 22428 40594
rect 22376 40530 22428 40536
rect 21732 40520 21784 40526
rect 21732 40462 21784 40468
rect 22112 40390 22140 40530
rect 22100 40384 22152 40390
rect 22100 40326 22152 40332
rect 21638 39264 21694 39273
rect 21638 39199 21694 39208
rect 21364 39092 21416 39098
rect 21364 39034 21416 39040
rect 21652 38894 21680 39199
rect 22008 39024 22060 39030
rect 22008 38966 22060 38972
rect 21640 38888 21692 38894
rect 21640 38830 21692 38836
rect 21180 38548 21232 38554
rect 21180 38490 21232 38496
rect 20996 38480 21048 38486
rect 20996 38422 21048 38428
rect 22020 38418 22048 38966
rect 22192 38548 22244 38554
rect 22192 38490 22244 38496
rect 21088 38412 21140 38418
rect 21732 38412 21784 38418
rect 21088 38354 21140 38360
rect 21652 38372 21732 38400
rect 20812 37800 20864 37806
rect 20812 37742 20864 37748
rect 20824 37466 20852 37742
rect 20720 37460 20772 37466
rect 20720 37402 20772 37408
rect 20812 37460 20864 37466
rect 20812 37402 20864 37408
rect 20824 37318 21036 37346
rect 21100 37330 21128 38354
rect 21178 37904 21234 37913
rect 21178 37839 21180 37848
rect 21232 37839 21234 37848
rect 21180 37810 21232 37816
rect 21652 37670 21680 38372
rect 21732 38354 21784 38360
rect 22008 38412 22060 38418
rect 22008 38354 22060 38360
rect 22204 37913 22232 38490
rect 22190 37904 22246 37913
rect 22190 37839 22246 37848
rect 21640 37664 21692 37670
rect 21640 37606 21692 37612
rect 21824 37664 21876 37670
rect 21824 37606 21876 37612
rect 21836 37330 21864 37606
rect 19984 37198 20036 37204
rect 20166 37224 20222 37233
rect 20824 37194 20852 37318
rect 20904 37256 20956 37262
rect 20904 37198 20956 37204
rect 20166 37159 20222 37168
rect 20812 37188 20864 37194
rect 20812 37130 20864 37136
rect 20916 37126 20944 37198
rect 21008 37126 21036 37318
rect 21088 37324 21140 37330
rect 21088 37266 21140 37272
rect 21824 37324 21876 37330
rect 21824 37266 21876 37272
rect 22284 37188 22336 37194
rect 22284 37130 22336 37136
rect 20904 37120 20956 37126
rect 20904 37062 20956 37068
rect 20996 37120 21048 37126
rect 20996 37062 21048 37068
rect 22296 36718 22324 37130
rect 22284 36712 22336 36718
rect 19340 36654 19392 36660
rect 19890 36680 19946 36689
rect 18970 36615 18972 36624
rect 19024 36615 19026 36624
rect 18972 36586 19024 36592
rect 18788 36100 18840 36106
rect 18788 36042 18840 36048
rect 18880 36100 18932 36106
rect 18880 36042 18932 36048
rect 18800 35698 18828 36042
rect 18788 35692 18840 35698
rect 18788 35634 18840 35640
rect 19076 35630 19104 36654
rect 19248 36032 19300 36038
rect 19248 35974 19300 35980
rect 19064 35624 19116 35630
rect 19064 35566 19116 35572
rect 19156 35556 19208 35562
rect 19156 35498 19208 35504
rect 19168 35290 19196 35498
rect 19156 35284 19208 35290
rect 19156 35226 19208 35232
rect 18788 34944 18840 34950
rect 18788 34886 18840 34892
rect 18800 34746 18828 34886
rect 18788 34740 18840 34746
rect 18788 34682 18840 34688
rect 19260 32774 19288 35974
rect 19352 35290 19380 36654
rect 22284 36654 22336 36660
rect 19890 36615 19946 36624
rect 20076 36644 20128 36650
rect 20076 36586 20128 36592
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19580 36400 19876 36420
rect 20088 36038 20116 36586
rect 20628 36576 20680 36582
rect 20628 36518 20680 36524
rect 20166 36272 20222 36281
rect 20166 36207 20222 36216
rect 20180 36106 20208 36207
rect 20168 36100 20220 36106
rect 20168 36042 20220 36048
rect 20076 36032 20128 36038
rect 20076 35974 20128 35980
rect 19984 35624 20036 35630
rect 19984 35566 20036 35572
rect 19996 35494 20024 35566
rect 19432 35488 19484 35494
rect 19432 35430 19484 35436
rect 19984 35488 20036 35494
rect 19984 35430 20036 35436
rect 19340 35284 19392 35290
rect 19340 35226 19392 35232
rect 19444 34746 19472 35430
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 19708 35216 19760 35222
rect 19706 35184 19708 35193
rect 19760 35184 19762 35193
rect 19706 35119 19762 35128
rect 19432 34740 19484 34746
rect 19432 34682 19484 34688
rect 20074 34640 20130 34649
rect 20074 34575 20076 34584
rect 20128 34575 20130 34584
rect 20076 34546 20128 34552
rect 19984 34536 20036 34542
rect 19984 34478 20036 34484
rect 19996 34406 20024 34478
rect 19984 34400 20036 34406
rect 19984 34342 20036 34348
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 19996 33862 20024 34342
rect 20180 34066 20208 36042
rect 20640 35630 20668 36518
rect 20904 36236 20956 36242
rect 20904 36178 20956 36184
rect 20720 36168 20772 36174
rect 20720 36110 20772 36116
rect 20732 35766 20760 36110
rect 20916 35834 20944 36178
rect 20904 35828 20956 35834
rect 20904 35770 20956 35776
rect 20720 35760 20772 35766
rect 20720 35702 20772 35708
rect 20628 35624 20680 35630
rect 20628 35566 20680 35572
rect 20732 35290 20760 35702
rect 21824 35488 21876 35494
rect 21824 35430 21876 35436
rect 20720 35284 20772 35290
rect 20720 35226 20772 35232
rect 21836 35154 21864 35430
rect 22192 35284 22244 35290
rect 22192 35226 22244 35232
rect 21824 35148 21876 35154
rect 21876 35108 22048 35136
rect 21824 35090 21876 35096
rect 21270 34776 21326 34785
rect 21180 34740 21232 34746
rect 21270 34711 21326 34720
rect 21180 34682 21232 34688
rect 21192 34542 21220 34682
rect 21284 34542 21312 34711
rect 20352 34536 20404 34542
rect 20352 34478 20404 34484
rect 21180 34536 21232 34542
rect 21180 34478 21232 34484
rect 21272 34536 21324 34542
rect 21272 34478 21324 34484
rect 20364 34406 20392 34478
rect 21192 34406 21220 34478
rect 20352 34400 20404 34406
rect 20352 34342 20404 34348
rect 21180 34400 21232 34406
rect 21180 34342 21232 34348
rect 20168 34060 20220 34066
rect 20168 34002 20220 34008
rect 19984 33856 20036 33862
rect 19984 33798 20036 33804
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 19616 32972 19668 32978
rect 19616 32914 19668 32920
rect 19248 32768 19300 32774
rect 19248 32710 19300 32716
rect 19628 32434 19656 32914
rect 19892 32768 19944 32774
rect 19892 32710 19944 32716
rect 19904 32502 19932 32710
rect 19892 32496 19944 32502
rect 19892 32438 19944 32444
rect 19616 32428 19668 32434
rect 19616 32370 19668 32376
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 19340 29096 19392 29102
rect 19340 29038 19392 29044
rect 19352 28626 19380 29038
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 19892 28688 19944 28694
rect 19522 28656 19578 28665
rect 19340 28620 19392 28626
rect 19892 28630 19944 28636
rect 19522 28591 19524 28600
rect 19340 28562 19392 28568
rect 19576 28591 19578 28600
rect 19524 28562 19576 28568
rect 19248 26920 19300 26926
rect 19248 26862 19300 26868
rect 18696 26852 18748 26858
rect 18696 26794 18748 26800
rect 19260 26518 19288 26862
rect 19248 26512 19300 26518
rect 19248 26454 19300 26460
rect 19352 26450 19380 28562
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19580 27696 19876 27716
rect 19904 27062 19932 28630
rect 19892 27056 19944 27062
rect 19892 26998 19944 27004
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 19340 26444 19392 26450
rect 19340 26386 19392 26392
rect 19432 26376 19484 26382
rect 19432 26318 19484 26324
rect 18236 26240 18288 26246
rect 18236 26182 18288 26188
rect 19444 25838 19472 26318
rect 19432 25832 19484 25838
rect 19432 25774 19484 25780
rect 19892 25832 19944 25838
rect 19892 25774 19944 25780
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 19904 25430 19932 25774
rect 19892 25424 19944 25430
rect 19892 25366 19944 25372
rect 19340 24608 19392 24614
rect 19340 24550 19392 24556
rect 18328 24336 18380 24342
rect 18328 24278 18380 24284
rect 18340 22234 18368 24278
rect 18420 24268 18472 24274
rect 18420 24210 18472 24216
rect 18432 22506 18460 24210
rect 18880 24200 18932 24206
rect 18880 24142 18932 24148
rect 18788 23860 18840 23866
rect 18788 23802 18840 23808
rect 18604 23588 18656 23594
rect 18604 23530 18656 23536
rect 18420 22500 18472 22506
rect 18420 22442 18472 22448
rect 18328 22228 18380 22234
rect 18328 22170 18380 22176
rect 18432 22098 18460 22442
rect 18420 22092 18472 22098
rect 18420 22034 18472 22040
rect 18616 21486 18644 23530
rect 18696 22160 18748 22166
rect 18696 22102 18748 22108
rect 18604 21480 18656 21486
rect 18604 21422 18656 21428
rect 18156 19230 18368 19258
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 17960 18828 18012 18834
rect 17960 18770 18012 18776
rect 18052 18828 18104 18834
rect 18052 18770 18104 18776
rect 18064 18222 18092 18770
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 18064 17746 18092 18158
rect 18052 17740 18104 17746
rect 18052 17682 18104 17688
rect 18156 17202 18184 19110
rect 18236 18624 18288 18630
rect 18236 18566 18288 18572
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 18248 17134 18276 18566
rect 18340 17678 18368 19230
rect 18708 18426 18736 22102
rect 18800 21350 18828 23802
rect 18892 23662 18920 24142
rect 18880 23656 18932 23662
rect 18880 23598 18932 23604
rect 19248 23520 19300 23526
rect 19248 23462 19300 23468
rect 19260 23186 19288 23462
rect 19248 23180 19300 23186
rect 19248 23122 19300 23128
rect 19064 22024 19116 22030
rect 19064 21966 19116 21972
rect 19076 21486 19104 21966
rect 19156 21888 19208 21894
rect 19156 21830 19208 21836
rect 19168 21486 19196 21830
rect 19064 21480 19116 21486
rect 19064 21422 19116 21428
rect 19156 21480 19208 21486
rect 19156 21422 19208 21428
rect 18788 21344 18840 21350
rect 18788 21286 18840 21292
rect 18696 18420 18748 18426
rect 18696 18362 18748 18368
rect 18708 18154 18736 18362
rect 18696 18148 18748 18154
rect 18696 18090 18748 18096
rect 18328 17672 18380 17678
rect 18328 17614 18380 17620
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18236 17128 18288 17134
rect 18236 17070 18288 17076
rect 18052 16992 18104 16998
rect 18052 16934 18104 16940
rect 17960 16584 18012 16590
rect 17960 16526 18012 16532
rect 17868 15904 17920 15910
rect 17868 15846 17920 15852
rect 17776 14612 17828 14618
rect 17776 14554 17828 14560
rect 17316 12368 17368 12374
rect 17316 12310 17368 12316
rect 17328 11898 17356 12310
rect 16580 11892 16632 11898
rect 16580 11834 16632 11840
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 16396 11212 16448 11218
rect 16396 11154 16448 11160
rect 16212 11076 16264 11082
rect 16212 11018 16264 11024
rect 16224 10470 16252 11018
rect 16580 11008 16632 11014
rect 16580 10950 16632 10956
rect 16592 10742 16620 10950
rect 17788 10742 17816 14554
rect 16580 10736 16632 10742
rect 16580 10678 16632 10684
rect 17776 10736 17828 10742
rect 17776 10678 17828 10684
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16224 9926 16252 10406
rect 16212 9920 16264 9926
rect 16212 9862 16264 9868
rect 16212 8560 16264 8566
rect 16212 8502 16264 8508
rect 15476 7948 15528 7954
rect 15476 7890 15528 7896
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 15108 7540 15160 7546
rect 15108 7482 15160 7488
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15120 7002 15148 7482
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 15304 6934 15332 7278
rect 15292 6928 15344 6934
rect 15292 6870 15344 6876
rect 15108 6724 15160 6730
rect 15108 6666 15160 6672
rect 15120 6254 15148 6666
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 15120 5846 15148 6190
rect 15396 5914 15424 7482
rect 15488 6866 15516 7890
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 16224 6798 16252 8502
rect 17880 8090 17908 15846
rect 17972 12442 18000 16526
rect 18064 16114 18092 16934
rect 18328 16720 18380 16726
rect 18328 16662 18380 16668
rect 18052 16108 18104 16114
rect 18052 16050 18104 16056
rect 18340 14006 18368 16662
rect 18432 16046 18460 17478
rect 18604 17128 18656 17134
rect 18604 17070 18656 17076
rect 18510 16688 18566 16697
rect 18510 16623 18512 16632
rect 18564 16623 18566 16632
rect 18512 16594 18564 16600
rect 18616 16046 18644 17070
rect 18420 16040 18472 16046
rect 18420 15982 18472 15988
rect 18604 16040 18656 16046
rect 18604 15982 18656 15988
rect 18800 14278 18828 21286
rect 19154 17368 19210 17377
rect 19154 17303 19210 17312
rect 19168 17202 19196 17303
rect 19156 17196 19208 17202
rect 19156 17138 19208 17144
rect 19064 17128 19116 17134
rect 19064 17070 19116 17076
rect 18972 17060 19024 17066
rect 18972 17002 19024 17008
rect 18984 16658 19012 17002
rect 19076 16998 19104 17070
rect 19064 16992 19116 16998
rect 19064 16934 19116 16940
rect 18972 16652 19024 16658
rect 18972 16594 19024 16600
rect 18984 16046 19012 16594
rect 19076 16454 19104 16934
rect 19064 16448 19116 16454
rect 19064 16390 19116 16396
rect 18972 16040 19024 16046
rect 18972 15982 19024 15988
rect 18788 14272 18840 14278
rect 18788 14214 18840 14220
rect 19168 14074 19196 17138
rect 19352 14074 19380 24550
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 19616 23112 19668 23118
rect 19616 23054 19668 23060
rect 19628 22642 19656 23054
rect 19616 22636 19668 22642
rect 19616 22578 19668 22584
rect 19892 22568 19944 22574
rect 19892 22510 19944 22516
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 19904 21690 19932 22510
rect 19892 21684 19944 21690
rect 19892 21626 19944 21632
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 19996 20602 20024 33798
rect 20364 33522 20392 34342
rect 21180 34128 21232 34134
rect 21178 34096 21180 34105
rect 21232 34096 21234 34105
rect 21178 34031 21234 34040
rect 21284 34066 21496 34082
rect 21284 34060 21508 34066
rect 21284 34054 21456 34060
rect 21284 33998 21312 34054
rect 21456 34002 21508 34008
rect 22020 33998 22048 35108
rect 22100 35080 22152 35086
rect 22100 35022 22152 35028
rect 22112 34746 22140 35022
rect 22100 34740 22152 34746
rect 22100 34682 22152 34688
rect 22204 34678 22232 35226
rect 22376 35148 22428 35154
rect 22376 35090 22428 35096
rect 22284 35080 22336 35086
rect 22284 35022 22336 35028
rect 22296 34950 22324 35022
rect 22284 34944 22336 34950
rect 22284 34886 22336 34892
rect 22282 34776 22338 34785
rect 22282 34711 22284 34720
rect 22336 34711 22338 34720
rect 22284 34682 22336 34688
rect 22192 34672 22244 34678
rect 22192 34614 22244 34620
rect 21272 33992 21324 33998
rect 20442 33960 20498 33969
rect 21272 33934 21324 33940
rect 21364 33992 21416 33998
rect 21364 33934 21416 33940
rect 22008 33992 22060 33998
rect 22008 33934 22060 33940
rect 20442 33895 20444 33904
rect 20496 33895 20498 33904
rect 20444 33866 20496 33872
rect 21270 33552 21326 33561
rect 20352 33516 20404 33522
rect 21270 33487 21326 33496
rect 20352 33458 20404 33464
rect 20364 33386 20392 33458
rect 21284 33454 21312 33487
rect 20996 33448 21048 33454
rect 20994 33416 20996 33425
rect 21272 33448 21324 33454
rect 21048 33416 21050 33425
rect 20352 33380 20404 33386
rect 20352 33322 20404 33328
rect 20812 33380 20864 33386
rect 21272 33390 21324 33396
rect 20994 33351 21050 33360
rect 20812 33322 20864 33328
rect 20260 32224 20312 32230
rect 20260 32166 20312 32172
rect 20272 32026 20300 32166
rect 20260 32020 20312 32026
rect 20260 31962 20312 31968
rect 20076 31340 20128 31346
rect 20076 31282 20128 31288
rect 20088 22234 20116 31282
rect 20168 31272 20220 31278
rect 20168 31214 20220 31220
rect 20180 30938 20208 31214
rect 20168 30932 20220 30938
rect 20168 30874 20220 30880
rect 20180 28694 20208 30874
rect 20272 30054 20300 31962
rect 20260 30048 20312 30054
rect 20260 29990 20312 29996
rect 20168 28688 20220 28694
rect 20168 28630 20220 28636
rect 20272 28540 20300 29990
rect 20364 28694 20392 33322
rect 20824 32502 20852 33322
rect 21376 33318 21404 33934
rect 21732 33856 21784 33862
rect 21732 33798 21784 33804
rect 21640 33652 21692 33658
rect 21640 33594 21692 33600
rect 21652 33522 21680 33594
rect 21640 33516 21692 33522
rect 21640 33458 21692 33464
rect 21548 33448 21600 33454
rect 21548 33390 21600 33396
rect 21272 33312 21324 33318
rect 21272 33254 21324 33260
rect 21364 33312 21416 33318
rect 21364 33254 21416 33260
rect 21284 33130 21312 33254
rect 21560 33130 21588 33390
rect 21744 33386 21772 33798
rect 22192 33652 22244 33658
rect 22192 33594 22244 33600
rect 22204 33561 22232 33594
rect 22190 33552 22246 33561
rect 22190 33487 22246 33496
rect 22388 33425 22416 35090
rect 22848 35086 22876 41958
rect 23124 41478 23152 42502
rect 23112 41472 23164 41478
rect 23112 41414 23164 41420
rect 23860 40186 23888 42774
rect 24768 42764 24820 42770
rect 24768 42706 24820 42712
rect 24780 42566 24808 42706
rect 24032 42560 24084 42566
rect 24032 42502 24084 42508
rect 24768 42560 24820 42566
rect 24768 42502 24820 42508
rect 24044 42158 24072 42502
rect 26068 42158 26096 42842
rect 26252 42702 26280 43658
rect 27160 43308 27212 43314
rect 27160 43250 27212 43256
rect 26700 43104 26752 43110
rect 26700 43046 26752 43052
rect 26712 42702 26740 43046
rect 26240 42696 26292 42702
rect 26240 42638 26292 42644
rect 26700 42696 26752 42702
rect 26700 42638 26752 42644
rect 24032 42152 24084 42158
rect 24032 42094 24084 42100
rect 26056 42152 26108 42158
rect 26056 42094 26108 42100
rect 23848 40180 23900 40186
rect 23848 40122 23900 40128
rect 24044 38214 24072 42094
rect 25688 42016 25740 42022
rect 25688 41958 25740 41964
rect 25780 42016 25832 42022
rect 25780 41958 25832 41964
rect 25700 41682 25728 41958
rect 25792 41750 25820 41958
rect 25780 41744 25832 41750
rect 25780 41686 25832 41692
rect 25044 41676 25096 41682
rect 25044 41618 25096 41624
rect 25688 41676 25740 41682
rect 25688 41618 25740 41624
rect 24860 41064 24912 41070
rect 24860 41006 24912 41012
rect 24872 40934 24900 41006
rect 25056 40934 25084 41618
rect 26068 41206 26096 42094
rect 26252 41834 26280 42638
rect 27172 42226 27200 43250
rect 28276 42906 28304 43794
rect 43628 43784 43680 43790
rect 43628 43726 43680 43732
rect 44456 43784 44508 43790
rect 44508 43744 44588 43772
rect 44456 43726 44508 43732
rect 34940 43548 35236 43568
rect 34996 43546 35020 43548
rect 35076 43546 35100 43548
rect 35156 43546 35180 43548
rect 35018 43494 35020 43546
rect 35082 43494 35094 43546
rect 35156 43494 35158 43546
rect 34996 43492 35020 43494
rect 35076 43492 35100 43494
rect 35156 43492 35180 43494
rect 34940 43472 35236 43492
rect 38844 43308 38896 43314
rect 38844 43250 38896 43256
rect 40040 43308 40092 43314
rect 40040 43250 40092 43256
rect 33232 43240 33284 43246
rect 33232 43182 33284 43188
rect 33968 43240 34020 43246
rect 33968 43182 34020 43188
rect 29184 43172 29236 43178
rect 29184 43114 29236 43120
rect 28448 43104 28500 43110
rect 28448 43046 28500 43052
rect 28264 42900 28316 42906
rect 28264 42842 28316 42848
rect 27896 42628 27948 42634
rect 27896 42570 27948 42576
rect 27160 42220 27212 42226
rect 27160 42162 27212 42168
rect 26608 42152 26660 42158
rect 26608 42094 26660 42100
rect 26700 42152 26752 42158
rect 26700 42094 26752 42100
rect 26620 42022 26648 42094
rect 26608 42016 26660 42022
rect 26608 41958 26660 41964
rect 26252 41806 26372 41834
rect 26148 41676 26200 41682
rect 26148 41618 26200 41624
rect 26056 41200 26108 41206
rect 26056 41142 26108 41148
rect 26160 41070 26188 41618
rect 26344 41614 26372 41806
rect 26712 41750 26740 42094
rect 27908 41818 27936 42570
rect 28460 42566 28488 43046
rect 29196 42770 29224 43114
rect 33244 43110 33272 43182
rect 31944 43104 31996 43110
rect 31944 43046 31996 43052
rect 32312 43104 32364 43110
rect 32312 43046 32364 43052
rect 33232 43104 33284 43110
rect 33232 43046 33284 43052
rect 29368 42900 29420 42906
rect 29368 42842 29420 42848
rect 29380 42809 29408 42842
rect 29366 42800 29422 42809
rect 29184 42764 29236 42770
rect 29184 42706 29236 42712
rect 29276 42764 29328 42770
rect 29366 42735 29422 42744
rect 29276 42706 29328 42712
rect 28448 42560 28500 42566
rect 28448 42502 28500 42508
rect 28170 42256 28226 42265
rect 28170 42191 28226 42200
rect 27896 41812 27948 41818
rect 27896 41754 27948 41760
rect 26700 41744 26752 41750
rect 26700 41686 26752 41692
rect 27908 41682 27936 41754
rect 28184 41750 28212 42191
rect 28172 41744 28224 41750
rect 28172 41686 28224 41692
rect 27344 41676 27396 41682
rect 27344 41618 27396 41624
rect 27896 41676 27948 41682
rect 27896 41618 27948 41624
rect 26332 41608 26384 41614
rect 26332 41550 26384 41556
rect 26240 41540 26292 41546
rect 26240 41482 26292 41488
rect 27160 41540 27212 41546
rect 27356 41528 27384 41618
rect 27212 41500 27384 41528
rect 27160 41482 27212 41488
rect 26252 41206 26280 41482
rect 26240 41200 26292 41206
rect 26240 41142 26292 41148
rect 26712 41138 27016 41154
rect 26700 41132 27028 41138
rect 26752 41126 26976 41132
rect 26700 41074 26752 41080
rect 26976 41074 27028 41080
rect 27264 41070 27292 41500
rect 27804 41200 27856 41206
rect 27540 41126 27752 41154
rect 27804 41142 27856 41148
rect 26148 41064 26200 41070
rect 26148 41006 26200 41012
rect 27252 41064 27304 41070
rect 27252 41006 27304 41012
rect 26160 40934 26188 41006
rect 24860 40928 24912 40934
rect 24860 40870 24912 40876
rect 25044 40928 25096 40934
rect 25044 40870 25096 40876
rect 26148 40928 26200 40934
rect 26148 40870 26200 40876
rect 26332 40928 26384 40934
rect 26332 40870 26384 40876
rect 26424 40928 26476 40934
rect 26424 40870 26476 40876
rect 27436 40928 27488 40934
rect 27540 40916 27568 41126
rect 27724 41070 27752 41126
rect 27620 41064 27672 41070
rect 27620 41006 27672 41012
rect 27712 41064 27764 41070
rect 27712 41006 27764 41012
rect 27632 40934 27660 41006
rect 27816 40934 27844 41142
rect 27488 40888 27568 40916
rect 27620 40928 27672 40934
rect 27436 40870 27488 40876
rect 27620 40870 27672 40876
rect 27804 40928 27856 40934
rect 27804 40870 27856 40876
rect 24124 39636 24176 39642
rect 24124 39578 24176 39584
rect 24136 38962 24164 39578
rect 24124 38956 24176 38962
rect 24124 38898 24176 38904
rect 24308 38412 24360 38418
rect 24308 38354 24360 38360
rect 24032 38208 24084 38214
rect 24032 38150 24084 38156
rect 23400 37806 23428 37837
rect 23388 37800 23440 37806
rect 23386 37768 23388 37777
rect 23440 37768 23442 37777
rect 23386 37703 23442 37712
rect 23400 37466 23428 37703
rect 23388 37460 23440 37466
rect 23388 37402 23440 37408
rect 24320 36718 24348 38354
rect 24872 38282 24900 40870
rect 24952 40724 25004 40730
rect 24952 40666 25004 40672
rect 24492 38276 24544 38282
rect 24492 38218 24544 38224
rect 24860 38276 24912 38282
rect 24860 38218 24912 38224
rect 24504 37466 24532 38218
rect 24492 37460 24544 37466
rect 24492 37402 24544 37408
rect 24768 37324 24820 37330
rect 24768 37266 24820 37272
rect 24308 36712 24360 36718
rect 24308 36654 24360 36660
rect 24492 36576 24544 36582
rect 24492 36518 24544 36524
rect 24504 36378 24532 36518
rect 24780 36378 24808 37266
rect 24492 36372 24544 36378
rect 24492 36314 24544 36320
rect 24768 36372 24820 36378
rect 24768 36314 24820 36320
rect 24400 36304 24452 36310
rect 24136 36252 24400 36258
rect 24872 36281 24900 38218
rect 24964 37262 24992 40666
rect 25056 40458 25084 40870
rect 26344 40662 26372 40870
rect 26436 40730 26464 40870
rect 26424 40724 26476 40730
rect 26424 40666 26476 40672
rect 26332 40656 26384 40662
rect 26332 40598 26384 40604
rect 27528 40656 27580 40662
rect 27528 40598 27580 40604
rect 26516 40520 26568 40526
rect 26516 40462 26568 40468
rect 26792 40520 26844 40526
rect 26792 40462 26844 40468
rect 25044 40452 25096 40458
rect 25044 40394 25096 40400
rect 26528 40118 26556 40462
rect 26804 40186 26832 40462
rect 27540 40390 27568 40598
rect 27632 40458 27660 40870
rect 27816 40730 27844 40870
rect 27804 40724 27856 40730
rect 27804 40666 27856 40672
rect 27620 40452 27672 40458
rect 27620 40394 27672 40400
rect 27528 40384 27580 40390
rect 27528 40326 27580 40332
rect 27896 40384 27948 40390
rect 27896 40326 27948 40332
rect 28264 40384 28316 40390
rect 28460 40372 28488 42502
rect 29288 41818 29316 42706
rect 29380 42022 29408 42735
rect 31956 42702 31984 43046
rect 32220 42764 32272 42770
rect 32220 42706 32272 42712
rect 31944 42696 31996 42702
rect 31944 42638 31996 42644
rect 32232 42226 32260 42706
rect 32324 42702 32352 43046
rect 33244 42838 33272 43046
rect 33232 42832 33284 42838
rect 33232 42774 33284 42780
rect 32312 42696 32364 42702
rect 32312 42638 32364 42644
rect 32220 42220 32272 42226
rect 32220 42162 32272 42168
rect 30748 42084 30800 42090
rect 30748 42026 30800 42032
rect 29368 42016 29420 42022
rect 29368 41958 29420 41964
rect 29276 41812 29328 41818
rect 29276 41754 29328 41760
rect 30760 41546 30788 42026
rect 32128 42016 32180 42022
rect 32128 41958 32180 41964
rect 31576 41812 31628 41818
rect 31576 41754 31628 41760
rect 30932 41676 30984 41682
rect 30932 41618 30984 41624
rect 30748 41540 30800 41546
rect 30748 41482 30800 41488
rect 30944 41206 30972 41618
rect 31484 41472 31536 41478
rect 31484 41414 31536 41420
rect 30932 41200 30984 41206
rect 30932 41142 30984 41148
rect 30288 40928 30340 40934
rect 30288 40870 30340 40876
rect 28998 40488 29054 40497
rect 28998 40423 29054 40432
rect 28316 40344 28488 40372
rect 28264 40326 28316 40332
rect 26792 40180 26844 40186
rect 26792 40122 26844 40128
rect 27344 40180 27396 40186
rect 27344 40122 27396 40128
rect 26516 40112 26568 40118
rect 26516 40054 26568 40060
rect 27356 39982 27384 40122
rect 27908 39982 27936 40326
rect 27988 40180 28040 40186
rect 27988 40122 28040 40128
rect 25412 39976 25464 39982
rect 25412 39918 25464 39924
rect 25780 39976 25832 39982
rect 25780 39918 25832 39924
rect 25964 39976 26016 39982
rect 26148 39976 26200 39982
rect 25964 39918 26016 39924
rect 26068 39936 26148 39964
rect 25424 39574 25452 39918
rect 25412 39568 25464 39574
rect 25412 39510 25464 39516
rect 25424 38486 25452 39510
rect 25596 39500 25648 39506
rect 25596 39442 25648 39448
rect 25412 38480 25464 38486
rect 25412 38422 25464 38428
rect 25608 38418 25636 39442
rect 25596 38412 25648 38418
rect 25596 38354 25648 38360
rect 25792 37806 25820 39918
rect 25976 39574 26004 39918
rect 25964 39568 26016 39574
rect 25964 39510 26016 39516
rect 25780 37800 25832 37806
rect 25700 37760 25780 37788
rect 25044 37324 25096 37330
rect 25044 37266 25096 37272
rect 25412 37324 25464 37330
rect 25412 37266 25464 37272
rect 24952 37256 25004 37262
rect 24952 37198 25004 37204
rect 24964 36786 24992 37198
rect 24952 36780 25004 36786
rect 24952 36722 25004 36728
rect 25056 36718 25084 37266
rect 25424 36718 25452 37266
rect 25044 36712 25096 36718
rect 25044 36654 25096 36660
rect 25412 36712 25464 36718
rect 25412 36654 25464 36660
rect 24136 36246 24452 36252
rect 24858 36272 24914 36281
rect 24136 36242 24440 36246
rect 24124 36236 24440 36242
rect 23860 36196 24124 36224
rect 23860 36106 23888 36196
rect 24176 36230 24440 36236
rect 25056 36242 25084 36654
rect 25136 36576 25188 36582
rect 25136 36518 25188 36524
rect 24858 36207 24914 36216
rect 25044 36236 25096 36242
rect 24124 36178 24176 36184
rect 25044 36178 25096 36184
rect 23848 36100 23900 36106
rect 23848 36042 23900 36048
rect 24122 35728 24178 35737
rect 24122 35663 24124 35672
rect 24176 35663 24178 35672
rect 24124 35634 24176 35640
rect 25056 35494 25084 36178
rect 25148 36174 25176 36518
rect 25424 36242 25452 36654
rect 25412 36236 25464 36242
rect 25412 36178 25464 36184
rect 25136 36168 25188 36174
rect 25136 36110 25188 36116
rect 25424 36106 25452 36178
rect 25412 36100 25464 36106
rect 25412 36042 25464 36048
rect 25424 35834 25452 36042
rect 25412 35828 25464 35834
rect 25412 35770 25464 35776
rect 25504 35828 25556 35834
rect 25504 35770 25556 35776
rect 25136 35760 25188 35766
rect 25136 35702 25188 35708
rect 25148 35630 25176 35702
rect 25136 35624 25188 35630
rect 25136 35566 25188 35572
rect 25044 35488 25096 35494
rect 25044 35430 25096 35436
rect 24308 35148 24360 35154
rect 24308 35090 24360 35096
rect 22836 35080 22888 35086
rect 22836 35022 22888 35028
rect 22928 35080 22980 35086
rect 22928 35022 22980 35028
rect 22940 34649 22968 35022
rect 23388 34944 23440 34950
rect 23388 34886 23440 34892
rect 23664 34944 23716 34950
rect 23664 34886 23716 34892
rect 22926 34640 22982 34649
rect 23400 34610 23428 34886
rect 22926 34575 22982 34584
rect 23388 34604 23440 34610
rect 23388 34546 23440 34552
rect 23112 34060 23164 34066
rect 23112 34002 23164 34008
rect 22468 33924 22520 33930
rect 22468 33866 22520 33872
rect 22374 33416 22430 33425
rect 21732 33380 21784 33386
rect 22374 33351 22430 33360
rect 21732 33322 21784 33328
rect 22388 33318 22416 33351
rect 22376 33312 22428 33318
rect 22376 33254 22428 33260
rect 21284 33102 21588 33130
rect 21732 32904 21784 32910
rect 21732 32846 21784 32852
rect 22192 32904 22244 32910
rect 22192 32846 22244 32852
rect 21744 32774 21772 32846
rect 21732 32768 21784 32774
rect 21732 32710 21784 32716
rect 20812 32496 20864 32502
rect 20812 32438 20864 32444
rect 20904 32496 20956 32502
rect 20904 32438 20956 32444
rect 20720 31272 20772 31278
rect 20720 31214 20772 31220
rect 20732 30938 20760 31214
rect 20720 30932 20772 30938
rect 20720 30874 20772 30880
rect 20824 30802 20852 32438
rect 20916 31822 20944 32438
rect 21548 32428 21600 32434
rect 21548 32370 21600 32376
rect 20904 31816 20956 31822
rect 20904 31758 20956 31764
rect 21560 31414 21588 32370
rect 21744 32026 21772 32710
rect 21824 32292 21876 32298
rect 21824 32234 21876 32240
rect 21836 32026 21864 32234
rect 21732 32020 21784 32026
rect 21732 31962 21784 31968
rect 21824 32020 21876 32026
rect 21824 31962 21876 31968
rect 21640 31952 21692 31958
rect 21638 31920 21640 31929
rect 21692 31920 21694 31929
rect 21638 31855 21694 31864
rect 22008 31884 22060 31890
rect 22008 31826 22060 31832
rect 21548 31408 21600 31414
rect 21548 31350 21600 31356
rect 22020 31362 22048 31826
rect 22020 31334 22140 31362
rect 20996 31136 21048 31142
rect 20996 31078 21048 31084
rect 20812 30796 20864 30802
rect 20812 30738 20864 30744
rect 20824 29714 20852 30738
rect 21008 30598 21036 31078
rect 22112 30938 22140 31334
rect 22204 31142 22232 32846
rect 22282 31920 22338 31929
rect 22282 31855 22284 31864
rect 22336 31855 22338 31864
rect 22284 31826 22336 31832
rect 22192 31136 22244 31142
rect 22192 31078 22244 31084
rect 22100 30932 22152 30938
rect 22100 30874 22152 30880
rect 20996 30592 21048 30598
rect 20996 30534 21048 30540
rect 20812 29708 20864 29714
rect 20812 29650 20864 29656
rect 20812 29504 20864 29510
rect 20812 29446 20864 29452
rect 20720 29028 20772 29034
rect 20720 28970 20772 28976
rect 20352 28688 20404 28694
rect 20352 28630 20404 28636
rect 20536 28688 20588 28694
rect 20536 28630 20588 28636
rect 20352 28552 20404 28558
rect 20272 28512 20352 28540
rect 20352 28494 20404 28500
rect 20364 28422 20392 28494
rect 20352 28416 20404 28422
rect 20352 28358 20404 28364
rect 20364 28014 20392 28358
rect 20352 28008 20404 28014
rect 20352 27950 20404 27956
rect 20168 26852 20220 26858
rect 20168 26794 20220 26800
rect 20180 24410 20208 26794
rect 20548 26568 20576 28630
rect 20732 28082 20760 28970
rect 20720 28076 20772 28082
rect 20720 28018 20772 28024
rect 20824 27962 20852 29446
rect 20732 27934 20852 27962
rect 20628 27056 20680 27062
rect 20628 26998 20680 27004
rect 20640 26926 20668 26998
rect 20628 26920 20680 26926
rect 20628 26862 20680 26868
rect 20732 26790 20760 27934
rect 20812 27872 20864 27878
rect 20812 27814 20864 27820
rect 20824 27334 20852 27814
rect 20812 27328 20864 27334
rect 20812 27270 20864 27276
rect 20720 26784 20772 26790
rect 20720 26726 20772 26732
rect 20364 26540 20576 26568
rect 20168 24404 20220 24410
rect 20168 24346 20220 24352
rect 20168 23656 20220 23662
rect 20168 23598 20220 23604
rect 20180 23526 20208 23598
rect 20168 23520 20220 23526
rect 20166 23488 20168 23497
rect 20220 23488 20222 23497
rect 20166 23423 20222 23432
rect 20180 23254 20208 23423
rect 20168 23248 20220 23254
rect 20168 23190 20220 23196
rect 20076 22228 20128 22234
rect 20076 22170 20128 22176
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 19996 20398 20024 20538
rect 19984 20392 20036 20398
rect 19984 20334 20036 20340
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 19444 19854 19472 20198
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19996 19514 20024 20334
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 20168 18352 20220 18358
rect 20168 18294 20220 18300
rect 19432 18080 19484 18086
rect 19432 18022 19484 18028
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 19444 17746 19472 18022
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 19890 17368 19946 17377
rect 19996 17338 20024 18022
rect 20180 17338 20208 18294
rect 19890 17303 19946 17312
rect 19984 17332 20036 17338
rect 19904 17270 19932 17303
rect 19984 17274 20036 17280
rect 20168 17332 20220 17338
rect 20168 17274 20220 17280
rect 19892 17264 19944 17270
rect 19892 17206 19944 17212
rect 19432 17128 19484 17134
rect 19432 17070 19484 17076
rect 19444 15570 19472 17070
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 19892 15972 19944 15978
rect 19892 15914 19944 15920
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 19904 15570 19932 15914
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 19892 15564 19944 15570
rect 19892 15506 19944 15512
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19444 14482 19472 15302
rect 20364 15162 20392 26540
rect 20536 26444 20588 26450
rect 20536 26386 20588 26392
rect 20548 24614 20576 26386
rect 20628 25356 20680 25362
rect 20628 25298 20680 25304
rect 20536 24608 20588 24614
rect 20536 24550 20588 24556
rect 20640 24410 20668 25298
rect 20732 25294 20760 26726
rect 20824 25702 20852 27270
rect 20812 25696 20864 25702
rect 20812 25638 20864 25644
rect 20904 25696 20956 25702
rect 20904 25638 20956 25644
rect 20720 25288 20772 25294
rect 20720 25230 20772 25236
rect 20732 25158 20760 25230
rect 20720 25152 20772 25158
rect 20720 25094 20772 25100
rect 20628 24404 20680 24410
rect 20628 24346 20680 24352
rect 20732 23798 20760 25094
rect 20824 24614 20852 25638
rect 20812 24608 20864 24614
rect 20812 24550 20864 24556
rect 20720 23792 20772 23798
rect 20720 23734 20772 23740
rect 20824 23118 20852 24550
rect 20916 24274 20944 25638
rect 20904 24268 20956 24274
rect 20904 24210 20956 24216
rect 21008 23866 21036 30534
rect 22100 30184 22152 30190
rect 22100 30126 22152 30132
rect 22112 29850 22140 30126
rect 22100 29844 22152 29850
rect 22100 29786 22152 29792
rect 21824 29096 21876 29102
rect 21824 29038 21876 29044
rect 21836 28218 21864 29038
rect 21824 28212 21876 28218
rect 21824 28154 21876 28160
rect 21364 27872 21416 27878
rect 21364 27814 21416 27820
rect 21376 27538 21404 27814
rect 21364 27532 21416 27538
rect 21364 27474 21416 27480
rect 21456 27464 21508 27470
rect 21456 27406 21508 27412
rect 21916 27464 21968 27470
rect 21916 27406 21968 27412
rect 21468 27334 21496 27406
rect 21456 27328 21508 27334
rect 21456 27270 21508 27276
rect 21928 26994 21956 27406
rect 21916 26988 21968 26994
rect 21916 26930 21968 26936
rect 21088 26240 21140 26246
rect 21088 26182 21140 26188
rect 21100 25498 21128 26182
rect 21088 25492 21140 25498
rect 21088 25434 21140 25440
rect 21100 25362 21128 25434
rect 21088 25356 21140 25362
rect 21088 25298 21140 25304
rect 21548 25356 21600 25362
rect 21548 25298 21600 25304
rect 21824 25356 21876 25362
rect 21824 25298 21876 25304
rect 20996 23860 21048 23866
rect 20996 23802 21048 23808
rect 21560 23662 21588 25298
rect 21836 24410 21864 25298
rect 22008 25220 22060 25226
rect 22008 25162 22060 25168
rect 21824 24404 21876 24410
rect 21824 24346 21876 24352
rect 21548 23656 21600 23662
rect 21548 23598 21600 23604
rect 20812 23112 20864 23118
rect 20812 23054 20864 23060
rect 21640 23112 21692 23118
rect 21640 23054 21692 23060
rect 21272 22500 21324 22506
rect 21272 22442 21324 22448
rect 21284 22166 21312 22442
rect 21272 22160 21324 22166
rect 21270 22128 21272 22137
rect 21324 22128 21326 22137
rect 21270 22063 21326 22072
rect 21180 21480 21232 21486
rect 21180 21422 21232 21428
rect 20812 20392 20864 20398
rect 20812 20334 20864 20340
rect 20824 20262 20852 20334
rect 20628 20256 20680 20262
rect 20628 20198 20680 20204
rect 20812 20256 20864 20262
rect 20812 20198 20864 20204
rect 20640 16250 20668 20198
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20732 18222 20760 19110
rect 20720 18216 20772 18222
rect 20720 18158 20772 18164
rect 20732 18086 20760 18158
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 20628 16244 20680 16250
rect 20628 16186 20680 16192
rect 20640 16130 20668 16186
rect 20548 16102 20668 16130
rect 20352 15156 20404 15162
rect 20352 15098 20404 15104
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19156 14068 19208 14074
rect 19156 14010 19208 14016
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 18328 14000 18380 14006
rect 18328 13942 18380 13948
rect 18236 13864 18288 13870
rect 18236 13806 18288 13812
rect 18248 13462 18276 13806
rect 18236 13456 18288 13462
rect 18236 13398 18288 13404
rect 17960 12436 18012 12442
rect 17960 12378 18012 12384
rect 18340 12306 18368 13942
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 20548 12986 20576 16102
rect 20628 14952 20680 14958
rect 20628 14894 20680 14900
rect 20640 14550 20668 14894
rect 20628 14544 20680 14550
rect 20628 14486 20680 14492
rect 20732 14074 20760 18022
rect 20824 17202 20852 20198
rect 20996 19848 21048 19854
rect 20996 19790 21048 19796
rect 20812 17196 20864 17202
rect 20812 17138 20864 17144
rect 21008 15706 21036 19790
rect 21192 18358 21220 21422
rect 21652 21010 21680 23054
rect 21640 21004 21692 21010
rect 21640 20946 21692 20952
rect 21916 20936 21968 20942
rect 21916 20878 21968 20884
rect 21272 20256 21324 20262
rect 21272 20198 21324 20204
rect 21284 19922 21312 20198
rect 21272 19916 21324 19922
rect 21272 19858 21324 19864
rect 21928 19514 21956 20878
rect 21916 19508 21968 19514
rect 21916 19450 21968 19456
rect 21732 18760 21784 18766
rect 21732 18702 21784 18708
rect 21180 18352 21232 18358
rect 21180 18294 21232 18300
rect 21192 18222 21220 18294
rect 21180 18216 21232 18222
rect 21180 18158 21232 18164
rect 21640 18216 21692 18222
rect 21640 18158 21692 18164
rect 21192 17082 21220 18158
rect 21652 17882 21680 18158
rect 21640 17876 21692 17882
rect 21640 17818 21692 17824
rect 21100 17054 21220 17082
rect 21548 17128 21600 17134
rect 21548 17070 21600 17076
rect 21100 16046 21128 17054
rect 21560 16794 21588 17070
rect 21548 16788 21600 16794
rect 21548 16730 21600 16736
rect 21560 16046 21588 16730
rect 21088 16040 21140 16046
rect 21088 15982 21140 15988
rect 21548 16040 21600 16046
rect 21548 15982 21600 15988
rect 20996 15700 21048 15706
rect 20996 15642 21048 15648
rect 21008 15026 21036 15642
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 20720 14068 20772 14074
rect 20720 14010 20772 14016
rect 20812 13864 20864 13870
rect 20812 13806 20864 13812
rect 20536 12980 20588 12986
rect 20536 12922 20588 12928
rect 20824 12782 20852 13806
rect 21744 13530 21772 18702
rect 21824 18352 21876 18358
rect 21824 18294 21876 18300
rect 21836 18222 21864 18294
rect 21824 18216 21876 18222
rect 21824 18158 21876 18164
rect 21824 17264 21876 17270
rect 21824 17206 21876 17212
rect 21836 16726 21864 17206
rect 21824 16720 21876 16726
rect 21824 16662 21876 16668
rect 21928 15366 21956 15397
rect 21916 15360 21968 15366
rect 21914 15328 21916 15337
rect 21968 15328 21970 15337
rect 21914 15263 21970 15272
rect 21928 15162 21956 15263
rect 21916 15156 21968 15162
rect 21916 15098 21968 15104
rect 21824 14272 21876 14278
rect 21824 14214 21876 14220
rect 21836 13870 21864 14214
rect 21824 13864 21876 13870
rect 21824 13806 21876 13812
rect 22020 13546 22048 25162
rect 22100 25152 22152 25158
rect 22100 25094 22152 25100
rect 22112 24818 22140 25094
rect 22100 24812 22152 24818
rect 22100 24754 22152 24760
rect 22284 24064 22336 24070
rect 22284 24006 22336 24012
rect 22296 23662 22324 24006
rect 22284 23656 22336 23662
rect 22284 23598 22336 23604
rect 22376 21548 22428 21554
rect 22376 21490 22428 21496
rect 22284 21344 22336 21350
rect 22284 21286 22336 21292
rect 22296 19310 22324 21286
rect 22388 21146 22416 21490
rect 22480 21486 22508 33866
rect 22652 33312 22704 33318
rect 22652 33254 22704 33260
rect 22560 31272 22612 31278
rect 22560 31214 22612 31220
rect 22572 30870 22600 31214
rect 22560 30864 22612 30870
rect 22560 30806 22612 30812
rect 22664 30326 22692 33254
rect 23020 31884 23072 31890
rect 23020 31826 23072 31832
rect 22744 31408 22796 31414
rect 22744 31350 22796 31356
rect 22756 30938 22784 31350
rect 22744 30932 22796 30938
rect 22744 30874 22796 30880
rect 22836 30728 22888 30734
rect 22836 30670 22888 30676
rect 22744 30388 22796 30394
rect 22744 30330 22796 30336
rect 22652 30320 22704 30326
rect 22652 30262 22704 30268
rect 22664 29850 22692 30262
rect 22652 29844 22704 29850
rect 22652 29786 22704 29792
rect 22664 29714 22692 29786
rect 22652 29708 22704 29714
rect 22652 29650 22704 29656
rect 22560 29096 22612 29102
rect 22560 29038 22612 29044
rect 22572 28558 22600 29038
rect 22652 28960 22704 28966
rect 22652 28902 22704 28908
rect 22664 28665 22692 28902
rect 22650 28656 22706 28665
rect 22650 28591 22706 28600
rect 22560 28552 22612 28558
rect 22560 28494 22612 28500
rect 22756 26738 22784 30330
rect 22664 26710 22784 26738
rect 22560 23520 22612 23526
rect 22560 23462 22612 23468
rect 22572 23186 22600 23462
rect 22560 23180 22612 23186
rect 22560 23122 22612 23128
rect 22468 21480 22520 21486
rect 22468 21422 22520 21428
rect 22560 21344 22612 21350
rect 22560 21286 22612 21292
rect 22572 21146 22600 21286
rect 22376 21140 22428 21146
rect 22376 21082 22428 21088
rect 22560 21140 22612 21146
rect 22560 21082 22612 21088
rect 22560 20392 22612 20398
rect 22560 20334 22612 20340
rect 22572 20058 22600 20334
rect 22560 20052 22612 20058
rect 22560 19994 22612 20000
rect 22284 19304 22336 19310
rect 22284 19246 22336 19252
rect 22192 18760 22244 18766
rect 22192 18702 22244 18708
rect 22204 18426 22232 18702
rect 22192 18420 22244 18426
rect 22192 18362 22244 18368
rect 22296 18154 22324 19246
rect 22284 18148 22336 18154
rect 22284 18090 22336 18096
rect 22664 16658 22692 26710
rect 22848 18970 22876 30670
rect 22928 27464 22980 27470
rect 22928 27406 22980 27412
rect 22940 21554 22968 27406
rect 23032 23322 23060 31826
rect 23020 23316 23072 23322
rect 23020 23258 23072 23264
rect 22928 21548 22980 21554
rect 22928 21490 22980 21496
rect 23124 20602 23152 34002
rect 23676 33998 23704 34886
rect 23848 34400 23900 34406
rect 23848 34342 23900 34348
rect 23664 33992 23716 33998
rect 23664 33934 23716 33940
rect 23204 33856 23256 33862
rect 23204 33798 23256 33804
rect 23216 27470 23244 33798
rect 23860 33658 23888 34342
rect 24320 34134 24348 35090
rect 25056 35018 25084 35430
rect 25320 35284 25372 35290
rect 25320 35226 25372 35232
rect 25332 35154 25360 35226
rect 25516 35193 25544 35770
rect 25502 35184 25558 35193
rect 25320 35148 25372 35154
rect 25502 35119 25558 35128
rect 25320 35090 25372 35096
rect 25044 35012 25096 35018
rect 25044 34954 25096 34960
rect 25332 34678 25360 35090
rect 25320 34672 25372 34678
rect 25320 34614 25372 34620
rect 24308 34128 24360 34134
rect 24308 34070 24360 34076
rect 24400 34128 24452 34134
rect 24400 34070 24452 34076
rect 24858 34096 24914 34105
rect 24412 33930 24440 34070
rect 24858 34031 24914 34040
rect 24582 33960 24638 33969
rect 24400 33924 24452 33930
rect 24582 33895 24638 33904
rect 24400 33866 24452 33872
rect 24596 33862 24624 33895
rect 24584 33856 24636 33862
rect 24584 33798 24636 33804
rect 24768 33788 24820 33794
rect 24768 33730 24820 33736
rect 23848 33652 23900 33658
rect 23848 33594 23900 33600
rect 24400 33652 24452 33658
rect 24400 33594 24452 33600
rect 24584 33652 24636 33658
rect 24780 33640 24808 33730
rect 24872 33658 24900 34031
rect 24636 33612 24808 33640
rect 24860 33652 24912 33658
rect 24584 33594 24636 33600
rect 24860 33594 24912 33600
rect 23296 31680 23348 31686
rect 23296 31622 23348 31628
rect 23308 31414 23336 31622
rect 23296 31408 23348 31414
rect 23296 31350 23348 31356
rect 23388 31408 23440 31414
rect 23388 31350 23440 31356
rect 23400 30394 23428 31350
rect 24214 30832 24270 30841
rect 24214 30767 24270 30776
rect 23388 30388 23440 30394
rect 23388 30330 23440 30336
rect 23478 30152 23534 30161
rect 23478 30087 23534 30096
rect 23492 29102 23520 30087
rect 23480 29096 23532 29102
rect 23480 29038 23532 29044
rect 23386 28112 23442 28121
rect 23386 28047 23442 28056
rect 23204 27464 23256 27470
rect 23204 27406 23256 27412
rect 23204 27328 23256 27334
rect 23204 27270 23256 27276
rect 23216 26450 23244 27270
rect 23296 26784 23348 26790
rect 23296 26726 23348 26732
rect 23308 26450 23336 26726
rect 23400 26518 23428 28047
rect 23388 26512 23440 26518
rect 23388 26454 23440 26460
rect 23204 26444 23256 26450
rect 23204 26386 23256 26392
rect 23296 26444 23348 26450
rect 23296 26386 23348 26392
rect 23572 24676 23624 24682
rect 23572 24618 23624 24624
rect 23584 24342 23612 24618
rect 23572 24336 23624 24342
rect 23572 24278 23624 24284
rect 23480 24268 23532 24274
rect 23480 24210 23532 24216
rect 23492 22982 23520 24210
rect 23584 24177 23612 24278
rect 24124 24200 24176 24206
rect 23570 24168 23626 24177
rect 24124 24142 24176 24148
rect 23570 24103 23626 24112
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23492 22817 23520 22918
rect 23478 22808 23534 22817
rect 23478 22743 23534 22752
rect 24136 21894 24164 24142
rect 24124 21888 24176 21894
rect 24124 21830 24176 21836
rect 23112 20596 23164 20602
rect 23112 20538 23164 20544
rect 23478 20088 23534 20097
rect 23478 20023 23534 20032
rect 22836 18964 22888 18970
rect 22836 18906 22888 18912
rect 22652 16652 22704 16658
rect 22652 16594 22704 16600
rect 22192 15972 22244 15978
rect 22192 15914 22244 15920
rect 22204 15570 22232 15914
rect 22192 15564 22244 15570
rect 22192 15506 22244 15512
rect 23386 14784 23442 14793
rect 23386 14719 23442 14728
rect 22192 13796 22244 13802
rect 22192 13738 22244 13744
rect 21732 13524 21784 13530
rect 21732 13466 21784 13472
rect 21836 13518 22048 13546
rect 21836 13410 21864 13518
rect 21744 13382 21864 13410
rect 22204 13394 22232 13738
rect 22008 13388 22060 13394
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 18328 12300 18380 12306
rect 18328 12242 18380 12248
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 19352 11218 19380 12038
rect 19892 11892 19944 11898
rect 19892 11834 19944 11840
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 19432 11348 19484 11354
rect 19432 11290 19484 11296
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 18328 11008 18380 11014
rect 18328 10950 18380 10956
rect 18340 10674 18368 10950
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 19444 9178 19472 11290
rect 19904 11082 19932 11834
rect 20824 11762 20852 12718
rect 21364 12300 21416 12306
rect 21364 12242 21416 12248
rect 21376 11898 21404 12242
rect 21364 11892 21416 11898
rect 21364 11834 21416 11840
rect 20812 11756 20864 11762
rect 20812 11698 20864 11704
rect 20904 11552 20956 11558
rect 20904 11494 20956 11500
rect 19892 11076 19944 11082
rect 19892 11018 19944 11024
rect 19904 10810 19932 11018
rect 19892 10804 19944 10810
rect 19892 10746 19944 10752
rect 20916 10674 20944 11494
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 20904 10668 20956 10674
rect 20904 10610 20956 10616
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 20548 10266 20576 10610
rect 21456 10464 21508 10470
rect 21456 10406 21508 10412
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 20548 9722 20576 10202
rect 21468 10130 21496 10406
rect 21456 10124 21508 10130
rect 21456 10066 21508 10072
rect 20536 9716 20588 9722
rect 20536 9658 20588 9664
rect 20076 9512 20128 9518
rect 20076 9454 20128 9460
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 19352 8430 19380 8774
rect 20088 8634 20116 9454
rect 20548 9382 20576 9658
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20548 9178 20576 9318
rect 20536 9172 20588 9178
rect 20536 9114 20588 9120
rect 20548 8634 20576 9114
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 20536 8628 20588 8634
rect 20536 8570 20588 8576
rect 20720 8560 20772 8566
rect 20720 8502 20772 8508
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 17868 8084 17920 8090
rect 17868 8026 17920 8032
rect 19352 7410 19380 8366
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 20732 7546 20760 8502
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 19340 7404 19392 7410
rect 19340 7346 19392 7352
rect 19984 7200 20036 7206
rect 19984 7142 20036 7148
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 19996 6866 20024 7142
rect 20732 7002 20760 7482
rect 20720 6996 20772 7002
rect 20720 6938 20772 6944
rect 16304 6860 16356 6866
rect 16304 6802 16356 6808
rect 19984 6860 20036 6866
rect 19984 6802 20036 6808
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 15672 6254 15700 6734
rect 16224 6254 16252 6734
rect 16316 6458 16344 6802
rect 20732 6798 20760 6938
rect 20720 6792 20772 6798
rect 20720 6734 20772 6740
rect 19892 6656 19944 6662
rect 19892 6598 19944 6604
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 15660 6248 15712 6254
rect 15660 6190 15712 6196
rect 16212 6248 16264 6254
rect 16212 6190 16264 6196
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15200 5908 15252 5914
rect 15200 5850 15252 5856
rect 15384 5908 15436 5914
rect 15384 5850 15436 5856
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 15108 5840 15160 5846
rect 15108 5782 15160 5788
rect 15212 5710 15240 5850
rect 15580 5778 15608 6054
rect 15672 5914 15700 6190
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 16224 5710 16252 6190
rect 16856 6180 16908 6186
rect 16856 6122 16908 6128
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 16212 5704 16264 5710
rect 16212 5646 16264 5652
rect 15212 5370 15240 5646
rect 16868 5370 16896 6122
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 19904 5778 19932 6598
rect 20732 6322 20760 6734
rect 20720 6316 20772 6322
rect 20720 6258 20772 6264
rect 20732 5914 20760 6258
rect 20904 6248 20956 6254
rect 20904 6190 20956 6196
rect 20720 5908 20772 5914
rect 20720 5850 20772 5856
rect 19892 5772 19944 5778
rect 19892 5714 19944 5720
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 16856 5364 16908 5370
rect 16856 5306 16908 5312
rect 16672 5160 16724 5166
rect 16672 5102 16724 5108
rect 16684 4826 16712 5102
rect 16672 4820 16724 4826
rect 16672 4762 16724 4768
rect 19352 4690 19380 5510
rect 19904 5234 19932 5714
rect 19892 5228 19944 5234
rect 19892 5170 19944 5176
rect 20732 5166 20760 5850
rect 20916 5370 20944 6190
rect 21744 5914 21772 13382
rect 22008 13330 22060 13336
rect 22192 13388 22244 13394
rect 22192 13330 22244 13336
rect 21824 12640 21876 12646
rect 21824 12582 21876 12588
rect 21836 12306 21864 12582
rect 22020 12442 22048 13330
rect 22284 12776 22336 12782
rect 22284 12718 22336 12724
rect 22008 12436 22060 12442
rect 22008 12378 22060 12384
rect 21824 12300 21876 12306
rect 21824 12242 21876 12248
rect 22296 11898 22324 12718
rect 23400 12374 23428 14719
rect 23492 14482 23520 20023
rect 24136 17134 24164 21830
rect 24124 17128 24176 17134
rect 24124 17070 24176 17076
rect 23572 16652 23624 16658
rect 23572 16594 23624 16600
rect 23584 15638 23612 16594
rect 23572 15632 23624 15638
rect 23572 15574 23624 15580
rect 23480 14476 23532 14482
rect 23480 14418 23532 14424
rect 23492 13530 23520 14418
rect 23480 13524 23532 13530
rect 23480 13466 23532 13472
rect 23388 12368 23440 12374
rect 23388 12310 23440 12316
rect 22284 11892 22336 11898
rect 22284 11834 22336 11840
rect 23400 11694 23428 12310
rect 23388 11688 23440 11694
rect 23388 11630 23440 11636
rect 24228 11354 24256 30767
rect 24412 27878 24440 33594
rect 24860 32428 24912 32434
rect 24860 32370 24912 32376
rect 24492 30252 24544 30258
rect 24492 30194 24544 30200
rect 24400 27872 24452 27878
rect 24400 27814 24452 27820
rect 24306 26752 24362 26761
rect 24306 26687 24362 26696
rect 24320 26586 24348 26687
rect 24308 26580 24360 26586
rect 24308 26522 24360 26528
rect 24504 22098 24532 30194
rect 24766 29472 24822 29481
rect 24766 29407 24822 29416
rect 24780 29170 24808 29407
rect 24768 29164 24820 29170
rect 24768 29106 24820 29112
rect 24872 26450 24900 32370
rect 25700 27130 25728 37760
rect 25780 37742 25832 37748
rect 26068 37262 26096 39936
rect 26148 39918 26200 39924
rect 27344 39976 27396 39982
rect 27344 39918 27396 39924
rect 27896 39976 27948 39982
rect 27896 39918 27948 39924
rect 27620 39500 27672 39506
rect 27620 39442 27672 39448
rect 26332 38956 26384 38962
rect 26332 38898 26384 38904
rect 26240 38208 26292 38214
rect 26240 38150 26292 38156
rect 26148 37800 26200 37806
rect 26252 37788 26280 38150
rect 26344 37942 26372 38898
rect 26424 38888 26476 38894
rect 26424 38830 26476 38836
rect 26436 37942 26464 38830
rect 27160 38820 27212 38826
rect 27160 38762 27212 38768
rect 27172 38214 27200 38762
rect 27344 38344 27396 38350
rect 27344 38286 27396 38292
rect 27356 38214 27384 38286
rect 27160 38208 27212 38214
rect 27160 38150 27212 38156
rect 27344 38208 27396 38214
rect 27344 38150 27396 38156
rect 27172 37942 27200 38150
rect 26332 37936 26384 37942
rect 26332 37878 26384 37884
rect 26424 37936 26476 37942
rect 26424 37878 26476 37884
rect 27160 37936 27212 37942
rect 27160 37878 27212 37884
rect 26200 37760 26280 37788
rect 26148 37742 26200 37748
rect 26252 37466 26280 37760
rect 26240 37460 26292 37466
rect 26240 37402 26292 37408
rect 26252 37330 26280 37402
rect 27356 37330 27384 38150
rect 26240 37324 26292 37330
rect 26240 37266 26292 37272
rect 27344 37324 27396 37330
rect 27344 37266 27396 37272
rect 26056 37256 26108 37262
rect 26056 37198 26108 37204
rect 26792 36780 26844 36786
rect 26792 36722 26844 36728
rect 26424 36644 26476 36650
rect 26424 36586 26476 36592
rect 26240 36372 26292 36378
rect 26240 36314 26292 36320
rect 26056 34944 26108 34950
rect 26056 34886 26108 34892
rect 26068 34474 26096 34886
rect 26252 34474 26280 36314
rect 26056 34468 26108 34474
rect 26056 34410 26108 34416
rect 26240 34468 26292 34474
rect 26240 34410 26292 34416
rect 26436 29782 26464 36586
rect 26804 35630 26832 36722
rect 27160 36712 27212 36718
rect 27160 36654 27212 36660
rect 26976 36372 27028 36378
rect 26976 36314 27028 36320
rect 26988 36242 27016 36314
rect 26976 36236 27028 36242
rect 26976 36178 27028 36184
rect 27172 36106 27200 36654
rect 27160 36100 27212 36106
rect 27160 36042 27212 36048
rect 26974 35728 27030 35737
rect 26974 35663 26976 35672
rect 27028 35663 27030 35672
rect 26976 35634 27028 35640
rect 27172 35630 27200 36042
rect 26792 35624 26844 35630
rect 26792 35566 26844 35572
rect 27160 35624 27212 35630
rect 27160 35566 27212 35572
rect 26516 35488 26568 35494
rect 26516 35430 26568 35436
rect 26608 35488 26660 35494
rect 26608 35430 26660 35436
rect 26424 29776 26476 29782
rect 26424 29718 26476 29724
rect 26528 28422 26556 35430
rect 26620 34785 26648 35430
rect 26606 34776 26662 34785
rect 26606 34711 26662 34720
rect 26620 34406 26648 34711
rect 26700 34536 26752 34542
rect 26700 34478 26752 34484
rect 26608 34400 26660 34406
rect 26608 34342 26660 34348
rect 26712 30258 26740 34478
rect 26976 31544 27028 31550
rect 26976 31486 27028 31492
rect 26792 31068 26844 31074
rect 26792 31010 26844 31016
rect 26700 30252 26752 30258
rect 26700 30194 26752 30200
rect 26516 28416 26568 28422
rect 26516 28358 26568 28364
rect 25688 27124 25740 27130
rect 25688 27066 25740 27072
rect 24860 26444 24912 26450
rect 24860 26386 24912 26392
rect 24768 25696 24820 25702
rect 24768 25638 24820 25644
rect 24780 25537 24808 25638
rect 24766 25528 24822 25537
rect 24766 25463 24822 25472
rect 26804 24750 26832 31010
rect 26884 30932 26936 30938
rect 26884 30874 26936 30880
rect 26792 24744 26844 24750
rect 26792 24686 26844 24692
rect 24492 22092 24544 22098
rect 24492 22034 24544 22040
rect 26896 16522 26924 30874
rect 26988 17950 27016 31486
rect 27068 31000 27120 31006
rect 27068 30942 27120 30948
rect 26976 17944 27028 17950
rect 26976 17886 27028 17892
rect 27080 17338 27108 30942
rect 27356 28966 27384 37266
rect 27632 34950 27660 39442
rect 27712 39432 27764 39438
rect 27804 39432 27856 39438
rect 27764 39380 27804 39386
rect 27712 39374 27856 39380
rect 27724 39358 27844 39374
rect 28000 39302 28028 40122
rect 28276 40118 28304 40326
rect 28264 40112 28316 40118
rect 28264 40054 28316 40060
rect 28080 39976 28132 39982
rect 28080 39918 28132 39924
rect 27804 39296 27856 39302
rect 27804 39238 27856 39244
rect 27988 39296 28040 39302
rect 28092 39273 28120 39918
rect 27988 39238 28040 39244
rect 28078 39264 28134 39273
rect 27816 38486 27844 39238
rect 28078 39199 28134 39208
rect 28276 38758 28304 40054
rect 29012 39982 29040 40423
rect 29000 39976 29052 39982
rect 29000 39918 29052 39924
rect 30300 39846 30328 40870
rect 30944 40594 30972 41142
rect 31496 41070 31524 41414
rect 31588 41070 31616 41754
rect 31760 41608 31812 41614
rect 31760 41550 31812 41556
rect 31484 41064 31536 41070
rect 31484 41006 31536 41012
rect 31576 41064 31628 41070
rect 31576 41006 31628 41012
rect 30932 40588 30984 40594
rect 30932 40530 30984 40536
rect 31588 40526 31616 41006
rect 31772 40934 31800 41550
rect 32140 41138 32168 41958
rect 32220 41540 32272 41546
rect 32220 41482 32272 41488
rect 32128 41132 32180 41138
rect 32128 41074 32180 41080
rect 31944 41064 31996 41070
rect 31944 41006 31996 41012
rect 31760 40928 31812 40934
rect 31760 40870 31812 40876
rect 31760 40724 31812 40730
rect 31760 40666 31812 40672
rect 31576 40520 31628 40526
rect 31576 40462 31628 40468
rect 31666 40488 31722 40497
rect 31666 40423 31722 40432
rect 31680 40118 31708 40423
rect 31772 40186 31800 40666
rect 31956 40526 31984 41006
rect 32036 40656 32088 40662
rect 32036 40598 32088 40604
rect 31944 40520 31996 40526
rect 31944 40462 31996 40468
rect 31760 40180 31812 40186
rect 31760 40122 31812 40128
rect 32048 40118 32076 40598
rect 32232 40458 32260 41482
rect 32220 40452 32272 40458
rect 32220 40394 32272 40400
rect 31668 40112 31720 40118
rect 31668 40054 31720 40060
rect 32036 40112 32088 40118
rect 32036 40054 32088 40060
rect 31574 39944 31630 39953
rect 31574 39879 31576 39888
rect 31628 39879 31630 39888
rect 31576 39850 31628 39856
rect 30288 39840 30340 39846
rect 30288 39782 30340 39788
rect 31588 39574 31616 39850
rect 32324 39846 32352 42638
rect 33876 42560 33928 42566
rect 33876 42502 33928 42508
rect 33888 42242 33916 42502
rect 32588 42220 32640 42226
rect 32588 42162 32640 42168
rect 33152 42214 33916 42242
rect 32600 42022 32628 42162
rect 33152 42090 33180 42214
rect 33508 42152 33560 42158
rect 33508 42094 33560 42100
rect 33140 42084 33192 42090
rect 33140 42026 33192 42032
rect 32588 42016 32640 42022
rect 32588 41958 32640 41964
rect 32404 41676 32456 41682
rect 32404 41618 32456 41624
rect 32680 41676 32732 41682
rect 32680 41618 32732 41624
rect 32416 41585 32444 41618
rect 32402 41576 32458 41585
rect 32402 41511 32458 41520
rect 32692 41478 32720 41618
rect 32864 41540 32916 41546
rect 32864 41482 32916 41488
rect 32680 41472 32732 41478
rect 32680 41414 32732 41420
rect 32692 41070 32720 41414
rect 32404 41064 32456 41070
rect 32496 41064 32548 41070
rect 32404 41006 32456 41012
rect 32494 41032 32496 41041
rect 32680 41064 32732 41070
rect 32548 41032 32550 41041
rect 32416 40934 32444 41006
rect 32680 41006 32732 41012
rect 32494 40967 32550 40976
rect 32404 40928 32456 40934
rect 32404 40870 32456 40876
rect 32772 40588 32824 40594
rect 32772 40530 32824 40536
rect 32784 40497 32812 40530
rect 32770 40488 32826 40497
rect 32770 40423 32826 40432
rect 32404 39976 32456 39982
rect 32402 39944 32404 39953
rect 32456 39944 32458 39953
rect 32402 39879 32458 39888
rect 32678 39944 32734 39953
rect 32678 39879 32734 39888
rect 32312 39840 32364 39846
rect 32312 39782 32364 39788
rect 32220 39636 32272 39642
rect 32220 39578 32272 39584
rect 31576 39568 31628 39574
rect 31576 39510 31628 39516
rect 31760 39568 31812 39574
rect 31760 39510 31812 39516
rect 31772 39438 31800 39510
rect 31760 39432 31812 39438
rect 31760 39374 31812 39380
rect 28264 38752 28316 38758
rect 28264 38694 28316 38700
rect 31484 38548 31536 38554
rect 31484 38490 31536 38496
rect 27804 38480 27856 38486
rect 27804 38422 27856 38428
rect 28816 38480 28868 38486
rect 28816 38422 28868 38428
rect 27816 37330 27844 38422
rect 27896 38412 27948 38418
rect 27896 38354 27948 38360
rect 28632 38412 28684 38418
rect 28632 38354 28684 38360
rect 27908 37806 27936 38354
rect 27896 37800 27948 37806
rect 27896 37742 27948 37748
rect 27804 37324 27856 37330
rect 27804 37266 27856 37272
rect 28644 36786 28672 38354
rect 28828 37466 28856 38422
rect 28908 38208 28960 38214
rect 28908 38150 28960 38156
rect 28920 37874 28948 38150
rect 31496 37942 31524 38490
rect 31484 37936 31536 37942
rect 31484 37878 31536 37884
rect 31944 37936 31996 37942
rect 31944 37878 31996 37884
rect 28908 37868 28960 37874
rect 28908 37810 28960 37816
rect 31956 37806 31984 37878
rect 31852 37800 31904 37806
rect 31852 37742 31904 37748
rect 31944 37800 31996 37806
rect 31996 37760 32076 37788
rect 31944 37742 31996 37748
rect 31864 37466 31892 37742
rect 32048 37670 32076 37760
rect 32036 37664 32088 37670
rect 32036 37606 32088 37612
rect 28816 37460 28868 37466
rect 28816 37402 28868 37408
rect 31852 37460 31904 37466
rect 31852 37402 31904 37408
rect 28828 37346 28856 37402
rect 28736 37330 28856 37346
rect 28724 37324 28856 37330
rect 28776 37318 28856 37324
rect 28724 37266 28776 37272
rect 28632 36780 28684 36786
rect 28632 36722 28684 36728
rect 28736 36718 28764 37266
rect 28816 37256 28868 37262
rect 28816 37198 28868 37204
rect 28828 36922 28856 37198
rect 31760 37120 31812 37126
rect 31760 37062 31812 37068
rect 28816 36916 28868 36922
rect 28816 36858 28868 36864
rect 28724 36712 28776 36718
rect 28724 36654 28776 36660
rect 30380 36712 30432 36718
rect 30380 36654 30432 36660
rect 29092 36372 29144 36378
rect 29092 36314 29144 36320
rect 29644 36372 29696 36378
rect 29644 36314 29696 36320
rect 29104 36122 29132 36314
rect 29550 36272 29606 36281
rect 29368 36236 29420 36242
rect 29420 36216 29550 36224
rect 29420 36196 29552 36216
rect 29368 36178 29420 36184
rect 29604 36207 29606 36216
rect 29552 36178 29604 36184
rect 28920 36094 29132 36122
rect 29656 36106 29684 36314
rect 29644 36100 29696 36106
rect 28448 36032 28500 36038
rect 28448 35974 28500 35980
rect 28460 35154 28488 35974
rect 28920 35630 28948 36094
rect 29644 36042 29696 36048
rect 30104 36100 30156 36106
rect 30104 36042 30156 36048
rect 28908 35624 28960 35630
rect 28908 35566 28960 35572
rect 29092 35624 29144 35630
rect 29092 35566 29144 35572
rect 28080 35148 28132 35154
rect 28080 35090 28132 35096
rect 28448 35148 28500 35154
rect 28448 35090 28500 35096
rect 28092 34950 28120 35090
rect 28460 34950 28488 35090
rect 29104 35018 29132 35566
rect 30116 35562 30144 36042
rect 30288 35760 30340 35766
rect 30288 35702 30340 35708
rect 30194 35592 30250 35601
rect 30104 35556 30156 35562
rect 30194 35527 30250 35536
rect 30104 35498 30156 35504
rect 30116 35154 30144 35498
rect 30208 35494 30236 35527
rect 30196 35488 30248 35494
rect 30196 35430 30248 35436
rect 30300 35154 30328 35702
rect 30392 35290 30420 36654
rect 31772 36174 31800 37062
rect 31864 36718 31892 37402
rect 31944 37120 31996 37126
rect 31944 37062 31996 37068
rect 31852 36712 31904 36718
rect 31852 36654 31904 36660
rect 31956 36242 31984 37062
rect 32048 36854 32076 37606
rect 32036 36848 32088 36854
rect 32036 36790 32088 36796
rect 32128 36780 32180 36786
rect 32128 36722 32180 36728
rect 32140 36242 32168 36722
rect 31944 36236 31996 36242
rect 31944 36178 31996 36184
rect 32128 36236 32180 36242
rect 32128 36178 32180 36184
rect 31760 36168 31812 36174
rect 31760 36110 31812 36116
rect 30564 36032 30616 36038
rect 30564 35974 30616 35980
rect 30576 35698 30604 35974
rect 30564 35692 30616 35698
rect 30564 35634 30616 35640
rect 31300 35624 31352 35630
rect 31300 35566 31352 35572
rect 30380 35284 30432 35290
rect 30380 35226 30432 35232
rect 30472 35284 30524 35290
rect 30472 35226 30524 35232
rect 30104 35148 30156 35154
rect 30104 35090 30156 35096
rect 30288 35148 30340 35154
rect 30288 35090 30340 35096
rect 29092 35012 29144 35018
rect 29092 34954 29144 34960
rect 27620 34944 27672 34950
rect 27620 34886 27672 34892
rect 28080 34944 28132 34950
rect 28080 34886 28132 34892
rect 28448 34944 28500 34950
rect 28448 34886 28500 34892
rect 27528 34196 27580 34202
rect 27528 34138 27580 34144
rect 27540 33833 27568 34138
rect 27526 33824 27582 33833
rect 27526 33759 27582 33768
rect 28356 32632 28408 32638
rect 28356 32574 28408 32580
rect 27344 28960 27396 28966
rect 27344 28902 27396 28908
rect 28368 27402 28396 32574
rect 28356 27396 28408 27402
rect 28356 27338 28408 27344
rect 28460 21962 28488 34886
rect 30484 34678 30512 35226
rect 31312 35222 31340 35566
rect 31956 35494 31984 36178
rect 32128 35760 32180 35766
rect 32128 35702 32180 35708
rect 31760 35488 31812 35494
rect 31760 35430 31812 35436
rect 31944 35488 31996 35494
rect 31944 35430 31996 35436
rect 31772 35306 31800 35430
rect 32140 35306 32168 35702
rect 31772 35278 32168 35306
rect 31300 35216 31352 35222
rect 30562 35184 30618 35193
rect 31300 35158 31352 35164
rect 30562 35119 30618 35128
rect 30472 34672 30524 34678
rect 30472 34614 30524 34620
rect 30576 34542 30604 35119
rect 31668 35080 31720 35086
rect 31668 35022 31720 35028
rect 31760 35080 31812 35086
rect 31760 35022 31812 35028
rect 31680 34950 31708 35022
rect 31668 34944 31720 34950
rect 31668 34886 31720 34892
rect 30564 34536 30616 34542
rect 30564 34478 30616 34484
rect 30748 34536 30800 34542
rect 30748 34478 30800 34484
rect 30932 34536 30984 34542
rect 30932 34478 30984 34484
rect 30760 33522 30788 34478
rect 30748 33516 30800 33522
rect 30748 33458 30800 33464
rect 30944 33046 30972 34478
rect 30932 33040 30984 33046
rect 30932 32982 30984 32988
rect 31772 32910 31800 35022
rect 32232 34610 32260 39578
rect 32312 39500 32364 39506
rect 32312 39442 32364 39448
rect 32324 38758 32352 39442
rect 32312 38752 32364 38758
rect 32312 38694 32364 38700
rect 32692 37126 32720 39879
rect 32772 39500 32824 39506
rect 32772 39442 32824 39448
rect 32784 39030 32812 39442
rect 32772 39024 32824 39030
rect 32772 38966 32824 38972
rect 32876 38418 32904 41482
rect 33520 41478 33548 42094
rect 33980 41682 34008 43182
rect 35256 43172 35308 43178
rect 35256 43114 35308 43120
rect 34152 43104 34204 43110
rect 34152 43046 34204 43052
rect 34164 42226 34192 43046
rect 35268 42770 35296 43114
rect 38198 42800 38254 42809
rect 35256 42764 35308 42770
rect 38198 42735 38254 42744
rect 35256 42706 35308 42712
rect 38212 42702 38240 42735
rect 34980 42696 35032 42702
rect 34978 42664 34980 42673
rect 37740 42696 37792 42702
rect 35032 42664 35034 42673
rect 34978 42599 35034 42608
rect 37738 42664 37740 42673
rect 38200 42696 38252 42702
rect 37792 42664 37794 42673
rect 38200 42638 38252 42644
rect 37738 42599 37794 42608
rect 34940 42460 35236 42480
rect 34996 42458 35020 42460
rect 35076 42458 35100 42460
rect 35156 42458 35180 42460
rect 35018 42406 35020 42458
rect 35082 42406 35094 42458
rect 35156 42406 35158 42458
rect 34996 42404 35020 42406
rect 35076 42404 35100 42406
rect 35156 42404 35180 42406
rect 34940 42384 35236 42404
rect 38660 42356 38712 42362
rect 38660 42298 38712 42304
rect 37372 42288 37424 42294
rect 37094 42256 37150 42265
rect 34152 42220 34204 42226
rect 37372 42230 37424 42236
rect 37094 42191 37096 42200
rect 34152 42162 34204 42168
rect 37148 42191 37150 42200
rect 37096 42162 37148 42168
rect 37384 42158 37412 42230
rect 34428 42152 34480 42158
rect 34428 42094 34480 42100
rect 37372 42152 37424 42158
rect 37372 42094 37424 42100
rect 34336 42016 34388 42022
rect 34336 41958 34388 41964
rect 34060 41744 34112 41750
rect 34060 41686 34112 41692
rect 33876 41676 33928 41682
rect 33876 41618 33928 41624
rect 33968 41676 34020 41682
rect 33968 41618 34020 41624
rect 33690 41576 33746 41585
rect 33690 41511 33692 41520
rect 33744 41511 33746 41520
rect 33692 41482 33744 41488
rect 33508 41472 33560 41478
rect 33508 41414 33560 41420
rect 33416 41132 33468 41138
rect 33416 41074 33468 41080
rect 33322 41032 33378 41041
rect 33428 41002 33456 41074
rect 33322 40967 33378 40976
rect 33416 40996 33468 41002
rect 33336 40934 33364 40967
rect 33416 40938 33468 40944
rect 33140 40928 33192 40934
rect 33140 40870 33192 40876
rect 33324 40928 33376 40934
rect 33324 40870 33376 40876
rect 33508 40928 33560 40934
rect 33508 40870 33560 40876
rect 33046 39808 33102 39817
rect 33046 39743 33102 39752
rect 33060 39506 33088 39743
rect 33048 39500 33100 39506
rect 33048 39442 33100 39448
rect 33060 39302 33088 39442
rect 33048 39296 33100 39302
rect 33048 39238 33100 39244
rect 32864 38412 32916 38418
rect 32864 38354 32916 38360
rect 32772 38276 32824 38282
rect 32772 38218 32824 38224
rect 32784 37330 32812 38218
rect 33152 38214 33180 40870
rect 33336 40458 33364 40870
rect 33232 40452 33284 40458
rect 33232 40394 33284 40400
rect 33324 40452 33376 40458
rect 33324 40394 33376 40400
rect 33244 40338 33272 40394
rect 33520 40390 33548 40870
rect 33704 40662 33732 41482
rect 33888 41478 33916 41618
rect 34072 41478 34100 41686
rect 34348 41682 34376 41958
rect 34336 41676 34388 41682
rect 34336 41618 34388 41624
rect 33876 41472 33928 41478
rect 33876 41414 33928 41420
rect 34060 41472 34112 41478
rect 34060 41414 34112 41420
rect 33692 40656 33744 40662
rect 33692 40598 33744 40604
rect 33508 40384 33560 40390
rect 33428 40344 33508 40372
rect 33428 40338 33456 40344
rect 33244 40310 33456 40338
rect 33508 40326 33560 40332
rect 33704 39982 33732 40598
rect 33888 40118 33916 41414
rect 34440 41206 34468 42094
rect 35532 42016 35584 42022
rect 35532 41958 35584 41964
rect 35544 41818 35572 41958
rect 35532 41812 35584 41818
rect 35532 41754 35584 41760
rect 38016 41812 38068 41818
rect 38016 41754 38068 41760
rect 34704 41744 34756 41750
rect 34704 41686 34756 41692
rect 34428 41200 34480 41206
rect 34428 41142 34480 41148
rect 34612 40520 34664 40526
rect 34612 40462 34664 40468
rect 33876 40112 33928 40118
rect 33876 40054 33928 40060
rect 34428 40044 34480 40050
rect 34428 39986 34480 39992
rect 33692 39976 33744 39982
rect 34440 39953 34468 39986
rect 33692 39918 33744 39924
rect 34426 39944 34482 39953
rect 34336 39908 34388 39914
rect 34426 39879 34482 39888
rect 34336 39850 34388 39856
rect 33968 39636 34020 39642
rect 33968 39578 34020 39584
rect 33508 39432 33560 39438
rect 33508 39374 33560 39380
rect 33232 39296 33284 39302
rect 33232 39238 33284 39244
rect 33244 38350 33272 39238
rect 33520 38826 33548 39374
rect 33980 39302 34008 39578
rect 34348 39506 34376 39850
rect 34336 39500 34388 39506
rect 34336 39442 34388 39448
rect 34520 39432 34572 39438
rect 34520 39374 34572 39380
rect 33876 39296 33928 39302
rect 33876 39238 33928 39244
rect 33968 39296 34020 39302
rect 33968 39238 34020 39244
rect 33888 38962 33916 39238
rect 34532 39030 34560 39374
rect 34624 39302 34652 40462
rect 34716 40186 34744 41686
rect 38028 41682 38056 41754
rect 38672 41750 38700 42298
rect 38660 41744 38712 41750
rect 38660 41686 38712 41692
rect 38016 41676 38068 41682
rect 38016 41618 38068 41624
rect 38568 41676 38620 41682
rect 38568 41618 38620 41624
rect 37924 41608 37976 41614
rect 38580 41562 38608 41618
rect 37924 41550 37976 41556
rect 34940 41372 35236 41392
rect 34996 41370 35020 41372
rect 35076 41370 35100 41372
rect 35156 41370 35180 41372
rect 35018 41318 35020 41370
rect 35082 41318 35094 41370
rect 35156 41318 35158 41370
rect 34996 41316 35020 41318
rect 35076 41316 35100 41318
rect 35156 41316 35180 41318
rect 34940 41296 35236 41316
rect 34796 41064 34848 41070
rect 34796 41006 34848 41012
rect 37372 41064 37424 41070
rect 37372 41006 37424 41012
rect 37648 41064 37700 41070
rect 37936 41052 37964 41550
rect 38488 41534 38608 41562
rect 37700 41024 37964 41052
rect 38108 41064 38160 41070
rect 37648 41006 37700 41012
rect 34704 40180 34756 40186
rect 34704 40122 34756 40128
rect 34808 39302 34836 41006
rect 34940 40284 35236 40304
rect 34996 40282 35020 40284
rect 35076 40282 35100 40284
rect 35156 40282 35180 40284
rect 35018 40230 35020 40282
rect 35082 40230 35094 40282
rect 35156 40230 35158 40282
rect 34996 40228 35020 40230
rect 35076 40228 35100 40230
rect 35156 40228 35180 40230
rect 34940 40208 35236 40228
rect 37384 40118 37412 41006
rect 37648 40724 37700 40730
rect 37648 40666 37700 40672
rect 37660 40390 37688 40666
rect 37648 40384 37700 40390
rect 37648 40326 37700 40332
rect 37372 40112 37424 40118
rect 37372 40054 37424 40060
rect 37384 39982 37412 40054
rect 37372 39976 37424 39982
rect 37372 39918 37424 39924
rect 37556 39976 37608 39982
rect 37608 39936 37780 39964
rect 37556 39918 37608 39924
rect 37752 39846 37780 39936
rect 37740 39840 37792 39846
rect 37740 39782 37792 39788
rect 34612 39296 34664 39302
rect 34612 39238 34664 39244
rect 34796 39296 34848 39302
rect 34796 39238 34848 39244
rect 34520 39024 34572 39030
rect 34520 38966 34572 38972
rect 33876 38956 33928 38962
rect 33876 38898 33928 38904
rect 33508 38820 33560 38826
rect 33508 38762 33560 38768
rect 33232 38344 33284 38350
rect 33232 38286 33284 38292
rect 33324 38276 33376 38282
rect 33324 38218 33376 38224
rect 33140 38208 33192 38214
rect 33140 38150 33192 38156
rect 32772 37324 32824 37330
rect 32772 37266 32824 37272
rect 32680 37120 32732 37126
rect 32680 37062 32732 37068
rect 32772 36576 32824 36582
rect 32772 36518 32824 36524
rect 32784 35766 32812 36518
rect 32772 35760 32824 35766
rect 32772 35702 32824 35708
rect 33336 35154 33364 38218
rect 33600 37800 33652 37806
rect 33598 37768 33600 37777
rect 33652 37768 33654 37777
rect 33598 37703 33654 37712
rect 34808 37482 34836 39238
rect 34940 39196 35236 39216
rect 34996 39194 35020 39196
rect 35076 39194 35100 39196
rect 35156 39194 35180 39196
rect 35018 39142 35020 39194
rect 35082 39142 35094 39194
rect 35156 39142 35158 39194
rect 34996 39140 35020 39142
rect 35076 39140 35100 39142
rect 35156 39140 35180 39142
rect 34940 39120 35236 39140
rect 34940 38108 35236 38128
rect 34996 38106 35020 38108
rect 35076 38106 35100 38108
rect 35156 38106 35180 38108
rect 35018 38054 35020 38106
rect 35082 38054 35094 38106
rect 35156 38054 35158 38106
rect 34996 38052 35020 38054
rect 35076 38052 35100 38054
rect 35156 38052 35180 38054
rect 34940 38032 35236 38052
rect 37004 37868 37056 37874
rect 37004 37810 37056 37816
rect 35992 37732 36044 37738
rect 35992 37674 36044 37680
rect 34716 37454 34836 37482
rect 34716 37330 34744 37454
rect 34704 37324 34756 37330
rect 34704 37266 34756 37272
rect 34796 37324 34848 37330
rect 34796 37266 34848 37272
rect 35716 37324 35768 37330
rect 35716 37266 35768 37272
rect 34808 36922 34836 37266
rect 35440 37256 35492 37262
rect 35440 37198 35492 37204
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 35452 36922 35480 37198
rect 34796 36916 34848 36922
rect 34796 36858 34848 36864
rect 35440 36916 35492 36922
rect 35440 36858 35492 36864
rect 35728 36854 35756 37266
rect 36004 37126 36032 37674
rect 36176 37324 36228 37330
rect 36176 37266 36228 37272
rect 35992 37120 36044 37126
rect 35992 37062 36044 37068
rect 35716 36848 35768 36854
rect 35716 36790 35768 36796
rect 36004 36718 36032 37062
rect 35992 36712 36044 36718
rect 35992 36654 36044 36660
rect 35622 36272 35678 36281
rect 35622 36207 35624 36216
rect 35676 36207 35678 36216
rect 35624 36178 35676 36184
rect 35348 36168 35400 36174
rect 35348 36110 35400 36116
rect 35360 36038 35388 36110
rect 35348 36032 35400 36038
rect 35348 35974 35400 35980
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 35360 35698 35388 35974
rect 35348 35692 35400 35698
rect 35348 35634 35400 35640
rect 35360 35494 35388 35634
rect 36188 35630 36216 37266
rect 37016 36922 37044 37810
rect 37556 37800 37608 37806
rect 37556 37742 37608 37748
rect 37568 37670 37596 37742
rect 37556 37664 37608 37670
rect 37556 37606 37608 37612
rect 37740 37664 37792 37670
rect 37740 37606 37792 37612
rect 37568 37262 37596 37606
rect 37752 37398 37780 37606
rect 37740 37392 37792 37398
rect 37740 37334 37792 37340
rect 37556 37256 37608 37262
rect 37740 37256 37792 37262
rect 37608 37216 37740 37244
rect 37556 37198 37608 37204
rect 37740 37198 37792 37204
rect 37004 36916 37056 36922
rect 37004 36858 37056 36864
rect 36452 36712 36504 36718
rect 36452 36654 36504 36660
rect 36728 36712 36780 36718
rect 36728 36654 36780 36660
rect 36464 36310 36492 36654
rect 36452 36304 36504 36310
rect 36452 36246 36504 36252
rect 36176 35624 36228 35630
rect 36452 35624 36504 35630
rect 36176 35566 36228 35572
rect 36450 35592 36452 35601
rect 36504 35592 36506 35601
rect 36450 35527 36506 35536
rect 34612 35488 34664 35494
rect 34612 35430 34664 35436
rect 35348 35488 35400 35494
rect 35348 35430 35400 35436
rect 36268 35488 36320 35494
rect 36268 35430 36320 35436
rect 32312 35148 32364 35154
rect 32312 35090 32364 35096
rect 32864 35148 32916 35154
rect 32864 35090 32916 35096
rect 33324 35148 33376 35154
rect 33324 35090 33376 35096
rect 32220 34604 32272 34610
rect 32220 34546 32272 34552
rect 32324 34406 32352 35090
rect 32876 34610 32904 35090
rect 33876 35080 33928 35086
rect 33876 35022 33928 35028
rect 33508 34944 33560 34950
rect 33508 34886 33560 34892
rect 33600 34944 33652 34950
rect 33600 34886 33652 34892
rect 33520 34678 33548 34886
rect 33508 34672 33560 34678
rect 33508 34614 33560 34620
rect 32864 34604 32916 34610
rect 32864 34546 32916 34552
rect 33324 34536 33376 34542
rect 33612 34490 33640 34886
rect 33888 34649 33916 35022
rect 33874 34640 33930 34649
rect 33874 34575 33930 34584
rect 33376 34484 33640 34490
rect 33324 34478 33640 34484
rect 33336 34462 33640 34478
rect 32312 34400 32364 34406
rect 32312 34342 32364 34348
rect 31760 32904 31812 32910
rect 31760 32846 31812 32852
rect 34624 32842 34652 35430
rect 36280 35154 36308 35430
rect 36740 35154 36768 36654
rect 37844 36582 37872 41024
rect 38108 41006 38160 41012
rect 38120 40594 38148 41006
rect 38488 40730 38516 41534
rect 38752 41132 38804 41138
rect 38752 41074 38804 41080
rect 38476 40724 38528 40730
rect 38476 40666 38528 40672
rect 38108 40588 38160 40594
rect 38108 40530 38160 40536
rect 38016 40520 38068 40526
rect 38016 40462 38068 40468
rect 38028 40066 38056 40462
rect 38120 40186 38148 40530
rect 38108 40180 38160 40186
rect 38108 40122 38160 40128
rect 37936 40038 38056 40066
rect 37936 39982 37964 40038
rect 38120 39982 38148 40122
rect 38660 40044 38712 40050
rect 38660 39986 38712 39992
rect 37924 39976 37976 39982
rect 37924 39918 37976 39924
rect 38108 39976 38160 39982
rect 38672 39930 38700 39986
rect 38108 39918 38160 39924
rect 38580 39902 38700 39930
rect 38580 39817 38608 39902
rect 38566 39808 38622 39817
rect 38566 39743 38622 39752
rect 38566 39672 38622 39681
rect 38566 39607 38622 39616
rect 38580 39409 38608 39607
rect 38566 39400 38622 39409
rect 38566 39335 38622 39344
rect 38658 39128 38714 39137
rect 38658 39063 38660 39072
rect 38712 39063 38714 39072
rect 38660 39034 38712 39040
rect 38764 38962 38792 41074
rect 38752 38956 38804 38962
rect 38752 38898 38804 38904
rect 38856 38894 38884 43250
rect 39028 43104 39080 43110
rect 39028 43046 39080 43052
rect 39040 42634 39068 43046
rect 39028 42628 39080 42634
rect 39028 42570 39080 42576
rect 39040 42362 39068 42570
rect 39304 42560 39356 42566
rect 39304 42502 39356 42508
rect 39580 42560 39632 42566
rect 39580 42502 39632 42508
rect 39672 42560 39724 42566
rect 39672 42502 39724 42508
rect 39028 42356 39080 42362
rect 39028 42298 39080 42304
rect 39120 42356 39172 42362
rect 39120 42298 39172 42304
rect 39132 42265 39160 42298
rect 39118 42256 39174 42265
rect 39118 42191 39174 42200
rect 39316 42158 39344 42502
rect 39396 42288 39448 42294
rect 39396 42230 39448 42236
rect 39304 42152 39356 42158
rect 39304 42094 39356 42100
rect 39316 41970 39344 42094
rect 39224 41942 39344 41970
rect 39028 41608 39080 41614
rect 39028 41550 39080 41556
rect 39118 41576 39174 41585
rect 38936 41472 38988 41478
rect 38934 41440 38936 41449
rect 38988 41440 38990 41449
rect 38934 41375 38990 41384
rect 38936 40928 38988 40934
rect 38936 40870 38988 40876
rect 38948 40118 38976 40870
rect 38936 40112 38988 40118
rect 38936 40054 38988 40060
rect 38948 39846 38976 40054
rect 38936 39840 38988 39846
rect 38936 39782 38988 39788
rect 39040 39030 39068 41550
rect 39118 41511 39120 41520
rect 39172 41511 39174 41520
rect 39120 41482 39172 41488
rect 39120 39500 39172 39506
rect 39120 39442 39172 39448
rect 39028 39024 39080 39030
rect 39028 38966 39080 38972
rect 38844 38888 38896 38894
rect 38844 38830 38896 38836
rect 39132 38418 39160 39442
rect 39224 38418 39252 41942
rect 39408 41818 39436 42230
rect 39592 42158 39620 42502
rect 39580 42152 39632 42158
rect 39580 42094 39632 42100
rect 39684 41818 39712 42502
rect 39856 42152 39908 42158
rect 39856 42094 39908 42100
rect 39396 41812 39448 41818
rect 39396 41754 39448 41760
rect 39672 41812 39724 41818
rect 39672 41754 39724 41760
rect 39684 41682 39712 41754
rect 39672 41676 39724 41682
rect 39672 41618 39724 41624
rect 39304 40384 39356 40390
rect 39302 40352 39304 40361
rect 39356 40352 39358 40361
rect 39302 40287 39358 40296
rect 39316 40186 39344 40287
rect 39304 40180 39356 40186
rect 39304 40122 39356 40128
rect 39868 39506 39896 42094
rect 40052 42022 40080 43250
rect 40960 43104 41012 43110
rect 40960 43046 41012 43052
rect 42616 43104 42668 43110
rect 42616 43046 42668 43052
rect 40132 42764 40184 42770
rect 40132 42706 40184 42712
rect 40500 42764 40552 42770
rect 40500 42706 40552 42712
rect 40144 42022 40172 42706
rect 40408 42220 40460 42226
rect 40408 42162 40460 42168
rect 40040 42016 40092 42022
rect 40040 41958 40092 41964
rect 40132 42016 40184 42022
rect 40132 41958 40184 41964
rect 40420 39982 40448 42162
rect 40512 40118 40540 42706
rect 40972 42673 41000 43046
rect 40958 42664 41014 42673
rect 40958 42599 41014 42608
rect 40972 42362 41000 42599
rect 40960 42356 41012 42362
rect 40960 42298 41012 42304
rect 41880 42288 41932 42294
rect 41880 42230 41932 42236
rect 41892 42022 41920 42230
rect 41984 42226 42288 42242
rect 41972 42220 42300 42226
rect 42024 42214 42248 42220
rect 41972 42162 42024 42168
rect 42248 42162 42300 42168
rect 40592 42016 40644 42022
rect 40592 41958 40644 41964
rect 41880 42016 41932 42022
rect 41880 41958 41932 41964
rect 40604 41750 40632 41958
rect 40592 41744 40644 41750
rect 40592 41686 40644 41692
rect 42628 41682 42656 43046
rect 43536 42628 43588 42634
rect 43536 42570 43588 42576
rect 43548 42362 43576 42570
rect 43536 42356 43588 42362
rect 43536 42298 43588 42304
rect 43168 41812 43220 41818
rect 43168 41754 43220 41760
rect 42616 41676 42668 41682
rect 42616 41618 42668 41624
rect 42340 41608 42392 41614
rect 42340 41550 42392 41556
rect 42352 41478 42380 41550
rect 42340 41472 42392 41478
rect 42340 41414 42392 41420
rect 43180 40730 43208 41754
rect 43640 41750 43668 43726
rect 44560 43654 44588 43744
rect 45940 43654 45968 43862
rect 48780 43852 48832 43858
rect 48780 43794 48832 43800
rect 48320 43716 48372 43722
rect 48320 43658 48372 43664
rect 44548 43648 44600 43654
rect 44548 43590 44600 43596
rect 45652 43648 45704 43654
rect 45652 43590 45704 43596
rect 45928 43648 45980 43654
rect 45928 43590 45980 43596
rect 43720 42560 43772 42566
rect 43720 42502 43772 42508
rect 43628 41744 43680 41750
rect 43628 41686 43680 41692
rect 43536 41676 43588 41682
rect 43536 41618 43588 41624
rect 43444 41472 43496 41478
rect 43442 41440 43444 41449
rect 43496 41440 43498 41449
rect 43442 41375 43498 41384
rect 43168 40724 43220 40730
rect 43168 40666 43220 40672
rect 43444 40724 43496 40730
rect 43444 40666 43496 40672
rect 42708 40588 42760 40594
rect 42708 40530 42760 40536
rect 40592 40520 40644 40526
rect 40592 40462 40644 40468
rect 40500 40112 40552 40118
rect 40500 40054 40552 40060
rect 40604 40050 40632 40462
rect 40592 40044 40644 40050
rect 40592 39986 40644 39992
rect 40408 39976 40460 39982
rect 40408 39918 40460 39924
rect 40960 39976 41012 39982
rect 40960 39918 41012 39924
rect 40972 39846 41000 39918
rect 40316 39840 40368 39846
rect 40316 39782 40368 39788
rect 40960 39840 41012 39846
rect 40960 39782 41012 39788
rect 41144 39840 41196 39846
rect 41144 39782 41196 39788
rect 39488 39500 39540 39506
rect 39488 39442 39540 39448
rect 39856 39500 39908 39506
rect 39856 39442 39908 39448
rect 39948 39500 40000 39506
rect 39948 39442 40000 39448
rect 39120 38412 39172 38418
rect 39120 38354 39172 38360
rect 39212 38412 39264 38418
rect 39212 38354 39264 38360
rect 38936 38344 38988 38350
rect 38936 38286 38988 38292
rect 38948 37670 38976 38286
rect 39132 38214 39160 38354
rect 39120 38208 39172 38214
rect 39120 38150 39172 38156
rect 39028 37936 39080 37942
rect 39028 37878 39080 37884
rect 38936 37664 38988 37670
rect 38936 37606 38988 37612
rect 38108 36780 38160 36786
rect 38108 36722 38160 36728
rect 37832 36576 37884 36582
rect 37832 36518 37884 36524
rect 38120 36242 38148 36722
rect 38580 36650 38700 36666
rect 38568 36644 38700 36650
rect 38620 36638 38700 36644
rect 38568 36586 38620 36592
rect 38672 36582 38700 36638
rect 38660 36576 38712 36582
rect 38660 36518 38712 36524
rect 38108 36236 38160 36242
rect 38108 36178 38160 36184
rect 38948 36174 38976 37606
rect 38936 36168 38988 36174
rect 38936 36110 38988 36116
rect 38948 35290 38976 36110
rect 38936 35284 38988 35290
rect 38936 35226 38988 35232
rect 36820 35216 36872 35222
rect 36818 35184 36820 35193
rect 36872 35184 36874 35193
rect 36268 35148 36320 35154
rect 36268 35090 36320 35096
rect 36636 35148 36688 35154
rect 36636 35090 36688 35096
rect 36728 35148 36780 35154
rect 36818 35119 36874 35128
rect 37280 35148 37332 35154
rect 36728 35090 36780 35096
rect 37280 35090 37332 35096
rect 38016 35148 38068 35154
rect 38016 35090 38068 35096
rect 38660 35148 38712 35154
rect 38660 35090 38712 35096
rect 35624 35080 35676 35086
rect 35624 35022 35676 35028
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 34612 32836 34664 32842
rect 34612 32778 34664 32784
rect 35636 31958 35664 35022
rect 36648 34746 36676 35090
rect 37004 35080 37056 35086
rect 37004 35022 37056 35028
rect 37016 34746 37044 35022
rect 37292 34950 37320 35090
rect 37096 34944 37148 34950
rect 37096 34886 37148 34892
rect 37280 34944 37332 34950
rect 37280 34886 37332 34892
rect 36636 34740 36688 34746
rect 36636 34682 36688 34688
rect 37004 34740 37056 34746
rect 37004 34682 37056 34688
rect 37108 34406 37136 34886
rect 37096 34400 37148 34406
rect 37096 34342 37148 34348
rect 37292 32978 37320 34886
rect 38028 34542 38056 35090
rect 38672 34542 38700 35090
rect 38752 35012 38804 35018
rect 38752 34954 38804 34960
rect 38764 34921 38792 34954
rect 38750 34912 38806 34921
rect 38750 34847 38806 34856
rect 38842 34776 38898 34785
rect 39040 34746 39068 37878
rect 39304 37868 39356 37874
rect 39304 37810 39356 37816
rect 39316 36718 39344 37810
rect 39396 37732 39448 37738
rect 39396 37674 39448 37680
rect 39408 37398 39436 37674
rect 39396 37392 39448 37398
rect 39396 37334 39448 37340
rect 39304 36712 39356 36718
rect 39304 36654 39356 36660
rect 39408 36242 39436 37334
rect 39500 36922 39528 39442
rect 39580 39432 39632 39438
rect 39580 39374 39632 39380
rect 39592 38962 39620 39374
rect 39580 38956 39632 38962
rect 39580 38898 39632 38904
rect 39960 38418 39988 39442
rect 40328 39302 40356 39782
rect 40868 39432 40920 39438
rect 40868 39374 40920 39380
rect 40316 39296 40368 39302
rect 40316 39238 40368 39244
rect 40684 39296 40736 39302
rect 40684 39238 40736 39244
rect 40224 38820 40276 38826
rect 40224 38762 40276 38768
rect 39948 38412 40000 38418
rect 39948 38354 40000 38360
rect 39946 38312 40002 38321
rect 39946 38247 40002 38256
rect 39960 37874 39988 38247
rect 39948 37868 40000 37874
rect 39948 37810 40000 37816
rect 40132 37868 40184 37874
rect 40132 37810 40184 37816
rect 40144 37670 40172 37810
rect 40132 37664 40184 37670
rect 40132 37606 40184 37612
rect 39488 36916 39540 36922
rect 39488 36858 39540 36864
rect 39396 36236 39448 36242
rect 39396 36178 39448 36184
rect 40144 36145 40172 37606
rect 40236 37398 40264 38762
rect 40592 38412 40644 38418
rect 40592 38354 40644 38360
rect 40500 38344 40552 38350
rect 40498 38312 40500 38321
rect 40552 38312 40554 38321
rect 40498 38247 40554 38256
rect 40408 37800 40460 37806
rect 40408 37742 40460 37748
rect 40420 37641 40448 37742
rect 40406 37632 40462 37641
rect 40406 37567 40462 37576
rect 40316 37460 40368 37466
rect 40316 37402 40368 37408
rect 40224 37392 40276 37398
rect 40224 37334 40276 37340
rect 40328 37126 40356 37402
rect 40604 37262 40632 38354
rect 40696 38026 40724 39238
rect 40880 38214 40908 39374
rect 40960 39296 41012 39302
rect 40960 39238 41012 39244
rect 40972 38894 41000 39238
rect 40960 38888 41012 38894
rect 40960 38830 41012 38836
rect 40868 38208 40920 38214
rect 40868 38150 40920 38156
rect 40696 37998 40908 38026
rect 40880 37874 40908 37998
rect 40868 37868 40920 37874
rect 40868 37810 40920 37816
rect 41156 37806 41184 39782
rect 42720 39302 42748 40530
rect 43456 40526 43484 40666
rect 42892 40520 42944 40526
rect 42892 40462 42944 40468
rect 43444 40520 43496 40526
rect 43444 40462 43496 40468
rect 42904 40390 42932 40462
rect 42892 40384 42944 40390
rect 42892 40326 42944 40332
rect 42800 39908 42852 39914
rect 42800 39850 42852 39856
rect 42812 39438 42840 39850
rect 42800 39432 42852 39438
rect 42800 39374 42852 39380
rect 42708 39296 42760 39302
rect 42708 39238 42760 39244
rect 42904 38758 42932 40326
rect 43548 40050 43576 41618
rect 43732 41614 43760 42502
rect 43904 42152 43956 42158
rect 43904 42094 43956 42100
rect 43720 41608 43772 41614
rect 43720 41550 43772 41556
rect 43916 41138 43944 42094
rect 44180 42016 44232 42022
rect 44180 41958 44232 41964
rect 44192 41206 44220 41958
rect 44560 41682 44588 43590
rect 44916 42764 44968 42770
rect 44916 42706 44968 42712
rect 44928 42158 44956 42706
rect 44916 42152 44968 42158
rect 44916 42094 44968 42100
rect 45192 42016 45244 42022
rect 45192 41958 45244 41964
rect 44824 41812 44876 41818
rect 44824 41754 44876 41760
rect 44836 41682 44864 41754
rect 44548 41676 44600 41682
rect 44548 41618 44600 41624
rect 44824 41676 44876 41682
rect 44824 41618 44876 41624
rect 44560 41478 44588 41618
rect 44548 41472 44600 41478
rect 44548 41414 44600 41420
rect 44180 41200 44232 41206
rect 44180 41142 44232 41148
rect 43904 41132 43956 41138
rect 43904 41074 43956 41080
rect 45100 41132 45152 41138
rect 45100 41074 45152 41080
rect 43996 41064 44048 41070
rect 43996 41006 44048 41012
rect 44088 41064 44140 41070
rect 44088 41006 44140 41012
rect 44008 40390 44036 41006
rect 43996 40384 44048 40390
rect 43996 40326 44048 40332
rect 44008 40202 44036 40326
rect 43916 40174 44036 40202
rect 43536 40044 43588 40050
rect 43536 39986 43588 39992
rect 43916 39982 43944 40174
rect 44100 40066 44128 41006
rect 44180 40724 44232 40730
rect 44180 40666 44232 40672
rect 44192 40594 44220 40666
rect 44180 40588 44232 40594
rect 44180 40530 44232 40536
rect 44008 40038 44128 40066
rect 43904 39976 43956 39982
rect 43904 39918 43956 39924
rect 43628 39636 43680 39642
rect 43628 39578 43680 39584
rect 43444 39296 43496 39302
rect 43444 39238 43496 39244
rect 42892 38752 42944 38758
rect 42892 38694 42944 38700
rect 43260 38752 43312 38758
rect 43260 38694 43312 38700
rect 42982 38584 43038 38593
rect 42892 38548 42944 38554
rect 42982 38519 43038 38528
rect 42892 38490 42944 38496
rect 41234 37904 41290 37913
rect 41234 37839 41236 37848
rect 41288 37839 41290 37848
rect 41236 37810 41288 37816
rect 41144 37800 41196 37806
rect 41144 37742 41196 37748
rect 42904 37738 42932 38490
rect 42996 38486 43024 38519
rect 42984 38480 43036 38486
rect 42984 38422 43036 38428
rect 42892 37732 42944 37738
rect 42892 37674 42944 37680
rect 42800 37664 42852 37670
rect 42800 37606 42852 37612
rect 40866 37496 40922 37505
rect 41420 37460 41472 37466
rect 40866 37431 40868 37440
rect 40920 37431 40922 37440
rect 40868 37402 40920 37408
rect 41248 37420 41420 37448
rect 40592 37256 40644 37262
rect 40592 37198 40644 37204
rect 40316 37120 40368 37126
rect 40316 37062 40368 37068
rect 40500 37120 40552 37126
rect 40500 37062 40552 37068
rect 40130 36136 40186 36145
rect 40130 36071 40186 36080
rect 39672 35624 39724 35630
rect 39672 35566 39724 35572
rect 39578 35184 39634 35193
rect 39578 35119 39580 35128
rect 39632 35119 39634 35128
rect 39580 35090 39632 35096
rect 39592 34746 39620 35090
rect 39684 34746 39712 35566
rect 40512 35290 40540 37062
rect 41248 35562 41276 37420
rect 41420 37402 41472 37408
rect 42812 36394 42840 37606
rect 43168 36848 43220 36854
rect 43166 36816 43168 36825
rect 43220 36816 43222 36825
rect 43166 36751 43222 36760
rect 43272 36582 43300 38694
rect 43352 36644 43404 36650
rect 43352 36586 43404 36592
rect 43260 36576 43312 36582
rect 43260 36518 43312 36524
rect 42628 36366 42840 36394
rect 42628 35698 42656 36366
rect 43364 36242 43392 36586
rect 43456 36310 43484 39238
rect 43640 38978 43668 39578
rect 43904 39500 43956 39506
rect 43904 39442 43956 39448
rect 43916 39302 43944 39442
rect 43904 39296 43956 39302
rect 43904 39238 43956 39244
rect 43640 38950 43944 38978
rect 43812 38888 43864 38894
rect 43812 38830 43864 38836
rect 43824 38758 43852 38830
rect 43916 38758 43944 38950
rect 43812 38752 43864 38758
rect 43812 38694 43864 38700
rect 43904 38752 43956 38758
rect 43904 38694 43956 38700
rect 44008 37262 44036 40038
rect 45112 39982 45140 41074
rect 45204 41070 45232 41958
rect 45664 41750 45692 43590
rect 45940 41818 45968 43590
rect 48332 43450 48360 43658
rect 48320 43444 48372 43450
rect 48320 43386 48372 43392
rect 48792 43246 48820 43794
rect 49608 43784 49660 43790
rect 49608 43726 49660 43732
rect 48780 43240 48832 43246
rect 48780 43182 48832 43188
rect 46572 43172 46624 43178
rect 46572 43114 46624 43120
rect 46584 42770 46612 43114
rect 46572 42764 46624 42770
rect 46572 42706 46624 42712
rect 46020 42696 46072 42702
rect 46020 42638 46072 42644
rect 46112 42696 46164 42702
rect 46112 42638 46164 42644
rect 45928 41812 45980 41818
rect 45928 41754 45980 41760
rect 45652 41744 45704 41750
rect 45652 41686 45704 41692
rect 45560 41676 45612 41682
rect 45560 41618 45612 41624
rect 45192 41064 45244 41070
rect 45192 41006 45244 41012
rect 45468 41064 45520 41070
rect 45468 41006 45520 41012
rect 45192 40928 45244 40934
rect 45192 40870 45244 40876
rect 45376 40928 45428 40934
rect 45376 40870 45428 40876
rect 45204 40594 45232 40870
rect 45192 40588 45244 40594
rect 45192 40530 45244 40536
rect 45388 40390 45416 40870
rect 45376 40384 45428 40390
rect 45376 40326 45428 40332
rect 44180 39976 44232 39982
rect 45100 39976 45152 39982
rect 44180 39918 44232 39924
rect 45098 39944 45100 39953
rect 45152 39944 45154 39953
rect 44088 39296 44140 39302
rect 44088 39238 44140 39244
rect 44100 38894 44128 39238
rect 44088 38888 44140 38894
rect 44088 38830 44140 38836
rect 44088 38208 44140 38214
rect 44088 38150 44140 38156
rect 44100 37806 44128 38150
rect 44088 37800 44140 37806
rect 44088 37742 44140 37748
rect 44088 37664 44140 37670
rect 44088 37606 44140 37612
rect 44100 37262 44128 37606
rect 43996 37256 44048 37262
rect 43996 37198 44048 37204
rect 44088 37256 44140 37262
rect 44088 37198 44140 37204
rect 43444 36304 43496 36310
rect 43444 36246 43496 36252
rect 42800 36236 42852 36242
rect 42800 36178 42852 36184
rect 43352 36236 43404 36242
rect 43352 36178 43404 36184
rect 42812 35766 42840 36178
rect 43628 36168 43680 36174
rect 43628 36110 43680 36116
rect 42800 35760 42852 35766
rect 42800 35702 42852 35708
rect 42892 35760 42944 35766
rect 42892 35702 42944 35708
rect 42616 35692 42668 35698
rect 42616 35634 42668 35640
rect 42812 35630 42840 35702
rect 42800 35624 42852 35630
rect 42800 35566 42852 35572
rect 41236 35556 41288 35562
rect 41236 35498 41288 35504
rect 42064 35556 42116 35562
rect 42064 35498 42116 35504
rect 41786 35320 41842 35329
rect 40500 35284 40552 35290
rect 41786 35255 41842 35264
rect 40500 35226 40552 35232
rect 41696 35216 41748 35222
rect 41696 35158 41748 35164
rect 40592 35148 40644 35154
rect 40592 35090 40644 35096
rect 40604 34785 40632 35090
rect 40960 35080 41012 35086
rect 40960 35022 41012 35028
rect 40590 34776 40646 34785
rect 38842 34711 38844 34720
rect 38896 34711 38898 34720
rect 39028 34740 39080 34746
rect 38844 34682 38896 34688
rect 39028 34682 39080 34688
rect 39580 34740 39632 34746
rect 39580 34682 39632 34688
rect 39672 34740 39724 34746
rect 40590 34711 40646 34720
rect 39672 34682 39724 34688
rect 40972 34542 41000 35022
rect 41708 34746 41736 35158
rect 41800 35154 41828 35255
rect 41788 35148 41840 35154
rect 41788 35090 41840 35096
rect 41512 34740 41564 34746
rect 41512 34682 41564 34688
rect 41696 34740 41748 34746
rect 41696 34682 41748 34688
rect 37464 34536 37516 34542
rect 37464 34478 37516 34484
rect 38016 34536 38068 34542
rect 38016 34478 38068 34484
rect 38660 34536 38712 34542
rect 38660 34478 38712 34484
rect 40040 34536 40092 34542
rect 40040 34478 40092 34484
rect 40960 34536 41012 34542
rect 40960 34478 41012 34484
rect 37280 32972 37332 32978
rect 37280 32914 37332 32920
rect 37476 32774 37504 34478
rect 40052 33114 40080 34478
rect 41524 34474 41552 34682
rect 42076 34678 42104 35498
rect 42904 35290 42932 35702
rect 42984 35488 43036 35494
rect 42984 35430 43036 35436
rect 42892 35284 42944 35290
rect 42892 35226 42944 35232
rect 42996 35222 43024 35430
rect 42984 35216 43036 35222
rect 42984 35158 43036 35164
rect 43444 35080 43496 35086
rect 43444 35022 43496 35028
rect 42892 34740 42944 34746
rect 42892 34682 42944 34688
rect 42064 34672 42116 34678
rect 42064 34614 42116 34620
rect 42904 34626 42932 34682
rect 42904 34610 43024 34626
rect 42904 34604 43036 34610
rect 42904 34598 42984 34604
rect 42984 34546 43036 34552
rect 41512 34468 41564 34474
rect 41512 34410 41564 34416
rect 40040 33108 40092 33114
rect 40040 33050 40092 33056
rect 37464 32768 37516 32774
rect 37464 32710 37516 32716
rect 35624 31952 35676 31958
rect 35624 31894 35676 31900
rect 43456 31278 43484 35022
rect 43640 34746 43668 36110
rect 44008 35290 44036 37198
rect 44192 36854 44220 39918
rect 45098 39879 45154 39888
rect 44272 39840 44324 39846
rect 44272 39782 44324 39788
rect 45100 39840 45152 39846
rect 45100 39782 45152 39788
rect 44284 38865 44312 39782
rect 44364 39500 44416 39506
rect 44364 39442 44416 39448
rect 44916 39500 44968 39506
rect 44916 39442 44968 39448
rect 44376 39302 44404 39442
rect 44928 39302 44956 39442
rect 44364 39296 44416 39302
rect 44364 39238 44416 39244
rect 44916 39296 44968 39302
rect 44916 39238 44968 39244
rect 44928 38894 44956 39238
rect 45112 38962 45140 39782
rect 45100 38956 45152 38962
rect 45100 38898 45152 38904
rect 44916 38888 44968 38894
rect 44270 38856 44326 38865
rect 44916 38830 44968 38836
rect 44270 38791 44326 38800
rect 44916 38412 44968 38418
rect 44916 38354 44968 38360
rect 45376 38412 45428 38418
rect 45376 38354 45428 38360
rect 44456 37800 44508 37806
rect 44456 37742 44508 37748
rect 44180 36848 44232 36854
rect 44180 36790 44232 36796
rect 44088 35692 44140 35698
rect 44088 35634 44140 35640
rect 43996 35284 44048 35290
rect 43996 35226 44048 35232
rect 43628 34740 43680 34746
rect 43628 34682 43680 34688
rect 44008 34542 44036 35226
rect 44100 35222 44128 35634
rect 44088 35216 44140 35222
rect 44088 35158 44140 35164
rect 44192 35086 44220 36790
rect 44468 36718 44496 37742
rect 44928 37346 44956 38354
rect 45388 37942 45416 38354
rect 45376 37936 45428 37942
rect 45376 37878 45428 37884
rect 45480 37720 45508 41006
rect 45572 40730 45600 41618
rect 46032 41614 46060 42638
rect 46124 42294 46152 42638
rect 48872 42356 48924 42362
rect 48872 42298 48924 42304
rect 46112 42288 46164 42294
rect 46112 42230 46164 42236
rect 48884 42242 48912 42298
rect 48884 42226 49188 42242
rect 48884 42220 49200 42226
rect 48884 42214 49148 42220
rect 49148 42162 49200 42168
rect 48320 42152 48372 42158
rect 48318 42120 48320 42129
rect 48596 42152 48648 42158
rect 48372 42120 48374 42129
rect 47768 42084 47820 42090
rect 48648 42112 48728 42140
rect 48596 42094 48648 42100
rect 48318 42055 48374 42064
rect 47768 42026 47820 42032
rect 47780 41750 47808 42026
rect 48504 42016 48556 42022
rect 48504 41958 48556 41964
rect 48228 41812 48280 41818
rect 48228 41754 48280 41760
rect 47768 41744 47820 41750
rect 47768 41686 47820 41692
rect 45836 41608 45888 41614
rect 45836 41550 45888 41556
rect 46020 41608 46072 41614
rect 46020 41550 46072 41556
rect 45560 40724 45612 40730
rect 45560 40666 45612 40672
rect 45848 39438 45876 41550
rect 45928 41472 45980 41478
rect 45928 41414 45980 41420
rect 46388 41472 46440 41478
rect 46388 41414 46440 41420
rect 46572 41472 46624 41478
rect 46572 41414 46624 41420
rect 45940 41274 45968 41414
rect 45928 41268 45980 41274
rect 45928 41210 45980 41216
rect 45928 40724 45980 40730
rect 45928 40666 45980 40672
rect 45836 39432 45888 39438
rect 45836 39374 45888 39380
rect 45940 39302 45968 40666
rect 46400 40662 46428 41414
rect 46388 40656 46440 40662
rect 46388 40598 46440 40604
rect 46112 39568 46164 39574
rect 46112 39510 46164 39516
rect 45928 39296 45980 39302
rect 45928 39238 45980 39244
rect 45940 38962 45968 39238
rect 45928 38956 45980 38962
rect 45928 38898 45980 38904
rect 46124 38894 46152 39510
rect 46204 39296 46256 39302
rect 46204 39238 46256 39244
rect 46216 39030 46244 39238
rect 46204 39024 46256 39030
rect 46204 38966 46256 38972
rect 46584 38894 46612 41414
rect 48240 41154 48268 41754
rect 48516 41682 48544 41958
rect 48596 41812 48648 41818
rect 48596 41754 48648 41760
rect 48608 41721 48636 41754
rect 48594 41712 48650 41721
rect 48504 41676 48556 41682
rect 48594 41647 48650 41656
rect 48504 41618 48556 41624
rect 48240 41126 48360 41154
rect 48332 41002 48360 41126
rect 48516 41070 48544 41618
rect 48700 41138 48728 42112
rect 49514 42120 49570 42129
rect 49514 42055 49570 42064
rect 49528 42022 49556 42055
rect 49620 42022 49648 43726
rect 53392 43314 53420 45440
rect 75552 44192 75604 44198
rect 75552 44134 75604 44140
rect 54576 43852 54628 43858
rect 54576 43794 54628 43800
rect 58532 43852 58584 43858
rect 58532 43794 58584 43800
rect 59544 43852 59596 43858
rect 59544 43794 59596 43800
rect 60004 43852 60056 43858
rect 60004 43794 60056 43800
rect 74080 43852 74132 43858
rect 74080 43794 74132 43800
rect 53840 43648 53892 43654
rect 53840 43590 53892 43596
rect 53852 43450 53880 43590
rect 54588 43450 54616 43794
rect 53840 43444 53892 43450
rect 53840 43386 53892 43392
rect 54576 43444 54628 43450
rect 54576 43386 54628 43392
rect 54668 43444 54720 43450
rect 54668 43386 54720 43392
rect 53380 43308 53432 43314
rect 53380 43250 53432 43256
rect 49792 43104 49844 43110
rect 49792 43046 49844 43052
rect 52276 43104 52328 43110
rect 52276 43046 52328 43052
rect 49700 42084 49752 42090
rect 49700 42026 49752 42032
rect 49516 42016 49568 42022
rect 49516 41958 49568 41964
rect 49608 42016 49660 42022
rect 49608 41958 49660 41964
rect 48964 41608 49016 41614
rect 48964 41550 49016 41556
rect 48976 41274 49004 41550
rect 48964 41268 49016 41274
rect 48964 41210 49016 41216
rect 49056 41268 49108 41274
rect 49056 41210 49108 41216
rect 48688 41132 48740 41138
rect 48688 41074 48740 41080
rect 48976 41070 49004 41210
rect 49068 41070 49096 41210
rect 49528 41138 49556 41958
rect 49620 41682 49648 41958
rect 49608 41676 49660 41682
rect 49608 41618 49660 41624
rect 49516 41132 49568 41138
rect 49516 41074 49568 41080
rect 48504 41064 48556 41070
rect 48504 41006 48556 41012
rect 48964 41064 49016 41070
rect 48964 41006 49016 41012
rect 49056 41064 49108 41070
rect 49056 41006 49108 41012
rect 48320 40996 48372 41002
rect 48320 40938 48372 40944
rect 49332 40928 49384 40934
rect 49332 40870 49384 40876
rect 48320 40384 48372 40390
rect 48226 40352 48282 40361
rect 48320 40326 48372 40332
rect 49146 40352 49202 40361
rect 48226 40287 48282 40296
rect 48240 40186 48268 40287
rect 48228 40180 48280 40186
rect 48228 40122 48280 40128
rect 48332 40050 48360 40326
rect 49146 40287 49202 40296
rect 49160 40118 49188 40287
rect 49238 40216 49294 40225
rect 49238 40151 49294 40160
rect 49148 40112 49200 40118
rect 49054 40080 49110 40089
rect 48320 40044 48372 40050
rect 49148 40054 49200 40060
rect 49054 40015 49110 40024
rect 48320 39986 48372 39992
rect 48792 39630 49004 39658
rect 49068 39642 49096 40015
rect 49252 39982 49280 40151
rect 49344 40050 49372 40870
rect 49528 40526 49556 41074
rect 49516 40520 49568 40526
rect 49516 40462 49568 40468
rect 49712 40390 49740 42026
rect 49804 40526 49832 43046
rect 50300 43004 50596 43024
rect 50356 43002 50380 43004
rect 50436 43002 50460 43004
rect 50516 43002 50540 43004
rect 50378 42950 50380 43002
rect 50442 42950 50454 43002
rect 50516 42950 50518 43002
rect 50356 42948 50380 42950
rect 50436 42948 50460 42950
rect 50516 42948 50540 42950
rect 50300 42928 50596 42948
rect 51356 42764 51408 42770
rect 51356 42706 51408 42712
rect 50804 42628 50856 42634
rect 50804 42570 50856 42576
rect 50816 42514 50844 42570
rect 50988 42560 51040 42566
rect 50816 42508 50988 42514
rect 50816 42502 51040 42508
rect 50816 42486 51028 42502
rect 50068 42152 50120 42158
rect 50068 42094 50120 42100
rect 49882 41712 49938 41721
rect 49882 41647 49884 41656
rect 49936 41647 49938 41656
rect 49884 41618 49936 41624
rect 50080 41206 50108 42094
rect 51080 42016 51132 42022
rect 51080 41958 51132 41964
rect 50300 41916 50596 41936
rect 50356 41914 50380 41916
rect 50436 41914 50460 41916
rect 50516 41914 50540 41916
rect 50378 41862 50380 41914
rect 50442 41862 50454 41914
rect 50516 41862 50518 41914
rect 50356 41860 50380 41862
rect 50436 41860 50460 41862
rect 50516 41860 50540 41862
rect 50300 41840 50596 41860
rect 50160 41472 50212 41478
rect 50160 41414 50212 41420
rect 50068 41200 50120 41206
rect 50068 41142 50120 41148
rect 50172 40662 50200 41414
rect 50300 40828 50596 40848
rect 50356 40826 50380 40828
rect 50436 40826 50460 40828
rect 50516 40826 50540 40828
rect 50378 40774 50380 40826
rect 50442 40774 50454 40826
rect 50516 40774 50518 40826
rect 50356 40772 50380 40774
rect 50436 40772 50460 40774
rect 50516 40772 50540 40774
rect 50300 40752 50596 40772
rect 50160 40656 50212 40662
rect 50160 40598 50212 40604
rect 49792 40520 49844 40526
rect 49792 40462 49844 40468
rect 49700 40384 49752 40390
rect 49700 40326 49752 40332
rect 49790 40352 49846 40361
rect 49790 40287 49846 40296
rect 49804 40118 49832 40287
rect 49792 40112 49844 40118
rect 51092 40089 51120 41958
rect 51264 41812 51316 41818
rect 51264 41754 51316 41760
rect 51276 41274 51304 41754
rect 51264 41268 51316 41274
rect 51264 41210 51316 41216
rect 49792 40054 49844 40060
rect 51078 40080 51134 40089
rect 49332 40044 49384 40050
rect 51078 40015 51134 40024
rect 49332 39986 49384 39992
rect 49240 39976 49292 39982
rect 49240 39918 49292 39924
rect 49332 39908 49384 39914
rect 49332 39850 49384 39856
rect 49344 39681 49372 39850
rect 49608 39840 49660 39846
rect 49608 39782 49660 39788
rect 50068 39840 50120 39846
rect 50068 39782 50120 39788
rect 49330 39672 49386 39681
rect 48792 39574 48820 39630
rect 48596 39568 48648 39574
rect 48596 39510 48648 39516
rect 48780 39568 48832 39574
rect 48780 39510 48832 39516
rect 48872 39568 48924 39574
rect 48872 39510 48924 39516
rect 48976 39522 49004 39630
rect 49056 39636 49108 39642
rect 49330 39607 49386 39616
rect 49056 39578 49108 39584
rect 49424 39568 49476 39574
rect 46756 39432 46808 39438
rect 46756 39374 46808 39380
rect 46112 38888 46164 38894
rect 46112 38830 46164 38836
rect 46572 38888 46624 38894
rect 46572 38830 46624 38836
rect 46664 38888 46716 38894
rect 46664 38830 46716 38836
rect 46676 38758 46704 38830
rect 46664 38752 46716 38758
rect 46664 38694 46716 38700
rect 46768 38350 46796 39374
rect 47032 39296 47084 39302
rect 47032 39238 47084 39244
rect 47044 38962 47072 39238
rect 48226 39128 48282 39137
rect 48282 39098 48360 39114
rect 48282 39092 48372 39098
rect 48282 39086 48320 39092
rect 48226 39063 48282 39072
rect 48320 39034 48372 39040
rect 47032 38956 47084 38962
rect 47032 38898 47084 38904
rect 48412 38752 48464 38758
rect 48412 38694 48464 38700
rect 48226 38584 48282 38593
rect 48282 38554 48360 38570
rect 48282 38548 48372 38554
rect 48282 38542 48320 38548
rect 48226 38519 48282 38528
rect 48320 38490 48372 38496
rect 46756 38344 46808 38350
rect 46756 38286 46808 38292
rect 45560 38208 45612 38214
rect 45560 38150 45612 38156
rect 48320 38208 48372 38214
rect 48320 38150 48372 38156
rect 45572 37874 45600 38150
rect 45560 37868 45612 37874
rect 45560 37810 45612 37816
rect 46664 37868 46716 37874
rect 46664 37810 46716 37816
rect 46204 37800 46256 37806
rect 46204 37742 46256 37748
rect 45560 37732 45612 37738
rect 45480 37692 45560 37720
rect 45560 37674 45612 37680
rect 45834 37632 45890 37641
rect 45834 37567 45890 37576
rect 45848 37398 45876 37567
rect 46216 37505 46244 37742
rect 46676 37670 46704 37810
rect 48332 37738 48360 38150
rect 48424 37738 48452 38694
rect 48320 37732 48372 37738
rect 48320 37674 48372 37680
rect 48412 37732 48464 37738
rect 48412 37674 48464 37680
rect 46664 37664 46716 37670
rect 46664 37606 46716 37612
rect 47860 37664 47912 37670
rect 47860 37606 47912 37612
rect 46202 37496 46258 37505
rect 46202 37431 46258 37440
rect 44744 37330 44956 37346
rect 45836 37392 45888 37398
rect 45836 37334 45888 37340
rect 47872 37330 47900 37606
rect 47952 37460 48004 37466
rect 47952 37402 48004 37408
rect 47964 37330 47992 37402
rect 48608 37330 48636 39510
rect 48884 38894 48912 39510
rect 48976 39506 49372 39522
rect 49424 39510 49476 39516
rect 48976 39500 49384 39506
rect 48976 39494 49332 39500
rect 49332 39442 49384 39448
rect 48964 39432 49016 39438
rect 48962 39400 48964 39409
rect 49016 39400 49018 39409
rect 48962 39335 49018 39344
rect 48962 39128 49018 39137
rect 48962 39063 49018 39072
rect 48976 38962 49004 39063
rect 48964 38956 49016 38962
rect 48964 38898 49016 38904
rect 49436 38894 49464 39510
rect 48872 38888 48924 38894
rect 48872 38830 48924 38836
rect 49424 38888 49476 38894
rect 49424 38830 49476 38836
rect 49516 38888 49568 38894
rect 49516 38830 49568 38836
rect 49528 38758 49556 38830
rect 49516 38752 49568 38758
rect 49516 38694 49568 38700
rect 49528 37856 49556 38694
rect 49620 37874 49648 39782
rect 49792 39636 49844 39642
rect 49792 39578 49844 39584
rect 49804 39506 49832 39578
rect 49792 39500 49844 39506
rect 49792 39442 49844 39448
rect 49884 39364 49936 39370
rect 49884 39306 49936 39312
rect 49896 39030 49924 39306
rect 50080 39137 50108 39782
rect 50300 39740 50596 39760
rect 50356 39738 50380 39740
rect 50436 39738 50460 39740
rect 50516 39738 50540 39740
rect 50378 39686 50380 39738
rect 50442 39686 50454 39738
rect 50516 39686 50518 39738
rect 50356 39684 50380 39686
rect 50436 39684 50460 39686
rect 50516 39684 50540 39686
rect 50158 39672 50214 39681
rect 50300 39664 50596 39684
rect 50710 39672 50766 39681
rect 50158 39607 50160 39616
rect 50212 39607 50214 39616
rect 50710 39607 50712 39616
rect 50160 39578 50212 39584
rect 50764 39607 50766 39616
rect 50804 39636 50856 39642
rect 50712 39578 50764 39584
rect 50804 39578 50856 39584
rect 50436 39568 50488 39574
rect 50436 39510 50488 39516
rect 50448 39438 50476 39510
rect 50724 39506 50752 39578
rect 50712 39500 50764 39506
rect 50712 39442 50764 39448
rect 50436 39432 50488 39438
rect 50436 39374 50488 39380
rect 50066 39128 50122 39137
rect 50066 39063 50122 39072
rect 50448 39030 50476 39374
rect 50724 39030 50752 39442
rect 50816 39409 50844 39578
rect 50802 39400 50858 39409
rect 50802 39335 50858 39344
rect 49884 39024 49936 39030
rect 49884 38966 49936 38972
rect 50436 39024 50488 39030
rect 50436 38966 50488 38972
rect 50712 39024 50764 39030
rect 50712 38966 50764 38972
rect 51080 38956 51132 38962
rect 51080 38898 51132 38904
rect 50300 38652 50596 38672
rect 50356 38650 50380 38652
rect 50436 38650 50460 38652
rect 50516 38650 50540 38652
rect 50378 38598 50380 38650
rect 50442 38598 50454 38650
rect 50516 38598 50518 38650
rect 50356 38596 50380 38598
rect 50436 38596 50460 38598
rect 50516 38596 50540 38598
rect 50300 38576 50596 38596
rect 50342 38448 50398 38457
rect 50068 38412 50120 38418
rect 50342 38383 50344 38392
rect 50068 38354 50120 38360
rect 50396 38383 50398 38392
rect 50344 38354 50396 38360
rect 49884 38344 49936 38350
rect 50080 38321 50108 38354
rect 50252 38344 50304 38350
rect 49884 38286 49936 38292
rect 50066 38312 50122 38321
rect 49792 38276 49844 38282
rect 49792 38218 49844 38224
rect 49804 38010 49832 38218
rect 49896 38010 49924 38286
rect 50252 38286 50304 38292
rect 50066 38247 50122 38256
rect 50264 38214 50292 38286
rect 50252 38208 50304 38214
rect 50252 38150 50304 38156
rect 50710 38040 50766 38049
rect 49792 38004 49844 38010
rect 49792 37946 49844 37952
rect 49884 38004 49936 38010
rect 50710 37975 50766 37984
rect 49884 37946 49936 37952
rect 49160 37828 49556 37856
rect 49608 37868 49660 37874
rect 48964 37392 49016 37398
rect 48964 37334 49016 37340
rect 44732 37324 44956 37330
rect 44784 37318 44956 37324
rect 44732 37266 44784 37272
rect 44456 36712 44508 36718
rect 44456 36654 44508 36660
rect 44468 35766 44496 36654
rect 44928 36310 44956 37318
rect 47860 37324 47912 37330
rect 47860 37266 47912 37272
rect 47952 37324 48004 37330
rect 47952 37266 48004 37272
rect 48596 37324 48648 37330
rect 48596 37266 48648 37272
rect 48688 37324 48740 37330
rect 48688 37266 48740 37272
rect 48504 37120 48556 37126
rect 48504 37062 48556 37068
rect 48044 36848 48096 36854
rect 48042 36816 48044 36825
rect 48096 36816 48098 36825
rect 48516 36786 48544 37062
rect 48700 36786 48728 37266
rect 48976 37233 49004 37334
rect 48962 37224 49018 37233
rect 48962 37159 49018 37168
rect 49160 37126 49188 37828
rect 49608 37810 49660 37816
rect 50724 37806 50752 37975
rect 50712 37800 50764 37806
rect 50712 37742 50764 37748
rect 50300 37564 50596 37584
rect 50356 37562 50380 37564
rect 50436 37562 50460 37564
rect 50516 37562 50540 37564
rect 50378 37510 50380 37562
rect 50442 37510 50454 37562
rect 50516 37510 50518 37562
rect 50356 37508 50380 37510
rect 50436 37508 50460 37510
rect 50516 37508 50540 37510
rect 50300 37488 50596 37508
rect 51092 37346 51120 38898
rect 51262 38312 51318 38321
rect 51262 38247 51318 38256
rect 51276 38010 51304 38247
rect 51172 38004 51224 38010
rect 51172 37946 51224 37952
rect 51264 38004 51316 38010
rect 51264 37946 51316 37952
rect 51184 37466 51212 37946
rect 51368 37874 51396 42706
rect 51448 40384 51500 40390
rect 51448 40326 51500 40332
rect 51460 39098 51488 40326
rect 51816 39976 51868 39982
rect 51816 39918 51868 39924
rect 52000 39976 52052 39982
rect 52052 39936 52132 39964
rect 52000 39918 52052 39924
rect 51538 39808 51594 39817
rect 51538 39743 51594 39752
rect 51552 39642 51580 39743
rect 51540 39636 51592 39642
rect 51540 39578 51592 39584
rect 51828 39522 51856 39918
rect 52104 39846 52132 39936
rect 52092 39840 52144 39846
rect 52092 39782 52144 39788
rect 51828 39494 52040 39522
rect 52104 39506 52132 39782
rect 51632 39432 51684 39438
rect 51630 39400 51632 39409
rect 51908 39432 51960 39438
rect 51684 39400 51686 39409
rect 51908 39374 51960 39380
rect 51630 39335 51686 39344
rect 51448 39092 51500 39098
rect 51448 39034 51500 39040
rect 51448 38752 51500 38758
rect 51920 38729 51948 39374
rect 52012 38944 52040 39494
rect 52092 39500 52144 39506
rect 52092 39442 52144 39448
rect 52184 39432 52236 39438
rect 52184 39374 52236 39380
rect 52196 39098 52224 39374
rect 52184 39092 52236 39098
rect 52184 39034 52236 39040
rect 52092 38956 52144 38962
rect 52012 38916 52092 38944
rect 52092 38898 52144 38904
rect 51448 38694 51500 38700
rect 51906 38720 51962 38729
rect 51460 38486 51488 38694
rect 51906 38655 51962 38664
rect 51448 38480 51500 38486
rect 51448 38422 51500 38428
rect 51814 38448 51870 38457
rect 51814 38383 51870 38392
rect 51448 38208 51500 38214
rect 51448 38150 51500 38156
rect 51356 37868 51408 37874
rect 51356 37810 51408 37816
rect 51172 37460 51224 37466
rect 51172 37402 51224 37408
rect 50068 37324 50120 37330
rect 50068 37266 50120 37272
rect 50804 37324 50856 37330
rect 51092 37318 51212 37346
rect 50804 37266 50856 37272
rect 49148 37120 49200 37126
rect 49148 37062 49200 37068
rect 49240 37120 49292 37126
rect 49240 37062 49292 37068
rect 48042 36751 48098 36760
rect 48504 36780 48556 36786
rect 48504 36722 48556 36728
rect 48688 36780 48740 36786
rect 48688 36722 48740 36728
rect 49252 36718 49280 37062
rect 49792 36916 49844 36922
rect 49792 36858 49844 36864
rect 47308 36712 47360 36718
rect 47308 36654 47360 36660
rect 49240 36712 49292 36718
rect 49240 36654 49292 36660
rect 47320 36378 47348 36654
rect 48320 36576 48372 36582
rect 48320 36518 48372 36524
rect 49148 36576 49200 36582
rect 49148 36518 49200 36524
rect 47308 36372 47360 36378
rect 47308 36314 47360 36320
rect 44916 36304 44968 36310
rect 44916 36246 44968 36252
rect 44456 35760 44508 35766
rect 44456 35702 44508 35708
rect 47766 35320 47822 35329
rect 48332 35306 48360 36518
rect 48780 36032 48832 36038
rect 48780 35974 48832 35980
rect 48792 35698 48820 35974
rect 48780 35692 48832 35698
rect 48780 35634 48832 35640
rect 48792 35494 48820 35634
rect 48872 35556 48924 35562
rect 48872 35498 48924 35504
rect 48780 35488 48832 35494
rect 48780 35430 48832 35436
rect 47766 35255 47822 35264
rect 48044 35284 48096 35290
rect 47780 35222 47808 35255
rect 48240 35278 48360 35306
rect 48240 35272 48268 35278
rect 48096 35244 48268 35272
rect 48044 35226 48096 35232
rect 46572 35216 46624 35222
rect 46572 35158 46624 35164
rect 47768 35216 47820 35222
rect 47768 35158 47820 35164
rect 44364 35148 44416 35154
rect 44284 35108 44364 35136
rect 44180 35080 44232 35086
rect 44180 35022 44232 35028
rect 44284 35018 44312 35108
rect 44416 35108 44588 35136
rect 44364 35090 44416 35096
rect 44272 35012 44324 35018
rect 44272 34954 44324 34960
rect 44560 34610 44588 35108
rect 46584 34950 46612 35158
rect 46756 35080 46808 35086
rect 46756 35022 46808 35028
rect 46768 34950 46796 35022
rect 46572 34944 46624 34950
rect 46572 34886 46624 34892
rect 46756 34944 46808 34950
rect 46848 34944 46900 34950
rect 46756 34886 46808 34892
rect 46846 34912 46848 34921
rect 46900 34912 46902 34921
rect 44548 34604 44600 34610
rect 44548 34546 44600 34552
rect 43996 34536 44048 34542
rect 43996 34478 44048 34484
rect 46584 33794 46612 34886
rect 46572 33788 46624 33794
rect 46572 33730 46624 33736
rect 46768 32298 46796 34886
rect 46846 34847 46902 34856
rect 48792 34134 48820 35430
rect 48884 35086 48912 35498
rect 48964 35488 49016 35494
rect 48964 35430 49016 35436
rect 48872 35080 48924 35086
rect 48872 35022 48924 35028
rect 48780 34128 48832 34134
rect 48780 34070 48832 34076
rect 48976 32638 49004 35430
rect 49160 35154 49188 36518
rect 49252 35630 49280 36654
rect 49516 36032 49568 36038
rect 49516 35974 49568 35980
rect 49240 35624 49292 35630
rect 49240 35566 49292 35572
rect 49422 35592 49478 35601
rect 49422 35527 49478 35536
rect 49148 35148 49200 35154
rect 49148 35090 49200 35096
rect 49436 34950 49464 35527
rect 49528 35170 49556 35974
rect 49804 35766 49832 36858
rect 49976 36236 50028 36242
rect 49976 36178 50028 36184
rect 49882 35864 49938 35873
rect 49882 35799 49938 35808
rect 49792 35760 49844 35766
rect 49792 35702 49844 35708
rect 49896 35290 49924 35799
rect 49988 35630 50016 36178
rect 49976 35624 50028 35630
rect 49976 35566 50028 35572
rect 50080 35476 50108 37266
rect 50816 37210 50844 37266
rect 50816 37182 51120 37210
rect 50804 37120 50856 37126
rect 50804 37062 50856 37068
rect 50436 36848 50488 36854
rect 50434 36816 50436 36825
rect 50712 36848 50764 36854
rect 50488 36816 50490 36825
rect 50712 36790 50764 36796
rect 50434 36751 50490 36760
rect 50300 36476 50596 36496
rect 50356 36474 50380 36476
rect 50436 36474 50460 36476
rect 50516 36474 50540 36476
rect 50378 36422 50380 36474
rect 50442 36422 50454 36474
rect 50516 36422 50518 36474
rect 50356 36420 50380 36422
rect 50436 36420 50460 36422
rect 50516 36420 50540 36422
rect 50300 36400 50596 36420
rect 50724 36310 50752 36790
rect 50816 36786 50844 37062
rect 50804 36780 50856 36786
rect 50804 36722 50856 36728
rect 50896 36644 50948 36650
rect 50896 36586 50948 36592
rect 50712 36304 50764 36310
rect 50712 36246 50764 36252
rect 50160 36236 50212 36242
rect 50160 36178 50212 36184
rect 50344 36236 50396 36242
rect 50344 36178 50396 36184
rect 49988 35448 50108 35476
rect 49988 35290 50016 35448
rect 49884 35284 49936 35290
rect 49884 35226 49936 35232
rect 49976 35284 50028 35290
rect 49976 35226 50028 35232
rect 49528 35154 49648 35170
rect 49528 35148 49660 35154
rect 49528 35142 49608 35148
rect 49608 35090 49660 35096
rect 49620 34950 49648 35090
rect 49988 35086 50016 35226
rect 50172 35136 50200 36178
rect 50356 36038 50384 36178
rect 50344 36032 50396 36038
rect 50344 35974 50396 35980
rect 50712 35624 50764 35630
rect 50712 35566 50764 35572
rect 50724 35494 50752 35566
rect 50908 35562 50936 36586
rect 51092 36310 51120 37182
rect 51184 36786 51212 37318
rect 51172 36780 51224 36786
rect 51172 36722 51224 36728
rect 51460 36718 51488 38150
rect 51828 37806 51856 38383
rect 52288 37890 52316 43046
rect 53852 42838 53880 43386
rect 54680 43246 54708 43386
rect 54668 43240 54720 43246
rect 54588 43200 54668 43228
rect 53840 42832 53892 42838
rect 53840 42774 53892 42780
rect 53748 42764 53800 42770
rect 53748 42706 53800 42712
rect 52368 42560 52420 42566
rect 52368 42502 52420 42508
rect 53104 42560 53156 42566
rect 53104 42502 53156 42508
rect 52380 42158 52408 42502
rect 52368 42152 52420 42158
rect 52368 42094 52420 42100
rect 53116 41682 53144 42502
rect 53760 42362 53788 42706
rect 53748 42356 53800 42362
rect 53748 42298 53800 42304
rect 54484 42152 54536 42158
rect 54220 42100 54484 42106
rect 54220 42094 54536 42100
rect 54220 42078 54524 42094
rect 54220 42022 54248 42078
rect 54208 42016 54260 42022
rect 54208 41958 54260 41964
rect 53104 41676 53156 41682
rect 53104 41618 53156 41624
rect 53288 41676 53340 41682
rect 53288 41618 53340 41624
rect 53300 41274 53328 41618
rect 53288 41268 53340 41274
rect 53288 41210 53340 41216
rect 52644 41064 52696 41070
rect 52644 41006 52696 41012
rect 52656 40526 52684 41006
rect 54588 40934 54616 43200
rect 54668 43182 54720 43188
rect 58440 43104 58492 43110
rect 58440 43046 58492 43052
rect 54668 42764 54720 42770
rect 54668 42706 54720 42712
rect 57152 42764 57204 42770
rect 57152 42706 57204 42712
rect 57336 42764 57388 42770
rect 57336 42706 57388 42712
rect 58348 42764 58400 42770
rect 58348 42706 58400 42712
rect 54680 42158 54708 42706
rect 54852 42696 54904 42702
rect 54852 42638 54904 42644
rect 54864 42158 54892 42638
rect 55680 42560 55732 42566
rect 55680 42502 55732 42508
rect 55692 42158 55720 42502
rect 57164 42158 57192 42706
rect 54668 42152 54720 42158
rect 54668 42094 54720 42100
rect 54852 42152 54904 42158
rect 54852 42094 54904 42100
rect 55680 42152 55732 42158
rect 55680 42094 55732 42100
rect 57152 42152 57204 42158
rect 57152 42094 57204 42100
rect 54668 42016 54720 42022
rect 54668 41958 54720 41964
rect 55956 42016 56008 42022
rect 55956 41958 56008 41964
rect 54576 40928 54628 40934
rect 54576 40870 54628 40876
rect 52644 40520 52696 40526
rect 52644 40462 52696 40468
rect 52920 40520 52972 40526
rect 52920 40462 52972 40468
rect 52368 39976 52420 39982
rect 52368 39918 52420 39924
rect 52380 39137 52408 39918
rect 52644 39908 52696 39914
rect 52644 39850 52696 39856
rect 52656 39681 52684 39850
rect 52826 39808 52882 39817
rect 52826 39743 52882 39752
rect 52642 39672 52698 39681
rect 52642 39607 52698 39616
rect 52656 39506 52684 39607
rect 52840 39506 52868 39743
rect 52644 39500 52696 39506
rect 52644 39442 52696 39448
rect 52828 39500 52880 39506
rect 52828 39442 52880 39448
rect 52366 39128 52422 39137
rect 52366 39063 52422 39072
rect 52552 39024 52604 39030
rect 52552 38966 52604 38972
rect 52460 38956 52512 38962
rect 52460 38898 52512 38904
rect 52472 38486 52500 38898
rect 52460 38480 52512 38486
rect 52460 38422 52512 38428
rect 52460 38344 52512 38350
rect 52460 38286 52512 38292
rect 52104 37862 52316 37890
rect 51540 37800 51592 37806
rect 51540 37742 51592 37748
rect 51816 37800 51868 37806
rect 51816 37742 51868 37748
rect 51552 37398 51580 37742
rect 51540 37392 51592 37398
rect 51540 37334 51592 37340
rect 51448 36712 51500 36718
rect 51448 36654 51500 36660
rect 51080 36304 51132 36310
rect 51080 36246 51132 36252
rect 51172 36032 51224 36038
rect 51172 35974 51224 35980
rect 50896 35556 50948 35562
rect 50896 35498 50948 35504
rect 50712 35488 50764 35494
rect 50908 35465 50936 35498
rect 51184 35494 51212 35974
rect 51356 35760 51408 35766
rect 51356 35702 51408 35708
rect 51172 35488 51224 35494
rect 50712 35430 50764 35436
rect 50894 35456 50950 35465
rect 50300 35388 50596 35408
rect 51172 35430 51224 35436
rect 50894 35391 50950 35400
rect 50356 35386 50380 35388
rect 50436 35386 50460 35388
rect 50516 35386 50540 35388
rect 50378 35334 50380 35386
rect 50442 35334 50454 35386
rect 50516 35334 50518 35386
rect 50356 35332 50380 35334
rect 50436 35332 50460 35334
rect 50516 35332 50540 35334
rect 50300 35312 50596 35332
rect 50252 35148 50304 35154
rect 50172 35108 50252 35136
rect 50252 35090 50304 35096
rect 51368 35086 51396 35702
rect 49976 35080 50028 35086
rect 49976 35022 50028 35028
rect 51356 35080 51408 35086
rect 51356 35022 51408 35028
rect 49424 34944 49476 34950
rect 49424 34886 49476 34892
rect 49608 34944 49660 34950
rect 49608 34886 49660 34892
rect 48964 32632 49016 32638
rect 48964 32574 49016 32580
rect 49620 32502 49648 34886
rect 49976 34400 50028 34406
rect 49976 34342 50028 34348
rect 49988 33862 50016 34342
rect 50300 34300 50596 34320
rect 50356 34298 50380 34300
rect 50436 34298 50460 34300
rect 50516 34298 50540 34300
rect 50378 34246 50380 34298
rect 50442 34246 50454 34298
rect 50516 34246 50518 34298
rect 50356 34244 50380 34246
rect 50436 34244 50460 34246
rect 50516 34244 50540 34246
rect 50300 34224 50596 34244
rect 49976 33856 50028 33862
rect 49976 33798 50028 33804
rect 49608 32496 49660 32502
rect 49608 32438 49660 32444
rect 46756 32292 46808 32298
rect 46756 32234 46808 32240
rect 51552 31890 51580 37334
rect 51632 37120 51684 37126
rect 51632 37062 51684 37068
rect 51644 36242 51672 37062
rect 51724 36576 51776 36582
rect 51724 36518 51776 36524
rect 51908 36576 51960 36582
rect 51908 36518 51960 36524
rect 51736 36417 51764 36518
rect 51722 36408 51778 36417
rect 51722 36343 51778 36352
rect 51816 36372 51868 36378
rect 51816 36314 51868 36320
rect 51632 36236 51684 36242
rect 51632 36178 51684 36184
rect 51644 35290 51672 36178
rect 51722 35864 51778 35873
rect 51722 35799 51778 35808
rect 51736 35562 51764 35799
rect 51724 35556 51776 35562
rect 51724 35498 51776 35504
rect 51632 35284 51684 35290
rect 51632 35226 51684 35232
rect 51828 35086 51856 36314
rect 51816 35080 51868 35086
rect 51816 35022 51868 35028
rect 51828 34921 51856 35022
rect 51814 34912 51870 34921
rect 51814 34847 51870 34856
rect 51920 34610 51948 36518
rect 52000 35488 52052 35494
rect 52000 35430 52052 35436
rect 52012 35290 52040 35430
rect 52000 35284 52052 35290
rect 52000 35226 52052 35232
rect 52000 35080 52052 35086
rect 52000 35022 52052 35028
rect 52012 34950 52040 35022
rect 52000 34944 52052 34950
rect 52000 34886 52052 34892
rect 51908 34604 51960 34610
rect 51908 34546 51960 34552
rect 51816 34536 51868 34542
rect 51814 34504 51816 34513
rect 51868 34504 51870 34513
rect 51814 34439 51870 34448
rect 52104 33454 52132 37862
rect 52472 37806 52500 38286
rect 52368 37800 52420 37806
rect 52368 37742 52420 37748
rect 52460 37800 52512 37806
rect 52460 37742 52512 37748
rect 52380 37398 52408 37742
rect 52460 37664 52512 37670
rect 52460 37606 52512 37612
rect 52368 37392 52420 37398
rect 52368 37334 52420 37340
rect 52472 36786 52500 37606
rect 52564 37330 52592 38966
rect 52734 38856 52790 38865
rect 52656 38814 52734 38842
rect 52552 37324 52604 37330
rect 52552 37266 52604 37272
rect 52460 36780 52512 36786
rect 52460 36722 52512 36728
rect 52460 36644 52512 36650
rect 52460 36586 52512 36592
rect 52472 35601 52500 36586
rect 52458 35592 52514 35601
rect 52458 35527 52514 35536
rect 52368 35488 52420 35494
rect 52368 35430 52420 35436
rect 52380 35222 52408 35430
rect 52368 35216 52420 35222
rect 52368 35158 52420 35164
rect 52656 34678 52684 38814
rect 52734 38791 52790 38800
rect 52932 38457 52960 40462
rect 53102 40216 53158 40225
rect 54588 40202 54616 40870
rect 54680 40662 54708 41958
rect 55968 41721 55996 41958
rect 55034 41712 55090 41721
rect 55954 41712 56010 41721
rect 55034 41647 55036 41656
rect 55088 41647 55090 41656
rect 55128 41676 55180 41682
rect 55036 41618 55088 41624
rect 57348 41682 57376 42706
rect 58360 42673 58388 42706
rect 58346 42664 58402 42673
rect 58452 42634 58480 43046
rect 58346 42599 58402 42608
rect 58440 42628 58492 42634
rect 58440 42570 58492 42576
rect 58544 42294 58572 43794
rect 59084 43648 59136 43654
rect 59084 43590 59136 43596
rect 59096 43314 59124 43590
rect 59084 43308 59136 43314
rect 59084 43250 59136 43256
rect 59360 43240 59412 43246
rect 59360 43182 59412 43188
rect 59372 42702 59400 43182
rect 59360 42696 59412 42702
rect 59556 42673 59584 43794
rect 59912 43104 59964 43110
rect 59912 43046 59964 43052
rect 59360 42638 59412 42644
rect 59542 42664 59598 42673
rect 58900 42628 58952 42634
rect 59542 42599 59598 42608
rect 59636 42628 59688 42634
rect 58900 42570 58952 42576
rect 59636 42570 59688 42576
rect 58532 42288 58584 42294
rect 58912 42276 58940 42570
rect 59176 42288 59228 42294
rect 58912 42248 59176 42276
rect 58532 42230 58584 42236
rect 59176 42230 59228 42236
rect 59188 41682 59216 42230
rect 59648 42158 59676 42570
rect 59636 42152 59688 42158
rect 59636 42094 59688 42100
rect 59924 41682 59952 43046
rect 60016 42838 60044 43794
rect 61016 43784 61068 43790
rect 61016 43726 61068 43732
rect 60004 42832 60056 42838
rect 60004 42774 60056 42780
rect 60016 42158 60044 42774
rect 61028 42770 61056 43726
rect 74092 43654 74120 43794
rect 74264 43716 74316 43722
rect 74264 43658 74316 43664
rect 74080 43648 74132 43654
rect 74080 43590 74132 43596
rect 65660 43548 65956 43568
rect 65716 43546 65740 43548
rect 65796 43546 65820 43548
rect 65876 43546 65900 43548
rect 65738 43494 65740 43546
rect 65802 43494 65814 43546
rect 65876 43494 65878 43546
rect 65716 43492 65740 43494
rect 65796 43492 65820 43494
rect 65876 43492 65900 43494
rect 65660 43472 65956 43492
rect 61108 43444 61160 43450
rect 61108 43386 61160 43392
rect 60464 42764 60516 42770
rect 60464 42706 60516 42712
rect 61016 42764 61068 42770
rect 61016 42706 61068 42712
rect 60186 42664 60242 42673
rect 60186 42599 60242 42608
rect 60096 42560 60148 42566
rect 60096 42502 60148 42508
rect 60004 42152 60056 42158
rect 60004 42094 60056 42100
rect 55954 41647 55956 41656
rect 55128 41618 55180 41624
rect 56008 41647 56010 41656
rect 57336 41676 57388 41682
rect 55956 41618 56008 41624
rect 57336 41618 57388 41624
rect 59176 41676 59228 41682
rect 59176 41618 59228 41624
rect 59912 41676 59964 41682
rect 59912 41618 59964 41624
rect 55036 41472 55088 41478
rect 55036 41414 55088 41420
rect 55048 41070 55076 41414
rect 55036 41064 55088 41070
rect 55036 41006 55088 41012
rect 54852 40928 54904 40934
rect 54852 40870 54904 40876
rect 54668 40656 54720 40662
rect 54668 40598 54720 40604
rect 54864 40594 54892 40870
rect 54852 40588 54904 40594
rect 54852 40530 54904 40536
rect 55140 40526 55168 41618
rect 55864 41608 55916 41614
rect 55968 41587 55996 41618
rect 60016 41596 60044 42094
rect 60108 42022 60136 42502
rect 60200 42158 60228 42599
rect 60188 42152 60240 42158
rect 60188 42094 60240 42100
rect 60476 42022 60504 42706
rect 61028 42158 61056 42706
rect 61120 42702 61148 43386
rect 73896 43308 73948 43314
rect 73896 43250 73948 43256
rect 63868 43240 63920 43246
rect 63868 43182 63920 43188
rect 66904 43240 66956 43246
rect 66904 43182 66956 43188
rect 67364 43240 67416 43246
rect 67364 43182 67416 43188
rect 70584 43240 70636 43246
rect 70584 43182 70636 43188
rect 63776 43104 63828 43110
rect 63776 43046 63828 43052
rect 63788 42770 63816 43046
rect 63776 42764 63828 42770
rect 63776 42706 63828 42712
rect 61108 42696 61160 42702
rect 61108 42638 61160 42644
rect 63592 42560 63644 42566
rect 63592 42502 63644 42508
rect 61200 42288 61252 42294
rect 61200 42230 61252 42236
rect 61212 42158 61240 42230
rect 60648 42152 60700 42158
rect 60648 42094 60700 42100
rect 61016 42152 61068 42158
rect 61016 42094 61068 42100
rect 61200 42152 61252 42158
rect 61200 42094 61252 42100
rect 60096 42016 60148 42022
rect 60096 41958 60148 41964
rect 60464 42016 60516 42022
rect 60464 41958 60516 41964
rect 60096 41608 60148 41614
rect 60016 41568 60096 41596
rect 55864 41550 55916 41556
rect 60660 41585 60688 42094
rect 60096 41550 60148 41556
rect 60646 41576 60702 41585
rect 55876 41274 55904 41550
rect 60646 41511 60702 41520
rect 55864 41268 55916 41274
rect 55864 41210 55916 41216
rect 63500 40928 63552 40934
rect 63500 40870 63552 40876
rect 57796 40588 57848 40594
rect 57796 40530 57848 40536
rect 58808 40588 58860 40594
rect 58808 40530 58860 40536
rect 62948 40588 63000 40594
rect 62948 40530 63000 40536
rect 55128 40520 55180 40526
rect 55128 40462 55180 40468
rect 57704 40384 57756 40390
rect 57704 40326 57756 40332
rect 54588 40174 54708 40202
rect 53102 40151 53158 40160
rect 53116 40050 53144 40151
rect 53104 40044 53156 40050
rect 53104 39986 53156 39992
rect 53288 39976 53340 39982
rect 53288 39918 53340 39924
rect 54576 39976 54628 39982
rect 54576 39918 54628 39924
rect 53300 39302 53328 39918
rect 53380 39840 53432 39846
rect 53380 39782 53432 39788
rect 53564 39840 53616 39846
rect 53564 39782 53616 39788
rect 53392 39302 53420 39782
rect 53576 39370 53604 39782
rect 53656 39636 53708 39642
rect 53656 39578 53708 39584
rect 53668 39409 53696 39578
rect 54300 39500 54352 39506
rect 54300 39442 54352 39448
rect 53654 39400 53710 39409
rect 53564 39364 53616 39370
rect 53654 39335 53710 39344
rect 53564 39306 53616 39312
rect 54312 39302 54340 39442
rect 53288 39296 53340 39302
rect 53288 39238 53340 39244
rect 53380 39296 53432 39302
rect 53380 39238 53432 39244
rect 54116 39296 54168 39302
rect 54300 39296 54352 39302
rect 54168 39256 54248 39284
rect 54116 39238 54168 39244
rect 54220 39030 54248 39256
rect 54300 39238 54352 39244
rect 54208 39024 54260 39030
rect 54312 39001 54340 39238
rect 54208 38966 54260 38972
rect 54298 38992 54354 39001
rect 54298 38927 54354 38936
rect 54208 38888 54260 38894
rect 54260 38836 54432 38842
rect 54208 38830 54432 38836
rect 54220 38814 54432 38830
rect 54404 38808 54432 38814
rect 54484 38820 54536 38826
rect 54404 38780 54484 38808
rect 54484 38762 54536 38768
rect 54588 38758 54616 39918
rect 54680 39846 54708 40174
rect 54668 39840 54720 39846
rect 54668 39782 54720 39788
rect 56784 39840 56836 39846
rect 56784 39782 56836 39788
rect 54680 39574 54708 39782
rect 54668 39568 54720 39574
rect 56796 39545 56824 39782
rect 54668 39510 54720 39516
rect 56782 39536 56838 39545
rect 54680 39438 54708 39510
rect 56782 39471 56838 39480
rect 54668 39432 54720 39438
rect 57716 39409 57744 40326
rect 57808 39794 57836 40530
rect 58072 39976 58124 39982
rect 58072 39918 58124 39924
rect 58624 39976 58676 39982
rect 58624 39918 58676 39924
rect 57888 39840 57940 39846
rect 57808 39788 57888 39794
rect 57808 39782 57940 39788
rect 57808 39766 57928 39782
rect 57808 39574 57836 39766
rect 57796 39568 57848 39574
rect 57796 39510 57848 39516
rect 58084 39506 58112 39918
rect 58072 39500 58124 39506
rect 58072 39442 58124 39448
rect 58164 39500 58216 39506
rect 58164 39442 58216 39448
rect 57980 39432 58032 39438
rect 54668 39374 54720 39380
rect 57702 39400 57758 39409
rect 56692 39364 56744 39370
rect 57980 39374 58032 39380
rect 57702 39335 57758 39344
rect 56692 39306 56744 39312
rect 54668 39296 54720 39302
rect 54668 39238 54720 39244
rect 54680 38962 54708 39238
rect 56230 39128 56286 39137
rect 56230 39063 56286 39072
rect 54668 38956 54720 38962
rect 54668 38898 54720 38904
rect 54208 38752 54260 38758
rect 54208 38694 54260 38700
rect 54576 38752 54628 38758
rect 54576 38694 54628 38700
rect 52918 38448 52974 38457
rect 52918 38383 52974 38392
rect 53196 38208 53248 38214
rect 53196 38150 53248 38156
rect 53288 38208 53340 38214
rect 53288 38150 53340 38156
rect 53208 38049 53236 38150
rect 53194 38040 53250 38049
rect 53194 37975 53250 37984
rect 52920 37664 52972 37670
rect 52920 37606 52972 37612
rect 52932 37398 52960 37606
rect 52920 37392 52972 37398
rect 52920 37334 52972 37340
rect 52736 36712 52788 36718
rect 52736 36654 52788 36660
rect 52748 36242 52776 36654
rect 52736 36236 52788 36242
rect 52736 36178 52788 36184
rect 53300 35154 53328 38150
rect 53380 37868 53432 37874
rect 53380 37810 53432 37816
rect 53392 37670 53420 37810
rect 54220 37670 54248 38694
rect 55034 38448 55090 38457
rect 55034 38383 55090 38392
rect 53380 37664 53432 37670
rect 53380 37606 53432 37612
rect 54208 37664 54260 37670
rect 54208 37606 54260 37612
rect 53392 36310 53420 37606
rect 53840 37256 53892 37262
rect 53840 37198 53892 37204
rect 53852 36718 53880 37198
rect 53840 36712 53892 36718
rect 53840 36654 53892 36660
rect 53748 36644 53800 36650
rect 53748 36586 53800 36592
rect 53380 36304 53432 36310
rect 53380 36246 53432 36252
rect 53760 35329 53788 36586
rect 54116 36576 54168 36582
rect 54116 36518 54168 36524
rect 54128 36242 54156 36518
rect 54116 36236 54168 36242
rect 54116 36178 54168 36184
rect 54220 36122 54248 37606
rect 54944 37256 54996 37262
rect 54944 37198 54996 37204
rect 54852 37120 54904 37126
rect 54852 37062 54904 37068
rect 54864 36378 54892 37062
rect 54956 36922 54984 37198
rect 54944 36916 54996 36922
rect 54944 36858 54996 36864
rect 55048 36786 55076 38383
rect 56244 38350 56272 39063
rect 56612 38758 56640 38789
rect 56600 38752 56652 38758
rect 56598 38720 56600 38729
rect 56652 38720 56654 38729
rect 56598 38655 56654 38664
rect 56612 38418 56640 38655
rect 56704 38486 56732 39306
rect 57992 39302 58020 39374
rect 57980 39296 58032 39302
rect 57980 39238 58032 39244
rect 57992 38894 58020 39238
rect 57980 38888 58032 38894
rect 57980 38830 58032 38836
rect 58176 38758 58204 39442
rect 58254 39400 58310 39409
rect 58254 39335 58310 39344
rect 58268 38894 58296 39335
rect 58636 38894 58664 39918
rect 58820 39914 58848 40530
rect 59176 40384 59228 40390
rect 59176 40326 59228 40332
rect 58808 39908 58860 39914
rect 58808 39850 58860 39856
rect 59188 39574 59216 40326
rect 62960 39982 62988 40530
rect 62948 39976 63000 39982
rect 62948 39918 63000 39924
rect 63512 39914 63540 40870
rect 63604 40390 63632 42502
rect 63880 42226 63908 43182
rect 66260 43172 66312 43178
rect 66260 43114 66312 43120
rect 66272 42770 66300 43114
rect 66916 42906 66944 43182
rect 66904 42900 66956 42906
rect 66904 42842 66956 42848
rect 67376 42770 67404 43182
rect 67916 43172 67968 43178
rect 67916 43114 67968 43120
rect 69204 43172 69256 43178
rect 69204 43114 69256 43120
rect 66260 42764 66312 42770
rect 66260 42706 66312 42712
rect 67364 42764 67416 42770
rect 67364 42706 67416 42712
rect 64236 42560 64288 42566
rect 64236 42502 64288 42508
rect 65524 42560 65576 42566
rect 65524 42502 65576 42508
rect 67272 42560 67324 42566
rect 67272 42502 67324 42508
rect 63868 42220 63920 42226
rect 63868 42162 63920 42168
rect 64248 41478 64276 42502
rect 64420 42220 64472 42226
rect 64420 42162 64472 42168
rect 64432 41750 64460 42162
rect 64512 42152 64564 42158
rect 64512 42094 64564 42100
rect 64880 42152 64932 42158
rect 64880 42094 64932 42100
rect 65064 42152 65116 42158
rect 65064 42094 65116 42100
rect 64420 41744 64472 41750
rect 64420 41686 64472 41692
rect 64328 41676 64380 41682
rect 64328 41618 64380 41624
rect 64236 41472 64288 41478
rect 64236 41414 64288 41420
rect 63776 41268 63828 41274
rect 63776 41210 63828 41216
rect 63788 40594 63816 41210
rect 64340 40934 64368 41618
rect 64524 41274 64552 42094
rect 64892 41750 64920 42094
rect 64880 41744 64932 41750
rect 64880 41686 64932 41692
rect 64512 41268 64564 41274
rect 64512 41210 64564 41216
rect 64892 41070 64920 41686
rect 65076 41682 65104 42094
rect 65064 41676 65116 41682
rect 65064 41618 65116 41624
rect 64880 41064 64932 41070
rect 64880 41006 64932 41012
rect 65076 41002 65104 41618
rect 65432 41608 65484 41614
rect 65432 41550 65484 41556
rect 65064 40996 65116 41002
rect 65064 40938 65116 40944
rect 64328 40928 64380 40934
rect 64328 40870 64380 40876
rect 64340 40594 64736 40610
rect 63776 40588 63828 40594
rect 63776 40530 63828 40536
rect 64328 40588 64748 40594
rect 64380 40582 64696 40588
rect 64328 40530 64380 40536
rect 64696 40530 64748 40536
rect 64604 40520 64656 40526
rect 64972 40520 65024 40526
rect 64604 40462 64656 40468
rect 64892 40480 64972 40508
rect 63592 40384 63644 40390
rect 63592 40326 63644 40332
rect 64616 39982 64644 40462
rect 64892 40186 64920 40480
rect 64972 40462 65024 40468
rect 65444 40390 65472 41550
rect 64972 40384 65024 40390
rect 64972 40326 65024 40332
rect 65432 40384 65484 40390
rect 65432 40326 65484 40332
rect 64984 40186 65012 40326
rect 64880 40180 64932 40186
rect 64880 40122 64932 40128
rect 64972 40180 65024 40186
rect 64972 40122 65024 40128
rect 64144 39976 64196 39982
rect 64604 39976 64656 39982
rect 64196 39924 64276 39930
rect 64144 39918 64276 39924
rect 64604 39918 64656 39924
rect 61200 39908 61252 39914
rect 61200 39850 61252 39856
rect 63500 39908 63552 39914
rect 64156 39902 64276 39918
rect 63500 39850 63552 39856
rect 59084 39568 59136 39574
rect 59084 39510 59136 39516
rect 59176 39568 59228 39574
rect 59176 39510 59228 39516
rect 59096 39370 59124 39510
rect 59084 39364 59136 39370
rect 59084 39306 59136 39312
rect 59188 39302 59216 39510
rect 61212 39506 61240 39850
rect 61660 39840 61712 39846
rect 61660 39782 61712 39788
rect 60924 39500 60976 39506
rect 60924 39442 60976 39448
rect 61200 39500 61252 39506
rect 61200 39442 61252 39448
rect 59452 39364 59504 39370
rect 59452 39306 59504 39312
rect 59176 39296 59228 39302
rect 59176 39238 59228 39244
rect 59360 39296 59412 39302
rect 59360 39238 59412 39244
rect 59372 38894 59400 39238
rect 58256 38888 58308 38894
rect 58256 38830 58308 38836
rect 58624 38888 58676 38894
rect 58624 38830 58676 38836
rect 59084 38888 59136 38894
rect 59084 38830 59136 38836
rect 59360 38888 59412 38894
rect 59360 38830 59412 38836
rect 58164 38752 58216 38758
rect 58164 38694 58216 38700
rect 56692 38480 56744 38486
rect 56692 38422 56744 38428
rect 58176 38418 58204 38694
rect 56600 38412 56652 38418
rect 56600 38354 56652 38360
rect 58164 38412 58216 38418
rect 58164 38354 58216 38360
rect 58992 38412 59044 38418
rect 58992 38354 59044 38360
rect 56232 38344 56284 38350
rect 56232 38286 56284 38292
rect 57428 38344 57480 38350
rect 57428 38286 57480 38292
rect 57980 38344 58032 38350
rect 57980 38286 58032 38292
rect 56244 37806 56272 38286
rect 57440 38214 57468 38286
rect 56692 38208 56744 38214
rect 56692 38150 56744 38156
rect 57428 38208 57480 38214
rect 57428 38150 57480 38156
rect 56324 37936 56376 37942
rect 56324 37878 56376 37884
rect 56232 37800 56284 37806
rect 56232 37742 56284 37748
rect 56336 37398 56364 37878
rect 56324 37392 56376 37398
rect 56324 37334 56376 37340
rect 55128 37324 55180 37330
rect 55128 37266 55180 37272
rect 55036 36780 55088 36786
rect 55036 36722 55088 36728
rect 54852 36372 54904 36378
rect 54852 36314 54904 36320
rect 54128 36094 54248 36122
rect 53746 35320 53802 35329
rect 53746 35255 53802 35264
rect 53288 35148 53340 35154
rect 53288 35090 53340 35096
rect 53840 35148 53892 35154
rect 53840 35090 53892 35096
rect 53012 34944 53064 34950
rect 53012 34886 53064 34892
rect 52644 34672 52696 34678
rect 52644 34614 52696 34620
rect 53024 34610 53052 34886
rect 53012 34604 53064 34610
rect 53012 34546 53064 34552
rect 52552 34468 52604 34474
rect 52552 34410 52604 34416
rect 52368 34400 52420 34406
rect 52368 34342 52420 34348
rect 52380 34134 52408 34342
rect 52368 34128 52420 34134
rect 52368 34070 52420 34076
rect 52092 33448 52144 33454
rect 52092 33390 52144 33396
rect 52092 33108 52144 33114
rect 52092 33050 52144 33056
rect 52104 32026 52132 33050
rect 52092 32020 52144 32026
rect 52092 31962 52144 31968
rect 51540 31884 51592 31890
rect 51540 31826 51592 31832
rect 51080 31680 51132 31686
rect 51080 31622 51132 31628
rect 43444 31272 43496 31278
rect 43444 31214 43496 31220
rect 51092 30841 51120 31622
rect 52000 31612 52052 31618
rect 52000 31554 52052 31560
rect 51078 30832 51134 30841
rect 51078 30767 51134 30776
rect 52012 25537 52040 31554
rect 51998 25528 52054 25537
rect 51998 25463 52054 25472
rect 28448 21956 28500 21962
rect 28448 21898 28500 21904
rect 27068 17332 27120 17338
rect 27068 17274 27120 17280
rect 26884 16516 26936 16522
rect 26884 16458 26936 16464
rect 24216 11348 24268 11354
rect 24216 11290 24268 11296
rect 22468 9920 22520 9926
rect 22468 9862 22520 9868
rect 22480 9042 22508 9862
rect 22468 9036 22520 9042
rect 22468 8978 22520 8984
rect 22284 8492 22336 8498
rect 22284 8434 22336 8440
rect 22296 7546 22324 8434
rect 22284 7540 22336 7546
rect 22284 7482 22336 7488
rect 22284 7336 22336 7342
rect 22284 7278 22336 7284
rect 22296 7002 22324 7278
rect 22284 6996 22336 7002
rect 22284 6938 22336 6944
rect 21732 5908 21784 5914
rect 21732 5850 21784 5856
rect 21364 5704 21416 5710
rect 21364 5646 21416 5652
rect 21376 5370 21404 5646
rect 23480 5568 23532 5574
rect 23480 5510 23532 5516
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 21364 5364 21416 5370
rect 21364 5306 21416 5312
rect 20720 5160 20772 5166
rect 20720 5102 20772 5108
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 23492 4865 23520 5510
rect 52104 4865 52132 31962
rect 52368 31408 52420 31414
rect 52368 31350 52420 31356
rect 52380 22817 52408 31350
rect 52366 22808 52422 22817
rect 52366 22743 52422 22752
rect 23478 4856 23534 4865
rect 23478 4791 23534 4800
rect 52090 4856 52146 4865
rect 52090 4791 52146 4800
rect 19340 4684 19392 4690
rect 19340 4626 19392 4632
rect 12992 4548 13044 4554
rect 12992 4490 13044 4496
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 13188 4146 13216 4422
rect 13176 4140 13228 4146
rect 13176 4082 13228 4088
rect 11336 4072 11388 4078
rect 11336 4014 11388 4020
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 10508 3188 10560 3194
rect 10508 3130 10560 3136
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 7564 2984 7616 2990
rect 7564 2926 7616 2932
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 10060 2650 10088 2790
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 52564 950 52592 34410
rect 53852 31482 53880 35090
rect 54024 34944 54076 34950
rect 54024 34886 54076 34892
rect 53932 34604 53984 34610
rect 53932 34546 53984 34552
rect 53840 31476 53892 31482
rect 53840 31418 53892 31424
rect 53840 31340 53892 31346
rect 53840 31282 53892 31288
rect 53852 30229 53880 31282
rect 53944 31074 53972 34546
rect 54036 31346 54064 34886
rect 54128 34785 54156 36094
rect 55140 35766 55168 37266
rect 56232 37256 56284 37262
rect 56230 37224 56232 37233
rect 56284 37224 56286 37233
rect 56230 37159 56286 37168
rect 56048 36848 56100 36854
rect 56048 36790 56100 36796
rect 55312 36780 55364 36786
rect 55312 36722 55364 36728
rect 54576 35760 54628 35766
rect 54576 35702 54628 35708
rect 55128 35760 55180 35766
rect 55128 35702 55180 35708
rect 55218 35728 55274 35737
rect 54484 35556 54536 35562
rect 54484 35498 54536 35504
rect 54208 34944 54260 34950
rect 54208 34886 54260 34892
rect 54114 34776 54170 34785
rect 54114 34711 54170 34720
rect 54128 34542 54156 34711
rect 54116 34536 54168 34542
rect 54116 34478 54168 34484
rect 54116 31476 54168 31482
rect 54116 31418 54168 31424
rect 54024 31340 54076 31346
rect 54024 31282 54076 31288
rect 53932 31068 53984 31074
rect 53932 31010 53984 31016
rect 53838 30220 53894 30229
rect 53838 30155 53894 30164
rect 53840 29504 53892 29510
rect 53838 29472 53840 29481
rect 53892 29472 53894 29481
rect 53838 29407 53894 29416
rect 53838 28180 53894 28189
rect 53944 28166 53972 31010
rect 54024 30524 54076 30530
rect 54024 30466 54076 30472
rect 53894 28138 53972 28166
rect 53838 28115 53894 28124
rect 53840 27600 53892 27606
rect 53840 27542 53892 27548
rect 53852 26761 53880 27542
rect 53838 26752 53894 26761
rect 53838 26687 53894 26696
rect 53840 24268 53892 24274
rect 53838 24236 53840 24245
rect 53892 24236 53894 24245
rect 53838 24171 53894 24180
rect 54036 24086 54064 30466
rect 54128 27606 54156 31418
rect 54220 29510 54248 34886
rect 54300 34536 54352 34542
rect 54300 34478 54352 34484
rect 54312 31550 54340 34478
rect 54392 34468 54444 34474
rect 54392 34410 54444 34416
rect 54404 33114 54432 34410
rect 54496 33590 54524 35498
rect 54588 35494 54616 35702
rect 54944 35692 54996 35698
rect 55218 35663 55274 35672
rect 54944 35634 54996 35640
rect 54576 35488 54628 35494
rect 54576 35430 54628 35436
rect 54588 34406 54616 35430
rect 54760 34944 54812 34950
rect 54760 34886 54812 34892
rect 54852 34944 54904 34950
rect 54852 34886 54904 34892
rect 54576 34400 54628 34406
rect 54576 34342 54628 34348
rect 54484 33584 54536 33590
rect 54484 33526 54536 33532
rect 54588 33386 54616 34342
rect 54576 33380 54628 33386
rect 54576 33322 54628 33328
rect 54392 33108 54444 33114
rect 54392 33050 54444 33056
rect 54300 31544 54352 31550
rect 54300 31486 54352 31492
rect 54208 29504 54260 29510
rect 54208 29446 54260 29452
rect 54312 28422 54340 31486
rect 54300 28416 54352 28422
rect 54300 28358 54352 28364
rect 54116 27600 54168 27606
rect 54116 27542 54168 27548
rect 54772 24274 54800 34886
rect 54864 34785 54892 34886
rect 54850 34776 54906 34785
rect 54850 34711 54906 34720
rect 54956 34542 54984 35634
rect 55232 35630 55260 35663
rect 55220 35624 55272 35630
rect 55220 35566 55272 35572
rect 54852 34536 54904 34542
rect 54852 34478 54904 34484
rect 54944 34536 54996 34542
rect 54944 34478 54996 34484
rect 54864 31686 54892 34478
rect 55220 34468 55272 34474
rect 55220 34410 55272 34416
rect 54852 31680 54904 31686
rect 54852 31622 54904 31628
rect 54864 30530 54892 31622
rect 55232 31618 55260 34410
rect 55324 31822 55352 36722
rect 55956 36032 56008 36038
rect 55956 35974 56008 35980
rect 55968 35873 55996 35974
rect 55954 35864 56010 35873
rect 55954 35799 56010 35808
rect 55772 35624 55824 35630
rect 55772 35566 55824 35572
rect 55784 35465 55812 35566
rect 55770 35456 55826 35465
rect 55770 35391 55826 35400
rect 55770 35320 55826 35329
rect 55770 35255 55826 35264
rect 55784 35154 55812 35255
rect 55772 35148 55824 35154
rect 55772 35090 55824 35096
rect 55404 34536 55456 34542
rect 55404 34478 55456 34484
rect 55312 31816 55364 31822
rect 55312 31758 55364 31764
rect 55220 31612 55272 31618
rect 55220 31554 55272 31560
rect 55416 31414 55444 34478
rect 55968 33658 55996 35799
rect 56060 34202 56088 36790
rect 56336 36718 56364 37334
rect 56600 37256 56652 37262
rect 56600 37198 56652 37204
rect 56612 37126 56640 37198
rect 56600 37120 56652 37126
rect 56600 37062 56652 37068
rect 56612 36854 56640 37062
rect 56600 36848 56652 36854
rect 56600 36790 56652 36796
rect 56704 36786 56732 38150
rect 57440 37806 57468 38150
rect 57428 37800 57480 37806
rect 57428 37742 57480 37748
rect 57440 37641 57468 37742
rect 57426 37632 57482 37641
rect 57426 37567 57482 37576
rect 57992 37466 58020 38286
rect 59004 38010 59032 38354
rect 59096 38350 59124 38830
rect 59464 38826 59492 39306
rect 59544 39296 59596 39302
rect 59544 39238 59596 39244
rect 59556 38865 59584 39238
rect 60648 39024 60700 39030
rect 60646 38992 60648 39001
rect 60740 39024 60792 39030
rect 60700 38992 60702 39001
rect 60740 38966 60792 38972
rect 60646 38927 60702 38936
rect 59542 38856 59598 38865
rect 59452 38820 59504 38826
rect 59542 38791 59598 38800
rect 59452 38762 59504 38768
rect 59728 38412 59780 38418
rect 59728 38354 59780 38360
rect 59084 38344 59136 38350
rect 59084 38286 59136 38292
rect 58992 38004 59044 38010
rect 58992 37946 59044 37952
rect 59740 37874 59768 38354
rect 60648 38004 60700 38010
rect 60648 37946 60700 37952
rect 59910 37904 59966 37913
rect 59728 37868 59780 37874
rect 60660 37890 60688 37946
rect 60752 37890 60780 38966
rect 59910 37839 59912 37848
rect 59728 37810 59780 37816
rect 59964 37839 59966 37848
rect 60464 37868 60516 37874
rect 59912 37810 59964 37816
rect 60660 37862 60780 37890
rect 60464 37810 60516 37816
rect 58256 37800 58308 37806
rect 58256 37742 58308 37748
rect 57980 37460 58032 37466
rect 57980 37402 58032 37408
rect 57336 37324 57388 37330
rect 57520 37324 57572 37330
rect 57388 37284 57520 37312
rect 57336 37266 57388 37272
rect 57520 37266 57572 37272
rect 58268 36854 58296 37742
rect 60476 37466 60504 37810
rect 60464 37460 60516 37466
rect 60464 37402 60516 37408
rect 60740 36916 60792 36922
rect 60740 36858 60792 36864
rect 58256 36848 58308 36854
rect 56782 36816 56838 36825
rect 56692 36780 56744 36786
rect 56782 36751 56838 36760
rect 57886 36816 57942 36825
rect 58532 36848 58584 36854
rect 58256 36790 58308 36796
rect 58452 36808 58532 36836
rect 57886 36751 57942 36760
rect 56692 36722 56744 36728
rect 56796 36718 56824 36751
rect 56324 36712 56376 36718
rect 56324 36654 56376 36660
rect 56784 36712 56836 36718
rect 56784 36654 56836 36660
rect 57900 36650 57928 36751
rect 57888 36644 57940 36650
rect 57888 36586 57940 36592
rect 58162 36408 58218 36417
rect 58162 36343 58218 36352
rect 56244 36242 56640 36258
rect 56244 36236 56652 36242
rect 56244 36230 56600 36236
rect 56244 36038 56272 36230
rect 56600 36178 56652 36184
rect 57796 36168 57848 36174
rect 57796 36110 57848 36116
rect 57978 36136 58034 36145
rect 56232 36032 56284 36038
rect 56232 35974 56284 35980
rect 56140 35556 56192 35562
rect 56140 35498 56192 35504
rect 56152 35290 56180 35498
rect 56140 35284 56192 35290
rect 56140 35226 56192 35232
rect 56244 35170 56272 35974
rect 56966 35864 57022 35873
rect 56966 35799 57022 35808
rect 56322 35728 56378 35737
rect 56980 35698 57008 35799
rect 57520 35760 57572 35766
rect 57520 35702 57572 35708
rect 56322 35663 56378 35672
rect 56600 35692 56652 35698
rect 56336 35290 56364 35663
rect 56600 35634 56652 35640
rect 56968 35692 57020 35698
rect 56968 35634 57020 35640
rect 56612 35465 56640 35634
rect 57532 35630 57560 35702
rect 57520 35624 57572 35630
rect 57520 35566 57572 35572
rect 56598 35456 56654 35465
rect 56598 35391 56654 35400
rect 56324 35284 56376 35290
rect 56324 35226 56376 35232
rect 56508 35284 56560 35290
rect 56508 35226 56560 35232
rect 56244 35142 56456 35170
rect 56428 35086 56456 35142
rect 56140 35080 56192 35086
rect 56140 35022 56192 35028
rect 56416 35080 56468 35086
rect 56416 35022 56468 35028
rect 56152 34610 56180 35022
rect 56428 34950 56456 35022
rect 56416 34944 56468 34950
rect 56416 34886 56468 34892
rect 56140 34604 56192 34610
rect 56140 34546 56192 34552
rect 56048 34196 56100 34202
rect 56048 34138 56100 34144
rect 56428 34066 56456 34886
rect 56520 34513 56548 35226
rect 56968 35148 57020 35154
rect 56968 35090 57020 35096
rect 56980 34950 57008 35090
rect 57808 34950 57836 36110
rect 57978 36071 58034 36080
rect 57992 35850 58020 36071
rect 57900 35834 58020 35850
rect 57888 35828 58020 35834
rect 57940 35822 58020 35828
rect 57888 35770 57940 35776
rect 57980 35216 58032 35222
rect 57980 35158 58032 35164
rect 57992 35086 58020 35158
rect 57980 35080 58032 35086
rect 57980 35022 58032 35028
rect 56968 34944 57020 34950
rect 56966 34912 56968 34921
rect 57796 34944 57848 34950
rect 57020 34912 57022 34921
rect 57796 34886 57848 34892
rect 56966 34847 57022 34856
rect 57520 34536 57572 34542
rect 56506 34504 56562 34513
rect 57520 34478 57572 34484
rect 57888 34536 57940 34542
rect 57980 34536 58032 34542
rect 57940 34496 57980 34524
rect 57888 34478 57940 34484
rect 58176 34513 58204 36343
rect 58452 36038 58480 36808
rect 58532 36790 58584 36796
rect 58624 36576 58676 36582
rect 58624 36518 58676 36524
rect 60752 36530 60780 36858
rect 58636 36242 58664 36518
rect 60752 36502 60872 36530
rect 60844 36378 60872 36502
rect 60740 36372 60792 36378
rect 60740 36314 60792 36320
rect 60832 36372 60884 36378
rect 60832 36314 60884 36320
rect 60752 36258 60780 36314
rect 60936 36258 60964 39442
rect 61108 39364 61160 39370
rect 61108 39306 61160 39312
rect 61120 39098 61148 39306
rect 61108 39092 61160 39098
rect 61108 39034 61160 39040
rect 61016 39024 61068 39030
rect 61016 38966 61068 38972
rect 61028 38894 61056 38966
rect 61672 38894 61700 39782
rect 63512 39438 63540 39850
rect 64248 39846 64276 39902
rect 64144 39840 64196 39846
rect 64144 39782 64196 39788
rect 64236 39840 64288 39846
rect 64236 39782 64288 39788
rect 61844 39432 61896 39438
rect 61844 39374 61896 39380
rect 63500 39432 63552 39438
rect 63500 39374 63552 39380
rect 61856 38894 61884 39374
rect 64156 39030 64184 39782
rect 65340 39296 65392 39302
rect 65340 39238 65392 39244
rect 64144 39024 64196 39030
rect 64144 38966 64196 38972
rect 61016 38888 61068 38894
rect 61016 38830 61068 38836
rect 61200 38888 61252 38894
rect 61200 38830 61252 38836
rect 61660 38888 61712 38894
rect 61660 38830 61712 38836
rect 61844 38888 61896 38894
rect 61844 38830 61896 38836
rect 61106 38584 61162 38593
rect 61106 38519 61108 38528
rect 61160 38519 61162 38528
rect 61108 38490 61160 38496
rect 58532 36236 58584 36242
rect 58532 36178 58584 36184
rect 58624 36236 58676 36242
rect 60752 36230 60964 36258
rect 58624 36178 58676 36184
rect 58440 36032 58492 36038
rect 58440 35974 58492 35980
rect 58452 35154 58480 35974
rect 58440 35148 58492 35154
rect 58440 35090 58492 35096
rect 57980 34478 58032 34484
rect 58162 34504 58218 34513
rect 56506 34439 56562 34448
rect 56784 34468 56836 34474
rect 56784 34410 56836 34416
rect 56416 34060 56468 34066
rect 56416 34002 56468 34008
rect 55956 33652 56008 33658
rect 55956 33594 56008 33600
rect 55404 31408 55456 31414
rect 55404 31350 55456 31356
rect 56796 31278 56824 34410
rect 57532 34406 57560 34478
rect 58162 34439 58218 34448
rect 58176 34406 58204 34439
rect 58544 34406 58572 36178
rect 59820 36168 59872 36174
rect 59820 36110 59872 36116
rect 58624 36032 58676 36038
rect 58624 35974 58676 35980
rect 58808 36032 58860 36038
rect 58808 35974 58860 35980
rect 58636 35698 58664 35974
rect 58624 35692 58676 35698
rect 58624 35634 58676 35640
rect 58622 35320 58678 35329
rect 58622 35255 58678 35264
rect 58636 35154 58664 35255
rect 58820 35222 58848 35974
rect 59084 35624 59136 35630
rect 59082 35592 59084 35601
rect 59136 35592 59138 35601
rect 59082 35527 59138 35536
rect 58900 35488 58952 35494
rect 58898 35456 58900 35465
rect 58952 35456 58954 35465
rect 58898 35391 58954 35400
rect 59832 35290 59860 36110
rect 59820 35284 59872 35290
rect 59820 35226 59872 35232
rect 58808 35216 58860 35222
rect 58808 35158 58860 35164
rect 58624 35148 58676 35154
rect 58624 35090 58676 35096
rect 58636 34950 58664 35090
rect 61212 35086 61240 38830
rect 63774 38584 63830 38593
rect 61292 38548 61344 38554
rect 63774 38519 63830 38528
rect 61292 38490 61344 38496
rect 61304 38457 61332 38490
rect 63788 38486 63816 38519
rect 63776 38480 63828 38486
rect 61290 38448 61346 38457
rect 63776 38422 63828 38428
rect 61290 38383 61346 38392
rect 62856 38412 62908 38418
rect 62856 38354 62908 38360
rect 63500 38412 63552 38418
rect 63500 38354 63552 38360
rect 61934 38312 61990 38321
rect 61934 38247 61990 38256
rect 61948 38214 61976 38247
rect 61936 38208 61988 38214
rect 61936 38150 61988 38156
rect 62120 38208 62172 38214
rect 62120 38150 62172 38156
rect 62580 38208 62632 38214
rect 62580 38150 62632 38156
rect 62132 38010 62160 38150
rect 62120 38004 62172 38010
rect 62120 37946 62172 37952
rect 62132 36650 62160 37946
rect 62592 37262 62620 38150
rect 62868 38010 62896 38354
rect 63512 38298 63540 38354
rect 63144 38270 63540 38298
rect 62856 38004 62908 38010
rect 62856 37946 62908 37952
rect 62580 37256 62632 37262
rect 62580 37198 62632 37204
rect 62592 37126 62620 37198
rect 62580 37120 62632 37126
rect 62580 37062 62632 37068
rect 62120 36644 62172 36650
rect 62120 36586 62172 36592
rect 62028 35488 62080 35494
rect 62028 35430 62080 35436
rect 61200 35080 61252 35086
rect 61200 35022 61252 35028
rect 62040 35018 62068 35430
rect 62028 35012 62080 35018
rect 62028 34954 62080 34960
rect 58624 34944 58676 34950
rect 58624 34886 58676 34892
rect 61752 34944 61804 34950
rect 61752 34886 61804 34892
rect 59084 34672 59136 34678
rect 59084 34614 59136 34620
rect 58992 34604 59044 34610
rect 58992 34546 59044 34552
rect 58900 34536 58952 34542
rect 58898 34504 58900 34513
rect 58952 34504 58954 34513
rect 58898 34439 58954 34448
rect 57520 34400 57572 34406
rect 57518 34368 57520 34377
rect 58164 34400 58216 34406
rect 57572 34368 57574 34377
rect 58164 34342 58216 34348
rect 58532 34400 58584 34406
rect 59004 34377 59032 34546
rect 59096 34542 59124 34614
rect 59084 34536 59136 34542
rect 59084 34478 59136 34484
rect 58532 34342 58584 34348
rect 58990 34368 59046 34377
rect 57518 34303 57574 34312
rect 58990 34303 59046 34312
rect 57532 34277 57560 34303
rect 61764 33998 61792 34886
rect 62488 34468 62540 34474
rect 62488 34410 62540 34416
rect 61752 33992 61804 33998
rect 61752 33934 61804 33940
rect 62500 33930 62528 34410
rect 62488 33924 62540 33930
rect 62488 33866 62540 33872
rect 62592 32434 62620 37062
rect 63144 36650 63172 38270
rect 65352 38214 65380 39238
rect 65444 38758 65472 40326
rect 65536 39030 65564 42502
rect 65660 42460 65956 42480
rect 65716 42458 65740 42460
rect 65796 42458 65820 42460
rect 65876 42458 65900 42460
rect 65738 42406 65740 42458
rect 65802 42406 65814 42458
rect 65876 42406 65878 42458
rect 65716 42404 65740 42406
rect 65796 42404 65820 42406
rect 65876 42404 65900 42406
rect 65660 42384 65956 42404
rect 66720 42288 66772 42294
rect 66720 42230 66772 42236
rect 66352 42016 66404 42022
rect 66352 41958 66404 41964
rect 66364 41750 66392 41958
rect 66352 41744 66404 41750
rect 66352 41686 66404 41692
rect 66352 41608 66404 41614
rect 66350 41576 66352 41585
rect 66404 41576 66406 41585
rect 66350 41511 66406 41520
rect 66732 41478 66760 42230
rect 67284 42158 67312 42502
rect 67376 42294 67404 42706
rect 67364 42288 67416 42294
rect 67364 42230 67416 42236
rect 67272 42152 67324 42158
rect 67272 42094 67324 42100
rect 67548 41676 67600 41682
rect 67548 41618 67600 41624
rect 66720 41472 66772 41478
rect 66720 41414 66772 41420
rect 65660 41372 65956 41392
rect 65716 41370 65740 41372
rect 65796 41370 65820 41372
rect 65876 41370 65900 41372
rect 65738 41318 65740 41370
rect 65802 41318 65814 41370
rect 65876 41318 65878 41370
rect 65716 41316 65740 41318
rect 65796 41316 65820 41318
rect 65876 41316 65900 41318
rect 65660 41296 65956 41316
rect 67560 41274 67588 41618
rect 67548 41268 67600 41274
rect 67548 41210 67600 41216
rect 66260 40928 66312 40934
rect 66180 40888 66260 40916
rect 66076 40588 66128 40594
rect 66180 40576 66208 40888
rect 66260 40870 66312 40876
rect 67364 40928 67416 40934
rect 67364 40870 67416 40876
rect 67376 40594 67404 40870
rect 67928 40594 67956 43114
rect 69216 42770 69244 43114
rect 69204 42764 69256 42770
rect 69204 42706 69256 42712
rect 70596 42226 70624 43182
rect 73252 43172 73304 43178
rect 73252 43114 73304 43120
rect 71780 43104 71832 43110
rect 71780 43046 71832 43052
rect 71228 42764 71280 42770
rect 71228 42706 71280 42712
rect 71240 42566 71268 42706
rect 71504 42628 71556 42634
rect 71504 42570 71556 42576
rect 71228 42560 71280 42566
rect 71228 42502 71280 42508
rect 70584 42220 70636 42226
rect 70584 42162 70636 42168
rect 71240 42158 71268 42502
rect 71516 42226 71544 42570
rect 71504 42220 71556 42226
rect 71504 42162 71556 42168
rect 71228 42152 71280 42158
rect 71228 42094 71280 42100
rect 69848 42084 69900 42090
rect 69848 42026 69900 42032
rect 69664 42016 69716 42022
rect 69664 41958 69716 41964
rect 69676 41818 69704 41958
rect 69664 41812 69716 41818
rect 69664 41754 69716 41760
rect 69860 41750 69888 42026
rect 71688 41812 71740 41818
rect 71688 41754 71740 41760
rect 69848 41744 69900 41750
rect 69848 41686 69900 41692
rect 71228 41268 71280 41274
rect 71228 41210 71280 41216
rect 71240 41041 71268 41210
rect 71700 41206 71728 41754
rect 71792 41682 71820 43046
rect 73264 42702 73292 43114
rect 73908 42770 73936 43250
rect 73896 42764 73948 42770
rect 73896 42706 73948 42712
rect 73252 42696 73304 42702
rect 73252 42638 73304 42644
rect 72700 42560 72752 42566
rect 72700 42502 72752 42508
rect 72712 42294 72740 42502
rect 72700 42288 72752 42294
rect 72700 42230 72752 42236
rect 73264 42226 73292 42638
rect 73436 42560 73488 42566
rect 73436 42502 73488 42508
rect 73252 42220 73304 42226
rect 73252 42162 73304 42168
rect 73252 42084 73304 42090
rect 73252 42026 73304 42032
rect 73264 41750 73292 42026
rect 73252 41744 73304 41750
rect 73252 41686 73304 41692
rect 71780 41676 71832 41682
rect 71780 41618 71832 41624
rect 73160 41676 73212 41682
rect 73160 41618 73212 41624
rect 72608 41472 72660 41478
rect 72608 41414 72660 41420
rect 71688 41200 71740 41206
rect 71688 41142 71740 41148
rect 71226 41032 71282 41041
rect 71226 40967 71282 40976
rect 72148 40928 72200 40934
rect 72148 40870 72200 40876
rect 66128 40548 66208 40576
rect 66260 40588 66312 40594
rect 66076 40530 66128 40536
rect 66260 40530 66312 40536
rect 66352 40588 66404 40594
rect 66352 40530 66404 40536
rect 67364 40588 67416 40594
rect 67364 40530 67416 40536
rect 67456 40588 67508 40594
rect 67456 40530 67508 40536
rect 67916 40588 67968 40594
rect 67916 40530 67968 40536
rect 65660 40284 65956 40304
rect 65716 40282 65740 40284
rect 65796 40282 65820 40284
rect 65876 40282 65900 40284
rect 65738 40230 65740 40282
rect 65802 40230 65814 40282
rect 65876 40230 65878 40282
rect 65716 40228 65740 40230
rect 65796 40228 65820 40230
rect 65876 40228 65900 40230
rect 65660 40208 65956 40228
rect 66272 40089 66300 40530
rect 66364 40390 66392 40530
rect 67270 40488 67326 40497
rect 67270 40423 67272 40432
rect 67324 40423 67326 40432
rect 67272 40394 67324 40400
rect 66352 40384 66404 40390
rect 66352 40326 66404 40332
rect 67364 40384 67416 40390
rect 67468 40372 67496 40530
rect 67416 40344 67496 40372
rect 67364 40326 67416 40332
rect 67548 40112 67600 40118
rect 66258 40080 66314 40089
rect 66258 40015 66314 40024
rect 66994 40080 67050 40089
rect 67548 40054 67600 40060
rect 66994 40015 67050 40024
rect 67008 39982 67036 40015
rect 66996 39976 67048 39982
rect 66996 39918 67048 39924
rect 67456 39908 67508 39914
rect 67456 39850 67508 39856
rect 65708 39840 65760 39846
rect 65708 39782 65760 39788
rect 65720 39574 65748 39782
rect 65708 39568 65760 39574
rect 65708 39510 65760 39516
rect 67468 39506 67496 39850
rect 67456 39500 67508 39506
rect 67456 39442 67508 39448
rect 67560 39370 67588 40054
rect 67928 39982 67956 40530
rect 71044 40520 71096 40526
rect 71044 40462 71096 40468
rect 70768 40112 70820 40118
rect 71056 40089 71084 40462
rect 71964 40384 72016 40390
rect 71964 40326 72016 40332
rect 70768 40054 70820 40060
rect 71042 40080 71098 40089
rect 67916 39976 67968 39982
rect 67916 39918 67968 39924
rect 70780 39846 70808 40054
rect 71042 40015 71098 40024
rect 71044 39976 71096 39982
rect 71044 39918 71096 39924
rect 67640 39840 67692 39846
rect 67640 39782 67692 39788
rect 70768 39840 70820 39846
rect 70768 39782 70820 39788
rect 67548 39364 67600 39370
rect 67548 39306 67600 39312
rect 66168 39296 66220 39302
rect 66168 39238 66220 39244
rect 65660 39196 65956 39216
rect 65716 39194 65740 39196
rect 65796 39194 65820 39196
rect 65876 39194 65900 39196
rect 65738 39142 65740 39194
rect 65802 39142 65814 39194
rect 65876 39142 65878 39194
rect 65716 39140 65740 39142
rect 65796 39140 65820 39142
rect 65876 39140 65900 39142
rect 65660 39120 65956 39140
rect 65524 39024 65576 39030
rect 65524 38966 65576 38972
rect 66180 38894 66208 39238
rect 67652 39030 67680 39782
rect 71056 39642 71084 39918
rect 71044 39636 71096 39642
rect 71044 39578 71096 39584
rect 71976 39506 72004 40326
rect 72160 40118 72188 40870
rect 72148 40112 72200 40118
rect 72148 40054 72200 40060
rect 72620 39642 72648 41414
rect 73068 41200 73120 41206
rect 73068 41142 73120 41148
rect 72976 40928 73028 40934
rect 72976 40870 73028 40876
rect 72988 40594 73016 40870
rect 73080 40746 73108 41142
rect 73172 40934 73200 41618
rect 73252 41608 73304 41614
rect 73252 41550 73304 41556
rect 73344 41608 73396 41614
rect 73344 41550 73396 41556
rect 73264 41070 73292 41550
rect 73356 41478 73384 41550
rect 73344 41472 73396 41478
rect 73344 41414 73396 41420
rect 73448 41154 73476 42502
rect 73528 41472 73580 41478
rect 73528 41414 73580 41420
rect 73540 41206 73568 41414
rect 73356 41126 73476 41154
rect 73528 41200 73580 41206
rect 73528 41142 73580 41148
rect 73252 41064 73304 41070
rect 73252 41006 73304 41012
rect 73160 40928 73212 40934
rect 73160 40870 73212 40876
rect 73080 40718 73200 40746
rect 72976 40588 73028 40594
rect 72976 40530 73028 40536
rect 73068 40588 73120 40594
rect 73068 40530 73120 40536
rect 72608 39636 72660 39642
rect 72608 39578 72660 39584
rect 71964 39500 72016 39506
rect 71964 39442 72016 39448
rect 72332 39500 72384 39506
rect 72332 39442 72384 39448
rect 67640 39024 67692 39030
rect 67546 38992 67602 39001
rect 67640 38966 67692 38972
rect 70214 38992 70270 39001
rect 67546 38927 67548 38936
rect 67600 38927 67602 38936
rect 70214 38927 70216 38936
rect 67548 38898 67600 38904
rect 70268 38927 70270 38936
rect 70216 38898 70268 38904
rect 72344 38894 72372 39442
rect 72424 39432 72476 39438
rect 72424 39374 72476 39380
rect 72436 38962 72464 39374
rect 72424 38956 72476 38962
rect 72424 38898 72476 38904
rect 65524 38888 65576 38894
rect 65524 38830 65576 38836
rect 66168 38888 66220 38894
rect 66168 38830 66220 38836
rect 69664 38888 69716 38894
rect 69664 38830 69716 38836
rect 70308 38888 70360 38894
rect 70308 38830 70360 38836
rect 71504 38888 71556 38894
rect 72332 38888 72384 38894
rect 71556 38848 71820 38876
rect 71504 38830 71556 38836
rect 65432 38752 65484 38758
rect 65432 38694 65484 38700
rect 64696 38208 64748 38214
rect 64696 38150 64748 38156
rect 65340 38208 65392 38214
rect 65340 38150 65392 38156
rect 64708 37874 64736 38150
rect 64236 37868 64288 37874
rect 64236 37810 64288 37816
rect 64696 37868 64748 37874
rect 64696 37810 64748 37816
rect 64248 37670 64276 37810
rect 64328 37800 64380 37806
rect 64328 37742 64380 37748
rect 64236 37664 64288 37670
rect 64234 37632 64236 37641
rect 64288 37632 64290 37641
rect 64234 37567 64290 37576
rect 63868 37324 63920 37330
rect 63868 37266 63920 37272
rect 63132 36644 63184 36650
rect 63132 36586 63184 36592
rect 63144 36174 63172 36586
rect 63316 36372 63368 36378
rect 63316 36314 63368 36320
rect 63328 36242 63356 36314
rect 63880 36242 63908 37266
rect 63316 36236 63368 36242
rect 63316 36178 63368 36184
rect 63868 36236 63920 36242
rect 63868 36178 63920 36184
rect 62672 36168 62724 36174
rect 62672 36110 62724 36116
rect 63132 36168 63184 36174
rect 63132 36110 63184 36116
rect 62580 32428 62632 32434
rect 62580 32370 62632 32376
rect 62684 31754 62712 36110
rect 63328 35630 63356 36178
rect 63500 36168 63552 36174
rect 63500 36110 63552 36116
rect 63512 35766 63540 36110
rect 63500 35760 63552 35766
rect 63500 35702 63552 35708
rect 63684 35760 63736 35766
rect 63684 35702 63736 35708
rect 63316 35624 63368 35630
rect 63316 35566 63368 35572
rect 62764 35148 62816 35154
rect 62764 35090 62816 35096
rect 63040 35148 63092 35154
rect 63092 35108 63172 35136
rect 63040 35090 63092 35096
rect 62776 34950 62804 35090
rect 63144 34950 63172 35108
rect 62764 34944 62816 34950
rect 62764 34886 62816 34892
rect 63132 34944 63184 34950
rect 63132 34886 63184 34892
rect 63144 34542 63172 34886
rect 63132 34536 63184 34542
rect 63132 34478 63184 34484
rect 63696 32230 63724 35702
rect 64340 35154 64368 37742
rect 65352 37670 65380 38150
rect 65432 37936 65484 37942
rect 65432 37878 65484 37884
rect 64420 37664 64472 37670
rect 64420 37606 64472 37612
rect 65340 37664 65392 37670
rect 65340 37606 65392 37612
rect 64432 36854 64460 37606
rect 64788 37120 64840 37126
rect 64788 37062 64840 37068
rect 64420 36848 64472 36854
rect 64420 36790 64472 36796
rect 64800 36786 64828 37062
rect 64788 36780 64840 36786
rect 64788 36722 64840 36728
rect 64420 36168 64472 36174
rect 64420 36110 64472 36116
rect 64432 35630 64460 36110
rect 64420 35624 64472 35630
rect 64420 35566 64472 35572
rect 64604 35624 64656 35630
rect 64604 35566 64656 35572
rect 64616 35222 64644 35566
rect 64604 35216 64656 35222
rect 64604 35158 64656 35164
rect 64328 35148 64380 35154
rect 64328 35090 64380 35096
rect 63868 34944 63920 34950
rect 63868 34886 63920 34892
rect 64512 34944 64564 34950
rect 64512 34886 64564 34892
rect 63880 34542 63908 34886
rect 63868 34536 63920 34542
rect 63868 34478 63920 34484
rect 64524 34406 64552 34886
rect 65352 34678 65380 37606
rect 65444 37398 65472 37878
rect 65432 37392 65484 37398
rect 65536 37369 65564 38830
rect 67732 38752 67784 38758
rect 67732 38694 67784 38700
rect 67744 38486 67772 38694
rect 69676 38486 69704 38830
rect 70320 38758 70348 38830
rect 70308 38752 70360 38758
rect 70308 38694 70360 38700
rect 70780 38554 71268 38570
rect 70768 38548 71280 38554
rect 70820 38542 71228 38548
rect 70768 38490 70820 38496
rect 71228 38490 71280 38496
rect 67732 38480 67784 38486
rect 67732 38422 67784 38428
rect 69664 38480 69716 38486
rect 69664 38422 69716 38428
rect 70124 38480 70176 38486
rect 70124 38422 70176 38428
rect 67824 38344 67876 38350
rect 67362 38312 67418 38321
rect 67362 38247 67364 38256
rect 67416 38247 67418 38256
rect 67468 38292 67824 38298
rect 67468 38286 67876 38292
rect 68928 38344 68980 38350
rect 68928 38286 68980 38292
rect 67468 38270 67864 38286
rect 67364 38218 67416 38224
rect 67468 38214 67496 38270
rect 67456 38208 67508 38214
rect 67456 38150 67508 38156
rect 65660 38108 65956 38128
rect 65716 38106 65740 38108
rect 65796 38106 65820 38108
rect 65876 38106 65900 38108
rect 65738 38054 65740 38106
rect 65802 38054 65814 38106
rect 65876 38054 65878 38106
rect 65716 38052 65740 38054
rect 65796 38052 65820 38054
rect 65876 38052 65900 38054
rect 65660 38032 65956 38052
rect 65432 37334 65484 37340
rect 65522 37360 65578 37369
rect 65522 37295 65578 37304
rect 67468 37194 67496 38150
rect 68940 37806 68968 38286
rect 68928 37800 68980 37806
rect 70136 37777 70164 38422
rect 71792 38350 71820 38848
rect 72332 38830 72384 38836
rect 72344 38418 72372 38830
rect 72424 38752 72476 38758
rect 72424 38694 72476 38700
rect 72332 38412 72384 38418
rect 72332 38354 72384 38360
rect 71780 38344 71832 38350
rect 71780 38286 71832 38292
rect 71596 38276 71648 38282
rect 71596 38218 71648 38224
rect 71608 37890 71636 38218
rect 71056 37874 71636 37890
rect 71056 37868 71648 37874
rect 71056 37862 71596 37868
rect 71056 37806 71084 37862
rect 71596 37810 71648 37816
rect 72436 37806 72464 38694
rect 72620 38350 72648 39578
rect 73080 38894 73108 40530
rect 73172 40526 73200 40718
rect 73160 40520 73212 40526
rect 73160 40462 73212 40468
rect 73172 40390 73200 40462
rect 73160 40384 73212 40390
rect 73160 40326 73212 40332
rect 73356 40050 73384 41126
rect 73436 41064 73488 41070
rect 73436 41006 73488 41012
rect 73448 40594 73476 41006
rect 73528 40996 73580 41002
rect 73528 40938 73580 40944
rect 73436 40588 73488 40594
rect 73436 40530 73488 40536
rect 73540 40526 73568 40938
rect 73528 40520 73580 40526
rect 73528 40462 73580 40468
rect 73344 40044 73396 40050
rect 73344 39986 73396 39992
rect 73908 39846 73936 42706
rect 74092 42566 74120 43590
rect 74172 43240 74224 43246
rect 74172 43182 74224 43188
rect 74080 42560 74132 42566
rect 74080 42502 74132 42508
rect 74184 41750 74212 43182
rect 74276 42158 74304 43658
rect 75564 43450 75592 44134
rect 81020 44092 81316 44112
rect 81076 44090 81100 44092
rect 81156 44090 81180 44092
rect 81236 44090 81260 44092
rect 81098 44038 81100 44090
rect 81162 44038 81174 44090
rect 81236 44038 81238 44090
rect 81076 44036 81100 44038
rect 81156 44036 81180 44038
rect 81236 44036 81260 44038
rect 81020 44016 81316 44036
rect 78588 43852 78640 43858
rect 78588 43794 78640 43800
rect 78864 43852 78916 43858
rect 78864 43794 78916 43800
rect 81440 43852 81492 43858
rect 81440 43794 81492 43800
rect 82360 43852 82412 43858
rect 82360 43794 82412 43800
rect 78496 43716 78548 43722
rect 78496 43658 78548 43664
rect 74632 43444 74684 43450
rect 74632 43386 74684 43392
rect 75552 43444 75604 43450
rect 75552 43386 75604 43392
rect 74540 43240 74592 43246
rect 74540 43182 74592 43188
rect 74552 42226 74580 43182
rect 74644 42770 74672 43386
rect 75564 43246 75592 43386
rect 78508 43314 78536 43658
rect 78496 43308 78548 43314
rect 78496 43250 78548 43256
rect 75552 43240 75604 43246
rect 75552 43182 75604 43188
rect 75564 42838 75592 43182
rect 75920 43104 75972 43110
rect 75920 43046 75972 43052
rect 75552 42832 75604 42838
rect 75552 42774 75604 42780
rect 74632 42764 74684 42770
rect 74632 42706 74684 42712
rect 75932 42226 75960 43046
rect 78600 42906 78628 43794
rect 78680 43784 78732 43790
rect 78680 43726 78732 43732
rect 78692 43246 78720 43726
rect 78772 43648 78824 43654
rect 78876 43602 78904 43794
rect 78824 43596 78904 43602
rect 78772 43590 78904 43596
rect 78784 43574 78904 43590
rect 78876 43246 78904 43574
rect 78680 43240 78732 43246
rect 78680 43182 78732 43188
rect 78864 43240 78916 43246
rect 78864 43182 78916 43188
rect 78772 43172 78824 43178
rect 78772 43114 78824 43120
rect 78588 42900 78640 42906
rect 78588 42842 78640 42848
rect 77668 42628 77720 42634
rect 77668 42570 77720 42576
rect 74356 42220 74408 42226
rect 74356 42162 74408 42168
rect 74540 42220 74592 42226
rect 74540 42162 74592 42168
rect 75920 42220 75972 42226
rect 75920 42162 75972 42168
rect 74264 42152 74316 42158
rect 74264 42094 74316 42100
rect 74368 42022 74396 42162
rect 74356 42016 74408 42022
rect 74356 41958 74408 41964
rect 74368 41818 74396 41958
rect 74356 41812 74408 41818
rect 74356 41754 74408 41760
rect 74172 41744 74224 41750
rect 74172 41686 74224 41692
rect 74184 40050 74212 41686
rect 74172 40044 74224 40050
rect 74172 39986 74224 39992
rect 73988 39976 74040 39982
rect 73988 39918 74040 39924
rect 73896 39840 73948 39846
rect 73896 39782 73948 39788
rect 73908 39438 73936 39782
rect 73896 39432 73948 39438
rect 73896 39374 73948 39380
rect 73160 39364 73212 39370
rect 73160 39306 73212 39312
rect 73068 38888 73120 38894
rect 73068 38830 73120 38836
rect 72608 38344 72660 38350
rect 72608 38286 72660 38292
rect 72792 38344 72844 38350
rect 72792 38286 72844 38292
rect 72700 38208 72752 38214
rect 72700 38150 72752 38156
rect 72712 37874 72740 38150
rect 72700 37868 72752 37874
rect 72700 37810 72752 37816
rect 70492 37800 70544 37806
rect 68928 37742 68980 37748
rect 70122 37768 70178 37777
rect 69296 37732 69348 37738
rect 69296 37674 69348 37680
rect 69572 37732 69624 37738
rect 70492 37742 70544 37748
rect 70768 37800 70820 37806
rect 70768 37742 70820 37748
rect 71044 37800 71096 37806
rect 71044 37742 71096 37748
rect 71228 37800 71280 37806
rect 71228 37742 71280 37748
rect 71320 37800 71372 37806
rect 71320 37742 71372 37748
rect 72240 37800 72292 37806
rect 72240 37742 72292 37748
rect 72424 37800 72476 37806
rect 72424 37742 72476 37748
rect 70122 37703 70178 37712
rect 69572 37674 69624 37680
rect 68928 37664 68980 37670
rect 69112 37664 69164 37670
rect 68980 37612 69060 37618
rect 68928 37606 69060 37612
rect 69112 37606 69164 37612
rect 68940 37590 69060 37606
rect 67456 37188 67508 37194
rect 67456 37130 67508 37136
rect 65660 37020 65956 37040
rect 65716 37018 65740 37020
rect 65796 37018 65820 37020
rect 65876 37018 65900 37020
rect 65738 36966 65740 37018
rect 65802 36966 65814 37018
rect 65876 36966 65878 37018
rect 65716 36964 65740 36966
rect 65796 36964 65820 36966
rect 65876 36964 65900 36966
rect 65660 36944 65956 36964
rect 69032 36786 69060 37590
rect 69124 37466 69152 37606
rect 69112 37460 69164 37466
rect 69112 37402 69164 37408
rect 69308 37194 69336 37674
rect 69584 37466 69612 37674
rect 69572 37460 69624 37466
rect 69572 37402 69624 37408
rect 69756 37256 69808 37262
rect 69756 37198 69808 37204
rect 69296 37188 69348 37194
rect 69296 37130 69348 37136
rect 69020 36780 69072 36786
rect 69020 36722 69072 36728
rect 69308 36718 69336 37130
rect 69296 36712 69348 36718
rect 69296 36654 69348 36660
rect 69768 36650 69796 37198
rect 70504 37126 70532 37742
rect 70780 37466 70808 37742
rect 71240 37670 71268 37742
rect 71228 37664 71280 37670
rect 71228 37606 71280 37612
rect 71240 37466 71268 37606
rect 70768 37460 70820 37466
rect 70768 37402 70820 37408
rect 71228 37460 71280 37466
rect 71228 37402 71280 37408
rect 70492 37120 70544 37126
rect 70492 37062 70544 37068
rect 69756 36644 69808 36650
rect 69756 36586 69808 36592
rect 66076 36576 66128 36582
rect 66076 36518 66128 36524
rect 66088 36242 66116 36518
rect 66076 36236 66128 36242
rect 66076 36178 66128 36184
rect 70504 36174 70532 37062
rect 71044 36780 71096 36786
rect 71044 36722 71096 36728
rect 70492 36168 70544 36174
rect 67454 36136 67510 36145
rect 70492 36110 70544 36116
rect 67454 36071 67510 36080
rect 65660 35932 65956 35952
rect 65716 35930 65740 35932
rect 65796 35930 65820 35932
rect 65876 35930 65900 35932
rect 65738 35878 65740 35930
rect 65802 35878 65814 35930
rect 65876 35878 65878 35930
rect 65716 35876 65740 35878
rect 65796 35876 65820 35878
rect 65876 35876 65900 35878
rect 65660 35856 65956 35876
rect 67468 35850 67496 36071
rect 70216 36032 70268 36038
rect 70216 35974 70268 35980
rect 67638 35864 67694 35873
rect 67468 35822 67638 35850
rect 67638 35799 67694 35808
rect 68744 35760 68796 35766
rect 68744 35702 68796 35708
rect 66260 35692 66312 35698
rect 66260 35634 66312 35640
rect 65984 35556 66036 35562
rect 65984 35498 66036 35504
rect 65660 34844 65956 34864
rect 65716 34842 65740 34844
rect 65796 34842 65820 34844
rect 65876 34842 65900 34844
rect 65738 34790 65740 34842
rect 65802 34790 65814 34842
rect 65876 34790 65878 34842
rect 65716 34788 65740 34790
rect 65796 34788 65820 34790
rect 65876 34788 65900 34790
rect 65660 34768 65956 34788
rect 65340 34672 65392 34678
rect 65340 34614 65392 34620
rect 65996 34406 66024 35498
rect 66076 35488 66128 35494
rect 66076 35430 66128 35436
rect 66168 35488 66220 35494
rect 66168 35430 66220 35436
rect 66088 35034 66116 35430
rect 66180 35329 66208 35430
rect 66166 35320 66222 35329
rect 66166 35255 66222 35264
rect 66272 35034 66300 35634
rect 68560 35624 68612 35630
rect 68560 35566 68612 35572
rect 66994 35456 67050 35465
rect 66994 35391 67050 35400
rect 66720 35148 66772 35154
rect 66720 35090 66772 35096
rect 66088 35006 66300 35034
rect 66352 35080 66404 35086
rect 66352 35022 66404 35028
rect 66180 34950 66208 35006
rect 66168 34944 66220 34950
rect 66168 34886 66220 34892
rect 64512 34400 64564 34406
rect 64512 34342 64564 34348
rect 65984 34400 66036 34406
rect 65984 34342 66036 34348
rect 66180 32570 66208 34886
rect 66364 34762 66392 35022
rect 66732 34950 66760 35090
rect 66720 34944 66772 34950
rect 66720 34886 66772 34892
rect 66272 34734 66392 34762
rect 66272 34610 66300 34734
rect 67008 34678 67036 35391
rect 67272 35216 67324 35222
rect 67272 35158 67324 35164
rect 67088 35148 67140 35154
rect 67088 35090 67140 35096
rect 67100 34950 67128 35090
rect 67284 35018 67312 35158
rect 68572 35086 68600 35566
rect 68652 35556 68704 35562
rect 68652 35498 68704 35504
rect 68664 35465 68692 35498
rect 68650 35456 68706 35465
rect 68650 35391 68706 35400
rect 68756 35154 68784 35702
rect 70228 35698 70256 35974
rect 71056 35834 71084 36722
rect 71332 36242 71360 37742
rect 72252 37466 72280 37742
rect 72804 37466 72832 38286
rect 73172 37466 73200 39306
rect 74000 38758 74028 39918
rect 74368 39914 74396 41754
rect 74724 41064 74776 41070
rect 74724 41006 74776 41012
rect 74814 41032 74870 41041
rect 74736 40594 74764 41006
rect 74814 40967 74870 40976
rect 74908 40996 74960 41002
rect 74828 40934 74856 40967
rect 74908 40938 74960 40944
rect 74816 40928 74868 40934
rect 74816 40870 74868 40876
rect 74920 40594 74948 40938
rect 74724 40588 74776 40594
rect 74724 40530 74776 40536
rect 74908 40588 74960 40594
rect 74908 40530 74960 40536
rect 75826 40488 75882 40497
rect 75826 40423 75828 40432
rect 75880 40423 75882 40432
rect 75828 40394 75880 40400
rect 74448 39976 74500 39982
rect 74448 39918 74500 39924
rect 74356 39908 74408 39914
rect 74356 39850 74408 39856
rect 74460 38962 74488 39918
rect 74908 39908 74960 39914
rect 74908 39850 74960 39856
rect 74920 39506 74948 39850
rect 74908 39500 74960 39506
rect 74908 39442 74960 39448
rect 74908 39296 74960 39302
rect 74908 39238 74960 39244
rect 74722 38992 74778 39001
rect 74448 38956 74500 38962
rect 74722 38927 74724 38936
rect 74448 38898 74500 38904
rect 74776 38927 74778 38936
rect 74724 38898 74776 38904
rect 74920 38894 74948 39238
rect 74908 38888 74960 38894
rect 74908 38830 74960 38836
rect 73988 38752 74040 38758
rect 73988 38694 74040 38700
rect 74000 38418 74028 38694
rect 73988 38412 74040 38418
rect 73988 38354 74040 38360
rect 74172 38208 74224 38214
rect 74172 38150 74224 38156
rect 72240 37460 72292 37466
rect 72240 37402 72292 37408
rect 72792 37460 72844 37466
rect 72792 37402 72844 37408
rect 73160 37460 73212 37466
rect 73160 37402 73212 37408
rect 71780 37392 71832 37398
rect 71780 37334 71832 37340
rect 71504 37324 71556 37330
rect 71504 37266 71556 37272
rect 71412 36712 71464 36718
rect 71412 36654 71464 36660
rect 71320 36236 71372 36242
rect 71320 36178 71372 36184
rect 70492 35828 70544 35834
rect 70492 35770 70544 35776
rect 71044 35828 71096 35834
rect 71044 35770 71096 35776
rect 70216 35692 70268 35698
rect 70216 35634 70268 35640
rect 69112 35624 69164 35630
rect 68848 35584 69112 35612
rect 68744 35148 68796 35154
rect 68744 35090 68796 35096
rect 68560 35080 68612 35086
rect 68560 35022 68612 35028
rect 67272 35012 67324 35018
rect 67272 34954 67324 34960
rect 68744 35012 68796 35018
rect 68848 35000 68876 35584
rect 69112 35566 69164 35572
rect 69938 35592 69994 35601
rect 69938 35527 69994 35536
rect 69848 35488 69900 35494
rect 69848 35430 69900 35436
rect 69204 35284 69256 35290
rect 69204 35226 69256 35232
rect 68928 35216 68980 35222
rect 69216 35170 69244 35226
rect 68980 35164 69244 35170
rect 68928 35158 69244 35164
rect 68940 35142 69244 35158
rect 68796 34972 68876 35000
rect 68744 34954 68796 34960
rect 69860 34950 69888 35430
rect 69952 34950 69980 35527
rect 70504 35494 70532 35770
rect 71424 35630 71452 36654
rect 71516 36378 71544 37266
rect 71792 36854 71820 37334
rect 72976 37324 73028 37330
rect 72976 37266 73028 37272
rect 72332 37256 72384 37262
rect 72332 37198 72384 37204
rect 71780 36848 71832 36854
rect 71780 36790 71832 36796
rect 71504 36372 71556 36378
rect 71504 36314 71556 36320
rect 71516 36038 71544 36314
rect 72344 36242 72372 37198
rect 72988 37126 73016 37266
rect 72976 37120 73028 37126
rect 72976 37062 73028 37068
rect 72988 36854 73016 37062
rect 72976 36848 73028 36854
rect 72976 36790 73028 36796
rect 71780 36236 71832 36242
rect 71780 36178 71832 36184
rect 72332 36236 72384 36242
rect 72332 36178 72384 36184
rect 73068 36236 73120 36242
rect 73068 36178 73120 36184
rect 71504 36032 71556 36038
rect 71504 35974 71556 35980
rect 71412 35624 71464 35630
rect 71412 35566 71464 35572
rect 70492 35488 70544 35494
rect 70492 35430 70544 35436
rect 70584 35488 70636 35494
rect 70584 35430 70636 35436
rect 70596 35086 70624 35430
rect 71792 35222 71820 36178
rect 73080 35873 73108 36178
rect 73172 36174 73200 37402
rect 73160 36168 73212 36174
rect 73160 36110 73212 36116
rect 73252 36032 73304 36038
rect 73252 35974 73304 35980
rect 73066 35864 73122 35873
rect 73066 35799 73068 35808
rect 73120 35799 73122 35808
rect 73068 35770 73120 35776
rect 73080 35739 73108 35770
rect 71780 35216 71832 35222
rect 71780 35158 71832 35164
rect 73264 35154 73292 35974
rect 74184 35154 74212 38150
rect 75932 37330 75960 42162
rect 77680 42158 77708 42570
rect 78312 42560 78364 42566
rect 78312 42502 78364 42508
rect 77668 42152 77720 42158
rect 77668 42094 77720 42100
rect 76748 42016 76800 42022
rect 76748 41958 76800 41964
rect 76760 41274 76788 41958
rect 76748 41268 76800 41274
rect 76748 41210 76800 41216
rect 76760 37874 76788 41210
rect 77208 40180 77260 40186
rect 77208 40122 77260 40128
rect 77220 40089 77248 40122
rect 77206 40080 77262 40089
rect 77206 40015 77262 40024
rect 77484 39976 77536 39982
rect 77484 39918 77536 39924
rect 77392 39840 77444 39846
rect 77392 39782 77444 39788
rect 77300 39500 77352 39506
rect 77300 39442 77352 39448
rect 77312 38758 77340 39442
rect 77404 38758 77432 39782
rect 77496 39642 77524 39918
rect 77576 39840 77628 39846
rect 77576 39782 77628 39788
rect 77484 39636 77536 39642
rect 77484 39578 77536 39584
rect 77300 38752 77352 38758
rect 77300 38694 77352 38700
rect 77392 38752 77444 38758
rect 77392 38694 77444 38700
rect 77404 38418 77432 38694
rect 77588 38554 77616 39782
rect 78324 39506 78352 42502
rect 78600 42294 78628 42842
rect 78784 42702 78812 43114
rect 78772 42696 78824 42702
rect 78772 42638 78824 42644
rect 78588 42288 78640 42294
rect 78588 42230 78640 42236
rect 78404 42152 78456 42158
rect 78404 42094 78456 42100
rect 78416 41070 78444 42094
rect 78680 41676 78732 41682
rect 78680 41618 78732 41624
rect 78692 41274 78720 41618
rect 78876 41546 78904 43182
rect 81020 43004 81316 43024
rect 81076 43002 81100 43004
rect 81156 43002 81180 43004
rect 81236 43002 81260 43004
rect 81098 42950 81100 43002
rect 81162 42950 81174 43002
rect 81236 42950 81238 43002
rect 81076 42948 81100 42950
rect 81156 42948 81180 42950
rect 81236 42948 81260 42950
rect 81020 42928 81316 42948
rect 81452 42906 81480 43794
rect 82084 43648 82136 43654
rect 82084 43590 82136 43596
rect 81992 43240 82044 43246
rect 81992 43182 82044 43188
rect 81532 43172 81584 43178
rect 81532 43114 81584 43120
rect 81440 42900 81492 42906
rect 81440 42842 81492 42848
rect 81544 42786 81572 43114
rect 81452 42770 81572 42786
rect 81440 42764 81572 42770
rect 81492 42758 81572 42764
rect 81440 42706 81492 42712
rect 79876 42560 79928 42566
rect 79876 42502 79928 42508
rect 79888 42158 79916 42502
rect 79876 42152 79928 42158
rect 79876 42094 79928 42100
rect 79968 42016 80020 42022
rect 79968 41958 80020 41964
rect 78864 41540 78916 41546
rect 78864 41482 78916 41488
rect 79980 41274 80008 41958
rect 81020 41916 81316 41936
rect 81076 41914 81100 41916
rect 81156 41914 81180 41916
rect 81236 41914 81260 41916
rect 81098 41862 81100 41914
rect 81162 41862 81174 41914
rect 81236 41862 81238 41914
rect 81076 41860 81100 41862
rect 81156 41860 81180 41862
rect 81236 41860 81260 41862
rect 81020 41840 81316 41860
rect 81176 41682 81388 41698
rect 81164 41676 81388 41682
rect 81216 41670 81388 41676
rect 81164 41618 81216 41624
rect 80888 41608 80940 41614
rect 80888 41550 80940 41556
rect 80900 41274 80928 41550
rect 78680 41268 78732 41274
rect 78680 41210 78732 41216
rect 79968 41268 80020 41274
rect 79968 41210 80020 41216
rect 80888 41268 80940 41274
rect 80888 41210 80940 41216
rect 78404 41064 78456 41070
rect 78404 41006 78456 41012
rect 78692 40458 78720 41210
rect 80796 41064 80848 41070
rect 80796 41006 80848 41012
rect 80808 40934 80836 41006
rect 79416 40928 79468 40934
rect 79416 40870 79468 40876
rect 80796 40928 80848 40934
rect 80796 40870 80848 40876
rect 78680 40452 78732 40458
rect 78680 40394 78732 40400
rect 79428 40050 79456 40870
rect 80808 40390 80836 40870
rect 81020 40828 81316 40848
rect 81076 40826 81100 40828
rect 81156 40826 81180 40828
rect 81236 40826 81260 40828
rect 81098 40774 81100 40826
rect 81162 40774 81174 40826
rect 81236 40774 81238 40826
rect 81076 40772 81100 40774
rect 81156 40772 81180 40774
rect 81236 40772 81260 40774
rect 81020 40752 81316 40772
rect 81360 40662 81388 41670
rect 81452 41206 81480 42706
rect 82004 42702 82032 43182
rect 81992 42696 82044 42702
rect 81992 42638 82044 42644
rect 82004 41750 82032 42638
rect 82096 42362 82124 43590
rect 82372 43314 82400 43794
rect 82820 43784 82872 43790
rect 82820 43726 82872 43732
rect 82360 43308 82412 43314
rect 82360 43250 82412 43256
rect 82832 42770 82860 43726
rect 96380 43548 96676 43568
rect 96436 43546 96460 43548
rect 96516 43546 96540 43548
rect 96596 43546 96620 43548
rect 96458 43494 96460 43546
rect 96522 43494 96534 43546
rect 96596 43494 96598 43546
rect 96436 43492 96460 43494
rect 96516 43492 96540 43494
rect 96596 43492 96620 43494
rect 96380 43472 96676 43492
rect 83832 43104 83884 43110
rect 83832 43046 83884 43052
rect 82820 42764 82872 42770
rect 82820 42706 82872 42712
rect 82728 42696 82780 42702
rect 82728 42638 82780 42644
rect 82084 42356 82136 42362
rect 82084 42298 82136 42304
rect 82360 42356 82412 42362
rect 82360 42298 82412 42304
rect 81992 41744 82044 41750
rect 81992 41686 82044 41692
rect 82372 41682 82400 42298
rect 82740 42158 82768 42638
rect 83844 42566 83872 43046
rect 85212 42900 85264 42906
rect 85212 42842 85264 42848
rect 83004 42560 83056 42566
rect 83004 42502 83056 42508
rect 83832 42560 83884 42566
rect 83832 42502 83884 42508
rect 82728 42152 82780 42158
rect 82728 42094 82780 42100
rect 82360 41676 82412 41682
rect 82360 41618 82412 41624
rect 82912 41676 82964 41682
rect 82912 41618 82964 41624
rect 81440 41200 81492 41206
rect 81440 41142 81492 41148
rect 81348 40656 81400 40662
rect 81348 40598 81400 40604
rect 80888 40588 80940 40594
rect 80888 40530 80940 40536
rect 80900 40390 80928 40530
rect 80796 40384 80848 40390
rect 80796 40326 80848 40332
rect 80888 40384 80940 40390
rect 80888 40326 80940 40332
rect 79876 40180 79928 40186
rect 79876 40122 79928 40128
rect 79888 40066 79916 40122
rect 80152 40112 80204 40118
rect 79888 40060 80152 40066
rect 79888 40054 80204 40060
rect 79416 40044 79468 40050
rect 79416 39986 79468 39992
rect 79508 40044 79560 40050
rect 79888 40038 80192 40054
rect 79508 39986 79560 39992
rect 78312 39500 78364 39506
rect 78312 39442 78364 39448
rect 79520 38894 79548 39986
rect 80808 39982 80836 40326
rect 80900 39982 80928 40326
rect 80336 39976 80388 39982
rect 80520 39976 80572 39982
rect 80388 39924 80520 39930
rect 80336 39918 80572 39924
rect 80796 39976 80848 39982
rect 80796 39918 80848 39924
rect 80888 39976 80940 39982
rect 80888 39918 80940 39924
rect 79876 39908 79928 39914
rect 80348 39902 80560 39918
rect 79876 39850 79928 39856
rect 79888 39506 79916 39850
rect 79876 39500 79928 39506
rect 79876 39442 79928 39448
rect 80532 39370 80560 39902
rect 80808 39846 80836 39918
rect 80900 39846 80928 39918
rect 80796 39840 80848 39846
rect 80796 39782 80848 39788
rect 80888 39840 80940 39846
rect 80888 39782 80940 39788
rect 80520 39364 80572 39370
rect 80520 39306 80572 39312
rect 80900 39030 80928 39782
rect 81020 39740 81316 39760
rect 81076 39738 81100 39740
rect 81156 39738 81180 39740
rect 81236 39738 81260 39740
rect 81098 39686 81100 39738
rect 81162 39686 81174 39738
rect 81236 39686 81238 39738
rect 81076 39684 81100 39686
rect 81156 39684 81180 39686
rect 81236 39684 81260 39686
rect 81020 39664 81316 39684
rect 81360 39506 81388 40598
rect 81440 40588 81492 40594
rect 81440 40530 81492 40536
rect 81452 39914 81480 40530
rect 82372 40050 82400 41618
rect 82728 40928 82780 40934
rect 82728 40870 82780 40876
rect 82740 40730 82768 40870
rect 82924 40730 82952 41618
rect 82728 40724 82780 40730
rect 82728 40666 82780 40672
rect 82912 40724 82964 40730
rect 82912 40666 82964 40672
rect 83016 40526 83044 42502
rect 83096 42152 83148 42158
rect 83096 42094 83148 42100
rect 83108 41478 83136 42094
rect 84108 42016 84160 42022
rect 84108 41958 84160 41964
rect 84120 41682 84148 41958
rect 83648 41676 83700 41682
rect 83648 41618 83700 41624
rect 84108 41676 84160 41682
rect 84108 41618 84160 41624
rect 83096 41472 83148 41478
rect 83096 41414 83148 41420
rect 83660 41070 83688 41618
rect 83648 41064 83700 41070
rect 83648 41006 83700 41012
rect 83004 40520 83056 40526
rect 83004 40462 83056 40468
rect 85224 40050 85252 42842
rect 96380 42460 96676 42480
rect 96436 42458 96460 42460
rect 96516 42458 96540 42460
rect 96596 42458 96620 42460
rect 96458 42406 96460 42458
rect 96522 42406 96534 42458
rect 96596 42406 96598 42458
rect 96436 42404 96460 42406
rect 96516 42404 96540 42406
rect 96596 42404 96620 42406
rect 96380 42384 96676 42404
rect 85764 42220 85816 42226
rect 85764 42162 85816 42168
rect 85776 40050 85804 42162
rect 87144 42084 87196 42090
rect 87144 42026 87196 42032
rect 87156 41274 87184 42026
rect 96380 41372 96676 41392
rect 96436 41370 96460 41372
rect 96516 41370 96540 41372
rect 96596 41370 96620 41372
rect 96458 41318 96460 41370
rect 96522 41318 96534 41370
rect 96596 41318 96598 41370
rect 96436 41316 96460 41318
rect 96516 41316 96540 41318
rect 96596 41316 96620 41318
rect 96380 41296 96676 41316
rect 87144 41268 87196 41274
rect 87144 41210 87196 41216
rect 88984 41132 89036 41138
rect 88984 41074 89036 41080
rect 87604 41064 87656 41070
rect 87604 41006 87656 41012
rect 87616 40662 87644 41006
rect 88524 40928 88576 40934
rect 88524 40870 88576 40876
rect 87604 40656 87656 40662
rect 87604 40598 87656 40604
rect 86500 40588 86552 40594
rect 86500 40530 86552 40536
rect 86224 40520 86276 40526
rect 86224 40462 86276 40468
rect 86236 40118 86264 40462
rect 86224 40112 86276 40118
rect 86224 40054 86276 40060
rect 82360 40044 82412 40050
rect 82360 39986 82412 39992
rect 84936 40044 84988 40050
rect 84936 39986 84988 39992
rect 85212 40044 85264 40050
rect 85212 39986 85264 39992
rect 85764 40044 85816 40050
rect 85764 39986 85816 39992
rect 82728 39976 82780 39982
rect 82728 39918 82780 39924
rect 84108 39976 84160 39982
rect 84108 39918 84160 39924
rect 81440 39908 81492 39914
rect 81440 39850 81492 39856
rect 81452 39642 81480 39850
rect 81440 39636 81492 39642
rect 81440 39578 81492 39584
rect 81348 39500 81400 39506
rect 81348 39442 81400 39448
rect 82360 39432 82412 39438
rect 82360 39374 82412 39380
rect 80888 39024 80940 39030
rect 80888 38966 80940 38972
rect 82372 38962 82400 39374
rect 82740 38962 82768 39918
rect 83004 39636 83056 39642
rect 83004 39578 83056 39584
rect 82360 38956 82412 38962
rect 82360 38898 82412 38904
rect 82728 38956 82780 38962
rect 82728 38898 82780 38904
rect 79508 38888 79560 38894
rect 79508 38830 79560 38836
rect 82820 38820 82872 38826
rect 82820 38762 82872 38768
rect 81532 38752 81584 38758
rect 81532 38694 81584 38700
rect 81020 38652 81316 38672
rect 81076 38650 81100 38652
rect 81156 38650 81180 38652
rect 81236 38650 81260 38652
rect 81098 38598 81100 38650
rect 81162 38598 81174 38650
rect 81236 38598 81238 38650
rect 81076 38596 81100 38598
rect 81156 38596 81180 38598
rect 81236 38596 81260 38598
rect 81020 38576 81316 38596
rect 77576 38548 77628 38554
rect 77576 38490 77628 38496
rect 77392 38412 77444 38418
rect 77392 38354 77444 38360
rect 81440 38412 81492 38418
rect 81440 38354 81492 38360
rect 77484 38208 77536 38214
rect 77484 38150 77536 38156
rect 77496 37942 77524 38150
rect 77484 37936 77536 37942
rect 77484 37878 77536 37884
rect 76748 37868 76800 37874
rect 76748 37810 76800 37816
rect 77484 37800 77536 37806
rect 77484 37742 77536 37748
rect 77668 37800 77720 37806
rect 77668 37742 77720 37748
rect 77300 37664 77352 37670
rect 77300 37606 77352 37612
rect 75920 37324 75972 37330
rect 75920 37266 75972 37272
rect 75932 36174 75960 37266
rect 76748 37120 76800 37126
rect 76748 37062 76800 37068
rect 75920 36168 75972 36174
rect 75920 36110 75972 36116
rect 75932 35630 75960 36110
rect 74264 35624 74316 35630
rect 74264 35566 74316 35572
rect 75920 35624 75972 35630
rect 75920 35566 75972 35572
rect 76288 35624 76340 35630
rect 76288 35566 76340 35572
rect 76656 35624 76708 35630
rect 76656 35566 76708 35572
rect 73252 35148 73304 35154
rect 73252 35090 73304 35096
rect 74172 35148 74224 35154
rect 74172 35090 74224 35096
rect 74276 35086 74304 35566
rect 76300 35222 76328 35566
rect 76564 35556 76616 35562
rect 76564 35498 76616 35504
rect 76288 35216 76340 35222
rect 75366 35184 75422 35193
rect 74632 35148 74684 35154
rect 76288 35158 76340 35164
rect 75366 35119 75368 35128
rect 74632 35090 74684 35096
rect 75420 35119 75422 35128
rect 75644 35148 75696 35154
rect 75368 35090 75420 35096
rect 75644 35090 75696 35096
rect 70584 35080 70636 35086
rect 74264 35080 74316 35086
rect 70584 35022 70636 35028
rect 74262 35048 74264 35057
rect 74316 35048 74318 35057
rect 74262 34983 74318 34992
rect 67088 34944 67140 34950
rect 67088 34886 67140 34892
rect 69848 34944 69900 34950
rect 69848 34886 69900 34892
rect 69940 34944 69992 34950
rect 69940 34886 69992 34892
rect 66996 34672 67048 34678
rect 66996 34614 67048 34620
rect 66260 34604 66312 34610
rect 66260 34546 66312 34552
rect 66352 34604 66404 34610
rect 66352 34546 66404 34552
rect 66364 34513 66392 34546
rect 66350 34504 66406 34513
rect 74644 34474 74672 35090
rect 75092 34944 75144 34950
rect 75092 34886 75144 34892
rect 75104 34610 75132 34886
rect 75656 34678 75684 35090
rect 76194 34912 76250 34921
rect 76194 34847 76250 34856
rect 75644 34672 75696 34678
rect 75644 34614 75696 34620
rect 75092 34604 75144 34610
rect 75092 34546 75144 34552
rect 76208 34542 76236 34847
rect 76576 34626 76604 35498
rect 76668 35465 76696 35566
rect 76654 35456 76710 35465
rect 76654 35391 76710 35400
rect 76760 34921 76788 37062
rect 77312 36786 77340 37606
rect 77392 37256 77444 37262
rect 77392 37198 77444 37204
rect 77300 36780 77352 36786
rect 77300 36722 77352 36728
rect 77404 36718 77432 37198
rect 77496 36786 77524 37742
rect 77484 36780 77536 36786
rect 77484 36722 77536 36728
rect 77392 36712 77444 36718
rect 77392 36654 77444 36660
rect 77300 36576 77352 36582
rect 77300 36518 77352 36524
rect 77312 35306 77340 36518
rect 77390 35864 77446 35873
rect 77390 35799 77446 35808
rect 77404 35630 77432 35799
rect 77496 35698 77524 36722
rect 77680 36718 77708 37742
rect 81452 37738 81480 38354
rect 81544 38214 81572 38694
rect 82832 38418 82860 38762
rect 82820 38412 82872 38418
rect 82820 38354 82872 38360
rect 82912 38412 82964 38418
rect 82912 38354 82964 38360
rect 81532 38208 81584 38214
rect 81532 38150 81584 38156
rect 81716 38208 81768 38214
rect 81716 38150 81768 38156
rect 81440 37732 81492 37738
rect 81440 37674 81492 37680
rect 81020 37564 81316 37584
rect 81076 37562 81100 37564
rect 81156 37562 81180 37564
rect 81236 37562 81260 37564
rect 81098 37510 81100 37562
rect 81162 37510 81174 37562
rect 81236 37510 81238 37562
rect 81076 37508 81100 37510
rect 81156 37508 81180 37510
rect 81236 37508 81260 37510
rect 81020 37488 81316 37508
rect 78404 37120 78456 37126
rect 78404 37062 78456 37068
rect 78416 36718 78444 37062
rect 79232 36780 79284 36786
rect 79232 36722 79284 36728
rect 77668 36712 77720 36718
rect 77668 36654 77720 36660
rect 78404 36712 78456 36718
rect 78404 36654 78456 36660
rect 78772 36712 78824 36718
rect 78772 36654 78824 36660
rect 77680 36310 77708 36654
rect 77668 36304 77720 36310
rect 77668 36246 77720 36252
rect 77850 36272 77906 36281
rect 77576 36236 77628 36242
rect 78784 36242 78812 36654
rect 79244 36281 79272 36722
rect 79784 36644 79836 36650
rect 79784 36586 79836 36592
rect 79230 36272 79286 36281
rect 77850 36207 77906 36216
rect 78772 36236 78824 36242
rect 77576 36178 77628 36184
rect 77588 36145 77616 36178
rect 77864 36174 77892 36207
rect 79230 36207 79232 36216
rect 78772 36178 78824 36184
rect 79284 36207 79286 36216
rect 79232 36178 79284 36184
rect 77852 36168 77904 36174
rect 77574 36136 77630 36145
rect 77852 36110 77904 36116
rect 78036 36168 78088 36174
rect 78312 36168 78364 36174
rect 78088 36128 78312 36156
rect 78036 36110 78088 36116
rect 78312 36110 78364 36116
rect 77574 36071 77630 36080
rect 77588 35766 77616 36071
rect 77944 36032 77996 36038
rect 77944 35974 77996 35980
rect 77956 35834 77984 35974
rect 77668 35828 77720 35834
rect 77668 35770 77720 35776
rect 77944 35828 77996 35834
rect 77944 35770 77996 35776
rect 77576 35760 77628 35766
rect 77576 35702 77628 35708
rect 77484 35692 77536 35698
rect 77484 35634 77536 35640
rect 77392 35624 77444 35630
rect 77392 35566 77444 35572
rect 77680 35578 77708 35770
rect 77944 35624 77996 35630
rect 77864 35584 77944 35612
rect 77864 35578 77892 35584
rect 77680 35562 77892 35578
rect 77944 35566 77996 35572
rect 78310 35592 78366 35601
rect 77668 35556 77892 35562
rect 77720 35550 77892 35556
rect 78784 35562 78812 36178
rect 79244 36147 79272 36178
rect 79796 36145 79824 36586
rect 81728 36582 81756 38150
rect 82544 37800 82596 37806
rect 82544 37742 82596 37748
rect 80060 36576 80112 36582
rect 80060 36518 80112 36524
rect 81716 36576 81768 36582
rect 81716 36518 81768 36524
rect 80072 36310 80100 36518
rect 81020 36476 81316 36496
rect 81076 36474 81100 36476
rect 81156 36474 81180 36476
rect 81236 36474 81260 36476
rect 81098 36422 81100 36474
rect 81162 36422 81174 36474
rect 81236 36422 81238 36474
rect 81076 36420 81100 36422
rect 81156 36420 81180 36422
rect 81236 36420 81260 36422
rect 81020 36400 81316 36420
rect 81728 36310 81756 36518
rect 80060 36304 80112 36310
rect 80060 36246 80112 36252
rect 81716 36304 81768 36310
rect 81716 36246 81768 36252
rect 79782 36136 79838 36145
rect 79782 36071 79838 36080
rect 79600 36032 79652 36038
rect 79600 35974 79652 35980
rect 78772 35556 78824 35562
rect 78310 35527 78366 35536
rect 77668 35498 77720 35504
rect 77036 35278 77340 35306
rect 77036 35018 77064 35278
rect 78324 35222 78352 35527
rect 78692 35516 78772 35544
rect 78312 35216 78364 35222
rect 78312 35158 78364 35164
rect 77116 35148 77168 35154
rect 77116 35090 77168 35096
rect 77024 35012 77076 35018
rect 77024 34954 77076 34960
rect 76746 34912 76802 34921
rect 76746 34847 76802 34856
rect 76484 34610 76604 34626
rect 76472 34604 76604 34610
rect 76524 34598 76604 34604
rect 76472 34546 76524 34552
rect 77128 34542 77156 35090
rect 77298 35048 77354 35057
rect 77298 34983 77354 34992
rect 77312 34950 77340 34983
rect 77300 34944 77352 34950
rect 78036 34944 78088 34950
rect 77300 34886 77352 34892
rect 78034 34912 78036 34921
rect 78088 34912 78090 34921
rect 78034 34847 78090 34856
rect 78494 34776 78550 34785
rect 78494 34711 78550 34720
rect 77760 34672 77812 34678
rect 77760 34614 77812 34620
rect 77772 34542 77800 34614
rect 78508 34610 78536 34711
rect 78586 34640 78642 34649
rect 78496 34604 78548 34610
rect 78586 34575 78642 34584
rect 78496 34546 78548 34552
rect 78600 34542 78628 34575
rect 76196 34536 76248 34542
rect 76196 34478 76248 34484
rect 77116 34536 77168 34542
rect 77116 34478 77168 34484
rect 77760 34536 77812 34542
rect 78588 34536 78640 34542
rect 77760 34478 77812 34484
rect 78494 34504 78550 34513
rect 66350 34439 66406 34448
rect 74632 34468 74684 34474
rect 78588 34478 78640 34484
rect 78494 34439 78496 34448
rect 74632 34410 74684 34416
rect 78548 34439 78550 34448
rect 78692 34456 78720 35516
rect 78772 35498 78824 35504
rect 79508 35488 79560 35494
rect 79508 35430 79560 35436
rect 79520 35193 79548 35430
rect 79506 35184 79562 35193
rect 79612 35154 79640 35974
rect 79796 35834 79824 36071
rect 82556 36038 82584 37742
rect 82832 37466 82860 38354
rect 82924 38010 82952 38354
rect 82912 38004 82964 38010
rect 82912 37946 82964 37952
rect 82820 37460 82872 37466
rect 82820 37402 82872 37408
rect 83016 37398 83044 39578
rect 83832 39500 83884 39506
rect 83832 39442 83884 39448
rect 83280 39364 83332 39370
rect 83280 39306 83332 39312
rect 83188 39024 83240 39030
rect 83186 38992 83188 39001
rect 83240 38992 83242 39001
rect 83186 38927 83242 38936
rect 83200 38282 83228 38927
rect 83188 38276 83240 38282
rect 83188 38218 83240 38224
rect 83096 38208 83148 38214
rect 83096 38150 83148 38156
rect 83108 37874 83136 38150
rect 83096 37868 83148 37874
rect 83096 37810 83148 37816
rect 83004 37392 83056 37398
rect 83004 37334 83056 37340
rect 83200 37330 83228 38218
rect 83188 37324 83240 37330
rect 83188 37266 83240 37272
rect 82544 36032 82596 36038
rect 82544 35974 82596 35980
rect 79784 35828 79836 35834
rect 79784 35770 79836 35776
rect 80150 35592 80206 35601
rect 79784 35556 79836 35562
rect 80150 35527 80206 35536
rect 79784 35498 79836 35504
rect 79506 35119 79562 35128
rect 79600 35148 79652 35154
rect 79600 35090 79652 35096
rect 78956 34944 79008 34950
rect 78956 34886 79008 34892
rect 78772 34672 78824 34678
rect 78824 34632 78904 34660
rect 78968 34649 78996 34886
rect 79796 34678 79824 35498
rect 80164 35494 80192 35527
rect 80152 35488 80204 35494
rect 80152 35430 80204 35436
rect 81020 35388 81316 35408
rect 81076 35386 81100 35388
rect 81156 35386 81180 35388
rect 81236 35386 81260 35388
rect 81098 35334 81100 35386
rect 81162 35334 81174 35386
rect 81236 35334 81238 35386
rect 81076 35332 81100 35334
rect 81156 35332 81180 35334
rect 81236 35332 81260 35334
rect 81020 35312 81316 35332
rect 81348 35148 81400 35154
rect 81348 35090 81400 35096
rect 81360 34746 81388 35090
rect 82268 35080 82320 35086
rect 82268 35022 82320 35028
rect 81808 34944 81860 34950
rect 81808 34886 81860 34892
rect 82084 34944 82136 34950
rect 82084 34886 82136 34892
rect 81438 34776 81494 34785
rect 81348 34740 81400 34746
rect 81438 34711 81440 34720
rect 81348 34682 81400 34688
rect 81492 34711 81494 34720
rect 81440 34682 81492 34688
rect 79784 34672 79836 34678
rect 78772 34614 78824 34620
rect 78876 34542 78904 34632
rect 78954 34640 79010 34649
rect 79784 34614 79836 34620
rect 81532 34672 81584 34678
rect 81532 34614 81584 34620
rect 78954 34575 78956 34584
rect 79008 34575 79010 34584
rect 81348 34604 81400 34610
rect 78956 34546 79008 34552
rect 81348 34546 81400 34552
rect 78864 34536 78916 34542
rect 80888 34536 80940 34542
rect 78864 34478 78916 34484
rect 79966 34504 80022 34513
rect 78772 34468 78824 34474
rect 78692 34428 78772 34456
rect 78496 34410 78548 34416
rect 80888 34478 80940 34484
rect 79966 34439 80022 34448
rect 78772 34410 78824 34416
rect 67364 34400 67416 34406
rect 67364 34342 67416 34348
rect 67376 34134 67404 34342
rect 67364 34128 67416 34134
rect 67364 34070 67416 34076
rect 66168 32564 66220 32570
rect 66168 32506 66220 32512
rect 63684 32224 63736 32230
rect 63684 32166 63736 32172
rect 62672 31748 62724 31754
rect 62672 31690 62724 31696
rect 56784 31272 56836 31278
rect 56784 31214 56836 31220
rect 54852 30524 54904 30530
rect 54852 30466 54904 30472
rect 54760 24268 54812 24274
rect 54760 24210 54812 24216
rect 53852 24058 54064 24086
rect 53852 20165 53880 24058
rect 53838 20156 53894 20165
rect 53838 20091 53894 20100
rect 54116 19372 54168 19378
rect 54116 19314 54168 19320
rect 54128 18170 54156 19314
rect 53852 18142 54156 18170
rect 53852 14861 53880 18142
rect 53838 14852 53894 14861
rect 53838 14787 53894 14796
rect 79980 4865 80008 34439
rect 80900 20097 80928 34478
rect 81020 34300 81316 34320
rect 81076 34298 81100 34300
rect 81156 34298 81180 34300
rect 81236 34298 81260 34300
rect 81098 34246 81100 34298
rect 81162 34246 81174 34298
rect 81236 34246 81238 34298
rect 81076 34244 81100 34246
rect 81156 34244 81180 34246
rect 81236 34244 81260 34246
rect 81020 34224 81316 34244
rect 81360 24245 81388 34546
rect 81440 34536 81492 34542
rect 81440 34478 81492 34484
rect 81452 31754 81480 34478
rect 81440 31748 81492 31754
rect 81440 31690 81492 31696
rect 81438 31648 81494 31657
rect 81438 31583 81494 31592
rect 81452 29549 81480 31583
rect 81544 30938 81572 34614
rect 81624 34604 81676 34610
rect 81624 34546 81676 34552
rect 81532 30932 81584 30938
rect 81532 30874 81584 30880
rect 81544 30229 81572 30874
rect 81530 30220 81586 30229
rect 81530 30155 81586 30164
rect 81438 29540 81494 29549
rect 81438 29475 81494 29484
rect 81636 28189 81664 34546
rect 81716 31748 81768 31754
rect 81716 31690 81768 31696
rect 81622 28180 81678 28189
rect 81622 28115 81678 28124
rect 81622 26820 81678 26829
rect 81728 26806 81756 31690
rect 81820 31006 81848 34886
rect 81990 34504 82046 34513
rect 81990 34439 81992 34448
rect 82044 34439 82046 34448
rect 81992 34410 82044 34416
rect 81808 31000 81860 31006
rect 81808 30942 81860 30948
rect 81678 26778 81756 26806
rect 81622 26755 81678 26764
rect 81622 25596 81678 25605
rect 81820 25582 81848 30942
rect 81678 25554 81848 25582
rect 81622 25531 81678 25540
rect 81346 24236 81402 24245
rect 81346 24171 81402 24180
rect 81624 22908 81676 22914
rect 81622 22876 81624 22885
rect 81676 22876 81678 22885
rect 81622 22811 81678 22820
rect 82096 21298 82124 34886
rect 82280 22914 82308 35022
rect 82556 35018 82584 35974
rect 83292 35154 83320 39306
rect 83740 39296 83792 39302
rect 83740 39238 83792 39244
rect 83752 39098 83780 39238
rect 83740 39092 83792 39098
rect 83740 39034 83792 39040
rect 83752 38962 83780 39034
rect 83372 38956 83424 38962
rect 83372 38898 83424 38904
rect 83740 38956 83792 38962
rect 83740 38898 83792 38904
rect 83384 38826 83412 38898
rect 83372 38820 83424 38826
rect 83372 38762 83424 38768
rect 83384 38729 83412 38762
rect 83370 38720 83426 38729
rect 83370 38655 83426 38664
rect 83844 37806 83872 39442
rect 84120 39438 84148 39918
rect 84200 39840 84252 39846
rect 84200 39782 84252 39788
rect 84568 39840 84620 39846
rect 84568 39782 84620 39788
rect 84108 39432 84160 39438
rect 84108 39374 84160 39380
rect 84212 39030 84240 39782
rect 84580 39506 84608 39782
rect 84568 39500 84620 39506
rect 84568 39442 84620 39448
rect 84580 39302 84608 39442
rect 84948 39438 84976 39986
rect 84844 39432 84896 39438
rect 84844 39374 84896 39380
rect 84936 39432 84988 39438
rect 84936 39374 84988 39380
rect 84568 39296 84620 39302
rect 84568 39238 84620 39244
rect 84580 39098 84608 39238
rect 84568 39092 84620 39098
rect 84568 39034 84620 39040
rect 84200 39024 84252 39030
rect 84106 38992 84162 39001
rect 84200 38966 84252 38972
rect 84106 38927 84108 38936
rect 84160 38927 84162 38936
rect 84108 38898 84160 38904
rect 84580 38894 84608 39034
rect 84568 38888 84620 38894
rect 84568 38830 84620 38836
rect 84856 38826 84884 39374
rect 84844 38820 84896 38826
rect 84844 38762 84896 38768
rect 84014 38720 84070 38729
rect 84014 38655 84070 38664
rect 84028 38554 84056 38655
rect 84016 38548 84068 38554
rect 84016 38490 84068 38496
rect 83832 37800 83884 37806
rect 83832 37742 83884 37748
rect 84476 37256 84528 37262
rect 84476 37198 84528 37204
rect 84292 37120 84344 37126
rect 84292 37062 84344 37068
rect 84304 36582 84332 37062
rect 84292 36576 84344 36582
rect 84292 36518 84344 36524
rect 83740 36372 83792 36378
rect 83740 36314 83792 36320
rect 83752 35630 83780 36314
rect 83740 35624 83792 35630
rect 83740 35566 83792 35572
rect 84304 35494 84332 36518
rect 84488 36242 84516 37198
rect 85224 36854 85252 39986
rect 85672 39636 85724 39642
rect 85672 39578 85724 39584
rect 85684 39098 85712 39578
rect 85776 39506 85804 39986
rect 86512 39982 86540 40530
rect 86684 40520 86736 40526
rect 86684 40462 86736 40468
rect 85948 39976 86000 39982
rect 85948 39918 86000 39924
rect 86500 39976 86552 39982
rect 86500 39918 86552 39924
rect 85960 39846 85988 39918
rect 86696 39846 86724 40462
rect 88432 40044 88484 40050
rect 88432 39986 88484 39992
rect 86866 39944 86922 39953
rect 86866 39879 86922 39888
rect 86880 39846 86908 39879
rect 85948 39840 86000 39846
rect 85948 39782 86000 39788
rect 86684 39840 86736 39846
rect 86684 39782 86736 39788
rect 86868 39840 86920 39846
rect 86868 39782 86920 39788
rect 85960 39642 85988 39782
rect 85948 39636 86000 39642
rect 85948 39578 86000 39584
rect 86880 39506 86908 39782
rect 85764 39500 85816 39506
rect 85764 39442 85816 39448
rect 86868 39500 86920 39506
rect 86868 39442 86920 39448
rect 86224 39296 86276 39302
rect 86224 39238 86276 39244
rect 85672 39092 85724 39098
rect 85672 39034 85724 39040
rect 86236 38418 86264 39238
rect 86868 38888 86920 38894
rect 86868 38830 86920 38836
rect 86960 38888 87012 38894
rect 86960 38830 87012 38836
rect 85672 38412 85724 38418
rect 85672 38354 85724 38360
rect 86224 38412 86276 38418
rect 86224 38354 86276 38360
rect 85684 37806 85712 38354
rect 85672 37800 85724 37806
rect 85672 37742 85724 37748
rect 85580 37392 85632 37398
rect 85580 37334 85632 37340
rect 85488 37120 85540 37126
rect 85488 37062 85540 37068
rect 85212 36848 85264 36854
rect 85212 36790 85264 36796
rect 85500 36718 85528 37062
rect 85592 36854 85620 37334
rect 86880 37330 86908 38830
rect 86972 38486 87000 38830
rect 88444 38486 88472 39986
rect 88536 39982 88564 40870
rect 88996 40730 89024 41074
rect 88984 40724 89036 40730
rect 88984 40666 89036 40672
rect 88996 40050 89024 40666
rect 89444 40520 89496 40526
rect 89444 40462 89496 40468
rect 88984 40044 89036 40050
rect 88984 39986 89036 39992
rect 88524 39976 88576 39982
rect 88524 39918 88576 39924
rect 89456 39642 89484 40462
rect 89904 40384 89956 40390
rect 89904 40326 89956 40332
rect 89444 39636 89496 39642
rect 89444 39578 89496 39584
rect 89916 39506 89944 40326
rect 96380 40284 96676 40304
rect 96436 40282 96460 40284
rect 96516 40282 96540 40284
rect 96596 40282 96620 40284
rect 96458 40230 96460 40282
rect 96522 40230 96534 40282
rect 96596 40230 96598 40282
rect 96436 40228 96460 40230
rect 96516 40228 96540 40230
rect 96596 40228 96620 40230
rect 96380 40208 96676 40228
rect 91100 39976 91152 39982
rect 91100 39918 91152 39924
rect 91112 39642 91140 39918
rect 91100 39636 91152 39642
rect 91100 39578 91152 39584
rect 89904 39500 89956 39506
rect 89904 39442 89956 39448
rect 91008 39500 91060 39506
rect 91008 39442 91060 39448
rect 88524 39432 88576 39438
rect 88524 39374 88576 39380
rect 88536 39302 88564 39374
rect 90088 39364 90140 39370
rect 90088 39306 90140 39312
rect 88524 39296 88576 39302
rect 88524 39238 88576 39244
rect 86960 38480 87012 38486
rect 86960 38422 87012 38428
rect 88432 38480 88484 38486
rect 88432 38422 88484 38428
rect 88536 38350 88564 39238
rect 89076 38888 89128 38894
rect 89076 38830 89128 38836
rect 89088 38554 89116 38830
rect 89904 38820 89956 38826
rect 89904 38762 89956 38768
rect 89076 38548 89128 38554
rect 89076 38490 89128 38496
rect 89444 38480 89496 38486
rect 89444 38422 89496 38428
rect 88524 38344 88576 38350
rect 88524 38286 88576 38292
rect 88708 38208 88760 38214
rect 88708 38150 88760 38156
rect 88720 37466 88748 38150
rect 89456 37942 89484 38422
rect 89628 38208 89680 38214
rect 89628 38150 89680 38156
rect 89720 38208 89772 38214
rect 89720 38150 89772 38156
rect 89444 37936 89496 37942
rect 89444 37878 89496 37884
rect 88708 37460 88760 37466
rect 88708 37402 88760 37408
rect 86224 37324 86276 37330
rect 86224 37266 86276 37272
rect 86868 37324 86920 37330
rect 89640 37312 89668 38150
rect 89732 37806 89760 38150
rect 89916 37874 89944 38762
rect 90100 38554 90128 39306
rect 90088 38548 90140 38554
rect 90088 38490 90140 38496
rect 90100 38350 90128 38490
rect 91020 38486 91048 39442
rect 96380 39196 96676 39216
rect 96436 39194 96460 39196
rect 96516 39194 96540 39196
rect 96596 39194 96620 39196
rect 96458 39142 96460 39194
rect 96522 39142 96534 39194
rect 96596 39142 96598 39194
rect 96436 39140 96460 39142
rect 96516 39140 96540 39142
rect 96596 39140 96620 39142
rect 96380 39120 96676 39140
rect 91560 38888 91612 38894
rect 91560 38830 91612 38836
rect 91100 38820 91152 38826
rect 91100 38762 91152 38768
rect 91008 38480 91060 38486
rect 91008 38422 91060 38428
rect 91112 38418 91140 38762
rect 91100 38412 91152 38418
rect 91100 38354 91152 38360
rect 90088 38344 90140 38350
rect 90088 38286 90140 38292
rect 90916 38344 90968 38350
rect 90916 38286 90968 38292
rect 89904 37868 89956 37874
rect 89904 37810 89956 37816
rect 89720 37800 89772 37806
rect 89720 37742 89772 37748
rect 90732 37664 90784 37670
rect 90732 37606 90784 37612
rect 89720 37324 89772 37330
rect 89640 37284 89720 37312
rect 86868 37266 86920 37272
rect 89720 37266 89772 37272
rect 85580 36848 85632 36854
rect 85580 36790 85632 36796
rect 86236 36786 86264 37266
rect 86224 36780 86276 36786
rect 86224 36722 86276 36728
rect 85488 36712 85540 36718
rect 85488 36654 85540 36660
rect 84476 36236 84528 36242
rect 84476 36178 84528 36184
rect 86224 36168 86276 36174
rect 86224 36110 86276 36116
rect 85854 35864 85910 35873
rect 85854 35799 85910 35808
rect 85868 35766 85896 35799
rect 84476 35760 84528 35766
rect 85856 35760 85908 35766
rect 84476 35702 84528 35708
rect 85486 35728 85542 35737
rect 84292 35488 84344 35494
rect 84292 35430 84344 35436
rect 84488 35222 84516 35702
rect 85856 35702 85908 35708
rect 85764 35692 85816 35698
rect 85542 35672 85764 35680
rect 85486 35663 85764 35672
rect 85500 35652 85764 35663
rect 85396 35556 85448 35562
rect 85396 35498 85448 35504
rect 84476 35216 84528 35222
rect 83554 35184 83610 35193
rect 83280 35148 83332 35154
rect 84476 35158 84528 35164
rect 84752 35216 84804 35222
rect 84752 35158 84804 35164
rect 83554 35119 83610 35128
rect 84384 35148 84436 35154
rect 83280 35090 83332 35096
rect 83568 35018 83596 35119
rect 84384 35090 84436 35096
rect 84396 35057 84424 35090
rect 84764 35057 84792 35158
rect 85408 35154 85436 35498
rect 85396 35148 85448 35154
rect 85396 35090 85448 35096
rect 84382 35048 84438 35057
rect 82544 35012 82596 35018
rect 82544 34954 82596 34960
rect 83464 35012 83516 35018
rect 83464 34954 83516 34960
rect 83556 35012 83608 35018
rect 84382 34983 84438 34992
rect 84750 35048 84806 35057
rect 84750 34983 84806 34992
rect 83556 34954 83608 34960
rect 82556 34678 82584 34954
rect 82544 34672 82596 34678
rect 82544 34614 82596 34620
rect 82556 34542 82584 34614
rect 83476 34542 83504 34954
rect 85500 34678 85528 35652
rect 85764 35634 85816 35640
rect 86236 35222 86264 36110
rect 86776 36032 86828 36038
rect 86776 35974 86828 35980
rect 86788 35630 86816 35974
rect 86880 35834 86908 37266
rect 89732 37126 89760 37266
rect 87420 37120 87472 37126
rect 87420 37062 87472 37068
rect 89720 37120 89772 37126
rect 89720 37062 89772 37068
rect 86868 35828 86920 35834
rect 86868 35770 86920 35776
rect 86776 35624 86828 35630
rect 86776 35566 86828 35572
rect 87432 35290 87460 37062
rect 88432 36780 88484 36786
rect 88432 36722 88484 36728
rect 88444 36310 88472 36722
rect 89168 36644 89220 36650
rect 89168 36586 89220 36592
rect 90180 36644 90232 36650
rect 90180 36586 90232 36592
rect 88432 36304 88484 36310
rect 88432 36246 88484 36252
rect 88444 35698 88472 36246
rect 88432 35692 88484 35698
rect 88432 35634 88484 35640
rect 88156 35624 88208 35630
rect 88156 35566 88208 35572
rect 88248 35624 88300 35630
rect 88248 35566 88300 35572
rect 87420 35284 87472 35290
rect 87420 35226 87472 35232
rect 86040 35216 86092 35222
rect 86040 35158 86092 35164
rect 86224 35216 86276 35222
rect 86224 35158 86276 35164
rect 85580 35148 85632 35154
rect 85580 35090 85632 35096
rect 85592 35057 85620 35090
rect 86052 35057 86080 35158
rect 85578 35048 85634 35057
rect 85578 34983 85634 34992
rect 86038 35048 86094 35057
rect 86038 34983 86094 34992
rect 85488 34672 85540 34678
rect 85488 34614 85540 34620
rect 85500 34542 85528 34614
rect 82360 34536 82412 34542
rect 82360 34478 82412 34484
rect 82544 34536 82596 34542
rect 82544 34478 82596 34484
rect 83464 34536 83516 34542
rect 83464 34478 83516 34484
rect 85488 34536 85540 34542
rect 85488 34478 85540 34484
rect 82372 31657 82400 34478
rect 85592 34406 85620 34983
rect 88168 34746 88196 35566
rect 88260 35154 88288 35566
rect 88984 35488 89036 35494
rect 88984 35430 89036 35436
rect 88432 35284 88484 35290
rect 88432 35226 88484 35232
rect 88248 35148 88300 35154
rect 88248 35090 88300 35096
rect 88156 34740 88208 34746
rect 88156 34682 88208 34688
rect 88260 34542 88288 35090
rect 88340 34944 88392 34950
rect 88340 34886 88392 34892
rect 88352 34610 88380 34886
rect 88444 34678 88472 35226
rect 88432 34672 88484 34678
rect 88432 34614 88484 34620
rect 88340 34604 88392 34610
rect 88340 34546 88392 34552
rect 88996 34542 89024 35430
rect 89180 35086 89208 36586
rect 89720 36236 89772 36242
rect 89720 36178 89772 36184
rect 89536 36032 89588 36038
rect 89536 35974 89588 35980
rect 89548 35154 89576 35974
rect 89732 35698 89760 36178
rect 89720 35692 89772 35698
rect 89720 35634 89772 35640
rect 89536 35148 89588 35154
rect 89536 35090 89588 35096
rect 89168 35080 89220 35086
rect 89168 35022 89220 35028
rect 90192 34950 90220 36586
rect 90744 36174 90772 37606
rect 90928 36582 90956 38286
rect 91008 38208 91060 38214
rect 91008 38150 91060 38156
rect 91020 37738 91048 38150
rect 91284 37936 91336 37942
rect 91284 37878 91336 37884
rect 91008 37732 91060 37738
rect 91008 37674 91060 37680
rect 91020 37398 91048 37674
rect 91296 37398 91324 37878
rect 91572 37874 91600 38830
rect 93492 38820 93544 38826
rect 93492 38762 93544 38768
rect 93400 38752 93452 38758
rect 93400 38694 93452 38700
rect 93412 38554 93440 38694
rect 93400 38548 93452 38554
rect 93400 38490 93452 38496
rect 91560 37868 91612 37874
rect 91560 37810 91612 37816
rect 91572 37398 91600 37810
rect 91008 37392 91060 37398
rect 91008 37334 91060 37340
rect 91284 37392 91336 37398
rect 91284 37334 91336 37340
rect 91560 37392 91612 37398
rect 91560 37334 91612 37340
rect 91296 36922 91324 37334
rect 93412 36922 93440 38490
rect 93504 37806 93532 38762
rect 94596 38344 94648 38350
rect 94596 38286 94648 38292
rect 94504 38208 94556 38214
rect 94504 38150 94556 38156
rect 93492 37800 93544 37806
rect 93492 37742 93544 37748
rect 93584 37800 93636 37806
rect 93584 37742 93636 37748
rect 94516 37754 94544 38150
rect 94608 37874 94636 38286
rect 96380 38108 96676 38128
rect 96436 38106 96460 38108
rect 96516 38106 96540 38108
rect 96596 38106 96620 38108
rect 96458 38054 96460 38106
rect 96522 38054 96534 38106
rect 96596 38054 96598 38106
rect 96436 38052 96460 38054
rect 96516 38052 96540 38054
rect 96596 38052 96620 38054
rect 96380 38032 96676 38052
rect 94596 37868 94648 37874
rect 94596 37810 94648 37816
rect 95240 37800 95292 37806
rect 93596 37262 93624 37742
rect 94516 37726 94636 37754
rect 95240 37742 95292 37748
rect 97080 37800 97132 37806
rect 97080 37742 97132 37748
rect 94608 37398 94636 37726
rect 94596 37392 94648 37398
rect 94596 37334 94648 37340
rect 93584 37256 93636 37262
rect 93584 37198 93636 37204
rect 93676 37120 93728 37126
rect 93676 37062 93728 37068
rect 91008 36916 91060 36922
rect 91008 36858 91060 36864
rect 91284 36916 91336 36922
rect 91284 36858 91336 36864
rect 93400 36916 93452 36922
rect 93400 36858 93452 36864
rect 91020 36825 91048 36858
rect 91006 36816 91062 36825
rect 91006 36751 91062 36760
rect 91284 36780 91336 36786
rect 91284 36722 91336 36728
rect 90916 36576 90968 36582
rect 90916 36518 90968 36524
rect 90732 36168 90784 36174
rect 90732 36110 90784 36116
rect 90640 36032 90692 36038
rect 90640 35974 90692 35980
rect 90180 34944 90232 34950
rect 90180 34886 90232 34892
rect 90652 34542 90680 35974
rect 90744 35698 90772 36110
rect 90732 35692 90784 35698
rect 90732 35634 90784 35640
rect 91296 35630 91324 36722
rect 92756 36644 92808 36650
rect 92756 36586 92808 36592
rect 92768 36242 92796 36586
rect 91744 36236 91796 36242
rect 91744 36178 91796 36184
rect 92756 36236 92808 36242
rect 92756 36178 92808 36184
rect 91284 35624 91336 35630
rect 91284 35566 91336 35572
rect 91284 35488 91336 35494
rect 91284 35430 91336 35436
rect 91296 34746 91324 35430
rect 91756 35154 91784 36178
rect 93688 35630 93716 37062
rect 94044 36916 94096 36922
rect 94044 36858 94096 36864
rect 93952 36032 94004 36038
rect 93952 35974 94004 35980
rect 93676 35624 93728 35630
rect 93964 35612 93992 35974
rect 94056 35766 94084 36858
rect 94608 36174 94636 37334
rect 95252 37262 95280 37742
rect 95332 37732 95384 37738
rect 95332 37674 95384 37680
rect 95700 37732 95752 37738
rect 95700 37674 95752 37680
rect 95240 37256 95292 37262
rect 95240 37198 95292 37204
rect 95148 37188 95200 37194
rect 95148 37130 95200 37136
rect 95056 37120 95108 37126
rect 95056 37062 95108 37068
rect 95160 37074 95188 37130
rect 95068 36718 95096 37062
rect 95160 37046 95280 37074
rect 95252 36786 95280 37046
rect 95344 36922 95372 37674
rect 95712 37330 95740 37674
rect 96712 37664 96764 37670
rect 96712 37606 96764 37612
rect 96724 37466 96752 37606
rect 96712 37460 96764 37466
rect 96712 37402 96764 37408
rect 95700 37324 95752 37330
rect 95700 37266 95752 37272
rect 97092 37126 97120 37742
rect 97080 37120 97132 37126
rect 97080 37062 97132 37068
rect 96380 37020 96676 37040
rect 96436 37018 96460 37020
rect 96516 37018 96540 37020
rect 96596 37018 96620 37020
rect 96458 36966 96460 37018
rect 96522 36966 96534 37018
rect 96596 36966 96598 37018
rect 96436 36964 96460 36966
rect 96516 36964 96540 36966
rect 96596 36964 96620 36966
rect 96380 36944 96676 36964
rect 95332 36916 95384 36922
rect 95332 36858 95384 36864
rect 95330 36816 95386 36825
rect 95240 36780 95292 36786
rect 95330 36751 95386 36760
rect 95240 36722 95292 36728
rect 94688 36712 94740 36718
rect 94688 36654 94740 36660
rect 94964 36712 95016 36718
rect 94964 36654 95016 36660
rect 95056 36712 95108 36718
rect 95056 36654 95108 36660
rect 94700 36582 94728 36654
rect 94688 36576 94740 36582
rect 94688 36518 94740 36524
rect 94596 36168 94648 36174
rect 94596 36110 94648 36116
rect 94044 35760 94096 35766
rect 94044 35702 94096 35708
rect 93676 35566 93728 35572
rect 93872 35584 93992 35612
rect 91744 35148 91796 35154
rect 91744 35090 91796 35096
rect 93872 35086 93900 35584
rect 94056 35494 94084 35702
rect 94976 35630 95004 36654
rect 94964 35624 95016 35630
rect 94964 35566 95016 35572
rect 95068 35562 95096 36654
rect 95252 35698 95280 36722
rect 95344 36718 95372 36751
rect 95332 36712 95384 36718
rect 95332 36654 95384 36660
rect 97092 36242 97120 37062
rect 97264 36712 97316 36718
rect 97264 36654 97316 36660
rect 97276 36378 97304 36654
rect 97264 36372 97316 36378
rect 97264 36314 97316 36320
rect 97080 36236 97132 36242
rect 97080 36178 97132 36184
rect 96712 36032 96764 36038
rect 96712 35974 96764 35980
rect 96380 35932 96676 35952
rect 96436 35930 96460 35932
rect 96516 35930 96540 35932
rect 96596 35930 96620 35932
rect 96458 35878 96460 35930
rect 96522 35878 96534 35930
rect 96596 35878 96598 35930
rect 96436 35876 96460 35878
rect 96516 35876 96540 35878
rect 96596 35876 96620 35878
rect 96380 35856 96676 35876
rect 95240 35692 95292 35698
rect 95240 35634 95292 35640
rect 96724 35630 96752 35974
rect 96712 35624 96764 35630
rect 96712 35566 96764 35572
rect 94136 35556 94188 35562
rect 94136 35498 94188 35504
rect 95056 35556 95108 35562
rect 95056 35498 95108 35504
rect 94044 35488 94096 35494
rect 94044 35430 94096 35436
rect 94148 35154 94176 35498
rect 94136 35148 94188 35154
rect 94136 35090 94188 35096
rect 93860 35080 93912 35086
rect 93860 35022 93912 35028
rect 96380 34844 96676 34864
rect 96436 34842 96460 34844
rect 96516 34842 96540 34844
rect 96596 34842 96620 34844
rect 96458 34790 96460 34842
rect 96522 34790 96534 34842
rect 96596 34790 96598 34842
rect 96436 34788 96460 34790
rect 96516 34788 96540 34790
rect 96596 34788 96620 34790
rect 96380 34768 96676 34788
rect 91284 34740 91336 34746
rect 91284 34682 91336 34688
rect 88248 34536 88300 34542
rect 88248 34478 88300 34484
rect 88984 34536 89036 34542
rect 88984 34478 89036 34484
rect 90640 34536 90692 34542
rect 90640 34478 90692 34484
rect 85580 34400 85632 34406
rect 85580 34342 85632 34348
rect 82358 31648 82414 31657
rect 82358 31583 82414 31592
rect 82268 22908 82320 22914
rect 82268 22850 82320 22856
rect 81636 21270 82124 21298
rect 80886 20088 80942 20097
rect 80886 20023 80942 20032
rect 81636 16017 81664 21270
rect 81622 16008 81678 16017
rect 81622 15943 81678 15952
rect 81636 14861 81664 15943
rect 81622 14852 81678 14861
rect 81622 14787 81678 14796
rect 79966 4856 80022 4865
rect 79966 4791 80022 4800
rect 52552 944 52604 950
rect 52552 886 52604 892
rect 53380 944 53432 950
rect 53380 886 53432 892
rect 53392 800 53420 886
rect 2780 468 2832 474
rect 2780 410 2832 416
rect 5356 468 5408 474
rect 5356 410 5408 416
rect 2792 377 2820 410
rect 2778 368 2834 377
rect 2778 303 2834 312
rect 53378 0 53434 800
<< via2 >>
rect 3606 45872 3662 45928
rect 2778 44648 2834 44704
rect 3514 44104 3570 44160
rect 1490 40568 1546 40624
rect 3330 40024 3386 40080
rect 3238 38800 3294 38856
rect 3238 34040 3294 34096
rect 3422 35264 3478 35320
rect 3054 31048 3110 31104
rect 2962 29824 3018 29880
rect 3054 28872 3110 28928
rect 2962 16904 3018 16960
rect 2870 2624 2926 2680
rect 4066 45328 4122 45384
rect 19580 44090 19636 44092
rect 19660 44090 19716 44092
rect 19740 44090 19796 44092
rect 19820 44090 19876 44092
rect 19580 44038 19606 44090
rect 19606 44038 19636 44090
rect 19660 44038 19670 44090
rect 19670 44038 19716 44090
rect 19740 44038 19786 44090
rect 19786 44038 19796 44090
rect 19820 44038 19850 44090
rect 19850 44038 19876 44090
rect 19580 44036 19636 44038
rect 19660 44036 19716 44038
rect 19740 44036 19796 44038
rect 19820 44036 19876 44038
rect 50300 44090 50356 44092
rect 50380 44090 50436 44092
rect 50460 44090 50516 44092
rect 50540 44090 50596 44092
rect 50300 44038 50326 44090
rect 50326 44038 50356 44090
rect 50380 44038 50390 44090
rect 50390 44038 50436 44090
rect 50460 44038 50506 44090
rect 50506 44038 50516 44090
rect 50540 44038 50570 44090
rect 50570 44038 50596 44090
rect 50300 44036 50356 44038
rect 50380 44036 50436 44038
rect 50460 44036 50516 44038
rect 50540 44036 50596 44038
rect 4220 43546 4276 43548
rect 4300 43546 4356 43548
rect 4380 43546 4436 43548
rect 4460 43546 4516 43548
rect 4220 43494 4246 43546
rect 4246 43494 4276 43546
rect 4300 43494 4310 43546
rect 4310 43494 4356 43546
rect 4380 43494 4426 43546
rect 4426 43494 4436 43546
rect 4460 43494 4490 43546
rect 4490 43494 4516 43546
rect 4220 43492 4276 43494
rect 4300 43492 4356 43494
rect 4380 43492 4436 43494
rect 4460 43492 4516 43494
rect 4220 42458 4276 42460
rect 4300 42458 4356 42460
rect 4380 42458 4436 42460
rect 4460 42458 4516 42460
rect 4220 42406 4246 42458
rect 4246 42406 4276 42458
rect 4300 42406 4310 42458
rect 4310 42406 4356 42458
rect 4380 42406 4426 42458
rect 4426 42406 4436 42458
rect 4460 42406 4490 42458
rect 4490 42406 4516 42458
rect 4220 42404 4276 42406
rect 4300 42404 4356 42406
rect 4380 42404 4436 42406
rect 4460 42404 4516 42406
rect 4220 41370 4276 41372
rect 4300 41370 4356 41372
rect 4380 41370 4436 41372
rect 4460 41370 4516 41372
rect 4220 41318 4246 41370
rect 4246 41318 4276 41370
rect 4300 41318 4310 41370
rect 4310 41318 4356 41370
rect 4380 41318 4426 41370
rect 4426 41318 4436 41370
rect 4460 41318 4490 41370
rect 4490 41318 4516 41370
rect 4220 41316 4276 41318
rect 4300 41316 4356 41318
rect 4380 41316 4436 41318
rect 4460 41316 4516 41318
rect 3882 41112 3938 41168
rect 4220 40282 4276 40284
rect 4300 40282 4356 40284
rect 4380 40282 4436 40284
rect 4460 40282 4516 40284
rect 4220 40230 4246 40282
rect 4246 40230 4276 40282
rect 4300 40230 4310 40282
rect 4310 40230 4356 40282
rect 4380 40230 4426 40282
rect 4426 40230 4436 40282
rect 4460 40230 4490 40282
rect 4490 40230 4516 40282
rect 4220 40228 4276 40230
rect 4300 40228 4356 40230
rect 4380 40228 4436 40230
rect 4460 40228 4516 40230
rect 3974 39344 4030 39400
rect 4220 39194 4276 39196
rect 4300 39194 4356 39196
rect 4380 39194 4436 39196
rect 4460 39194 4516 39196
rect 4220 39142 4246 39194
rect 4246 39142 4276 39194
rect 4300 39142 4310 39194
rect 4310 39142 4356 39194
rect 4380 39142 4426 39194
rect 4426 39142 4436 39194
rect 4460 39142 4490 39194
rect 4490 39142 4516 39194
rect 4220 39140 4276 39142
rect 4300 39140 4356 39142
rect 4380 39140 4436 39142
rect 4460 39140 4516 39142
rect 4066 38120 4122 38176
rect 4220 38106 4276 38108
rect 4300 38106 4356 38108
rect 4380 38106 4436 38108
rect 4460 38106 4516 38108
rect 4220 38054 4246 38106
rect 4246 38054 4276 38106
rect 4300 38054 4310 38106
rect 4310 38054 4356 38106
rect 4380 38054 4426 38106
rect 4426 38054 4436 38106
rect 4460 38054 4490 38106
rect 4490 38054 4516 38106
rect 4220 38052 4276 38054
rect 4300 38052 4356 38054
rect 4380 38052 4436 38054
rect 4460 38052 4516 38054
rect 3882 37576 3938 37632
rect 3974 37032 4030 37088
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 4066 36352 4122 36408
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 4066 35808 4122 35864
rect 3882 34584 3938 34640
rect 3422 31728 3478 31784
rect 3330 28872 3386 28928
rect 3882 32816 3938 32872
rect 3238 23432 3294 23488
rect 3330 20440 3386 20496
rect 3146 19760 3202 19816
rect 3330 19216 3386 19272
rect 3698 17992 3754 18048
rect 3698 16224 3754 16280
rect 3606 15680 3662 15736
rect 3882 30504 3938 30560
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 4066 33496 4122 33552
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 4066 29280 4122 29336
rect 4066 28736 4122 28792
rect 3882 28056 3938 28112
rect 3882 26968 3938 27024
rect 3882 25744 3938 25800
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 4066 27512 4122 27568
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 4066 26288 4122 26344
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 4066 25200 4122 25256
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 3882 24520 3938 24576
rect 4066 23976 4122 24032
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 4066 22752 4122 22808
rect 3882 22208 3938 22264
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 4066 20984 4122 21040
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 3882 18672 3938 18728
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 3882 17448 3938 17504
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 3882 15000 3938 15056
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 3882 13912 3938 13968
rect 4066 13232 4122 13288
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 3882 12688 3938 12744
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 3882 11500 3884 11520
rect 3884 11500 3936 11520
rect 3936 11500 3938 11520
rect 3882 11464 3938 11500
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 3882 10412 3884 10432
rect 3884 10412 3936 10432
rect 3936 10412 3938 10432
rect 3882 10376 3938 10412
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 3882 9152 3938 9208
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4066 8608 4122 8664
rect 3882 7928 3938 7984
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 4066 7384 4122 7440
rect 3882 6704 3938 6760
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4066 6160 4122 6216
rect 3882 5616 3938 5672
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 3882 4392 3938 4448
rect 4066 4936 4122 4992
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 3882 3168 3938 3224
rect 4066 3848 4122 3904
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 5906 32272 5962 32328
rect 7378 39380 7380 39400
rect 7380 39380 7432 39400
rect 7432 39380 7434 39400
rect 7378 39344 7434 39380
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 3514 2080 3570 2136
rect 2962 1400 3018 1456
rect 2778 856 2834 912
rect 7102 19236 7158 19272
rect 7102 19216 7104 19236
rect 7104 19216 7156 19236
rect 7156 19216 7158 19236
rect 7194 19080 7250 19136
rect 7838 39500 7894 39536
rect 7838 39480 7840 39500
rect 7840 39480 7892 39500
rect 7892 39480 7894 39500
rect 7746 39364 7802 39400
rect 7746 39344 7748 39364
rect 7748 39344 7800 39364
rect 7800 39344 7802 39364
rect 8298 39516 8300 39536
rect 8300 39516 8352 39536
rect 8352 39516 8354 39536
rect 8298 39480 8354 39516
rect 7470 26152 7526 26208
rect 8390 31864 8446 31920
rect 8482 27376 8538 27432
rect 7470 12180 7472 12200
rect 7472 12180 7524 12200
rect 7524 12180 7526 12200
rect 7470 12144 7526 12180
rect 8114 18672 8170 18728
rect 9954 31900 9956 31920
rect 9956 31900 10008 31920
rect 10008 31900 10010 31920
rect 9954 31864 10010 31900
rect 9678 31456 9734 31512
rect 8850 19216 8906 19272
rect 8482 19080 8538 19136
rect 8482 18672 8538 18728
rect 8022 10668 8078 10704
rect 8022 10648 8024 10668
rect 8024 10648 8076 10668
rect 8076 10648 8078 10668
rect 9126 18672 9182 18728
rect 9586 27512 9642 27568
rect 9770 27376 9826 27432
rect 9678 22772 9734 22808
rect 9678 22752 9680 22772
rect 9680 22752 9732 22772
rect 9732 22752 9734 22772
rect 9494 21528 9550 21584
rect 8666 14456 8722 14512
rect 8114 9968 8170 10024
rect 9494 18028 9496 18048
rect 9496 18028 9548 18048
rect 9548 18028 9550 18048
rect 9494 17992 9550 18028
rect 11794 37712 11850 37768
rect 12254 36760 12310 36816
rect 12346 36660 12348 36680
rect 12348 36660 12400 36680
rect 12400 36660 12402 36680
rect 12346 36624 12402 36660
rect 14278 39480 14334 39536
rect 14462 39244 14464 39264
rect 14464 39244 14516 39264
rect 14516 39244 14518 39264
rect 14462 39208 14518 39244
rect 14094 38936 14150 38992
rect 11794 31476 11850 31512
rect 11794 31456 11796 31476
rect 11796 31456 11848 31476
rect 11848 31456 11850 31476
rect 9770 7404 9826 7440
rect 9770 7384 9772 7404
rect 9772 7384 9824 7404
rect 9824 7384 9826 7404
rect 13174 36116 13176 36136
rect 13176 36116 13228 36136
rect 13228 36116 13230 36136
rect 13174 36080 13230 36116
rect 14554 37324 14610 37360
rect 14554 37304 14556 37324
rect 14556 37304 14608 37324
rect 14608 37304 14610 37324
rect 14094 36660 14096 36680
rect 14096 36660 14148 36680
rect 14148 36660 14150 36680
rect 14094 36624 14150 36660
rect 12438 27512 12494 27568
rect 12622 23432 12678 23488
rect 15474 37712 15530 37768
rect 14646 35028 14648 35048
rect 14648 35028 14700 35048
rect 14700 35028 14702 35048
rect 14646 34992 14702 35028
rect 19580 43002 19636 43004
rect 19660 43002 19716 43004
rect 19740 43002 19796 43004
rect 19820 43002 19876 43004
rect 19580 42950 19606 43002
rect 19606 42950 19636 43002
rect 19660 42950 19670 43002
rect 19670 42950 19716 43002
rect 19740 42950 19786 43002
rect 19786 42950 19796 43002
rect 19820 42950 19850 43002
rect 19850 42950 19876 43002
rect 19580 42948 19636 42950
rect 19660 42948 19716 42950
rect 19740 42948 19796 42950
rect 19820 42948 19876 42950
rect 19580 41914 19636 41916
rect 19660 41914 19716 41916
rect 19740 41914 19796 41916
rect 19820 41914 19876 41916
rect 19580 41862 19606 41914
rect 19606 41862 19636 41914
rect 19660 41862 19670 41914
rect 19670 41862 19716 41914
rect 19740 41862 19786 41914
rect 19786 41862 19796 41914
rect 19820 41862 19850 41914
rect 19850 41862 19876 41914
rect 19580 41860 19636 41862
rect 19660 41860 19716 41862
rect 19740 41860 19796 41862
rect 19820 41860 19876 41862
rect 19580 40826 19636 40828
rect 19660 40826 19716 40828
rect 19740 40826 19796 40828
rect 19820 40826 19876 40828
rect 19580 40774 19606 40826
rect 19606 40774 19636 40826
rect 19660 40774 19670 40826
rect 19670 40774 19716 40826
rect 19740 40774 19786 40826
rect 19786 40774 19796 40826
rect 19820 40774 19850 40826
rect 19850 40774 19876 40826
rect 19580 40772 19636 40774
rect 19660 40772 19716 40774
rect 19740 40772 19796 40774
rect 19820 40772 19876 40774
rect 19062 39208 19118 39264
rect 19246 39208 19302 39264
rect 19580 39738 19636 39740
rect 19660 39738 19716 39740
rect 19740 39738 19796 39740
rect 19820 39738 19876 39740
rect 19580 39686 19606 39738
rect 19606 39686 19636 39738
rect 19660 39686 19670 39738
rect 19670 39686 19716 39738
rect 19740 39686 19786 39738
rect 19786 39686 19796 39738
rect 19820 39686 19850 39738
rect 19850 39686 19876 39738
rect 19580 39684 19636 39686
rect 19660 39684 19716 39686
rect 19740 39684 19796 39686
rect 19820 39684 19876 39686
rect 19580 38650 19636 38652
rect 19660 38650 19716 38652
rect 19740 38650 19796 38652
rect 19820 38650 19876 38652
rect 19580 38598 19606 38650
rect 19606 38598 19636 38650
rect 19660 38598 19670 38650
rect 19670 38598 19716 38650
rect 19740 38598 19786 38650
rect 19786 38598 19796 38650
rect 19820 38598 19850 38650
rect 19850 38598 19876 38650
rect 19580 38596 19636 38598
rect 19660 38596 19716 38598
rect 19740 38596 19796 38598
rect 19820 38596 19876 38598
rect 18142 37748 18144 37768
rect 18144 37748 18196 37768
rect 18196 37748 18198 37768
rect 18142 37712 18198 37748
rect 13266 14592 13322 14648
rect 13634 7384 13690 7440
rect 16394 15952 16450 16008
rect 18050 33768 18106 33824
rect 19430 38392 19486 38448
rect 19430 38256 19486 38312
rect 19338 37712 19394 37768
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 19338 37168 19394 37224
rect 19246 36760 19302 36816
rect 18970 36644 19026 36680
rect 21822 42200 21878 42256
rect 21638 39208 21694 39264
rect 21178 37868 21234 37904
rect 21178 37848 21180 37868
rect 21180 37848 21232 37868
rect 21232 37848 21234 37868
rect 22190 37848 22246 37904
rect 20166 37168 20222 37224
rect 18970 36624 18972 36644
rect 18972 36624 19024 36644
rect 19024 36624 19026 36644
rect 19890 36624 19946 36680
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 20166 36216 20222 36272
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 19706 35164 19708 35184
rect 19708 35164 19760 35184
rect 19760 35164 19762 35184
rect 19706 35128 19762 35164
rect 20074 34604 20130 34640
rect 20074 34584 20076 34604
rect 20076 34584 20128 34604
rect 20128 34584 20130 34604
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 21270 34720 21326 34776
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 19522 28620 19578 28656
rect 19522 28600 19524 28620
rect 19524 28600 19576 28620
rect 19576 28600 19578 28620
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 18510 16652 18566 16688
rect 18510 16632 18512 16652
rect 18512 16632 18564 16652
rect 18564 16632 18566 16652
rect 19154 17312 19210 17368
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 21178 34076 21180 34096
rect 21180 34076 21232 34096
rect 21232 34076 21234 34096
rect 21178 34040 21234 34076
rect 22282 34740 22338 34776
rect 22282 34720 22284 34740
rect 22284 34720 22336 34740
rect 22336 34720 22338 34740
rect 20442 33924 20498 33960
rect 20442 33904 20444 33924
rect 20444 33904 20496 33924
rect 20496 33904 20498 33924
rect 21270 33496 21326 33552
rect 20994 33396 20996 33416
rect 20996 33396 21048 33416
rect 21048 33396 21050 33416
rect 20994 33360 21050 33396
rect 22190 33496 22246 33552
rect 34940 43546 34996 43548
rect 35020 43546 35076 43548
rect 35100 43546 35156 43548
rect 35180 43546 35236 43548
rect 34940 43494 34966 43546
rect 34966 43494 34996 43546
rect 35020 43494 35030 43546
rect 35030 43494 35076 43546
rect 35100 43494 35146 43546
rect 35146 43494 35156 43546
rect 35180 43494 35210 43546
rect 35210 43494 35236 43546
rect 34940 43492 34996 43494
rect 35020 43492 35076 43494
rect 35100 43492 35156 43494
rect 35180 43492 35236 43494
rect 29366 42744 29422 42800
rect 28170 42200 28226 42256
rect 23386 37748 23388 37768
rect 23388 37748 23440 37768
rect 23440 37748 23442 37768
rect 23386 37712 23442 37748
rect 28998 40432 29054 40488
rect 24858 36216 24914 36272
rect 24122 35692 24178 35728
rect 24122 35672 24124 35692
rect 24124 35672 24176 35692
rect 24176 35672 24178 35692
rect 22926 34584 22982 34640
rect 22374 33360 22430 33416
rect 21638 31900 21640 31920
rect 21640 31900 21692 31920
rect 21692 31900 21694 31920
rect 21638 31864 21694 31900
rect 22282 31884 22338 31920
rect 22282 31864 22284 31884
rect 22284 31864 22336 31884
rect 22336 31864 22338 31884
rect 20166 23468 20168 23488
rect 20168 23468 20220 23488
rect 20220 23468 20222 23488
rect 20166 23432 20222 23468
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 19890 17312 19946 17368
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 21270 22108 21272 22128
rect 21272 22108 21324 22128
rect 21324 22108 21326 22128
rect 21270 22072 21326 22108
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 21914 15308 21916 15328
rect 21916 15308 21968 15328
rect 21968 15308 21970 15328
rect 21914 15272 21970 15308
rect 22650 28600 22706 28656
rect 25502 35128 25558 35184
rect 24858 34040 24914 34096
rect 24582 33904 24638 33960
rect 24214 30776 24270 30832
rect 23478 30096 23534 30152
rect 23386 28056 23442 28112
rect 23570 24112 23626 24168
rect 23478 22752 23534 22808
rect 23478 20032 23534 20088
rect 23386 14728 23442 14784
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 24306 26696 24362 26752
rect 24766 29416 24822 29472
rect 26974 35692 27030 35728
rect 26974 35672 26976 35692
rect 26976 35672 27028 35692
rect 27028 35672 27030 35692
rect 26606 34720 26662 34776
rect 24766 25472 24822 25528
rect 28078 39208 28134 39264
rect 31666 40432 31722 40488
rect 31574 39908 31630 39944
rect 31574 39888 31576 39908
rect 31576 39888 31628 39908
rect 31628 39888 31630 39908
rect 32402 41520 32458 41576
rect 32494 41012 32496 41032
rect 32496 41012 32548 41032
rect 32548 41012 32550 41032
rect 32494 40976 32550 41012
rect 32770 40432 32826 40488
rect 32402 39924 32404 39944
rect 32404 39924 32456 39944
rect 32456 39924 32458 39944
rect 32402 39888 32458 39924
rect 32678 39888 32734 39944
rect 29550 36236 29606 36272
rect 29550 36216 29552 36236
rect 29552 36216 29604 36236
rect 29604 36216 29606 36236
rect 30194 35536 30250 35592
rect 27526 33768 27582 33824
rect 30562 35128 30618 35184
rect 38198 42744 38254 42800
rect 34978 42644 34980 42664
rect 34980 42644 35032 42664
rect 35032 42644 35034 42664
rect 34978 42608 35034 42644
rect 37738 42644 37740 42664
rect 37740 42644 37792 42664
rect 37792 42644 37794 42664
rect 37738 42608 37794 42644
rect 34940 42458 34996 42460
rect 35020 42458 35076 42460
rect 35100 42458 35156 42460
rect 35180 42458 35236 42460
rect 34940 42406 34966 42458
rect 34966 42406 34996 42458
rect 35020 42406 35030 42458
rect 35030 42406 35076 42458
rect 35100 42406 35146 42458
rect 35146 42406 35156 42458
rect 35180 42406 35210 42458
rect 35210 42406 35236 42458
rect 34940 42404 34996 42406
rect 35020 42404 35076 42406
rect 35100 42404 35156 42406
rect 35180 42404 35236 42406
rect 37094 42220 37150 42256
rect 37094 42200 37096 42220
rect 37096 42200 37148 42220
rect 37148 42200 37150 42220
rect 33690 41540 33746 41576
rect 33690 41520 33692 41540
rect 33692 41520 33744 41540
rect 33744 41520 33746 41540
rect 33322 40976 33378 41032
rect 33046 39752 33102 39808
rect 34426 39888 34482 39944
rect 34940 41370 34996 41372
rect 35020 41370 35076 41372
rect 35100 41370 35156 41372
rect 35180 41370 35236 41372
rect 34940 41318 34966 41370
rect 34966 41318 34996 41370
rect 35020 41318 35030 41370
rect 35030 41318 35076 41370
rect 35100 41318 35146 41370
rect 35146 41318 35156 41370
rect 35180 41318 35210 41370
rect 35210 41318 35236 41370
rect 34940 41316 34996 41318
rect 35020 41316 35076 41318
rect 35100 41316 35156 41318
rect 35180 41316 35236 41318
rect 34940 40282 34996 40284
rect 35020 40282 35076 40284
rect 35100 40282 35156 40284
rect 35180 40282 35236 40284
rect 34940 40230 34966 40282
rect 34966 40230 34996 40282
rect 35020 40230 35030 40282
rect 35030 40230 35076 40282
rect 35100 40230 35146 40282
rect 35146 40230 35156 40282
rect 35180 40230 35210 40282
rect 35210 40230 35236 40282
rect 34940 40228 34996 40230
rect 35020 40228 35076 40230
rect 35100 40228 35156 40230
rect 35180 40228 35236 40230
rect 33598 37748 33600 37768
rect 33600 37748 33652 37768
rect 33652 37748 33654 37768
rect 33598 37712 33654 37748
rect 34940 39194 34996 39196
rect 35020 39194 35076 39196
rect 35100 39194 35156 39196
rect 35180 39194 35236 39196
rect 34940 39142 34966 39194
rect 34966 39142 34996 39194
rect 35020 39142 35030 39194
rect 35030 39142 35076 39194
rect 35100 39142 35146 39194
rect 35146 39142 35156 39194
rect 35180 39142 35210 39194
rect 35210 39142 35236 39194
rect 34940 39140 34996 39142
rect 35020 39140 35076 39142
rect 35100 39140 35156 39142
rect 35180 39140 35236 39142
rect 34940 38106 34996 38108
rect 35020 38106 35076 38108
rect 35100 38106 35156 38108
rect 35180 38106 35236 38108
rect 34940 38054 34966 38106
rect 34966 38054 34996 38106
rect 35020 38054 35030 38106
rect 35030 38054 35076 38106
rect 35100 38054 35146 38106
rect 35146 38054 35156 38106
rect 35180 38054 35210 38106
rect 35210 38054 35236 38106
rect 34940 38052 34996 38054
rect 35020 38052 35076 38054
rect 35100 38052 35156 38054
rect 35180 38052 35236 38054
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 35622 36236 35678 36272
rect 35622 36216 35624 36236
rect 35624 36216 35676 36236
rect 35676 36216 35678 36236
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 36450 35572 36452 35592
rect 36452 35572 36504 35592
rect 36504 35572 36506 35592
rect 36450 35536 36506 35572
rect 33874 34584 33930 34640
rect 38566 39752 38622 39808
rect 38566 39616 38622 39672
rect 38566 39344 38622 39400
rect 38658 39092 38714 39128
rect 38658 39072 38660 39092
rect 38660 39072 38712 39092
rect 38712 39072 38714 39092
rect 39118 42200 39174 42256
rect 38934 41420 38936 41440
rect 38936 41420 38988 41440
rect 38988 41420 38990 41440
rect 38934 41384 38990 41420
rect 39118 41540 39174 41576
rect 39118 41520 39120 41540
rect 39120 41520 39172 41540
rect 39172 41520 39174 41540
rect 39302 40332 39304 40352
rect 39304 40332 39356 40352
rect 39356 40332 39358 40352
rect 39302 40296 39358 40332
rect 40958 42608 41014 42664
rect 43442 41420 43444 41440
rect 43444 41420 43496 41440
rect 43496 41420 43498 41440
rect 43442 41384 43498 41420
rect 36818 35164 36820 35184
rect 36820 35164 36872 35184
rect 36872 35164 36874 35184
rect 36818 35128 36874 35164
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 38750 34856 38806 34912
rect 38842 34740 38898 34776
rect 39946 38256 40002 38312
rect 40498 38292 40500 38312
rect 40500 38292 40552 38312
rect 40552 38292 40554 38312
rect 40498 38256 40554 38292
rect 40406 37576 40462 37632
rect 42982 38528 43038 38584
rect 41234 37868 41290 37904
rect 41234 37848 41236 37868
rect 41236 37848 41288 37868
rect 41288 37848 41290 37868
rect 40866 37460 40922 37496
rect 40866 37440 40868 37460
rect 40868 37440 40920 37460
rect 40920 37440 40922 37460
rect 40130 36080 40186 36136
rect 39578 35148 39634 35184
rect 39578 35128 39580 35148
rect 39580 35128 39632 35148
rect 39632 35128 39634 35148
rect 43166 36796 43168 36816
rect 43168 36796 43220 36816
rect 43220 36796 43222 36816
rect 43166 36760 43222 36796
rect 45098 39924 45100 39944
rect 45100 39924 45152 39944
rect 45152 39924 45154 39944
rect 41786 35264 41842 35320
rect 38842 34720 38844 34740
rect 38844 34720 38896 34740
rect 38896 34720 38898 34740
rect 40590 34720 40646 34776
rect 45098 39888 45154 39924
rect 44270 38800 44326 38856
rect 48318 42100 48320 42120
rect 48320 42100 48372 42120
rect 48372 42100 48374 42120
rect 48318 42064 48374 42100
rect 48594 41656 48650 41712
rect 49514 42064 49570 42120
rect 48226 40296 48282 40352
rect 49146 40296 49202 40352
rect 49238 40160 49294 40216
rect 49054 40024 49110 40080
rect 50300 43002 50356 43004
rect 50380 43002 50436 43004
rect 50460 43002 50516 43004
rect 50540 43002 50596 43004
rect 50300 42950 50326 43002
rect 50326 42950 50356 43002
rect 50380 42950 50390 43002
rect 50390 42950 50436 43002
rect 50460 42950 50506 43002
rect 50506 42950 50516 43002
rect 50540 42950 50570 43002
rect 50570 42950 50596 43002
rect 50300 42948 50356 42950
rect 50380 42948 50436 42950
rect 50460 42948 50516 42950
rect 50540 42948 50596 42950
rect 49882 41676 49938 41712
rect 49882 41656 49884 41676
rect 49884 41656 49936 41676
rect 49936 41656 49938 41676
rect 50300 41914 50356 41916
rect 50380 41914 50436 41916
rect 50460 41914 50516 41916
rect 50540 41914 50596 41916
rect 50300 41862 50326 41914
rect 50326 41862 50356 41914
rect 50380 41862 50390 41914
rect 50390 41862 50436 41914
rect 50460 41862 50506 41914
rect 50506 41862 50516 41914
rect 50540 41862 50570 41914
rect 50570 41862 50596 41914
rect 50300 41860 50356 41862
rect 50380 41860 50436 41862
rect 50460 41860 50516 41862
rect 50540 41860 50596 41862
rect 50300 40826 50356 40828
rect 50380 40826 50436 40828
rect 50460 40826 50516 40828
rect 50540 40826 50596 40828
rect 50300 40774 50326 40826
rect 50326 40774 50356 40826
rect 50380 40774 50390 40826
rect 50390 40774 50436 40826
rect 50460 40774 50506 40826
rect 50506 40774 50516 40826
rect 50540 40774 50570 40826
rect 50570 40774 50596 40826
rect 50300 40772 50356 40774
rect 50380 40772 50436 40774
rect 50460 40772 50516 40774
rect 50540 40772 50596 40774
rect 49790 40296 49846 40352
rect 51078 40024 51134 40080
rect 49330 39616 49386 39672
rect 48226 39072 48282 39128
rect 48226 38528 48282 38584
rect 45834 37576 45890 37632
rect 46202 37440 46258 37496
rect 48962 39380 48964 39400
rect 48964 39380 49016 39400
rect 49016 39380 49018 39400
rect 48962 39344 49018 39380
rect 48962 39072 49018 39128
rect 50300 39738 50356 39740
rect 50380 39738 50436 39740
rect 50460 39738 50516 39740
rect 50540 39738 50596 39740
rect 50300 39686 50326 39738
rect 50326 39686 50356 39738
rect 50380 39686 50390 39738
rect 50390 39686 50436 39738
rect 50460 39686 50506 39738
rect 50506 39686 50516 39738
rect 50540 39686 50570 39738
rect 50570 39686 50596 39738
rect 50300 39684 50356 39686
rect 50380 39684 50436 39686
rect 50460 39684 50516 39686
rect 50540 39684 50596 39686
rect 50158 39636 50214 39672
rect 50158 39616 50160 39636
rect 50160 39616 50212 39636
rect 50212 39616 50214 39636
rect 50710 39636 50766 39672
rect 50710 39616 50712 39636
rect 50712 39616 50764 39636
rect 50764 39616 50766 39636
rect 50066 39072 50122 39128
rect 50802 39344 50858 39400
rect 50300 38650 50356 38652
rect 50380 38650 50436 38652
rect 50460 38650 50516 38652
rect 50540 38650 50596 38652
rect 50300 38598 50326 38650
rect 50326 38598 50356 38650
rect 50380 38598 50390 38650
rect 50390 38598 50436 38650
rect 50460 38598 50506 38650
rect 50506 38598 50516 38650
rect 50540 38598 50570 38650
rect 50570 38598 50596 38650
rect 50300 38596 50356 38598
rect 50380 38596 50436 38598
rect 50460 38596 50516 38598
rect 50540 38596 50596 38598
rect 50342 38412 50398 38448
rect 50342 38392 50344 38412
rect 50344 38392 50396 38412
rect 50396 38392 50398 38412
rect 50066 38256 50122 38312
rect 50710 37984 50766 38040
rect 48042 36796 48044 36816
rect 48044 36796 48096 36816
rect 48096 36796 48098 36816
rect 48042 36760 48098 36796
rect 48962 37168 49018 37224
rect 50300 37562 50356 37564
rect 50380 37562 50436 37564
rect 50460 37562 50516 37564
rect 50540 37562 50596 37564
rect 50300 37510 50326 37562
rect 50326 37510 50356 37562
rect 50380 37510 50390 37562
rect 50390 37510 50436 37562
rect 50460 37510 50506 37562
rect 50506 37510 50516 37562
rect 50540 37510 50570 37562
rect 50570 37510 50596 37562
rect 50300 37508 50356 37510
rect 50380 37508 50436 37510
rect 50460 37508 50516 37510
rect 50540 37508 50596 37510
rect 51262 38256 51318 38312
rect 51538 39752 51594 39808
rect 51630 39380 51632 39400
rect 51632 39380 51684 39400
rect 51684 39380 51686 39400
rect 51630 39344 51686 39380
rect 51906 38664 51962 38720
rect 51814 38392 51870 38448
rect 47766 35264 47822 35320
rect 46846 34892 46848 34912
rect 46848 34892 46900 34912
rect 46900 34892 46902 34912
rect 46846 34856 46902 34892
rect 49422 35536 49478 35592
rect 49882 35808 49938 35864
rect 50434 36796 50436 36816
rect 50436 36796 50488 36816
rect 50488 36796 50490 36816
rect 50434 36760 50490 36796
rect 50300 36474 50356 36476
rect 50380 36474 50436 36476
rect 50460 36474 50516 36476
rect 50540 36474 50596 36476
rect 50300 36422 50326 36474
rect 50326 36422 50356 36474
rect 50380 36422 50390 36474
rect 50390 36422 50436 36474
rect 50460 36422 50506 36474
rect 50506 36422 50516 36474
rect 50540 36422 50570 36474
rect 50570 36422 50596 36474
rect 50300 36420 50356 36422
rect 50380 36420 50436 36422
rect 50460 36420 50516 36422
rect 50540 36420 50596 36422
rect 52826 39752 52882 39808
rect 52642 39616 52698 39672
rect 52366 39072 52422 39128
rect 50894 35400 50950 35456
rect 50300 35386 50356 35388
rect 50380 35386 50436 35388
rect 50460 35386 50516 35388
rect 50540 35386 50596 35388
rect 50300 35334 50326 35386
rect 50326 35334 50356 35386
rect 50380 35334 50390 35386
rect 50390 35334 50436 35386
rect 50460 35334 50506 35386
rect 50506 35334 50516 35386
rect 50540 35334 50570 35386
rect 50570 35334 50596 35386
rect 50300 35332 50356 35334
rect 50380 35332 50436 35334
rect 50460 35332 50516 35334
rect 50540 35332 50596 35334
rect 50300 34298 50356 34300
rect 50380 34298 50436 34300
rect 50460 34298 50516 34300
rect 50540 34298 50596 34300
rect 50300 34246 50326 34298
rect 50326 34246 50356 34298
rect 50380 34246 50390 34298
rect 50390 34246 50436 34298
rect 50460 34246 50506 34298
rect 50506 34246 50516 34298
rect 50540 34246 50570 34298
rect 50570 34246 50596 34298
rect 50300 34244 50356 34246
rect 50380 34244 50436 34246
rect 50460 34244 50516 34246
rect 50540 34244 50596 34246
rect 51722 36352 51778 36408
rect 51722 35808 51778 35864
rect 51814 34856 51870 34912
rect 51814 34484 51816 34504
rect 51816 34484 51868 34504
rect 51868 34484 51870 34504
rect 51814 34448 51870 34484
rect 52458 35536 52514 35592
rect 52734 38800 52790 38856
rect 53102 40160 53158 40216
rect 55034 41676 55090 41712
rect 55034 41656 55036 41676
rect 55036 41656 55088 41676
rect 55088 41656 55090 41676
rect 55954 41676 56010 41712
rect 58346 42608 58402 42664
rect 59542 42608 59598 42664
rect 65660 43546 65716 43548
rect 65740 43546 65796 43548
rect 65820 43546 65876 43548
rect 65900 43546 65956 43548
rect 65660 43494 65686 43546
rect 65686 43494 65716 43546
rect 65740 43494 65750 43546
rect 65750 43494 65796 43546
rect 65820 43494 65866 43546
rect 65866 43494 65876 43546
rect 65900 43494 65930 43546
rect 65930 43494 65956 43546
rect 65660 43492 65716 43494
rect 65740 43492 65796 43494
rect 65820 43492 65876 43494
rect 65900 43492 65956 43494
rect 60186 42608 60242 42664
rect 55954 41656 55956 41676
rect 55956 41656 56008 41676
rect 56008 41656 56010 41676
rect 60646 41520 60702 41576
rect 53654 39344 53710 39400
rect 54298 38936 54354 38992
rect 56782 39480 56838 39536
rect 57702 39344 57758 39400
rect 56230 39072 56286 39128
rect 52918 38392 52974 38448
rect 53194 37984 53250 38040
rect 55034 38392 55090 38448
rect 56598 38700 56600 38720
rect 56600 38700 56652 38720
rect 56652 38700 56654 38720
rect 56598 38664 56654 38700
rect 58254 39344 58310 39400
rect 53746 35264 53802 35320
rect 51078 30776 51134 30832
rect 51998 25472 52054 25528
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 52366 22752 52422 22808
rect 23478 4800 23534 4856
rect 52090 4800 52146 4856
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 56230 37204 56232 37224
rect 56232 37204 56284 37224
rect 56284 37204 56286 37224
rect 56230 37168 56286 37204
rect 54114 34720 54170 34776
rect 53838 30164 53894 30220
rect 53838 29452 53840 29472
rect 53840 29452 53892 29472
rect 53892 29452 53894 29472
rect 53838 29416 53894 29452
rect 53838 28124 53894 28180
rect 53838 26696 53894 26752
rect 53838 24216 53840 24236
rect 53840 24216 53892 24236
rect 53892 24216 53894 24236
rect 53838 24180 53894 24216
rect 55218 35672 55274 35728
rect 54850 34720 54906 34776
rect 55954 35808 56010 35864
rect 55770 35400 55826 35456
rect 55770 35264 55826 35320
rect 57426 37576 57482 37632
rect 60646 38972 60648 38992
rect 60648 38972 60700 38992
rect 60700 38972 60702 38992
rect 60646 38936 60702 38972
rect 59542 38800 59598 38856
rect 59910 37868 59966 37904
rect 59910 37848 59912 37868
rect 59912 37848 59964 37868
rect 59964 37848 59966 37868
rect 56782 36760 56838 36816
rect 57886 36760 57942 36816
rect 58162 36352 58218 36408
rect 56966 35808 57022 35864
rect 56322 35672 56378 35728
rect 56598 35400 56654 35456
rect 57978 36080 58034 36136
rect 56966 34892 56968 34912
rect 56968 34892 57020 34912
rect 57020 34892 57022 34912
rect 56966 34856 57022 34892
rect 56506 34448 56562 34504
rect 61106 38548 61162 38584
rect 61106 38528 61108 38548
rect 61108 38528 61160 38548
rect 61160 38528 61162 38548
rect 58162 34448 58218 34504
rect 58622 35264 58678 35320
rect 59082 35572 59084 35592
rect 59084 35572 59136 35592
rect 59136 35572 59138 35592
rect 59082 35536 59138 35572
rect 58898 35436 58900 35456
rect 58900 35436 58952 35456
rect 58952 35436 58954 35456
rect 58898 35400 58954 35436
rect 63774 38528 63830 38584
rect 61290 38392 61346 38448
rect 61934 38256 61990 38312
rect 58898 34484 58900 34504
rect 58900 34484 58952 34504
rect 58952 34484 58954 34504
rect 58898 34448 58954 34484
rect 57518 34348 57520 34368
rect 57520 34348 57572 34368
rect 57572 34348 57574 34368
rect 57518 34312 57574 34348
rect 58990 34312 59046 34368
rect 65660 42458 65716 42460
rect 65740 42458 65796 42460
rect 65820 42458 65876 42460
rect 65900 42458 65956 42460
rect 65660 42406 65686 42458
rect 65686 42406 65716 42458
rect 65740 42406 65750 42458
rect 65750 42406 65796 42458
rect 65820 42406 65866 42458
rect 65866 42406 65876 42458
rect 65900 42406 65930 42458
rect 65930 42406 65956 42458
rect 65660 42404 65716 42406
rect 65740 42404 65796 42406
rect 65820 42404 65876 42406
rect 65900 42404 65956 42406
rect 66350 41556 66352 41576
rect 66352 41556 66404 41576
rect 66404 41556 66406 41576
rect 66350 41520 66406 41556
rect 65660 41370 65716 41372
rect 65740 41370 65796 41372
rect 65820 41370 65876 41372
rect 65900 41370 65956 41372
rect 65660 41318 65686 41370
rect 65686 41318 65716 41370
rect 65740 41318 65750 41370
rect 65750 41318 65796 41370
rect 65820 41318 65866 41370
rect 65866 41318 65876 41370
rect 65900 41318 65930 41370
rect 65930 41318 65956 41370
rect 65660 41316 65716 41318
rect 65740 41316 65796 41318
rect 65820 41316 65876 41318
rect 65900 41316 65956 41318
rect 71226 40976 71282 41032
rect 65660 40282 65716 40284
rect 65740 40282 65796 40284
rect 65820 40282 65876 40284
rect 65900 40282 65956 40284
rect 65660 40230 65686 40282
rect 65686 40230 65716 40282
rect 65740 40230 65750 40282
rect 65750 40230 65796 40282
rect 65820 40230 65866 40282
rect 65866 40230 65876 40282
rect 65900 40230 65930 40282
rect 65930 40230 65956 40282
rect 65660 40228 65716 40230
rect 65740 40228 65796 40230
rect 65820 40228 65876 40230
rect 65900 40228 65956 40230
rect 67270 40452 67326 40488
rect 67270 40432 67272 40452
rect 67272 40432 67324 40452
rect 67324 40432 67326 40452
rect 66258 40024 66314 40080
rect 66994 40024 67050 40080
rect 71042 40024 71098 40080
rect 65660 39194 65716 39196
rect 65740 39194 65796 39196
rect 65820 39194 65876 39196
rect 65900 39194 65956 39196
rect 65660 39142 65686 39194
rect 65686 39142 65716 39194
rect 65740 39142 65750 39194
rect 65750 39142 65796 39194
rect 65820 39142 65866 39194
rect 65866 39142 65876 39194
rect 65900 39142 65930 39194
rect 65930 39142 65956 39194
rect 65660 39140 65716 39142
rect 65740 39140 65796 39142
rect 65820 39140 65876 39142
rect 65900 39140 65956 39142
rect 67546 38956 67602 38992
rect 67546 38936 67548 38956
rect 67548 38936 67600 38956
rect 67600 38936 67602 38956
rect 70214 38956 70270 38992
rect 70214 38936 70216 38956
rect 70216 38936 70268 38956
rect 70268 38936 70270 38956
rect 64234 37612 64236 37632
rect 64236 37612 64288 37632
rect 64288 37612 64290 37632
rect 64234 37576 64290 37612
rect 67362 38276 67418 38312
rect 67362 38256 67364 38276
rect 67364 38256 67416 38276
rect 67416 38256 67418 38276
rect 65660 38106 65716 38108
rect 65740 38106 65796 38108
rect 65820 38106 65876 38108
rect 65900 38106 65956 38108
rect 65660 38054 65686 38106
rect 65686 38054 65716 38106
rect 65740 38054 65750 38106
rect 65750 38054 65796 38106
rect 65820 38054 65866 38106
rect 65866 38054 65876 38106
rect 65900 38054 65930 38106
rect 65930 38054 65956 38106
rect 65660 38052 65716 38054
rect 65740 38052 65796 38054
rect 65820 38052 65876 38054
rect 65900 38052 65956 38054
rect 65522 37304 65578 37360
rect 81020 44090 81076 44092
rect 81100 44090 81156 44092
rect 81180 44090 81236 44092
rect 81260 44090 81316 44092
rect 81020 44038 81046 44090
rect 81046 44038 81076 44090
rect 81100 44038 81110 44090
rect 81110 44038 81156 44090
rect 81180 44038 81226 44090
rect 81226 44038 81236 44090
rect 81260 44038 81290 44090
rect 81290 44038 81316 44090
rect 81020 44036 81076 44038
rect 81100 44036 81156 44038
rect 81180 44036 81236 44038
rect 81260 44036 81316 44038
rect 70122 37712 70178 37768
rect 65660 37018 65716 37020
rect 65740 37018 65796 37020
rect 65820 37018 65876 37020
rect 65900 37018 65956 37020
rect 65660 36966 65686 37018
rect 65686 36966 65716 37018
rect 65740 36966 65750 37018
rect 65750 36966 65796 37018
rect 65820 36966 65866 37018
rect 65866 36966 65876 37018
rect 65900 36966 65930 37018
rect 65930 36966 65956 37018
rect 65660 36964 65716 36966
rect 65740 36964 65796 36966
rect 65820 36964 65876 36966
rect 65900 36964 65956 36966
rect 67454 36080 67510 36136
rect 65660 35930 65716 35932
rect 65740 35930 65796 35932
rect 65820 35930 65876 35932
rect 65900 35930 65956 35932
rect 65660 35878 65686 35930
rect 65686 35878 65716 35930
rect 65740 35878 65750 35930
rect 65750 35878 65796 35930
rect 65820 35878 65866 35930
rect 65866 35878 65876 35930
rect 65900 35878 65930 35930
rect 65930 35878 65956 35930
rect 65660 35876 65716 35878
rect 65740 35876 65796 35878
rect 65820 35876 65876 35878
rect 65900 35876 65956 35878
rect 67638 35808 67694 35864
rect 65660 34842 65716 34844
rect 65740 34842 65796 34844
rect 65820 34842 65876 34844
rect 65900 34842 65956 34844
rect 65660 34790 65686 34842
rect 65686 34790 65716 34842
rect 65740 34790 65750 34842
rect 65750 34790 65796 34842
rect 65820 34790 65866 34842
rect 65866 34790 65876 34842
rect 65900 34790 65930 34842
rect 65930 34790 65956 34842
rect 65660 34788 65716 34790
rect 65740 34788 65796 34790
rect 65820 34788 65876 34790
rect 65900 34788 65956 34790
rect 66166 35264 66222 35320
rect 66994 35400 67050 35456
rect 68650 35400 68706 35456
rect 74814 40976 74870 41032
rect 75826 40452 75882 40488
rect 75826 40432 75828 40452
rect 75828 40432 75880 40452
rect 75880 40432 75882 40452
rect 74722 38956 74778 38992
rect 74722 38936 74724 38956
rect 74724 38936 74776 38956
rect 74776 38936 74778 38956
rect 69938 35536 69994 35592
rect 73066 35828 73122 35864
rect 73066 35808 73068 35828
rect 73068 35808 73120 35828
rect 73120 35808 73122 35828
rect 77206 40024 77262 40080
rect 81020 43002 81076 43004
rect 81100 43002 81156 43004
rect 81180 43002 81236 43004
rect 81260 43002 81316 43004
rect 81020 42950 81046 43002
rect 81046 42950 81076 43002
rect 81100 42950 81110 43002
rect 81110 42950 81156 43002
rect 81180 42950 81226 43002
rect 81226 42950 81236 43002
rect 81260 42950 81290 43002
rect 81290 42950 81316 43002
rect 81020 42948 81076 42950
rect 81100 42948 81156 42950
rect 81180 42948 81236 42950
rect 81260 42948 81316 42950
rect 81020 41914 81076 41916
rect 81100 41914 81156 41916
rect 81180 41914 81236 41916
rect 81260 41914 81316 41916
rect 81020 41862 81046 41914
rect 81046 41862 81076 41914
rect 81100 41862 81110 41914
rect 81110 41862 81156 41914
rect 81180 41862 81226 41914
rect 81226 41862 81236 41914
rect 81260 41862 81290 41914
rect 81290 41862 81316 41914
rect 81020 41860 81076 41862
rect 81100 41860 81156 41862
rect 81180 41860 81236 41862
rect 81260 41860 81316 41862
rect 81020 40826 81076 40828
rect 81100 40826 81156 40828
rect 81180 40826 81236 40828
rect 81260 40826 81316 40828
rect 81020 40774 81046 40826
rect 81046 40774 81076 40826
rect 81100 40774 81110 40826
rect 81110 40774 81156 40826
rect 81180 40774 81226 40826
rect 81226 40774 81236 40826
rect 81260 40774 81290 40826
rect 81290 40774 81316 40826
rect 81020 40772 81076 40774
rect 81100 40772 81156 40774
rect 81180 40772 81236 40774
rect 81260 40772 81316 40774
rect 96380 43546 96436 43548
rect 96460 43546 96516 43548
rect 96540 43546 96596 43548
rect 96620 43546 96676 43548
rect 96380 43494 96406 43546
rect 96406 43494 96436 43546
rect 96460 43494 96470 43546
rect 96470 43494 96516 43546
rect 96540 43494 96586 43546
rect 96586 43494 96596 43546
rect 96620 43494 96650 43546
rect 96650 43494 96676 43546
rect 96380 43492 96436 43494
rect 96460 43492 96516 43494
rect 96540 43492 96596 43494
rect 96620 43492 96676 43494
rect 81020 39738 81076 39740
rect 81100 39738 81156 39740
rect 81180 39738 81236 39740
rect 81260 39738 81316 39740
rect 81020 39686 81046 39738
rect 81046 39686 81076 39738
rect 81100 39686 81110 39738
rect 81110 39686 81156 39738
rect 81180 39686 81226 39738
rect 81226 39686 81236 39738
rect 81260 39686 81290 39738
rect 81290 39686 81316 39738
rect 81020 39684 81076 39686
rect 81100 39684 81156 39686
rect 81180 39684 81236 39686
rect 81260 39684 81316 39686
rect 96380 42458 96436 42460
rect 96460 42458 96516 42460
rect 96540 42458 96596 42460
rect 96620 42458 96676 42460
rect 96380 42406 96406 42458
rect 96406 42406 96436 42458
rect 96460 42406 96470 42458
rect 96470 42406 96516 42458
rect 96540 42406 96586 42458
rect 96586 42406 96596 42458
rect 96620 42406 96650 42458
rect 96650 42406 96676 42458
rect 96380 42404 96436 42406
rect 96460 42404 96516 42406
rect 96540 42404 96596 42406
rect 96620 42404 96676 42406
rect 96380 41370 96436 41372
rect 96460 41370 96516 41372
rect 96540 41370 96596 41372
rect 96620 41370 96676 41372
rect 96380 41318 96406 41370
rect 96406 41318 96436 41370
rect 96460 41318 96470 41370
rect 96470 41318 96516 41370
rect 96540 41318 96586 41370
rect 96586 41318 96596 41370
rect 96620 41318 96650 41370
rect 96650 41318 96676 41370
rect 96380 41316 96436 41318
rect 96460 41316 96516 41318
rect 96540 41316 96596 41318
rect 96620 41316 96676 41318
rect 81020 38650 81076 38652
rect 81100 38650 81156 38652
rect 81180 38650 81236 38652
rect 81260 38650 81316 38652
rect 81020 38598 81046 38650
rect 81046 38598 81076 38650
rect 81100 38598 81110 38650
rect 81110 38598 81156 38650
rect 81180 38598 81226 38650
rect 81226 38598 81236 38650
rect 81260 38598 81290 38650
rect 81290 38598 81316 38650
rect 81020 38596 81076 38598
rect 81100 38596 81156 38598
rect 81180 38596 81236 38598
rect 81260 38596 81316 38598
rect 75366 35148 75422 35184
rect 75366 35128 75368 35148
rect 75368 35128 75420 35148
rect 75420 35128 75422 35148
rect 74262 35028 74264 35048
rect 74264 35028 74316 35048
rect 74316 35028 74318 35048
rect 74262 34992 74318 35028
rect 66350 34448 66406 34504
rect 76194 34856 76250 34912
rect 76654 35400 76710 35456
rect 77390 35808 77446 35864
rect 81020 37562 81076 37564
rect 81100 37562 81156 37564
rect 81180 37562 81236 37564
rect 81260 37562 81316 37564
rect 81020 37510 81046 37562
rect 81046 37510 81076 37562
rect 81100 37510 81110 37562
rect 81110 37510 81156 37562
rect 81180 37510 81226 37562
rect 81226 37510 81236 37562
rect 81260 37510 81290 37562
rect 81290 37510 81316 37562
rect 81020 37508 81076 37510
rect 81100 37508 81156 37510
rect 81180 37508 81236 37510
rect 81260 37508 81316 37510
rect 77850 36216 77906 36272
rect 79230 36236 79286 36272
rect 79230 36216 79232 36236
rect 79232 36216 79284 36236
rect 79284 36216 79286 36236
rect 77574 36080 77630 36136
rect 78310 35536 78366 35592
rect 81020 36474 81076 36476
rect 81100 36474 81156 36476
rect 81180 36474 81236 36476
rect 81260 36474 81316 36476
rect 81020 36422 81046 36474
rect 81046 36422 81076 36474
rect 81100 36422 81110 36474
rect 81110 36422 81156 36474
rect 81180 36422 81226 36474
rect 81226 36422 81236 36474
rect 81260 36422 81290 36474
rect 81290 36422 81316 36474
rect 81020 36420 81076 36422
rect 81100 36420 81156 36422
rect 81180 36420 81236 36422
rect 81260 36420 81316 36422
rect 79782 36080 79838 36136
rect 76746 34856 76802 34912
rect 77298 34992 77354 35048
rect 78034 34892 78036 34912
rect 78036 34892 78088 34912
rect 78088 34892 78090 34912
rect 78034 34856 78090 34892
rect 78494 34720 78550 34776
rect 78586 34584 78642 34640
rect 78494 34468 78550 34504
rect 78494 34448 78496 34468
rect 78496 34448 78548 34468
rect 78548 34448 78550 34468
rect 79506 35128 79562 35184
rect 83186 38972 83188 38992
rect 83188 38972 83240 38992
rect 83240 38972 83242 38992
rect 83186 38936 83242 38972
rect 80150 35536 80206 35592
rect 81020 35386 81076 35388
rect 81100 35386 81156 35388
rect 81180 35386 81236 35388
rect 81260 35386 81316 35388
rect 81020 35334 81046 35386
rect 81046 35334 81076 35386
rect 81100 35334 81110 35386
rect 81110 35334 81156 35386
rect 81180 35334 81226 35386
rect 81226 35334 81236 35386
rect 81260 35334 81290 35386
rect 81290 35334 81316 35386
rect 81020 35332 81076 35334
rect 81100 35332 81156 35334
rect 81180 35332 81236 35334
rect 81260 35332 81316 35334
rect 81438 34740 81494 34776
rect 81438 34720 81440 34740
rect 81440 34720 81492 34740
rect 81492 34720 81494 34740
rect 78954 34604 79010 34640
rect 78954 34584 78956 34604
rect 78956 34584 79008 34604
rect 79008 34584 79010 34604
rect 79966 34448 80022 34504
rect 53838 20100 53894 20156
rect 53838 14796 53894 14852
rect 81020 34298 81076 34300
rect 81100 34298 81156 34300
rect 81180 34298 81236 34300
rect 81260 34298 81316 34300
rect 81020 34246 81046 34298
rect 81046 34246 81076 34298
rect 81100 34246 81110 34298
rect 81110 34246 81156 34298
rect 81180 34246 81226 34298
rect 81226 34246 81236 34298
rect 81260 34246 81290 34298
rect 81290 34246 81316 34298
rect 81020 34244 81076 34246
rect 81100 34244 81156 34246
rect 81180 34244 81236 34246
rect 81260 34244 81316 34246
rect 81438 31592 81494 31648
rect 81530 30164 81586 30220
rect 81438 29484 81494 29540
rect 81622 28124 81678 28180
rect 81622 26764 81678 26820
rect 81990 34468 82046 34504
rect 81990 34448 81992 34468
rect 81992 34448 82044 34468
rect 82044 34448 82046 34468
rect 81622 25540 81678 25596
rect 81346 24180 81402 24236
rect 81622 22856 81624 22876
rect 81624 22856 81676 22876
rect 81676 22856 81678 22876
rect 81622 22820 81678 22856
rect 83370 38664 83426 38720
rect 84106 38956 84162 38992
rect 84106 38936 84108 38956
rect 84108 38936 84160 38956
rect 84160 38936 84162 38956
rect 84014 38664 84070 38720
rect 86866 39888 86922 39944
rect 96380 40282 96436 40284
rect 96460 40282 96516 40284
rect 96540 40282 96596 40284
rect 96620 40282 96676 40284
rect 96380 40230 96406 40282
rect 96406 40230 96436 40282
rect 96460 40230 96470 40282
rect 96470 40230 96516 40282
rect 96540 40230 96586 40282
rect 96586 40230 96596 40282
rect 96620 40230 96650 40282
rect 96650 40230 96676 40282
rect 96380 40228 96436 40230
rect 96460 40228 96516 40230
rect 96540 40228 96596 40230
rect 96620 40228 96676 40230
rect 96380 39194 96436 39196
rect 96460 39194 96516 39196
rect 96540 39194 96596 39196
rect 96620 39194 96676 39196
rect 96380 39142 96406 39194
rect 96406 39142 96436 39194
rect 96460 39142 96470 39194
rect 96470 39142 96516 39194
rect 96540 39142 96586 39194
rect 96586 39142 96596 39194
rect 96620 39142 96650 39194
rect 96650 39142 96676 39194
rect 96380 39140 96436 39142
rect 96460 39140 96516 39142
rect 96540 39140 96596 39142
rect 96620 39140 96676 39142
rect 85854 35808 85910 35864
rect 85486 35672 85542 35728
rect 83554 35128 83610 35184
rect 84382 34992 84438 35048
rect 84750 34992 84806 35048
rect 85578 34992 85634 35048
rect 86038 34992 86094 35048
rect 96380 38106 96436 38108
rect 96460 38106 96516 38108
rect 96540 38106 96596 38108
rect 96620 38106 96676 38108
rect 96380 38054 96406 38106
rect 96406 38054 96436 38106
rect 96460 38054 96470 38106
rect 96470 38054 96516 38106
rect 96540 38054 96586 38106
rect 96586 38054 96596 38106
rect 96620 38054 96650 38106
rect 96650 38054 96676 38106
rect 96380 38052 96436 38054
rect 96460 38052 96516 38054
rect 96540 38052 96596 38054
rect 96620 38052 96676 38054
rect 91006 36760 91062 36816
rect 96380 37018 96436 37020
rect 96460 37018 96516 37020
rect 96540 37018 96596 37020
rect 96620 37018 96676 37020
rect 96380 36966 96406 37018
rect 96406 36966 96436 37018
rect 96460 36966 96470 37018
rect 96470 36966 96516 37018
rect 96540 36966 96586 37018
rect 96586 36966 96596 37018
rect 96620 36966 96650 37018
rect 96650 36966 96676 37018
rect 96380 36964 96436 36966
rect 96460 36964 96516 36966
rect 96540 36964 96596 36966
rect 96620 36964 96676 36966
rect 95330 36760 95386 36816
rect 96380 35930 96436 35932
rect 96460 35930 96516 35932
rect 96540 35930 96596 35932
rect 96620 35930 96676 35932
rect 96380 35878 96406 35930
rect 96406 35878 96436 35930
rect 96460 35878 96470 35930
rect 96470 35878 96516 35930
rect 96540 35878 96586 35930
rect 96586 35878 96596 35930
rect 96620 35878 96650 35930
rect 96650 35878 96676 35930
rect 96380 35876 96436 35878
rect 96460 35876 96516 35878
rect 96540 35876 96596 35878
rect 96620 35876 96676 35878
rect 96380 34842 96436 34844
rect 96460 34842 96516 34844
rect 96540 34842 96596 34844
rect 96620 34842 96676 34844
rect 96380 34790 96406 34842
rect 96406 34790 96436 34842
rect 96460 34790 96470 34842
rect 96470 34790 96516 34842
rect 96540 34790 96586 34842
rect 96586 34790 96596 34842
rect 96620 34790 96650 34842
rect 96650 34790 96676 34842
rect 96380 34788 96436 34790
rect 96460 34788 96516 34790
rect 96540 34788 96596 34790
rect 96620 34788 96676 34790
rect 82358 31592 82414 31648
rect 80886 20032 80942 20088
rect 81622 15952 81678 16008
rect 81622 14796 81678 14852
rect 79966 4800 80022 4856
rect 2778 312 2834 368
<< metal3 >>
rect 0 45930 800 45960
rect 3601 45930 3667 45933
rect 0 45928 3667 45930
rect 0 45872 3606 45928
rect 3662 45872 3667 45928
rect 0 45870 3667 45872
rect 0 45840 800 45870
rect 3601 45867 3667 45870
rect 0 45386 800 45416
rect 4061 45386 4127 45389
rect 0 45384 4127 45386
rect 0 45328 4066 45384
rect 4122 45328 4127 45384
rect 0 45326 4127 45328
rect 0 45296 800 45326
rect 4061 45323 4127 45326
rect 0 44706 800 44736
rect 2773 44706 2839 44709
rect 0 44704 2839 44706
rect 0 44648 2778 44704
rect 2834 44648 2839 44704
rect 0 44646 2839 44648
rect 0 44616 800 44646
rect 2773 44643 2839 44646
rect 0 44162 800 44192
rect 3509 44162 3575 44165
rect 0 44160 3575 44162
rect 0 44104 3514 44160
rect 3570 44104 3575 44160
rect 0 44102 3575 44104
rect 0 44072 800 44102
rect 3509 44099 3575 44102
rect 19568 44096 19888 44097
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 44031 19888 44032
rect 50288 44096 50608 44097
rect 50288 44032 50296 44096
rect 50360 44032 50376 44096
rect 50440 44032 50456 44096
rect 50520 44032 50536 44096
rect 50600 44032 50608 44096
rect 50288 44031 50608 44032
rect 81008 44096 81328 44097
rect 81008 44032 81016 44096
rect 81080 44032 81096 44096
rect 81160 44032 81176 44096
rect 81240 44032 81256 44096
rect 81320 44032 81328 44096
rect 81008 44031 81328 44032
rect 0 43528 800 43648
rect 4208 43552 4528 43553
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 43487 4528 43488
rect 34928 43552 35248 43553
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 43487 35248 43488
rect 65648 43552 65968 43553
rect 65648 43488 65656 43552
rect 65720 43488 65736 43552
rect 65800 43488 65816 43552
rect 65880 43488 65896 43552
rect 65960 43488 65968 43552
rect 65648 43487 65968 43488
rect 96368 43552 96688 43553
rect 96368 43488 96376 43552
rect 96440 43488 96456 43552
rect 96520 43488 96536 43552
rect 96600 43488 96616 43552
rect 96680 43488 96688 43552
rect 96368 43487 96688 43488
rect 19568 43008 19888 43009
rect 0 42848 800 42968
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 42943 19888 42944
rect 50288 43008 50608 43009
rect 50288 42944 50296 43008
rect 50360 42944 50376 43008
rect 50440 42944 50456 43008
rect 50520 42944 50536 43008
rect 50600 42944 50608 43008
rect 50288 42943 50608 42944
rect 81008 43008 81328 43009
rect 81008 42944 81016 43008
rect 81080 42944 81096 43008
rect 81160 42944 81176 43008
rect 81240 42944 81256 43008
rect 81320 42944 81328 43008
rect 81008 42943 81328 42944
rect 29361 42802 29427 42805
rect 38193 42802 38259 42805
rect 29361 42800 38259 42802
rect 29361 42744 29366 42800
rect 29422 42744 38198 42800
rect 38254 42744 38259 42800
rect 29361 42742 38259 42744
rect 29361 42739 29427 42742
rect 38193 42739 38259 42742
rect 34973 42666 35039 42669
rect 37733 42666 37799 42669
rect 40953 42666 41019 42669
rect 34973 42664 41019 42666
rect 34973 42608 34978 42664
rect 35034 42608 37738 42664
rect 37794 42608 40958 42664
rect 41014 42608 41019 42664
rect 34973 42606 41019 42608
rect 34973 42603 35039 42606
rect 37733 42603 37799 42606
rect 40953 42603 41019 42606
rect 58341 42666 58407 42669
rect 59537 42666 59603 42669
rect 60181 42666 60247 42669
rect 58341 42664 60247 42666
rect 58341 42608 58346 42664
rect 58402 42608 59542 42664
rect 59598 42608 60186 42664
rect 60242 42608 60247 42664
rect 58341 42606 60247 42608
rect 58341 42603 58407 42606
rect 59537 42603 59603 42606
rect 60181 42603 60247 42606
rect 4208 42464 4528 42465
rect 0 42304 800 42424
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 42399 4528 42400
rect 34928 42464 35248 42465
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 42399 35248 42400
rect 65648 42464 65968 42465
rect 65648 42400 65656 42464
rect 65720 42400 65736 42464
rect 65800 42400 65816 42464
rect 65880 42400 65896 42464
rect 65960 42400 65968 42464
rect 65648 42399 65968 42400
rect 96368 42464 96688 42465
rect 96368 42400 96376 42464
rect 96440 42400 96456 42464
rect 96520 42400 96536 42464
rect 96600 42400 96616 42464
rect 96680 42400 96688 42464
rect 96368 42399 96688 42400
rect 21817 42258 21883 42261
rect 28165 42258 28231 42261
rect 21817 42256 28231 42258
rect 21817 42200 21822 42256
rect 21878 42200 28170 42256
rect 28226 42200 28231 42256
rect 21817 42198 28231 42200
rect 21817 42195 21883 42198
rect 28165 42195 28231 42198
rect 37089 42258 37155 42261
rect 39113 42258 39179 42261
rect 37089 42256 39179 42258
rect 37089 42200 37094 42256
rect 37150 42200 39118 42256
rect 39174 42200 39179 42256
rect 37089 42198 39179 42200
rect 37089 42195 37155 42198
rect 39113 42195 39179 42198
rect 48313 42122 48379 42125
rect 49509 42122 49575 42125
rect 48313 42120 49575 42122
rect 48313 42064 48318 42120
rect 48374 42064 49514 42120
rect 49570 42064 49575 42120
rect 48313 42062 49575 42064
rect 48313 42059 48379 42062
rect 49509 42059 49575 42062
rect 19568 41920 19888 41921
rect 0 41760 800 41880
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 41855 19888 41856
rect 50288 41920 50608 41921
rect 50288 41856 50296 41920
rect 50360 41856 50376 41920
rect 50440 41856 50456 41920
rect 50520 41856 50536 41920
rect 50600 41856 50608 41920
rect 50288 41855 50608 41856
rect 81008 41920 81328 41921
rect 81008 41856 81016 41920
rect 81080 41856 81096 41920
rect 81160 41856 81176 41920
rect 81240 41856 81256 41920
rect 81320 41856 81328 41920
rect 81008 41855 81328 41856
rect 48589 41714 48655 41717
rect 49877 41714 49943 41717
rect 48589 41712 49943 41714
rect 48589 41656 48594 41712
rect 48650 41656 49882 41712
rect 49938 41656 49943 41712
rect 48589 41654 49943 41656
rect 48589 41651 48655 41654
rect 49877 41651 49943 41654
rect 55029 41714 55095 41717
rect 55949 41714 56015 41717
rect 55029 41712 56015 41714
rect 55029 41656 55034 41712
rect 55090 41656 55954 41712
rect 56010 41656 56015 41712
rect 55029 41654 56015 41656
rect 55029 41651 55095 41654
rect 55949 41651 56015 41654
rect 32397 41578 32463 41581
rect 33685 41578 33751 41581
rect 39113 41578 39179 41581
rect 32397 41576 39179 41578
rect 32397 41520 32402 41576
rect 32458 41520 33690 41576
rect 33746 41520 39118 41576
rect 39174 41520 39179 41576
rect 32397 41518 39179 41520
rect 32397 41515 32463 41518
rect 33685 41515 33751 41518
rect 39113 41515 39179 41518
rect 60641 41578 60707 41581
rect 66345 41578 66411 41581
rect 60641 41576 66411 41578
rect 60641 41520 60646 41576
rect 60702 41520 66350 41576
rect 66406 41520 66411 41576
rect 60641 41518 66411 41520
rect 60641 41515 60707 41518
rect 66345 41515 66411 41518
rect 38929 41442 38995 41445
rect 43437 41442 43503 41445
rect 38929 41440 43503 41442
rect 38929 41384 38934 41440
rect 38990 41384 43442 41440
rect 43498 41384 43503 41440
rect 38929 41382 43503 41384
rect 38929 41379 38995 41382
rect 43437 41379 43503 41382
rect 4208 41376 4528 41377
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 41311 4528 41312
rect 34928 41376 35248 41377
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 41311 35248 41312
rect 65648 41376 65968 41377
rect 65648 41312 65656 41376
rect 65720 41312 65736 41376
rect 65800 41312 65816 41376
rect 65880 41312 65896 41376
rect 65960 41312 65968 41376
rect 65648 41311 65968 41312
rect 96368 41376 96688 41377
rect 96368 41312 96376 41376
rect 96440 41312 96456 41376
rect 96520 41312 96536 41376
rect 96600 41312 96616 41376
rect 96680 41312 96688 41376
rect 96368 41311 96688 41312
rect 0 41170 800 41200
rect 3877 41170 3943 41173
rect 0 41168 3943 41170
rect 0 41112 3882 41168
rect 3938 41112 3943 41168
rect 0 41110 3943 41112
rect 0 41080 800 41110
rect 3877 41107 3943 41110
rect 32489 41034 32555 41037
rect 33317 41034 33383 41037
rect 32489 41032 33383 41034
rect 32489 40976 32494 41032
rect 32550 40976 33322 41032
rect 33378 40976 33383 41032
rect 32489 40974 33383 40976
rect 32489 40971 32555 40974
rect 33317 40971 33383 40974
rect 71221 41034 71287 41037
rect 74809 41034 74875 41037
rect 71221 41032 74875 41034
rect 71221 40976 71226 41032
rect 71282 40976 74814 41032
rect 74870 40976 74875 41032
rect 71221 40974 74875 40976
rect 71221 40971 71287 40974
rect 74809 40971 74875 40974
rect 19568 40832 19888 40833
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 40767 19888 40768
rect 50288 40832 50608 40833
rect 50288 40768 50296 40832
rect 50360 40768 50376 40832
rect 50440 40768 50456 40832
rect 50520 40768 50536 40832
rect 50600 40768 50608 40832
rect 50288 40767 50608 40768
rect 81008 40832 81328 40833
rect 81008 40768 81016 40832
rect 81080 40768 81096 40832
rect 81160 40768 81176 40832
rect 81240 40768 81256 40832
rect 81320 40768 81328 40832
rect 81008 40767 81328 40768
rect 0 40626 800 40656
rect 1485 40626 1551 40629
rect 0 40624 1551 40626
rect 0 40568 1490 40624
rect 1546 40568 1551 40624
rect 0 40566 1551 40568
rect 0 40536 800 40566
rect 1485 40563 1551 40566
rect 28993 40490 29059 40493
rect 31661 40490 31727 40493
rect 32765 40490 32831 40493
rect 28993 40488 32831 40490
rect 28993 40432 28998 40488
rect 29054 40432 31666 40488
rect 31722 40432 32770 40488
rect 32826 40432 32831 40488
rect 28993 40430 32831 40432
rect 28993 40427 29059 40430
rect 31661 40427 31727 40430
rect 32765 40427 32831 40430
rect 67265 40490 67331 40493
rect 75821 40490 75887 40493
rect 67265 40488 75887 40490
rect 67265 40432 67270 40488
rect 67326 40432 75826 40488
rect 75882 40432 75887 40488
rect 67265 40430 75887 40432
rect 67265 40427 67331 40430
rect 75821 40427 75887 40430
rect 39297 40354 39363 40357
rect 48221 40354 48287 40357
rect 39297 40352 48287 40354
rect 39297 40296 39302 40352
rect 39358 40296 48226 40352
rect 48282 40296 48287 40352
rect 39297 40294 48287 40296
rect 39297 40291 39363 40294
rect 48221 40291 48287 40294
rect 49141 40354 49207 40357
rect 49785 40354 49851 40357
rect 49141 40352 49851 40354
rect 49141 40296 49146 40352
rect 49202 40296 49790 40352
rect 49846 40296 49851 40352
rect 49141 40294 49851 40296
rect 49141 40291 49207 40294
rect 49785 40291 49851 40294
rect 4208 40288 4528 40289
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 40223 4528 40224
rect 34928 40288 35248 40289
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 40223 35248 40224
rect 65648 40288 65968 40289
rect 65648 40224 65656 40288
rect 65720 40224 65736 40288
rect 65800 40224 65816 40288
rect 65880 40224 65896 40288
rect 65960 40224 65968 40288
rect 65648 40223 65968 40224
rect 96368 40288 96688 40289
rect 96368 40224 96376 40288
rect 96440 40224 96456 40288
rect 96520 40224 96536 40288
rect 96600 40224 96616 40288
rect 96680 40224 96688 40288
rect 96368 40223 96688 40224
rect 49233 40218 49299 40221
rect 53097 40218 53163 40221
rect 49233 40216 53163 40218
rect 49233 40160 49238 40216
rect 49294 40160 53102 40216
rect 53158 40160 53163 40216
rect 49233 40158 53163 40160
rect 49233 40155 49299 40158
rect 53097 40155 53163 40158
rect 0 40082 800 40112
rect 3325 40082 3391 40085
rect 0 40080 3391 40082
rect 0 40024 3330 40080
rect 3386 40024 3391 40080
rect 0 40022 3391 40024
rect 0 39992 800 40022
rect 3325 40019 3391 40022
rect 49049 40082 49115 40085
rect 51073 40082 51139 40085
rect 49049 40080 51139 40082
rect 49049 40024 49054 40080
rect 49110 40024 51078 40080
rect 51134 40024 51139 40080
rect 49049 40022 51139 40024
rect 49049 40019 49115 40022
rect 51073 40019 51139 40022
rect 66253 40082 66319 40085
rect 66989 40082 67055 40085
rect 66253 40080 67055 40082
rect 66253 40024 66258 40080
rect 66314 40024 66994 40080
rect 67050 40024 67055 40080
rect 66253 40022 67055 40024
rect 66253 40019 66319 40022
rect 66989 40019 67055 40022
rect 71037 40082 71103 40085
rect 77201 40082 77267 40085
rect 71037 40080 77267 40082
rect 71037 40024 71042 40080
rect 71098 40024 77206 40080
rect 77262 40024 77267 40080
rect 71037 40022 77267 40024
rect 71037 40019 71103 40022
rect 77201 40019 77267 40022
rect 31569 39946 31635 39949
rect 32397 39946 32463 39949
rect 31569 39944 32463 39946
rect 31569 39888 31574 39944
rect 31630 39888 32402 39944
rect 32458 39888 32463 39944
rect 31569 39886 32463 39888
rect 31569 39883 31635 39886
rect 32397 39883 32463 39886
rect 32673 39946 32739 39949
rect 34421 39946 34487 39949
rect 32673 39944 34487 39946
rect 32673 39888 32678 39944
rect 32734 39888 34426 39944
rect 34482 39888 34487 39944
rect 32673 39886 34487 39888
rect 32673 39883 32739 39886
rect 34421 39883 34487 39886
rect 45093 39946 45159 39949
rect 86861 39946 86927 39949
rect 45093 39944 86927 39946
rect 45093 39888 45098 39944
rect 45154 39888 86866 39944
rect 86922 39888 86927 39944
rect 45093 39886 86927 39888
rect 45093 39883 45159 39886
rect 86861 39883 86927 39886
rect 33041 39810 33107 39813
rect 38561 39810 38627 39813
rect 33041 39808 38627 39810
rect 33041 39752 33046 39808
rect 33102 39752 38566 39808
rect 38622 39752 38627 39808
rect 33041 39750 38627 39752
rect 33041 39747 33107 39750
rect 38561 39747 38627 39750
rect 51533 39810 51599 39813
rect 52821 39810 52887 39813
rect 51533 39808 52887 39810
rect 51533 39752 51538 39808
rect 51594 39752 52826 39808
rect 52882 39752 52887 39808
rect 51533 39750 52887 39752
rect 51533 39747 51599 39750
rect 52821 39747 52887 39750
rect 19568 39744 19888 39745
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 39679 19888 39680
rect 50288 39744 50608 39745
rect 50288 39680 50296 39744
rect 50360 39680 50376 39744
rect 50440 39680 50456 39744
rect 50520 39680 50536 39744
rect 50600 39680 50608 39744
rect 50288 39679 50608 39680
rect 81008 39744 81328 39745
rect 81008 39680 81016 39744
rect 81080 39680 81096 39744
rect 81160 39680 81176 39744
rect 81240 39680 81256 39744
rect 81320 39680 81328 39744
rect 81008 39679 81328 39680
rect 28942 39612 28948 39676
rect 29012 39674 29018 39676
rect 38561 39674 38627 39677
rect 29012 39672 38627 39674
rect 29012 39616 38566 39672
rect 38622 39616 38627 39672
rect 29012 39614 38627 39616
rect 29012 39612 29018 39614
rect 38561 39611 38627 39614
rect 49325 39674 49391 39677
rect 50153 39674 50219 39677
rect 49325 39672 50219 39674
rect 49325 39616 49330 39672
rect 49386 39616 50158 39672
rect 50214 39616 50219 39672
rect 49325 39614 50219 39616
rect 49325 39611 49391 39614
rect 50153 39611 50219 39614
rect 50705 39674 50771 39677
rect 52637 39674 52703 39677
rect 50705 39672 52703 39674
rect 50705 39616 50710 39672
rect 50766 39616 52642 39672
rect 52698 39616 52703 39672
rect 50705 39614 52703 39616
rect 50705 39611 50771 39614
rect 52637 39611 52703 39614
rect 7833 39538 7899 39541
rect 8293 39538 8359 39541
rect 7833 39536 8359 39538
rect 7833 39480 7838 39536
rect 7894 39480 8298 39536
rect 8354 39480 8359 39536
rect 7833 39478 8359 39480
rect 7833 39475 7899 39478
rect 8293 39475 8359 39478
rect 14273 39538 14339 39541
rect 56777 39538 56843 39541
rect 14273 39536 56843 39538
rect 14273 39480 14278 39536
rect 14334 39480 56782 39536
rect 56838 39480 56843 39536
rect 14273 39478 56843 39480
rect 14273 39475 14339 39478
rect 56777 39475 56843 39478
rect 0 39402 800 39432
rect 3969 39402 4035 39405
rect 0 39400 4035 39402
rect 0 39344 3974 39400
rect 4030 39344 4035 39400
rect 0 39342 4035 39344
rect 0 39312 800 39342
rect 3969 39339 4035 39342
rect 7373 39402 7439 39405
rect 7741 39402 7807 39405
rect 28942 39402 28948 39404
rect 7373 39400 7807 39402
rect 7373 39344 7378 39400
rect 7434 39344 7746 39400
rect 7802 39344 7807 39400
rect 7373 39342 7807 39344
rect 7373 39339 7439 39342
rect 7741 39339 7807 39342
rect 21406 39342 28948 39402
rect 14457 39266 14523 39269
rect 19057 39266 19123 39269
rect 14457 39264 19123 39266
rect 14457 39208 14462 39264
rect 14518 39208 19062 39264
rect 19118 39208 19123 39264
rect 14457 39206 19123 39208
rect 14457 39203 14523 39206
rect 19057 39203 19123 39206
rect 19241 39266 19307 39269
rect 21406 39266 21466 39342
rect 28942 39340 28948 39342
rect 29012 39340 29018 39404
rect 38561 39402 38627 39405
rect 48957 39402 49023 39405
rect 50797 39402 50863 39405
rect 38561 39400 48882 39402
rect 38561 39344 38566 39400
rect 38622 39344 48882 39400
rect 38561 39342 48882 39344
rect 38561 39339 38627 39342
rect 19241 39264 21466 39266
rect 19241 39208 19246 39264
rect 19302 39208 21466 39264
rect 19241 39206 21466 39208
rect 21633 39266 21699 39269
rect 28073 39266 28139 39269
rect 21633 39264 28139 39266
rect 21633 39208 21638 39264
rect 21694 39208 28078 39264
rect 28134 39208 28139 39264
rect 21633 39206 28139 39208
rect 48822 39266 48882 39342
rect 48957 39400 50863 39402
rect 48957 39344 48962 39400
rect 49018 39344 50802 39400
rect 50858 39344 50863 39400
rect 48957 39342 50863 39344
rect 48957 39339 49023 39342
rect 50797 39339 50863 39342
rect 51625 39402 51691 39405
rect 53649 39402 53715 39405
rect 57697 39402 57763 39405
rect 58249 39402 58315 39405
rect 51625 39400 53715 39402
rect 51625 39344 51630 39400
rect 51686 39344 53654 39400
rect 53710 39344 53715 39400
rect 51625 39342 53715 39344
rect 51625 39339 51691 39342
rect 53649 39339 53715 39342
rect 54710 39400 58315 39402
rect 54710 39344 57702 39400
rect 57758 39344 58254 39400
rect 58310 39344 58315 39400
rect 54710 39342 58315 39344
rect 54710 39266 54770 39342
rect 57697 39339 57763 39342
rect 58249 39339 58315 39342
rect 48822 39206 54770 39266
rect 19241 39203 19307 39206
rect 21633 39203 21699 39206
rect 28073 39203 28139 39206
rect 4208 39200 4528 39201
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 39135 4528 39136
rect 34928 39200 35248 39201
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 39135 35248 39136
rect 65648 39200 65968 39201
rect 65648 39136 65656 39200
rect 65720 39136 65736 39200
rect 65800 39136 65816 39200
rect 65880 39136 65896 39200
rect 65960 39136 65968 39200
rect 65648 39135 65968 39136
rect 96368 39200 96688 39201
rect 96368 39136 96376 39200
rect 96440 39136 96456 39200
rect 96520 39136 96536 39200
rect 96600 39136 96616 39200
rect 96680 39136 96688 39200
rect 96368 39135 96688 39136
rect 38653 39130 38719 39133
rect 48221 39130 48287 39133
rect 38653 39128 48287 39130
rect 38653 39072 38658 39128
rect 38714 39072 48226 39128
rect 48282 39072 48287 39128
rect 38653 39070 48287 39072
rect 38653 39067 38719 39070
rect 48221 39067 48287 39070
rect 48957 39130 49023 39133
rect 50061 39130 50127 39133
rect 48957 39128 50127 39130
rect 48957 39072 48962 39128
rect 49018 39072 50066 39128
rect 50122 39072 50127 39128
rect 48957 39070 50127 39072
rect 48957 39067 49023 39070
rect 50061 39067 50127 39070
rect 52361 39130 52427 39133
rect 56225 39130 56291 39133
rect 52361 39128 56291 39130
rect 52361 39072 52366 39128
rect 52422 39072 56230 39128
rect 56286 39072 56291 39128
rect 52361 39070 56291 39072
rect 52361 39067 52427 39070
rect 56225 39067 56291 39070
rect 14089 38994 14155 38997
rect 54293 38994 54359 38997
rect 14089 38992 54359 38994
rect 14089 38936 14094 38992
rect 14150 38936 54298 38992
rect 54354 38936 54359 38992
rect 14089 38934 54359 38936
rect 14089 38931 14155 38934
rect 54293 38931 54359 38934
rect 60641 38994 60707 38997
rect 67541 38994 67607 38997
rect 60641 38992 67607 38994
rect 60641 38936 60646 38992
rect 60702 38936 67546 38992
rect 67602 38936 67607 38992
rect 60641 38934 67607 38936
rect 60641 38931 60707 38934
rect 67541 38931 67607 38934
rect 70209 38994 70275 38997
rect 74717 38994 74783 38997
rect 70209 38992 74783 38994
rect 70209 38936 70214 38992
rect 70270 38936 74722 38992
rect 74778 38936 74783 38992
rect 70209 38934 74783 38936
rect 70209 38931 70275 38934
rect 74717 38931 74783 38934
rect 83181 38994 83247 38997
rect 84101 38994 84167 38997
rect 83181 38992 84167 38994
rect 83181 38936 83186 38992
rect 83242 38936 84106 38992
rect 84162 38936 84167 38992
rect 83181 38934 84167 38936
rect 83181 38931 83247 38934
rect 84101 38931 84167 38934
rect 0 38858 800 38888
rect 3233 38858 3299 38861
rect 0 38856 3299 38858
rect 0 38800 3238 38856
rect 3294 38800 3299 38856
rect 0 38798 3299 38800
rect 0 38768 800 38798
rect 3233 38795 3299 38798
rect 44265 38858 44331 38861
rect 52729 38858 52795 38861
rect 59537 38858 59603 38861
rect 44265 38856 59603 38858
rect 44265 38800 44270 38856
rect 44326 38800 52734 38856
rect 52790 38800 59542 38856
rect 59598 38800 59603 38856
rect 44265 38798 59603 38800
rect 44265 38795 44331 38798
rect 52729 38795 52795 38798
rect 59537 38795 59603 38798
rect 51901 38722 51967 38725
rect 56593 38722 56659 38725
rect 51901 38720 56659 38722
rect 51901 38664 51906 38720
rect 51962 38664 56598 38720
rect 56654 38664 56659 38720
rect 51901 38662 56659 38664
rect 51901 38659 51967 38662
rect 56593 38659 56659 38662
rect 83365 38722 83431 38725
rect 84009 38722 84075 38725
rect 83365 38720 84075 38722
rect 83365 38664 83370 38720
rect 83426 38664 84014 38720
rect 84070 38664 84075 38720
rect 83365 38662 84075 38664
rect 83365 38659 83431 38662
rect 84009 38659 84075 38662
rect 19568 38656 19888 38657
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 38591 19888 38592
rect 50288 38656 50608 38657
rect 50288 38592 50296 38656
rect 50360 38592 50376 38656
rect 50440 38592 50456 38656
rect 50520 38592 50536 38656
rect 50600 38592 50608 38656
rect 50288 38591 50608 38592
rect 81008 38656 81328 38657
rect 81008 38592 81016 38656
rect 81080 38592 81096 38656
rect 81160 38592 81176 38656
rect 81240 38592 81256 38656
rect 81320 38592 81328 38656
rect 81008 38591 81328 38592
rect 42977 38586 43043 38589
rect 48221 38586 48287 38589
rect 42977 38584 48287 38586
rect 42977 38528 42982 38584
rect 43038 38528 48226 38584
rect 48282 38528 48287 38584
rect 42977 38526 48287 38528
rect 42977 38523 43043 38526
rect 48221 38523 48287 38526
rect 61101 38586 61167 38589
rect 63769 38586 63835 38589
rect 61101 38584 63835 38586
rect 61101 38528 61106 38584
rect 61162 38528 63774 38584
rect 63830 38528 63835 38584
rect 61101 38526 63835 38528
rect 61101 38523 61167 38526
rect 63769 38523 63835 38526
rect 19425 38450 19491 38453
rect 19382 38448 19491 38450
rect 19382 38392 19430 38448
rect 19486 38392 19491 38448
rect 19382 38387 19491 38392
rect 50337 38450 50403 38453
rect 51809 38450 51875 38453
rect 52913 38450 52979 38453
rect 50337 38448 52979 38450
rect 50337 38392 50342 38448
rect 50398 38392 51814 38448
rect 51870 38392 52918 38448
rect 52974 38392 52979 38448
rect 50337 38390 52979 38392
rect 50337 38387 50403 38390
rect 51809 38387 51875 38390
rect 52913 38387 52979 38390
rect 55029 38450 55095 38453
rect 61285 38450 61351 38453
rect 55029 38448 61351 38450
rect 55029 38392 55034 38448
rect 55090 38392 61290 38448
rect 61346 38392 61351 38448
rect 55029 38390 61351 38392
rect 55029 38387 55095 38390
rect 61285 38387 61351 38390
rect 19382 38317 19442 38387
rect 19382 38312 19491 38317
rect 19382 38256 19430 38312
rect 19486 38256 19491 38312
rect 19382 38254 19491 38256
rect 19425 38251 19491 38254
rect 39941 38314 40007 38317
rect 40493 38314 40559 38317
rect 39941 38312 40559 38314
rect 39941 38256 39946 38312
rect 40002 38256 40498 38312
rect 40554 38256 40559 38312
rect 39941 38254 40559 38256
rect 39941 38251 40007 38254
rect 40493 38251 40559 38254
rect 50061 38314 50127 38317
rect 51257 38314 51323 38317
rect 50061 38312 51323 38314
rect 50061 38256 50066 38312
rect 50122 38256 51262 38312
rect 51318 38256 51323 38312
rect 50061 38254 51323 38256
rect 50061 38251 50127 38254
rect 51257 38251 51323 38254
rect 61929 38314 61995 38317
rect 67357 38314 67423 38317
rect 61929 38312 67423 38314
rect 61929 38256 61934 38312
rect 61990 38256 67362 38312
rect 67418 38256 67423 38312
rect 61929 38254 67423 38256
rect 61929 38251 61995 38254
rect 67357 38251 67423 38254
rect 0 38178 800 38208
rect 4061 38178 4127 38181
rect 0 38176 4127 38178
rect 0 38120 4066 38176
rect 4122 38120 4127 38176
rect 0 38118 4127 38120
rect 0 38088 800 38118
rect 4061 38115 4127 38118
rect 4208 38112 4528 38113
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 38047 4528 38048
rect 34928 38112 35248 38113
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 38047 35248 38048
rect 65648 38112 65968 38113
rect 65648 38048 65656 38112
rect 65720 38048 65736 38112
rect 65800 38048 65816 38112
rect 65880 38048 65896 38112
rect 65960 38048 65968 38112
rect 65648 38047 65968 38048
rect 96368 38112 96688 38113
rect 96368 38048 96376 38112
rect 96440 38048 96456 38112
rect 96520 38048 96536 38112
rect 96600 38048 96616 38112
rect 96680 38048 96688 38112
rect 96368 38047 96688 38048
rect 50705 38042 50771 38045
rect 53189 38042 53255 38045
rect 50705 38040 53255 38042
rect 50705 37984 50710 38040
rect 50766 37984 53194 38040
rect 53250 37984 53255 38040
rect 50705 37982 53255 37984
rect 50705 37979 50771 37982
rect 53189 37979 53255 37982
rect 21173 37906 21239 37909
rect 22185 37906 22251 37909
rect 21173 37904 22251 37906
rect 21173 37848 21178 37904
rect 21234 37848 22190 37904
rect 22246 37848 22251 37904
rect 21173 37846 22251 37848
rect 21173 37843 21239 37846
rect 22185 37843 22251 37846
rect 41229 37906 41295 37909
rect 59905 37906 59971 37909
rect 41229 37904 59971 37906
rect 41229 37848 41234 37904
rect 41290 37848 59910 37904
rect 59966 37848 59971 37904
rect 41229 37846 59971 37848
rect 41229 37843 41295 37846
rect 59905 37843 59971 37846
rect 11789 37770 11855 37773
rect 15469 37770 15535 37773
rect 18137 37770 18203 37773
rect 11789 37768 18203 37770
rect 11789 37712 11794 37768
rect 11850 37712 15474 37768
rect 15530 37712 18142 37768
rect 18198 37712 18203 37768
rect 11789 37710 18203 37712
rect 11789 37707 11855 37710
rect 15469 37707 15535 37710
rect 18137 37707 18203 37710
rect 19333 37770 19399 37773
rect 23381 37770 23447 37773
rect 19333 37768 23447 37770
rect 19333 37712 19338 37768
rect 19394 37712 23386 37768
rect 23442 37712 23447 37768
rect 19333 37710 23447 37712
rect 19333 37707 19399 37710
rect 23381 37707 23447 37710
rect 33593 37770 33659 37773
rect 70117 37770 70183 37773
rect 33593 37768 70183 37770
rect 33593 37712 33598 37768
rect 33654 37712 70122 37768
rect 70178 37712 70183 37768
rect 33593 37710 70183 37712
rect 33593 37707 33659 37710
rect 70117 37707 70183 37710
rect 0 37634 800 37664
rect 3877 37634 3943 37637
rect 0 37632 3943 37634
rect 0 37576 3882 37632
rect 3938 37576 3943 37632
rect 0 37574 3943 37576
rect 0 37544 800 37574
rect 3877 37571 3943 37574
rect 40401 37634 40467 37637
rect 45829 37634 45895 37637
rect 40401 37632 45895 37634
rect 40401 37576 40406 37632
rect 40462 37576 45834 37632
rect 45890 37576 45895 37632
rect 40401 37574 45895 37576
rect 40401 37571 40467 37574
rect 45829 37571 45895 37574
rect 57421 37634 57487 37637
rect 64229 37634 64295 37637
rect 57421 37632 64295 37634
rect 57421 37576 57426 37632
rect 57482 37576 64234 37632
rect 64290 37576 64295 37632
rect 57421 37574 64295 37576
rect 57421 37571 57487 37574
rect 64229 37571 64295 37574
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 50288 37568 50608 37569
rect 50288 37504 50296 37568
rect 50360 37504 50376 37568
rect 50440 37504 50456 37568
rect 50520 37504 50536 37568
rect 50600 37504 50608 37568
rect 50288 37503 50608 37504
rect 81008 37568 81328 37569
rect 81008 37504 81016 37568
rect 81080 37504 81096 37568
rect 81160 37504 81176 37568
rect 81240 37504 81256 37568
rect 81320 37504 81328 37568
rect 81008 37503 81328 37504
rect 40861 37498 40927 37501
rect 46197 37498 46263 37501
rect 40861 37496 46263 37498
rect 40861 37440 40866 37496
rect 40922 37440 46202 37496
rect 46258 37440 46263 37496
rect 40861 37438 46263 37440
rect 40861 37435 40927 37438
rect 46197 37435 46263 37438
rect 14549 37362 14615 37365
rect 65517 37362 65583 37365
rect 14549 37360 65583 37362
rect 14549 37304 14554 37360
rect 14610 37304 65522 37360
rect 65578 37304 65583 37360
rect 14549 37302 65583 37304
rect 14549 37299 14615 37302
rect 65517 37299 65583 37302
rect 19333 37226 19399 37229
rect 20161 37226 20227 37229
rect 19333 37224 20227 37226
rect 19333 37168 19338 37224
rect 19394 37168 20166 37224
rect 20222 37168 20227 37224
rect 19333 37166 20227 37168
rect 19333 37163 19399 37166
rect 20161 37163 20227 37166
rect 48957 37226 49023 37229
rect 56225 37226 56291 37229
rect 48957 37224 56291 37226
rect 48957 37168 48962 37224
rect 49018 37168 56230 37224
rect 56286 37168 56291 37224
rect 48957 37166 56291 37168
rect 48957 37163 49023 37166
rect 56225 37163 56291 37166
rect 0 37090 800 37120
rect 3969 37090 4035 37093
rect 0 37088 4035 37090
rect 0 37032 3974 37088
rect 4030 37032 4035 37088
rect 0 37030 4035 37032
rect 0 37000 800 37030
rect 3969 37027 4035 37030
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 65648 37024 65968 37025
rect 65648 36960 65656 37024
rect 65720 36960 65736 37024
rect 65800 36960 65816 37024
rect 65880 36960 65896 37024
rect 65960 36960 65968 37024
rect 65648 36959 65968 36960
rect 96368 37024 96688 37025
rect 96368 36960 96376 37024
rect 96440 36960 96456 37024
rect 96520 36960 96536 37024
rect 96600 36960 96616 37024
rect 96680 36960 96688 37024
rect 96368 36959 96688 36960
rect 12249 36818 12315 36821
rect 19241 36818 19307 36821
rect 12249 36816 19307 36818
rect 12249 36760 12254 36816
rect 12310 36760 19246 36816
rect 19302 36760 19307 36816
rect 12249 36758 19307 36760
rect 12249 36755 12315 36758
rect 19241 36755 19307 36758
rect 43161 36818 43227 36821
rect 48037 36818 48103 36821
rect 43161 36816 48103 36818
rect 43161 36760 43166 36816
rect 43222 36760 48042 36816
rect 48098 36760 48103 36816
rect 43161 36758 48103 36760
rect 43161 36755 43227 36758
rect 48037 36755 48103 36758
rect 50429 36818 50495 36821
rect 56777 36818 56843 36821
rect 57881 36818 57947 36821
rect 50429 36816 57947 36818
rect 50429 36760 50434 36816
rect 50490 36760 56782 36816
rect 56838 36760 57886 36816
rect 57942 36760 57947 36816
rect 50429 36758 57947 36760
rect 50429 36755 50495 36758
rect 56777 36755 56843 36758
rect 57881 36755 57947 36758
rect 91001 36818 91067 36821
rect 95325 36818 95391 36821
rect 91001 36816 95391 36818
rect 91001 36760 91006 36816
rect 91062 36760 95330 36816
rect 95386 36760 95391 36816
rect 91001 36758 95391 36760
rect 91001 36755 91067 36758
rect 95325 36755 95391 36758
rect 12341 36682 12407 36685
rect 14089 36682 14155 36685
rect 12341 36680 14155 36682
rect 12341 36624 12346 36680
rect 12402 36624 14094 36680
rect 14150 36624 14155 36680
rect 12341 36622 14155 36624
rect 12341 36619 12407 36622
rect 14089 36619 14155 36622
rect 18965 36682 19031 36685
rect 19885 36682 19951 36685
rect 18965 36680 19951 36682
rect 18965 36624 18970 36680
rect 19026 36624 19890 36680
rect 19946 36624 19951 36680
rect 18965 36622 19951 36624
rect 18965 36619 19031 36622
rect 19885 36619 19951 36622
rect 19568 36480 19888 36481
rect 0 36410 800 36440
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 50288 36480 50608 36481
rect 50288 36416 50296 36480
rect 50360 36416 50376 36480
rect 50440 36416 50456 36480
rect 50520 36416 50536 36480
rect 50600 36416 50608 36480
rect 50288 36415 50608 36416
rect 81008 36480 81328 36481
rect 81008 36416 81016 36480
rect 81080 36416 81096 36480
rect 81160 36416 81176 36480
rect 81240 36416 81256 36480
rect 81320 36416 81328 36480
rect 81008 36415 81328 36416
rect 4061 36410 4127 36413
rect 0 36408 4127 36410
rect 0 36352 4066 36408
rect 4122 36352 4127 36408
rect 0 36350 4127 36352
rect 0 36320 800 36350
rect 4061 36347 4127 36350
rect 51717 36410 51783 36413
rect 58157 36410 58223 36413
rect 51717 36408 58223 36410
rect 51717 36352 51722 36408
rect 51778 36352 58162 36408
rect 58218 36352 58223 36408
rect 51717 36350 58223 36352
rect 51717 36347 51783 36350
rect 58157 36347 58223 36350
rect 20161 36274 20227 36277
rect 24853 36274 24919 36277
rect 20161 36272 24919 36274
rect 20161 36216 20166 36272
rect 20222 36216 24858 36272
rect 24914 36216 24919 36272
rect 20161 36214 24919 36216
rect 20161 36211 20227 36214
rect 24853 36211 24919 36214
rect 29545 36274 29611 36277
rect 35617 36274 35683 36277
rect 29545 36272 35683 36274
rect 29545 36216 29550 36272
rect 29606 36216 35622 36272
rect 35678 36216 35683 36272
rect 29545 36214 35683 36216
rect 29545 36211 29611 36214
rect 35617 36211 35683 36214
rect 77845 36274 77911 36277
rect 79225 36274 79291 36277
rect 77845 36272 79291 36274
rect 77845 36216 77850 36272
rect 77906 36216 79230 36272
rect 79286 36216 79291 36272
rect 77845 36214 79291 36216
rect 77845 36211 77911 36214
rect 79225 36211 79291 36214
rect 13169 36138 13235 36141
rect 40125 36138 40191 36141
rect 13169 36136 40191 36138
rect 13169 36080 13174 36136
rect 13230 36080 40130 36136
rect 40186 36080 40191 36136
rect 13169 36078 40191 36080
rect 13169 36075 13235 36078
rect 40125 36075 40191 36078
rect 57973 36138 58039 36141
rect 67449 36138 67515 36141
rect 57973 36136 67515 36138
rect 57973 36080 57978 36136
rect 58034 36080 67454 36136
rect 67510 36080 67515 36136
rect 57973 36078 67515 36080
rect 57973 36075 58039 36078
rect 67449 36075 67515 36078
rect 77569 36138 77635 36141
rect 79777 36138 79843 36141
rect 77569 36136 79843 36138
rect 77569 36080 77574 36136
rect 77630 36080 79782 36136
rect 79838 36080 79843 36136
rect 77569 36078 79843 36080
rect 77569 36075 77635 36078
rect 79777 36075 79843 36078
rect 4208 35936 4528 35937
rect 0 35866 800 35896
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 35871 35248 35872
rect 65648 35936 65968 35937
rect 65648 35872 65656 35936
rect 65720 35872 65736 35936
rect 65800 35872 65816 35936
rect 65880 35872 65896 35936
rect 65960 35872 65968 35936
rect 65648 35871 65968 35872
rect 96368 35936 96688 35937
rect 96368 35872 96376 35936
rect 96440 35872 96456 35936
rect 96520 35872 96536 35936
rect 96600 35872 96616 35936
rect 96680 35872 96688 35936
rect 96368 35871 96688 35872
rect 4061 35866 4127 35869
rect 0 35864 4127 35866
rect 0 35808 4066 35864
rect 4122 35808 4127 35864
rect 0 35806 4127 35808
rect 0 35776 800 35806
rect 4061 35803 4127 35806
rect 49877 35866 49943 35869
rect 51717 35866 51783 35869
rect 49877 35864 51783 35866
rect 49877 35808 49882 35864
rect 49938 35808 51722 35864
rect 51778 35808 51783 35864
rect 49877 35806 51783 35808
rect 49877 35803 49943 35806
rect 51717 35803 51783 35806
rect 55949 35866 56015 35869
rect 56961 35866 57027 35869
rect 55949 35864 57027 35866
rect 55949 35808 55954 35864
rect 56010 35808 56966 35864
rect 57022 35808 57027 35864
rect 55949 35806 57027 35808
rect 55949 35803 56015 35806
rect 56961 35803 57027 35806
rect 67633 35866 67699 35869
rect 73061 35866 73127 35869
rect 67633 35864 73127 35866
rect 67633 35808 67638 35864
rect 67694 35808 73066 35864
rect 73122 35808 73127 35864
rect 67633 35806 73127 35808
rect 67633 35803 67699 35806
rect 73061 35803 73127 35806
rect 77385 35866 77451 35869
rect 85849 35866 85915 35869
rect 77385 35864 85915 35866
rect 77385 35808 77390 35864
rect 77446 35808 85854 35864
rect 85910 35808 85915 35864
rect 77385 35806 85915 35808
rect 77385 35803 77451 35806
rect 85849 35803 85915 35806
rect 24117 35730 24183 35733
rect 26969 35730 27035 35733
rect 24117 35728 27035 35730
rect 24117 35672 24122 35728
rect 24178 35672 26974 35728
rect 27030 35672 27035 35728
rect 24117 35670 27035 35672
rect 24117 35667 24183 35670
rect 26969 35667 27035 35670
rect 55213 35730 55279 35733
rect 56317 35730 56383 35733
rect 85481 35730 85547 35733
rect 55213 35728 85547 35730
rect 55213 35672 55218 35728
rect 55274 35672 56322 35728
rect 56378 35672 85486 35728
rect 85542 35672 85547 35728
rect 55213 35670 85547 35672
rect 55213 35667 55279 35670
rect 56317 35667 56383 35670
rect 85481 35667 85547 35670
rect 30189 35594 30255 35597
rect 36445 35594 36511 35597
rect 30189 35592 36511 35594
rect 30189 35536 30194 35592
rect 30250 35536 36450 35592
rect 36506 35536 36511 35592
rect 30189 35534 36511 35536
rect 30189 35531 30255 35534
rect 36445 35531 36511 35534
rect 49417 35594 49483 35597
rect 52453 35594 52519 35597
rect 49417 35592 52519 35594
rect 49417 35536 49422 35592
rect 49478 35536 52458 35592
rect 52514 35536 52519 35592
rect 49417 35534 52519 35536
rect 49417 35531 49483 35534
rect 52453 35531 52519 35534
rect 59077 35594 59143 35597
rect 69933 35594 69999 35597
rect 59077 35592 69999 35594
rect 59077 35536 59082 35592
rect 59138 35536 69938 35592
rect 69994 35536 69999 35592
rect 59077 35534 69999 35536
rect 59077 35531 59143 35534
rect 69933 35531 69999 35534
rect 78305 35594 78371 35597
rect 80145 35594 80211 35597
rect 78305 35592 80211 35594
rect 78305 35536 78310 35592
rect 78366 35536 80150 35592
rect 80206 35536 80211 35592
rect 78305 35534 80211 35536
rect 78305 35531 78371 35534
rect 80145 35531 80211 35534
rect 50889 35458 50955 35461
rect 55765 35458 55831 35461
rect 56593 35458 56659 35461
rect 50889 35456 56659 35458
rect 50889 35400 50894 35456
rect 50950 35400 55770 35456
rect 55826 35400 56598 35456
rect 56654 35400 56659 35456
rect 50889 35398 56659 35400
rect 50889 35395 50955 35398
rect 55765 35395 55831 35398
rect 56593 35395 56659 35398
rect 58893 35458 58959 35461
rect 66989 35458 67055 35461
rect 58893 35456 67055 35458
rect 58893 35400 58898 35456
rect 58954 35400 66994 35456
rect 67050 35400 67055 35456
rect 58893 35398 67055 35400
rect 58893 35395 58959 35398
rect 66989 35395 67055 35398
rect 68645 35458 68711 35461
rect 76649 35458 76715 35461
rect 68645 35456 76715 35458
rect 68645 35400 68650 35456
rect 68706 35400 76654 35456
rect 76710 35400 76715 35456
rect 68645 35398 76715 35400
rect 68645 35395 68711 35398
rect 76649 35395 76715 35398
rect 19568 35392 19888 35393
rect 0 35322 800 35352
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 35327 19888 35328
rect 50288 35392 50608 35393
rect 50288 35328 50296 35392
rect 50360 35328 50376 35392
rect 50440 35328 50456 35392
rect 50520 35328 50536 35392
rect 50600 35328 50608 35392
rect 50288 35327 50608 35328
rect 81008 35392 81328 35393
rect 81008 35328 81016 35392
rect 81080 35328 81096 35392
rect 81160 35328 81176 35392
rect 81240 35328 81256 35392
rect 81320 35328 81328 35392
rect 81008 35327 81328 35328
rect 3417 35322 3483 35325
rect 0 35320 3483 35322
rect 0 35264 3422 35320
rect 3478 35264 3483 35320
rect 0 35262 3483 35264
rect 0 35232 800 35262
rect 3417 35259 3483 35262
rect 41781 35322 41847 35325
rect 47761 35322 47827 35325
rect 41781 35320 47827 35322
rect 41781 35264 41786 35320
rect 41842 35264 47766 35320
rect 47822 35264 47827 35320
rect 41781 35262 47827 35264
rect 41781 35259 41847 35262
rect 47761 35259 47827 35262
rect 53741 35322 53807 35325
rect 55765 35322 55831 35325
rect 53741 35320 55831 35322
rect 53741 35264 53746 35320
rect 53802 35264 55770 35320
rect 55826 35264 55831 35320
rect 53741 35262 55831 35264
rect 53741 35259 53807 35262
rect 55765 35259 55831 35262
rect 58617 35322 58683 35325
rect 66161 35322 66227 35325
rect 58617 35320 66227 35322
rect 58617 35264 58622 35320
rect 58678 35264 66166 35320
rect 66222 35264 66227 35320
rect 58617 35262 66227 35264
rect 58617 35259 58683 35262
rect 66161 35259 66227 35262
rect 19701 35186 19767 35189
rect 25497 35186 25563 35189
rect 19701 35184 25563 35186
rect 19701 35128 19706 35184
rect 19762 35128 25502 35184
rect 25558 35128 25563 35184
rect 19701 35126 25563 35128
rect 19701 35123 19767 35126
rect 25497 35123 25563 35126
rect 30557 35186 30623 35189
rect 36813 35186 36879 35189
rect 30557 35184 36879 35186
rect 30557 35128 30562 35184
rect 30618 35128 36818 35184
rect 36874 35128 36879 35184
rect 30557 35126 36879 35128
rect 30557 35123 30623 35126
rect 36813 35123 36879 35126
rect 39573 35186 39639 35189
rect 75361 35186 75427 35189
rect 39573 35184 75427 35186
rect 39573 35128 39578 35184
rect 39634 35128 75366 35184
rect 75422 35128 75427 35184
rect 39573 35126 75427 35128
rect 39573 35123 39639 35126
rect 75361 35123 75427 35126
rect 79501 35186 79567 35189
rect 83549 35186 83615 35189
rect 79501 35184 83615 35186
rect 79501 35128 79506 35184
rect 79562 35128 83554 35184
rect 83610 35128 83615 35184
rect 79501 35126 83615 35128
rect 79501 35123 79567 35126
rect 83549 35123 83615 35126
rect 14641 35050 14707 35053
rect 74257 35050 74323 35053
rect 14641 35048 74323 35050
rect 14641 34992 14646 35048
rect 14702 34992 74262 35048
rect 74318 34992 74323 35048
rect 14641 34990 74323 34992
rect 14641 34987 14707 34990
rect 74257 34987 74323 34990
rect 77293 35050 77359 35053
rect 84377 35050 84443 35053
rect 84745 35050 84811 35053
rect 85573 35050 85639 35053
rect 86033 35050 86099 35053
rect 77293 35048 86099 35050
rect 77293 34992 77298 35048
rect 77354 34992 84382 35048
rect 84438 34992 84750 35048
rect 84806 34992 85578 35048
rect 85634 34992 86038 35048
rect 86094 34992 86099 35048
rect 77293 34990 86099 34992
rect 77293 34987 77359 34990
rect 84377 34987 84443 34990
rect 84745 34987 84811 34990
rect 85573 34987 85639 34990
rect 86033 34987 86099 34990
rect 38745 34914 38811 34917
rect 46841 34914 46907 34917
rect 38745 34912 46907 34914
rect 38745 34856 38750 34912
rect 38806 34856 46846 34912
rect 46902 34856 46907 34912
rect 38745 34854 46907 34856
rect 38745 34851 38811 34854
rect 46841 34851 46907 34854
rect 51809 34914 51875 34917
rect 56961 34914 57027 34917
rect 51809 34912 57027 34914
rect 51809 34856 51814 34912
rect 51870 34856 56966 34912
rect 57022 34856 57027 34912
rect 51809 34854 57027 34856
rect 51809 34851 51875 34854
rect 56961 34851 57027 34854
rect 76189 34914 76255 34917
rect 76741 34914 76807 34917
rect 78029 34914 78095 34917
rect 76189 34912 78095 34914
rect 76189 34856 76194 34912
rect 76250 34856 76746 34912
rect 76802 34856 78034 34912
rect 78090 34856 78095 34912
rect 76189 34854 78095 34856
rect 76189 34851 76255 34854
rect 76741 34851 76807 34854
rect 78029 34851 78095 34854
rect 4208 34848 4528 34849
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 65648 34848 65968 34849
rect 65648 34784 65656 34848
rect 65720 34784 65736 34848
rect 65800 34784 65816 34848
rect 65880 34784 65896 34848
rect 65960 34784 65968 34848
rect 65648 34783 65968 34784
rect 96368 34848 96688 34849
rect 96368 34784 96376 34848
rect 96440 34784 96456 34848
rect 96520 34784 96536 34848
rect 96600 34784 96616 34848
rect 96680 34784 96688 34848
rect 96368 34783 96688 34784
rect 21265 34778 21331 34781
rect 22277 34778 22343 34781
rect 26601 34778 26667 34781
rect 21265 34776 26667 34778
rect 21265 34720 21270 34776
rect 21326 34720 22282 34776
rect 22338 34720 26606 34776
rect 26662 34720 26667 34776
rect 21265 34718 26667 34720
rect 21265 34715 21331 34718
rect 22277 34715 22343 34718
rect 26601 34715 26667 34718
rect 38837 34778 38903 34781
rect 40585 34778 40651 34781
rect 38837 34776 40651 34778
rect 38837 34720 38842 34776
rect 38898 34720 40590 34776
rect 40646 34720 40651 34776
rect 38837 34718 40651 34720
rect 38837 34715 38903 34718
rect 40585 34715 40651 34718
rect 54109 34778 54175 34781
rect 54845 34778 54911 34781
rect 54109 34776 54911 34778
rect 54109 34720 54114 34776
rect 54170 34720 54850 34776
rect 54906 34720 54911 34776
rect 54109 34718 54911 34720
rect 54109 34715 54175 34718
rect 54845 34715 54911 34718
rect 78489 34778 78555 34781
rect 81433 34778 81499 34781
rect 78489 34776 81499 34778
rect 78489 34720 78494 34776
rect 78550 34720 81438 34776
rect 81494 34720 81499 34776
rect 78489 34718 81499 34720
rect 78489 34715 78555 34718
rect 81433 34715 81499 34718
rect 0 34642 800 34672
rect 3877 34642 3943 34645
rect 0 34640 3943 34642
rect 0 34584 3882 34640
rect 3938 34584 3943 34640
rect 0 34582 3943 34584
rect 0 34552 800 34582
rect 3877 34579 3943 34582
rect 20069 34642 20135 34645
rect 22921 34642 22987 34645
rect 20069 34640 22987 34642
rect 20069 34584 20074 34640
rect 20130 34584 22926 34640
rect 22982 34584 22987 34640
rect 20069 34582 22987 34584
rect 20069 34579 20135 34582
rect 22921 34579 22987 34582
rect 33869 34642 33935 34645
rect 78581 34642 78647 34645
rect 78949 34642 79015 34645
rect 33869 34640 79015 34642
rect 33869 34584 33874 34640
rect 33930 34584 78586 34640
rect 78642 34584 78954 34640
rect 79010 34584 79015 34640
rect 33869 34582 79015 34584
rect 33869 34579 33935 34582
rect 78581 34579 78647 34582
rect 78949 34579 79015 34582
rect 51809 34506 51875 34509
rect 56501 34506 56567 34509
rect 51809 34504 56567 34506
rect 51809 34448 51814 34504
rect 51870 34448 56506 34504
rect 56562 34448 56567 34504
rect 51809 34446 56567 34448
rect 51809 34443 51875 34446
rect 56501 34443 56567 34446
rect 58157 34506 58223 34509
rect 58893 34506 58959 34509
rect 66345 34506 66411 34509
rect 58157 34504 66411 34506
rect 58157 34448 58162 34504
rect 58218 34448 58898 34504
rect 58954 34448 66350 34504
rect 66406 34448 66411 34504
rect 58157 34446 66411 34448
rect 58157 34443 58223 34446
rect 58893 34443 58959 34446
rect 66345 34443 66411 34446
rect 78489 34506 78555 34509
rect 79961 34506 80027 34509
rect 81985 34506 82051 34509
rect 78489 34504 82051 34506
rect 78489 34448 78494 34504
rect 78550 34448 79966 34504
rect 80022 34448 81990 34504
rect 82046 34448 82051 34504
rect 78489 34446 82051 34448
rect 78489 34443 78555 34446
rect 79961 34443 80027 34446
rect 81985 34443 82051 34446
rect 57513 34370 57579 34373
rect 58985 34370 59051 34373
rect 57513 34368 59051 34370
rect 57513 34312 57518 34368
rect 57574 34312 58990 34368
rect 59046 34312 59051 34368
rect 57513 34310 59051 34312
rect 57513 34307 57579 34310
rect 58985 34307 59051 34310
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 50288 34304 50608 34305
rect 50288 34240 50296 34304
rect 50360 34240 50376 34304
rect 50440 34240 50456 34304
rect 50520 34240 50536 34304
rect 50600 34240 50608 34304
rect 50288 34239 50608 34240
rect 81008 34304 81328 34305
rect 81008 34240 81016 34304
rect 81080 34240 81096 34304
rect 81160 34240 81176 34304
rect 81240 34240 81256 34304
rect 81320 34240 81328 34304
rect 81008 34239 81328 34240
rect 0 34098 800 34128
rect 3233 34098 3299 34101
rect 0 34096 3299 34098
rect 0 34040 3238 34096
rect 3294 34040 3299 34096
rect 0 34038 3299 34040
rect 0 34008 800 34038
rect 3233 34035 3299 34038
rect 21173 34098 21239 34101
rect 24853 34098 24919 34101
rect 21173 34096 24919 34098
rect 21173 34040 21178 34096
rect 21234 34040 24858 34096
rect 24914 34040 24919 34096
rect 21173 34038 24919 34040
rect 21173 34035 21239 34038
rect 24853 34035 24919 34038
rect 20437 33962 20503 33965
rect 24577 33962 24643 33965
rect 20437 33960 24643 33962
rect 20437 33904 20442 33960
rect 20498 33904 24582 33960
rect 24638 33904 24643 33960
rect 20437 33902 24643 33904
rect 20437 33899 20503 33902
rect 24577 33899 24643 33902
rect 18045 33826 18111 33829
rect 27521 33826 27587 33829
rect 18045 33824 27587 33826
rect 18045 33768 18050 33824
rect 18106 33768 27526 33824
rect 27582 33768 27587 33824
rect 18045 33766 27587 33768
rect 18045 33763 18111 33766
rect 27521 33763 27587 33766
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 0 33554 800 33584
rect 4061 33554 4127 33557
rect 0 33552 4127 33554
rect 0 33496 4066 33552
rect 4122 33496 4127 33552
rect 0 33494 4127 33496
rect 0 33464 800 33494
rect 4061 33491 4127 33494
rect 21265 33554 21331 33557
rect 22185 33554 22251 33557
rect 21265 33552 22251 33554
rect 21265 33496 21270 33552
rect 21326 33496 22190 33552
rect 22246 33496 22251 33552
rect 21265 33494 22251 33496
rect 21265 33491 21331 33494
rect 22185 33491 22251 33494
rect 20989 33418 21055 33421
rect 22369 33418 22435 33421
rect 20989 33416 22435 33418
rect 20989 33360 20994 33416
rect 21050 33360 22374 33416
rect 22430 33360 22435 33416
rect 20989 33358 22435 33360
rect 20989 33355 21055 33358
rect 22369 33355 22435 33358
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 33151 19888 33152
rect 0 32874 800 32904
rect 3877 32874 3943 32877
rect 0 32872 3943 32874
rect 0 32816 3882 32872
rect 3938 32816 3943 32872
rect 0 32814 3943 32816
rect 0 32784 800 32814
rect 3877 32811 3943 32814
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 0 32330 800 32360
rect 5901 32330 5967 32333
rect 0 32328 5967 32330
rect 0 32272 5906 32328
rect 5962 32272 5967 32328
rect 0 32270 5967 32272
rect 0 32240 800 32270
rect 5901 32267 5967 32270
rect 19568 32128 19888 32129
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 8385 31922 8451 31925
rect 9949 31922 10015 31925
rect 8385 31920 10015 31922
rect 8385 31864 8390 31920
rect 8446 31864 9954 31920
rect 10010 31864 10015 31920
rect 8385 31862 10015 31864
rect 8385 31859 8451 31862
rect 9949 31859 10015 31862
rect 21633 31922 21699 31925
rect 22277 31922 22343 31925
rect 21633 31920 22343 31922
rect 21633 31864 21638 31920
rect 21694 31864 22282 31920
rect 22338 31864 22343 31920
rect 21633 31862 22343 31864
rect 21633 31859 21699 31862
rect 22277 31859 22343 31862
rect 0 31786 800 31816
rect 3417 31786 3483 31789
rect 0 31784 3483 31786
rect 0 31728 3422 31784
rect 3478 31728 3483 31784
rect 0 31726 3483 31728
rect 0 31696 800 31726
rect 3417 31723 3483 31726
rect 81433 31650 81499 31653
rect 82353 31650 82419 31653
rect 79918 31648 82419 31650
rect 79918 31592 81438 31648
rect 81494 31592 82358 31648
rect 82414 31592 82419 31648
rect 79918 31590 82419 31592
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 9673 31514 9739 31517
rect 11789 31514 11855 31517
rect 9673 31512 11855 31514
rect 9673 31456 9678 31512
rect 9734 31456 11794 31512
rect 11850 31456 11855 31512
rect 9673 31454 11855 31456
rect 9673 31451 9739 31454
rect 11789 31451 11855 31454
rect 29494 31452 29500 31516
rect 29564 31514 29570 31516
rect 29564 31454 72434 31514
rect 29564 31452 29570 31454
rect 72374 31378 72434 31454
rect 79918 31378 79978 31590
rect 81433 31587 81499 31590
rect 82353 31587 82419 31590
rect 102726 31514 102732 31516
rect 81758 31454 102732 31514
rect 81758 31378 81818 31454
rect 102726 31452 102732 31454
rect 102796 31452 102802 31516
rect 72374 31318 79978 31378
rect 81574 31318 81818 31378
rect 0 31106 800 31136
rect 3049 31106 3115 31109
rect 0 31104 3115 31106
rect 0 31048 3054 31104
rect 3110 31048 3115 31104
rect 0 31046 3115 31048
rect 0 31016 800 31046
rect 3049 31043 3115 31046
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 81574 30902 81634 31318
rect 81574 30842 81788 30902
rect 24209 30834 24275 30837
rect 51073 30834 51139 30837
rect 24209 30832 27508 30834
rect 24209 30776 24214 30832
rect 24270 30776 27508 30832
rect 24209 30774 27508 30776
rect 51073 30832 54004 30834
rect 51073 30776 51078 30832
rect 51134 30776 54004 30832
rect 51073 30774 54004 30776
rect 24209 30771 24275 30774
rect 51073 30771 51139 30774
rect 0 30562 800 30592
rect 3877 30562 3943 30565
rect 0 30560 3943 30562
rect 0 30504 3882 30560
rect 3938 30504 3943 30560
rect 0 30502 3943 30504
rect 0 30472 800 30502
rect 3877 30499 3943 30502
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 53833 30222 53899 30225
rect 81525 30222 81591 30225
rect 53833 30220 54004 30222
rect 53833 30164 53838 30220
rect 53894 30164 54004 30220
rect 53833 30162 54004 30164
rect 81525 30220 81788 30222
rect 81525 30164 81530 30220
rect 81586 30164 81788 30220
rect 81525 30162 81788 30164
rect 53833 30159 53899 30162
rect 81525 30159 81591 30162
rect 23473 30154 23539 30157
rect 23473 30152 27508 30154
rect 23473 30096 23478 30152
rect 23534 30096 27508 30152
rect 23473 30094 27508 30096
rect 23473 30091 23539 30094
rect 19568 29952 19888 29953
rect 0 29882 800 29912
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 2957 29882 3023 29885
rect 0 29880 3023 29882
rect 0 29824 2962 29880
rect 3018 29824 3023 29880
rect 0 29822 3023 29824
rect 0 29792 800 29822
rect 2957 29819 3023 29822
rect 81433 29542 81499 29545
rect 81433 29540 81788 29542
rect 81433 29484 81438 29540
rect 81494 29484 81788 29540
rect 81433 29482 81788 29484
rect 81433 29479 81499 29482
rect 24761 29474 24827 29477
rect 24761 29472 27508 29474
rect 24761 29416 24766 29472
rect 24822 29416 27508 29472
rect 24761 29414 27508 29416
rect 24761 29411 24827 29414
rect 51574 29412 51580 29476
rect 51644 29474 51650 29476
rect 53833 29474 53899 29477
rect 51644 29472 54004 29474
rect 51644 29416 53838 29472
rect 53894 29416 54004 29472
rect 51644 29414 54004 29416
rect 51644 29412 51650 29414
rect 53833 29411 53899 29414
rect 4208 29408 4528 29409
rect 0 29338 800 29368
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 4061 29338 4127 29341
rect 0 29336 4127 29338
rect 0 29280 4066 29336
rect 4122 29280 4127 29336
rect 0 29278 4127 29280
rect 0 29248 800 29278
rect 4061 29275 4127 29278
rect 3049 28930 3115 28933
rect 3325 28930 3391 28933
rect 3049 28928 3391 28930
rect 3049 28872 3054 28928
rect 3110 28872 3330 28928
rect 3386 28872 3391 28928
rect 3049 28870 3391 28872
rect 3049 28867 3115 28870
rect 3325 28867 3391 28870
rect 19568 28864 19888 28865
rect 0 28794 800 28824
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 4061 28794 4127 28797
rect 0 28792 4127 28794
rect 0 28736 4066 28792
rect 4122 28736 4127 28792
rect 0 28734 4127 28736
rect 0 28704 800 28734
rect 4061 28731 4127 28734
rect 19517 28658 19583 28661
rect 22645 28658 22711 28661
rect 19517 28656 22711 28658
rect 19517 28600 19522 28656
rect 19578 28600 22650 28656
rect 22706 28600 22711 28656
rect 19517 28598 22711 28600
rect 19517 28595 19583 28598
rect 22645 28595 22711 28598
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 53833 28182 53899 28185
rect 81617 28182 81683 28185
rect 53833 28180 54004 28182
rect 0 28114 800 28144
rect 53833 28124 53838 28180
rect 53894 28124 54004 28180
rect 53833 28122 54004 28124
rect 81206 28180 81788 28182
rect 81206 28124 81622 28180
rect 81678 28124 81788 28180
rect 81206 28122 81788 28124
rect 53833 28119 53899 28122
rect 3877 28114 3943 28117
rect 0 28112 3943 28114
rect 0 28056 3882 28112
rect 3938 28056 3943 28112
rect 0 28054 3943 28056
rect 0 28024 800 28054
rect 3877 28051 3943 28054
rect 23381 28114 23447 28117
rect 23381 28112 27508 28114
rect 23381 28056 23386 28112
rect 23442 28056 27508 28112
rect 23381 28054 27508 28056
rect 23381 28051 23447 28054
rect 79174 28052 79180 28116
rect 79244 28114 79250 28116
rect 81206 28114 81266 28122
rect 81617 28119 81683 28122
rect 79244 28054 81266 28114
rect 79244 28052 79250 28054
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 0 27570 800 27600
rect 4061 27570 4127 27573
rect 0 27568 4127 27570
rect 0 27512 4066 27568
rect 4122 27512 4127 27568
rect 0 27510 4127 27512
rect 0 27480 800 27510
rect 4061 27507 4127 27510
rect 9581 27570 9647 27573
rect 12433 27570 12499 27573
rect 9581 27568 12499 27570
rect 9581 27512 9586 27568
rect 9642 27512 12438 27568
rect 12494 27512 12499 27568
rect 9581 27510 12499 27512
rect 9581 27507 9647 27510
rect 12433 27507 12499 27510
rect 8477 27434 8543 27437
rect 9765 27434 9831 27437
rect 8477 27432 9831 27434
rect 8477 27376 8482 27432
rect 8538 27376 9770 27432
rect 9826 27376 9831 27432
rect 8477 27374 9831 27376
rect 8477 27371 8543 27374
rect 9765 27371 9831 27374
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 0 27026 800 27056
rect 3877 27026 3943 27029
rect 0 27024 3943 27026
rect 0 26968 3882 27024
rect 3938 26968 3943 27024
rect 0 26966 3943 26968
rect 0 26936 800 26966
rect 3877 26963 3943 26966
rect 81617 26822 81683 26825
rect 81206 26820 81788 26822
rect 81206 26764 81622 26820
rect 81678 26764 81788 26820
rect 81206 26762 81788 26764
rect 24301 26754 24367 26757
rect 24301 26752 27508 26754
rect 24301 26696 24306 26752
rect 24362 26696 27508 26752
rect 24301 26694 27508 26696
rect 24301 26691 24367 26694
rect 52310 26692 52316 26756
rect 52380 26754 52386 26756
rect 53833 26754 53899 26757
rect 52380 26752 54004 26754
rect 52380 26696 53838 26752
rect 53894 26696 54004 26752
rect 52380 26694 54004 26696
rect 52380 26692 52386 26694
rect 53833 26691 53899 26694
rect 79542 26692 79548 26756
rect 79612 26754 79618 26756
rect 81206 26754 81266 26762
rect 81617 26759 81683 26762
rect 79612 26694 81266 26754
rect 79612 26692 79618 26694
rect 19568 26688 19888 26689
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 0 26346 800 26376
rect 4061 26346 4127 26349
rect 0 26344 4127 26346
rect 0 26288 4066 26344
rect 4122 26288 4127 26344
rect 0 26286 4127 26288
rect 0 26256 800 26286
rect 4061 26283 4127 26286
rect 7465 26210 7531 26213
rect 7598 26210 7604 26212
rect 7465 26208 7604 26210
rect 7465 26152 7470 26208
rect 7526 26152 7604 26208
rect 7465 26150 7604 26152
rect 7465 26147 7531 26150
rect 7598 26148 7604 26150
rect 7668 26148 7674 26212
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 0 25802 800 25832
rect 3877 25802 3943 25805
rect 0 25800 3943 25802
rect 0 25744 3882 25800
rect 3938 25744 3943 25800
rect 0 25742 3943 25744
rect 0 25712 800 25742
rect 3877 25739 3943 25742
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 81617 25598 81683 25601
rect 81617 25596 81788 25598
rect 81617 25540 81622 25596
rect 81678 25540 81788 25596
rect 81617 25538 81788 25540
rect 81617 25535 81683 25538
rect 24761 25530 24827 25533
rect 51993 25530 52059 25533
rect 52310 25530 52316 25532
rect 24761 25528 27508 25530
rect 24761 25472 24766 25528
rect 24822 25472 27508 25528
rect 24761 25470 27508 25472
rect 51993 25528 52316 25530
rect 51993 25472 51998 25528
rect 52054 25472 52316 25528
rect 51993 25470 52316 25472
rect 24761 25467 24827 25470
rect 51993 25467 52059 25470
rect 52310 25468 52316 25470
rect 52380 25530 52386 25532
rect 52380 25470 54004 25530
rect 52380 25468 52386 25470
rect 0 25258 800 25288
rect 4061 25258 4127 25261
rect 0 25256 4127 25258
rect 0 25200 4066 25256
rect 4122 25200 4127 25256
rect 0 25198 4127 25200
rect 0 25168 800 25198
rect 4061 25195 4127 25198
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 0 24578 800 24608
rect 3877 24578 3943 24581
rect 0 24576 3943 24578
rect 0 24520 3882 24576
rect 3938 24520 3943 24576
rect 0 24518 3943 24520
rect 0 24488 800 24518
rect 3877 24515 3943 24518
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 53833 24238 53899 24241
rect 81341 24238 81407 24241
rect 53422 24236 54004 24238
rect 53422 24180 53838 24236
rect 53894 24180 54004 24236
rect 53422 24178 54004 24180
rect 81206 24236 81788 24238
rect 81206 24180 81346 24236
rect 81402 24180 81788 24236
rect 81206 24178 81788 24180
rect 23565 24170 23631 24173
rect 23565 24168 27508 24170
rect 23565 24112 23570 24168
rect 23626 24112 27508 24168
rect 23565 24110 27508 24112
rect 23565 24107 23631 24110
rect 51942 24108 51948 24172
rect 52012 24170 52018 24172
rect 53422 24170 53482 24178
rect 53833 24175 53899 24178
rect 52012 24110 53482 24170
rect 52012 24108 52018 24110
rect 79726 24108 79732 24172
rect 79796 24170 79802 24172
rect 81206 24170 81266 24178
rect 81341 24175 81407 24178
rect 79796 24110 81266 24170
rect 79796 24108 79802 24110
rect 0 24034 800 24064
rect 4061 24034 4127 24037
rect 0 24032 4127 24034
rect 0 23976 4066 24032
rect 4122 23976 4127 24032
rect 0 23974 4127 23976
rect 0 23944 800 23974
rect 4061 23971 4127 23974
rect 4208 23968 4528 23969
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 0 23490 800 23520
rect 3233 23490 3299 23493
rect 0 23488 3299 23490
rect 0 23432 3238 23488
rect 3294 23432 3299 23488
rect 0 23430 3299 23432
rect 0 23400 800 23430
rect 3233 23427 3299 23430
rect 12617 23490 12683 23493
rect 12750 23490 12756 23492
rect 12617 23488 12756 23490
rect 12617 23432 12622 23488
rect 12678 23432 12756 23488
rect 12617 23430 12756 23432
rect 12617 23427 12683 23430
rect 12750 23428 12756 23430
rect 12820 23428 12826 23492
rect 20161 23490 20227 23493
rect 26366 23490 26372 23492
rect 20161 23488 26372 23490
rect 20161 23432 20166 23488
rect 20222 23432 26372 23488
rect 20161 23430 26372 23432
rect 20161 23427 20227 23430
rect 26366 23428 26372 23430
rect 26436 23428 26442 23492
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 102726 23156 102732 23220
rect 102796 23218 102802 23220
rect 105920 23218 106720 23248
rect 102796 23158 106720 23218
rect 102796 23156 102802 23158
rect 105920 23128 106720 23158
rect 4208 22880 4528 22881
rect 0 22810 800 22840
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 81617 22878 81683 22881
rect 4208 22815 4528 22816
rect 81390 22876 81788 22878
rect 81390 22820 81622 22876
rect 81678 22820 81788 22876
rect 81390 22818 81788 22820
rect 4061 22810 4127 22813
rect 0 22808 4127 22810
rect 0 22752 4066 22808
rect 4122 22752 4127 22808
rect 0 22750 4127 22752
rect 0 22720 800 22750
rect 4061 22747 4127 22750
rect 9673 22810 9739 22813
rect 9806 22810 9812 22812
rect 9673 22808 9812 22810
rect 9673 22752 9678 22808
rect 9734 22752 9812 22808
rect 9673 22750 9812 22752
rect 9673 22747 9739 22750
rect 9806 22748 9812 22750
rect 9876 22748 9882 22812
rect 23473 22810 23539 22813
rect 52361 22812 52427 22813
rect 52310 22810 52316 22812
rect 23473 22808 27508 22810
rect 23473 22752 23478 22808
rect 23534 22752 27508 22808
rect 23473 22750 27508 22752
rect 52234 22750 52316 22810
rect 52380 22810 52427 22812
rect 52380 22808 54004 22810
rect 52422 22752 54004 22808
rect 23473 22747 23539 22750
rect 52310 22748 52316 22750
rect 52380 22750 54004 22752
rect 52380 22748 52427 22750
rect 78622 22748 78628 22812
rect 78692 22810 78698 22812
rect 81390 22810 81450 22818
rect 81617 22815 81683 22818
rect 78692 22750 81450 22810
rect 78692 22748 78698 22750
rect 52361 22747 52427 22748
rect 19568 22336 19888 22337
rect 0 22266 800 22296
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 3877 22266 3943 22269
rect 0 22264 3943 22266
rect 0 22208 3882 22264
rect 3938 22208 3943 22264
rect 0 22206 3943 22208
rect 0 22176 800 22206
rect 3877 22203 3943 22206
rect 21265 22130 21331 22133
rect 21398 22130 21404 22132
rect 21265 22128 21404 22130
rect 21265 22072 21270 22128
rect 21326 22072 21404 22128
rect 21265 22070 21404 22072
rect 21265 22067 21331 22070
rect 21398 22068 21404 22070
rect 21468 22068 21474 22132
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 0 21586 800 21616
rect 9489 21586 9555 21589
rect 0 21584 9555 21586
rect 0 21528 9494 21584
rect 9550 21528 9555 21584
rect 0 21526 9555 21528
rect 0 21496 800 21526
rect 9489 21523 9555 21526
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 0 21042 800 21072
rect 4061 21042 4127 21045
rect 0 21040 4127 21042
rect 0 20984 4066 21040
rect 4122 20984 4127 21040
rect 0 20982 4127 20984
rect 0 20952 800 20982
rect 4061 20979 4127 20982
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 0 20498 800 20528
rect 3325 20498 3391 20501
rect 0 20496 3391 20498
rect 0 20440 3330 20496
rect 3386 20440 3391 20496
rect 0 20438 3391 20440
rect 0 20408 800 20438
rect 3325 20435 3391 20438
rect 19568 20160 19888 20161
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 53833 20158 53899 20161
rect 53833 20156 54004 20158
rect 53833 20100 53838 20156
rect 53894 20100 54004 20156
rect 53833 20098 54004 20100
rect 53833 20095 53899 20098
rect 23473 20090 23539 20093
rect 23473 20088 27508 20090
rect 23473 20032 23478 20088
rect 23534 20032 27508 20088
rect 23473 20030 27508 20032
rect 23473 20027 23539 20030
rect 78806 20028 78812 20092
rect 78876 20090 78882 20092
rect 80881 20090 80947 20093
rect 78876 20088 81788 20090
rect 78876 20032 80886 20088
rect 80942 20032 81788 20088
rect 78876 20030 81788 20032
rect 78876 20028 78882 20030
rect 80881 20027 80947 20030
rect 0 19818 800 19848
rect 3141 19818 3207 19821
rect 0 19816 3207 19818
rect 0 19760 3146 19816
rect 3202 19760 3207 19816
rect 0 19758 3207 19760
rect 0 19728 800 19758
rect 3141 19755 3207 19758
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 0 19274 800 19304
rect 3325 19274 3391 19277
rect 0 19272 3391 19274
rect 0 19216 3330 19272
rect 3386 19216 3391 19272
rect 0 19214 3391 19216
rect 0 19184 800 19214
rect 3325 19211 3391 19214
rect 7097 19274 7163 19277
rect 8845 19274 8911 19277
rect 7097 19272 8911 19274
rect 7097 19216 7102 19272
rect 7158 19216 8850 19272
rect 8906 19216 8911 19272
rect 7097 19214 8911 19216
rect 7097 19211 7163 19214
rect 8845 19211 8911 19214
rect 7189 19138 7255 19141
rect 8477 19138 8543 19141
rect 7189 19136 8543 19138
rect 7189 19080 7194 19136
rect 7250 19080 8482 19136
rect 8538 19080 8543 19136
rect 7189 19078 8543 19080
rect 7189 19075 7255 19078
rect 8477 19075 8543 19078
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 19007 19888 19008
rect 0 18730 800 18760
rect 3877 18730 3943 18733
rect 0 18728 3943 18730
rect 0 18672 3882 18728
rect 3938 18672 3943 18728
rect 0 18670 3943 18672
rect 0 18640 800 18670
rect 3877 18667 3943 18670
rect 8109 18730 8175 18733
rect 8477 18730 8543 18733
rect 9121 18730 9187 18733
rect 9254 18730 9260 18732
rect 8109 18728 9260 18730
rect 8109 18672 8114 18728
rect 8170 18672 8482 18728
rect 8538 18672 9126 18728
rect 9182 18672 9260 18728
rect 8109 18670 9260 18672
rect 8109 18667 8175 18670
rect 8477 18667 8543 18670
rect 9121 18667 9187 18670
rect 9254 18668 9260 18670
rect 9324 18668 9330 18732
rect 78254 18668 78260 18732
rect 78324 18730 78330 18732
rect 79542 18730 79548 18732
rect 78324 18670 79548 18730
rect 78324 18668 78330 18670
rect 79542 18668 79548 18670
rect 79612 18668 79618 18732
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 0 18050 800 18080
rect 3693 18050 3759 18053
rect 9489 18052 9555 18053
rect 0 18048 3759 18050
rect 0 17992 3698 18048
rect 3754 17992 3759 18048
rect 0 17990 3759 17992
rect 0 17960 800 17990
rect 3693 17987 3759 17990
rect 9438 17988 9444 18052
rect 9508 18050 9555 18052
rect 9508 18048 9600 18050
rect 9550 17992 9600 18048
rect 9508 17990 9600 17992
rect 9508 17988 9555 17990
rect 9489 17987 9555 17988
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 78622 17716 78628 17780
rect 78692 17778 78698 17780
rect 79174 17778 79180 17780
rect 78692 17718 79180 17778
rect 78692 17716 78698 17718
rect 79174 17716 79180 17718
rect 79244 17716 79250 17780
rect 0 17506 800 17536
rect 3877 17506 3943 17509
rect 0 17504 3943 17506
rect 0 17448 3882 17504
rect 3938 17448 3943 17504
rect 0 17446 3943 17448
rect 0 17416 800 17446
rect 3877 17443 3943 17446
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 19149 17370 19215 17373
rect 19885 17370 19951 17373
rect 20110 17370 20116 17372
rect 19149 17368 20116 17370
rect 19149 17312 19154 17368
rect 19210 17312 19890 17368
rect 19946 17312 20116 17368
rect 19149 17310 20116 17312
rect 19149 17307 19215 17310
rect 19885 17307 19951 17310
rect 20110 17308 20116 17310
rect 20180 17308 20186 17372
rect 0 16962 800 16992
rect 2957 16962 3023 16965
rect 0 16960 3023 16962
rect 0 16904 2962 16960
rect 3018 16904 3023 16960
rect 0 16902 3023 16904
rect 0 16872 800 16902
rect 2957 16899 3023 16902
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 18505 16690 18571 16693
rect 18638 16690 18644 16692
rect 18505 16688 18644 16690
rect 18505 16632 18510 16688
rect 18566 16632 18644 16688
rect 18505 16630 18644 16632
rect 18505 16627 18571 16630
rect 18638 16628 18644 16630
rect 18708 16628 18714 16692
rect 4208 16352 4528 16353
rect 0 16282 800 16312
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 3693 16282 3759 16285
rect 0 16280 3759 16282
rect 0 16224 3698 16280
rect 3754 16224 3759 16280
rect 0 16222 3759 16224
rect 0 16192 800 16222
rect 3693 16219 3759 16222
rect 16389 16012 16455 16013
rect 16389 16010 16436 16012
rect 16344 16008 16436 16010
rect 16344 15952 16394 16008
rect 16344 15950 16436 15952
rect 16389 15948 16436 15950
rect 16500 15948 16506 16012
rect 79910 15948 79916 16012
rect 79980 16010 79986 16012
rect 81617 16010 81683 16013
rect 79980 16008 81683 16010
rect 79980 15952 81622 16008
rect 81678 15952 81683 16008
rect 79980 15950 81683 15952
rect 79980 15948 79986 15950
rect 16389 15947 16455 15948
rect 81617 15947 81683 15950
rect 19568 15808 19888 15809
rect 0 15738 800 15768
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 3601 15738 3667 15741
rect 0 15736 3667 15738
rect 0 15680 3606 15736
rect 3662 15680 3667 15736
rect 0 15678 3667 15680
rect 0 15648 800 15678
rect 3601 15675 3667 15678
rect 21909 15332 21975 15333
rect 21909 15330 21956 15332
rect 21864 15328 21956 15330
rect 21864 15272 21914 15328
rect 21864 15270 21956 15272
rect 21909 15268 21956 15270
rect 22020 15268 22026 15332
rect 21909 15267 21975 15268
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 0 15058 800 15088
rect 3877 15058 3943 15061
rect 0 15056 3943 15058
rect 0 15000 3882 15056
rect 3938 15000 3943 15056
rect 0 14998 3943 15000
rect 0 14968 800 14998
rect 3877 14995 3943 14998
rect 53833 14854 53899 14857
rect 81617 14854 81683 14857
rect 53833 14852 54004 14854
rect 53833 14796 53838 14852
rect 53894 14796 54004 14852
rect 53833 14794 54004 14796
rect 81617 14852 81788 14854
rect 81617 14796 81622 14852
rect 81678 14796 81788 14852
rect 81617 14794 81788 14796
rect 53833 14791 53899 14794
rect 81617 14791 81683 14794
rect 23381 14786 23447 14789
rect 23381 14784 27508 14786
rect 23381 14728 23386 14784
rect 23442 14728 27508 14784
rect 23381 14726 27508 14728
rect 23381 14723 23447 14726
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 13261 14650 13327 14653
rect 13670 14650 13676 14652
rect 13261 14648 13676 14650
rect 13261 14592 13266 14648
rect 13322 14592 13676 14648
rect 13261 14590 13676 14592
rect 13261 14587 13327 14590
rect 13670 14588 13676 14590
rect 13740 14588 13746 14652
rect 0 14514 800 14544
rect 8661 14514 8727 14517
rect 0 14512 8727 14514
rect 0 14456 8666 14512
rect 8722 14456 8727 14512
rect 0 14454 8727 14456
rect 0 14424 800 14454
rect 8661 14451 8727 14454
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 0 13970 800 14000
rect 3877 13970 3943 13973
rect 0 13968 3943 13970
rect 0 13912 3882 13968
rect 3938 13912 3943 13968
rect 0 13910 3943 13912
rect 0 13880 800 13910
rect 3877 13907 3943 13910
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 13567 19888 13568
rect 0 13290 800 13320
rect 4061 13290 4127 13293
rect 0 13288 4127 13290
rect 0 13232 4066 13288
rect 4122 13232 4127 13288
rect 0 13230 4127 13232
rect 0 13200 800 13230
rect 4061 13227 4127 13230
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 0 12746 800 12776
rect 3877 12746 3943 12749
rect 0 12744 3943 12746
rect 0 12688 3882 12744
rect 3938 12688 3943 12744
rect 0 12686 3943 12688
rect 0 12656 800 12686
rect 3877 12683 3943 12686
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 0 12202 800 12232
rect 7465 12202 7531 12205
rect 0 12200 7531 12202
rect 0 12144 7470 12200
rect 7526 12144 7531 12200
rect 0 12142 7531 12144
rect 0 12112 800 12142
rect 7465 12139 7531 12142
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 0 11522 800 11552
rect 3877 11522 3943 11525
rect 0 11520 3943 11522
rect 0 11464 3882 11520
rect 3938 11464 3943 11520
rect 0 11462 3943 11464
rect 0 11432 800 11462
rect 3877 11459 3943 11462
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 0 10978 800 11008
rect 0 10918 4124 10978
rect 0 10888 800 10918
rect 4064 10706 4124 10918
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 8017 10706 8083 10709
rect 4064 10704 8083 10706
rect 4064 10648 8022 10704
rect 8078 10648 8083 10704
rect 4064 10646 8083 10648
rect 8017 10643 8083 10646
rect 0 10434 800 10464
rect 3877 10434 3943 10437
rect 0 10432 3943 10434
rect 0 10376 3882 10432
rect 3938 10376 3943 10432
rect 0 10374 3943 10376
rect 0 10344 800 10374
rect 3877 10371 3943 10374
rect 19568 10368 19888 10369
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 8109 10026 8175 10029
rect 4064 10024 8175 10026
rect 4064 9968 8114 10024
rect 8170 9968 8175 10024
rect 4064 9966 8175 9968
rect 0 9754 800 9784
rect 4064 9754 4124 9966
rect 8109 9963 8175 9966
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 0 9694 4124 9754
rect 0 9664 800 9694
rect 19568 9280 19888 9281
rect 0 9210 800 9240
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 3877 9210 3943 9213
rect 0 9208 3943 9210
rect 0 9152 3882 9208
rect 3938 9152 3943 9208
rect 0 9150 3943 9152
rect 0 9120 800 9150
rect 3877 9147 3943 9150
rect 4208 8736 4528 8737
rect 0 8666 800 8696
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 4061 8666 4127 8669
rect 0 8664 4127 8666
rect 0 8608 4066 8664
rect 4122 8608 4127 8664
rect 0 8606 4127 8608
rect 0 8576 800 8606
rect 4061 8603 4127 8606
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 0 7986 800 8016
rect 3877 7986 3943 7989
rect 0 7984 3943 7986
rect 0 7928 3882 7984
rect 3938 7928 3943 7984
rect 0 7926 3943 7928
rect 0 7896 800 7926
rect 3877 7923 3943 7926
rect 4208 7648 4528 7649
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 0 7442 800 7472
rect 4061 7442 4127 7445
rect 0 7440 4127 7442
rect 0 7384 4066 7440
rect 4122 7384 4127 7440
rect 0 7382 4127 7384
rect 0 7352 800 7382
rect 4061 7379 4127 7382
rect 9765 7442 9831 7445
rect 13629 7442 13695 7445
rect 9765 7440 13695 7442
rect 9765 7384 9770 7440
rect 9826 7384 13634 7440
rect 13690 7384 13695 7440
rect 9765 7382 13695 7384
rect 9765 7379 9831 7382
rect 13629 7379 13695 7382
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 0 6762 800 6792
rect 3877 6762 3943 6765
rect 0 6760 3943 6762
rect 0 6704 3882 6760
rect 3938 6704 3943 6760
rect 0 6702 3943 6704
rect 0 6672 800 6702
rect 3877 6699 3943 6702
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 0 6218 800 6248
rect 4061 6218 4127 6221
rect 0 6216 4127 6218
rect 0 6160 4066 6216
rect 4122 6160 4127 6216
rect 0 6158 4127 6160
rect 0 6128 800 6158
rect 4061 6155 4127 6158
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 0 5674 800 5704
rect 3877 5674 3943 5677
rect 0 5672 3943 5674
rect 0 5616 3882 5672
rect 3938 5616 3943 5672
rect 0 5614 3943 5616
rect 0 5584 800 5614
rect 3877 5611 3943 5614
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 0 4994 800 5024
rect 4061 4994 4127 4997
rect 0 4992 4127 4994
rect 0 4936 4066 4992
rect 4122 4936 4127 4992
rect 0 4934 4127 4936
rect 0 4904 800 4934
rect 4061 4931 4127 4934
rect 19568 4928 19888 4929
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 23473 4858 23539 4861
rect 52085 4858 52151 4861
rect 79961 4858 80027 4861
rect 23473 4856 27508 4858
rect 23473 4800 23478 4856
rect 23534 4800 27508 4856
rect 23473 4798 27508 4800
rect 52085 4856 54004 4858
rect 52085 4800 52090 4856
rect 52146 4800 54004 4856
rect 52085 4798 54004 4800
rect 79961 4856 81788 4858
rect 79961 4800 79966 4856
rect 80022 4800 81788 4856
rect 79961 4798 81788 4800
rect 23473 4795 23539 4798
rect 52085 4795 52151 4798
rect 79961 4795 80027 4798
rect 0 4450 800 4480
rect 3877 4450 3943 4453
rect 0 4448 3943 4450
rect 0 4392 3882 4448
rect 3938 4392 3943 4448
rect 0 4390 3943 4392
rect 0 4360 800 4390
rect 3877 4387 3943 4390
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 0 3906 800 3936
rect 4061 3906 4127 3909
rect 0 3904 4127 3906
rect 0 3848 4066 3904
rect 4122 3848 4127 3904
rect 0 3846 4127 3848
rect 0 3816 800 3846
rect 4061 3843 4127 3846
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 4208 3296 4528 3297
rect 0 3226 800 3256
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 3877 3226 3943 3229
rect 0 3224 3943 3226
rect 0 3168 3882 3224
rect 3938 3168 3943 3224
rect 0 3166 3943 3168
rect 0 3136 800 3166
rect 3877 3163 3943 3166
rect 19568 2752 19888 2753
rect 0 2682 800 2712
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 2865 2682 2931 2685
rect 0 2680 2931 2682
rect 0 2624 2870 2680
rect 2926 2624 2931 2680
rect 0 2622 2931 2624
rect 0 2592 800 2622
rect 2865 2619 2931 2622
rect 4208 2208 4528 2209
rect 0 2138 800 2168
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 3509 2138 3575 2141
rect 0 2136 3575 2138
rect 0 2080 3514 2136
rect 3570 2080 3575 2136
rect 0 2078 3575 2080
rect 0 2048 800 2078
rect 3509 2075 3575 2078
rect 0 1458 800 1488
rect 2957 1458 3023 1461
rect 0 1456 3023 1458
rect 0 1400 2962 1456
rect 3018 1400 3023 1456
rect 0 1398 3023 1400
rect 0 1368 800 1398
rect 2957 1395 3023 1398
rect 0 914 800 944
rect 2773 914 2839 917
rect 0 912 2839 914
rect 0 856 2778 912
rect 2834 856 2839 912
rect 0 854 2839 856
rect 0 824 800 854
rect 2773 851 2839 854
rect 0 370 800 400
rect 2773 370 2839 373
rect 0 368 2839 370
rect 0 312 2778 368
rect 2834 312 2839 368
rect 0 310 2839 312
rect 0 280 800 310
rect 2773 307 2839 310
<< via3 >>
rect 19576 44092 19640 44096
rect 19576 44036 19580 44092
rect 19580 44036 19636 44092
rect 19636 44036 19640 44092
rect 19576 44032 19640 44036
rect 19656 44092 19720 44096
rect 19656 44036 19660 44092
rect 19660 44036 19716 44092
rect 19716 44036 19720 44092
rect 19656 44032 19720 44036
rect 19736 44092 19800 44096
rect 19736 44036 19740 44092
rect 19740 44036 19796 44092
rect 19796 44036 19800 44092
rect 19736 44032 19800 44036
rect 19816 44092 19880 44096
rect 19816 44036 19820 44092
rect 19820 44036 19876 44092
rect 19876 44036 19880 44092
rect 19816 44032 19880 44036
rect 50296 44092 50360 44096
rect 50296 44036 50300 44092
rect 50300 44036 50356 44092
rect 50356 44036 50360 44092
rect 50296 44032 50360 44036
rect 50376 44092 50440 44096
rect 50376 44036 50380 44092
rect 50380 44036 50436 44092
rect 50436 44036 50440 44092
rect 50376 44032 50440 44036
rect 50456 44092 50520 44096
rect 50456 44036 50460 44092
rect 50460 44036 50516 44092
rect 50516 44036 50520 44092
rect 50456 44032 50520 44036
rect 50536 44092 50600 44096
rect 50536 44036 50540 44092
rect 50540 44036 50596 44092
rect 50596 44036 50600 44092
rect 50536 44032 50600 44036
rect 81016 44092 81080 44096
rect 81016 44036 81020 44092
rect 81020 44036 81076 44092
rect 81076 44036 81080 44092
rect 81016 44032 81080 44036
rect 81096 44092 81160 44096
rect 81096 44036 81100 44092
rect 81100 44036 81156 44092
rect 81156 44036 81160 44092
rect 81096 44032 81160 44036
rect 81176 44092 81240 44096
rect 81176 44036 81180 44092
rect 81180 44036 81236 44092
rect 81236 44036 81240 44092
rect 81176 44032 81240 44036
rect 81256 44092 81320 44096
rect 81256 44036 81260 44092
rect 81260 44036 81316 44092
rect 81316 44036 81320 44092
rect 81256 44032 81320 44036
rect 4216 43548 4280 43552
rect 4216 43492 4220 43548
rect 4220 43492 4276 43548
rect 4276 43492 4280 43548
rect 4216 43488 4280 43492
rect 4296 43548 4360 43552
rect 4296 43492 4300 43548
rect 4300 43492 4356 43548
rect 4356 43492 4360 43548
rect 4296 43488 4360 43492
rect 4376 43548 4440 43552
rect 4376 43492 4380 43548
rect 4380 43492 4436 43548
rect 4436 43492 4440 43548
rect 4376 43488 4440 43492
rect 4456 43548 4520 43552
rect 4456 43492 4460 43548
rect 4460 43492 4516 43548
rect 4516 43492 4520 43548
rect 4456 43488 4520 43492
rect 34936 43548 35000 43552
rect 34936 43492 34940 43548
rect 34940 43492 34996 43548
rect 34996 43492 35000 43548
rect 34936 43488 35000 43492
rect 35016 43548 35080 43552
rect 35016 43492 35020 43548
rect 35020 43492 35076 43548
rect 35076 43492 35080 43548
rect 35016 43488 35080 43492
rect 35096 43548 35160 43552
rect 35096 43492 35100 43548
rect 35100 43492 35156 43548
rect 35156 43492 35160 43548
rect 35096 43488 35160 43492
rect 35176 43548 35240 43552
rect 35176 43492 35180 43548
rect 35180 43492 35236 43548
rect 35236 43492 35240 43548
rect 35176 43488 35240 43492
rect 65656 43548 65720 43552
rect 65656 43492 65660 43548
rect 65660 43492 65716 43548
rect 65716 43492 65720 43548
rect 65656 43488 65720 43492
rect 65736 43548 65800 43552
rect 65736 43492 65740 43548
rect 65740 43492 65796 43548
rect 65796 43492 65800 43548
rect 65736 43488 65800 43492
rect 65816 43548 65880 43552
rect 65816 43492 65820 43548
rect 65820 43492 65876 43548
rect 65876 43492 65880 43548
rect 65816 43488 65880 43492
rect 65896 43548 65960 43552
rect 65896 43492 65900 43548
rect 65900 43492 65956 43548
rect 65956 43492 65960 43548
rect 65896 43488 65960 43492
rect 96376 43548 96440 43552
rect 96376 43492 96380 43548
rect 96380 43492 96436 43548
rect 96436 43492 96440 43548
rect 96376 43488 96440 43492
rect 96456 43548 96520 43552
rect 96456 43492 96460 43548
rect 96460 43492 96516 43548
rect 96516 43492 96520 43548
rect 96456 43488 96520 43492
rect 96536 43548 96600 43552
rect 96536 43492 96540 43548
rect 96540 43492 96596 43548
rect 96596 43492 96600 43548
rect 96536 43488 96600 43492
rect 96616 43548 96680 43552
rect 96616 43492 96620 43548
rect 96620 43492 96676 43548
rect 96676 43492 96680 43548
rect 96616 43488 96680 43492
rect 19576 43004 19640 43008
rect 19576 42948 19580 43004
rect 19580 42948 19636 43004
rect 19636 42948 19640 43004
rect 19576 42944 19640 42948
rect 19656 43004 19720 43008
rect 19656 42948 19660 43004
rect 19660 42948 19716 43004
rect 19716 42948 19720 43004
rect 19656 42944 19720 42948
rect 19736 43004 19800 43008
rect 19736 42948 19740 43004
rect 19740 42948 19796 43004
rect 19796 42948 19800 43004
rect 19736 42944 19800 42948
rect 19816 43004 19880 43008
rect 19816 42948 19820 43004
rect 19820 42948 19876 43004
rect 19876 42948 19880 43004
rect 19816 42944 19880 42948
rect 50296 43004 50360 43008
rect 50296 42948 50300 43004
rect 50300 42948 50356 43004
rect 50356 42948 50360 43004
rect 50296 42944 50360 42948
rect 50376 43004 50440 43008
rect 50376 42948 50380 43004
rect 50380 42948 50436 43004
rect 50436 42948 50440 43004
rect 50376 42944 50440 42948
rect 50456 43004 50520 43008
rect 50456 42948 50460 43004
rect 50460 42948 50516 43004
rect 50516 42948 50520 43004
rect 50456 42944 50520 42948
rect 50536 43004 50600 43008
rect 50536 42948 50540 43004
rect 50540 42948 50596 43004
rect 50596 42948 50600 43004
rect 50536 42944 50600 42948
rect 81016 43004 81080 43008
rect 81016 42948 81020 43004
rect 81020 42948 81076 43004
rect 81076 42948 81080 43004
rect 81016 42944 81080 42948
rect 81096 43004 81160 43008
rect 81096 42948 81100 43004
rect 81100 42948 81156 43004
rect 81156 42948 81160 43004
rect 81096 42944 81160 42948
rect 81176 43004 81240 43008
rect 81176 42948 81180 43004
rect 81180 42948 81236 43004
rect 81236 42948 81240 43004
rect 81176 42944 81240 42948
rect 81256 43004 81320 43008
rect 81256 42948 81260 43004
rect 81260 42948 81316 43004
rect 81316 42948 81320 43004
rect 81256 42944 81320 42948
rect 4216 42460 4280 42464
rect 4216 42404 4220 42460
rect 4220 42404 4276 42460
rect 4276 42404 4280 42460
rect 4216 42400 4280 42404
rect 4296 42460 4360 42464
rect 4296 42404 4300 42460
rect 4300 42404 4356 42460
rect 4356 42404 4360 42460
rect 4296 42400 4360 42404
rect 4376 42460 4440 42464
rect 4376 42404 4380 42460
rect 4380 42404 4436 42460
rect 4436 42404 4440 42460
rect 4376 42400 4440 42404
rect 4456 42460 4520 42464
rect 4456 42404 4460 42460
rect 4460 42404 4516 42460
rect 4516 42404 4520 42460
rect 4456 42400 4520 42404
rect 34936 42460 35000 42464
rect 34936 42404 34940 42460
rect 34940 42404 34996 42460
rect 34996 42404 35000 42460
rect 34936 42400 35000 42404
rect 35016 42460 35080 42464
rect 35016 42404 35020 42460
rect 35020 42404 35076 42460
rect 35076 42404 35080 42460
rect 35016 42400 35080 42404
rect 35096 42460 35160 42464
rect 35096 42404 35100 42460
rect 35100 42404 35156 42460
rect 35156 42404 35160 42460
rect 35096 42400 35160 42404
rect 35176 42460 35240 42464
rect 35176 42404 35180 42460
rect 35180 42404 35236 42460
rect 35236 42404 35240 42460
rect 35176 42400 35240 42404
rect 65656 42460 65720 42464
rect 65656 42404 65660 42460
rect 65660 42404 65716 42460
rect 65716 42404 65720 42460
rect 65656 42400 65720 42404
rect 65736 42460 65800 42464
rect 65736 42404 65740 42460
rect 65740 42404 65796 42460
rect 65796 42404 65800 42460
rect 65736 42400 65800 42404
rect 65816 42460 65880 42464
rect 65816 42404 65820 42460
rect 65820 42404 65876 42460
rect 65876 42404 65880 42460
rect 65816 42400 65880 42404
rect 65896 42460 65960 42464
rect 65896 42404 65900 42460
rect 65900 42404 65956 42460
rect 65956 42404 65960 42460
rect 65896 42400 65960 42404
rect 96376 42460 96440 42464
rect 96376 42404 96380 42460
rect 96380 42404 96436 42460
rect 96436 42404 96440 42460
rect 96376 42400 96440 42404
rect 96456 42460 96520 42464
rect 96456 42404 96460 42460
rect 96460 42404 96516 42460
rect 96516 42404 96520 42460
rect 96456 42400 96520 42404
rect 96536 42460 96600 42464
rect 96536 42404 96540 42460
rect 96540 42404 96596 42460
rect 96596 42404 96600 42460
rect 96536 42400 96600 42404
rect 96616 42460 96680 42464
rect 96616 42404 96620 42460
rect 96620 42404 96676 42460
rect 96676 42404 96680 42460
rect 96616 42400 96680 42404
rect 19576 41916 19640 41920
rect 19576 41860 19580 41916
rect 19580 41860 19636 41916
rect 19636 41860 19640 41916
rect 19576 41856 19640 41860
rect 19656 41916 19720 41920
rect 19656 41860 19660 41916
rect 19660 41860 19716 41916
rect 19716 41860 19720 41916
rect 19656 41856 19720 41860
rect 19736 41916 19800 41920
rect 19736 41860 19740 41916
rect 19740 41860 19796 41916
rect 19796 41860 19800 41916
rect 19736 41856 19800 41860
rect 19816 41916 19880 41920
rect 19816 41860 19820 41916
rect 19820 41860 19876 41916
rect 19876 41860 19880 41916
rect 19816 41856 19880 41860
rect 50296 41916 50360 41920
rect 50296 41860 50300 41916
rect 50300 41860 50356 41916
rect 50356 41860 50360 41916
rect 50296 41856 50360 41860
rect 50376 41916 50440 41920
rect 50376 41860 50380 41916
rect 50380 41860 50436 41916
rect 50436 41860 50440 41916
rect 50376 41856 50440 41860
rect 50456 41916 50520 41920
rect 50456 41860 50460 41916
rect 50460 41860 50516 41916
rect 50516 41860 50520 41916
rect 50456 41856 50520 41860
rect 50536 41916 50600 41920
rect 50536 41860 50540 41916
rect 50540 41860 50596 41916
rect 50596 41860 50600 41916
rect 50536 41856 50600 41860
rect 81016 41916 81080 41920
rect 81016 41860 81020 41916
rect 81020 41860 81076 41916
rect 81076 41860 81080 41916
rect 81016 41856 81080 41860
rect 81096 41916 81160 41920
rect 81096 41860 81100 41916
rect 81100 41860 81156 41916
rect 81156 41860 81160 41916
rect 81096 41856 81160 41860
rect 81176 41916 81240 41920
rect 81176 41860 81180 41916
rect 81180 41860 81236 41916
rect 81236 41860 81240 41916
rect 81176 41856 81240 41860
rect 81256 41916 81320 41920
rect 81256 41860 81260 41916
rect 81260 41860 81316 41916
rect 81316 41860 81320 41916
rect 81256 41856 81320 41860
rect 4216 41372 4280 41376
rect 4216 41316 4220 41372
rect 4220 41316 4276 41372
rect 4276 41316 4280 41372
rect 4216 41312 4280 41316
rect 4296 41372 4360 41376
rect 4296 41316 4300 41372
rect 4300 41316 4356 41372
rect 4356 41316 4360 41372
rect 4296 41312 4360 41316
rect 4376 41372 4440 41376
rect 4376 41316 4380 41372
rect 4380 41316 4436 41372
rect 4436 41316 4440 41372
rect 4376 41312 4440 41316
rect 4456 41372 4520 41376
rect 4456 41316 4460 41372
rect 4460 41316 4516 41372
rect 4516 41316 4520 41372
rect 4456 41312 4520 41316
rect 34936 41372 35000 41376
rect 34936 41316 34940 41372
rect 34940 41316 34996 41372
rect 34996 41316 35000 41372
rect 34936 41312 35000 41316
rect 35016 41372 35080 41376
rect 35016 41316 35020 41372
rect 35020 41316 35076 41372
rect 35076 41316 35080 41372
rect 35016 41312 35080 41316
rect 35096 41372 35160 41376
rect 35096 41316 35100 41372
rect 35100 41316 35156 41372
rect 35156 41316 35160 41372
rect 35096 41312 35160 41316
rect 35176 41372 35240 41376
rect 35176 41316 35180 41372
rect 35180 41316 35236 41372
rect 35236 41316 35240 41372
rect 35176 41312 35240 41316
rect 65656 41372 65720 41376
rect 65656 41316 65660 41372
rect 65660 41316 65716 41372
rect 65716 41316 65720 41372
rect 65656 41312 65720 41316
rect 65736 41372 65800 41376
rect 65736 41316 65740 41372
rect 65740 41316 65796 41372
rect 65796 41316 65800 41372
rect 65736 41312 65800 41316
rect 65816 41372 65880 41376
rect 65816 41316 65820 41372
rect 65820 41316 65876 41372
rect 65876 41316 65880 41372
rect 65816 41312 65880 41316
rect 65896 41372 65960 41376
rect 65896 41316 65900 41372
rect 65900 41316 65956 41372
rect 65956 41316 65960 41372
rect 65896 41312 65960 41316
rect 96376 41372 96440 41376
rect 96376 41316 96380 41372
rect 96380 41316 96436 41372
rect 96436 41316 96440 41372
rect 96376 41312 96440 41316
rect 96456 41372 96520 41376
rect 96456 41316 96460 41372
rect 96460 41316 96516 41372
rect 96516 41316 96520 41372
rect 96456 41312 96520 41316
rect 96536 41372 96600 41376
rect 96536 41316 96540 41372
rect 96540 41316 96596 41372
rect 96596 41316 96600 41372
rect 96536 41312 96600 41316
rect 96616 41372 96680 41376
rect 96616 41316 96620 41372
rect 96620 41316 96676 41372
rect 96676 41316 96680 41372
rect 96616 41312 96680 41316
rect 19576 40828 19640 40832
rect 19576 40772 19580 40828
rect 19580 40772 19636 40828
rect 19636 40772 19640 40828
rect 19576 40768 19640 40772
rect 19656 40828 19720 40832
rect 19656 40772 19660 40828
rect 19660 40772 19716 40828
rect 19716 40772 19720 40828
rect 19656 40768 19720 40772
rect 19736 40828 19800 40832
rect 19736 40772 19740 40828
rect 19740 40772 19796 40828
rect 19796 40772 19800 40828
rect 19736 40768 19800 40772
rect 19816 40828 19880 40832
rect 19816 40772 19820 40828
rect 19820 40772 19876 40828
rect 19876 40772 19880 40828
rect 19816 40768 19880 40772
rect 50296 40828 50360 40832
rect 50296 40772 50300 40828
rect 50300 40772 50356 40828
rect 50356 40772 50360 40828
rect 50296 40768 50360 40772
rect 50376 40828 50440 40832
rect 50376 40772 50380 40828
rect 50380 40772 50436 40828
rect 50436 40772 50440 40828
rect 50376 40768 50440 40772
rect 50456 40828 50520 40832
rect 50456 40772 50460 40828
rect 50460 40772 50516 40828
rect 50516 40772 50520 40828
rect 50456 40768 50520 40772
rect 50536 40828 50600 40832
rect 50536 40772 50540 40828
rect 50540 40772 50596 40828
rect 50596 40772 50600 40828
rect 50536 40768 50600 40772
rect 81016 40828 81080 40832
rect 81016 40772 81020 40828
rect 81020 40772 81076 40828
rect 81076 40772 81080 40828
rect 81016 40768 81080 40772
rect 81096 40828 81160 40832
rect 81096 40772 81100 40828
rect 81100 40772 81156 40828
rect 81156 40772 81160 40828
rect 81096 40768 81160 40772
rect 81176 40828 81240 40832
rect 81176 40772 81180 40828
rect 81180 40772 81236 40828
rect 81236 40772 81240 40828
rect 81176 40768 81240 40772
rect 81256 40828 81320 40832
rect 81256 40772 81260 40828
rect 81260 40772 81316 40828
rect 81316 40772 81320 40828
rect 81256 40768 81320 40772
rect 4216 40284 4280 40288
rect 4216 40228 4220 40284
rect 4220 40228 4276 40284
rect 4276 40228 4280 40284
rect 4216 40224 4280 40228
rect 4296 40284 4360 40288
rect 4296 40228 4300 40284
rect 4300 40228 4356 40284
rect 4356 40228 4360 40284
rect 4296 40224 4360 40228
rect 4376 40284 4440 40288
rect 4376 40228 4380 40284
rect 4380 40228 4436 40284
rect 4436 40228 4440 40284
rect 4376 40224 4440 40228
rect 4456 40284 4520 40288
rect 4456 40228 4460 40284
rect 4460 40228 4516 40284
rect 4516 40228 4520 40284
rect 4456 40224 4520 40228
rect 34936 40284 35000 40288
rect 34936 40228 34940 40284
rect 34940 40228 34996 40284
rect 34996 40228 35000 40284
rect 34936 40224 35000 40228
rect 35016 40284 35080 40288
rect 35016 40228 35020 40284
rect 35020 40228 35076 40284
rect 35076 40228 35080 40284
rect 35016 40224 35080 40228
rect 35096 40284 35160 40288
rect 35096 40228 35100 40284
rect 35100 40228 35156 40284
rect 35156 40228 35160 40284
rect 35096 40224 35160 40228
rect 35176 40284 35240 40288
rect 35176 40228 35180 40284
rect 35180 40228 35236 40284
rect 35236 40228 35240 40284
rect 35176 40224 35240 40228
rect 65656 40284 65720 40288
rect 65656 40228 65660 40284
rect 65660 40228 65716 40284
rect 65716 40228 65720 40284
rect 65656 40224 65720 40228
rect 65736 40284 65800 40288
rect 65736 40228 65740 40284
rect 65740 40228 65796 40284
rect 65796 40228 65800 40284
rect 65736 40224 65800 40228
rect 65816 40284 65880 40288
rect 65816 40228 65820 40284
rect 65820 40228 65876 40284
rect 65876 40228 65880 40284
rect 65816 40224 65880 40228
rect 65896 40284 65960 40288
rect 65896 40228 65900 40284
rect 65900 40228 65956 40284
rect 65956 40228 65960 40284
rect 65896 40224 65960 40228
rect 96376 40284 96440 40288
rect 96376 40228 96380 40284
rect 96380 40228 96436 40284
rect 96436 40228 96440 40284
rect 96376 40224 96440 40228
rect 96456 40284 96520 40288
rect 96456 40228 96460 40284
rect 96460 40228 96516 40284
rect 96516 40228 96520 40284
rect 96456 40224 96520 40228
rect 96536 40284 96600 40288
rect 96536 40228 96540 40284
rect 96540 40228 96596 40284
rect 96596 40228 96600 40284
rect 96536 40224 96600 40228
rect 96616 40284 96680 40288
rect 96616 40228 96620 40284
rect 96620 40228 96676 40284
rect 96676 40228 96680 40284
rect 96616 40224 96680 40228
rect 19576 39740 19640 39744
rect 19576 39684 19580 39740
rect 19580 39684 19636 39740
rect 19636 39684 19640 39740
rect 19576 39680 19640 39684
rect 19656 39740 19720 39744
rect 19656 39684 19660 39740
rect 19660 39684 19716 39740
rect 19716 39684 19720 39740
rect 19656 39680 19720 39684
rect 19736 39740 19800 39744
rect 19736 39684 19740 39740
rect 19740 39684 19796 39740
rect 19796 39684 19800 39740
rect 19736 39680 19800 39684
rect 19816 39740 19880 39744
rect 19816 39684 19820 39740
rect 19820 39684 19876 39740
rect 19876 39684 19880 39740
rect 19816 39680 19880 39684
rect 50296 39740 50360 39744
rect 50296 39684 50300 39740
rect 50300 39684 50356 39740
rect 50356 39684 50360 39740
rect 50296 39680 50360 39684
rect 50376 39740 50440 39744
rect 50376 39684 50380 39740
rect 50380 39684 50436 39740
rect 50436 39684 50440 39740
rect 50376 39680 50440 39684
rect 50456 39740 50520 39744
rect 50456 39684 50460 39740
rect 50460 39684 50516 39740
rect 50516 39684 50520 39740
rect 50456 39680 50520 39684
rect 50536 39740 50600 39744
rect 50536 39684 50540 39740
rect 50540 39684 50596 39740
rect 50596 39684 50600 39740
rect 50536 39680 50600 39684
rect 81016 39740 81080 39744
rect 81016 39684 81020 39740
rect 81020 39684 81076 39740
rect 81076 39684 81080 39740
rect 81016 39680 81080 39684
rect 81096 39740 81160 39744
rect 81096 39684 81100 39740
rect 81100 39684 81156 39740
rect 81156 39684 81160 39740
rect 81096 39680 81160 39684
rect 81176 39740 81240 39744
rect 81176 39684 81180 39740
rect 81180 39684 81236 39740
rect 81236 39684 81240 39740
rect 81176 39680 81240 39684
rect 81256 39740 81320 39744
rect 81256 39684 81260 39740
rect 81260 39684 81316 39740
rect 81316 39684 81320 39740
rect 81256 39680 81320 39684
rect 28948 39612 29012 39676
rect 28948 39340 29012 39404
rect 4216 39196 4280 39200
rect 4216 39140 4220 39196
rect 4220 39140 4276 39196
rect 4276 39140 4280 39196
rect 4216 39136 4280 39140
rect 4296 39196 4360 39200
rect 4296 39140 4300 39196
rect 4300 39140 4356 39196
rect 4356 39140 4360 39196
rect 4296 39136 4360 39140
rect 4376 39196 4440 39200
rect 4376 39140 4380 39196
rect 4380 39140 4436 39196
rect 4436 39140 4440 39196
rect 4376 39136 4440 39140
rect 4456 39196 4520 39200
rect 4456 39140 4460 39196
rect 4460 39140 4516 39196
rect 4516 39140 4520 39196
rect 4456 39136 4520 39140
rect 34936 39196 35000 39200
rect 34936 39140 34940 39196
rect 34940 39140 34996 39196
rect 34996 39140 35000 39196
rect 34936 39136 35000 39140
rect 35016 39196 35080 39200
rect 35016 39140 35020 39196
rect 35020 39140 35076 39196
rect 35076 39140 35080 39196
rect 35016 39136 35080 39140
rect 35096 39196 35160 39200
rect 35096 39140 35100 39196
rect 35100 39140 35156 39196
rect 35156 39140 35160 39196
rect 35096 39136 35160 39140
rect 35176 39196 35240 39200
rect 35176 39140 35180 39196
rect 35180 39140 35236 39196
rect 35236 39140 35240 39196
rect 35176 39136 35240 39140
rect 65656 39196 65720 39200
rect 65656 39140 65660 39196
rect 65660 39140 65716 39196
rect 65716 39140 65720 39196
rect 65656 39136 65720 39140
rect 65736 39196 65800 39200
rect 65736 39140 65740 39196
rect 65740 39140 65796 39196
rect 65796 39140 65800 39196
rect 65736 39136 65800 39140
rect 65816 39196 65880 39200
rect 65816 39140 65820 39196
rect 65820 39140 65876 39196
rect 65876 39140 65880 39196
rect 65816 39136 65880 39140
rect 65896 39196 65960 39200
rect 65896 39140 65900 39196
rect 65900 39140 65956 39196
rect 65956 39140 65960 39196
rect 65896 39136 65960 39140
rect 96376 39196 96440 39200
rect 96376 39140 96380 39196
rect 96380 39140 96436 39196
rect 96436 39140 96440 39196
rect 96376 39136 96440 39140
rect 96456 39196 96520 39200
rect 96456 39140 96460 39196
rect 96460 39140 96516 39196
rect 96516 39140 96520 39196
rect 96456 39136 96520 39140
rect 96536 39196 96600 39200
rect 96536 39140 96540 39196
rect 96540 39140 96596 39196
rect 96596 39140 96600 39196
rect 96536 39136 96600 39140
rect 96616 39196 96680 39200
rect 96616 39140 96620 39196
rect 96620 39140 96676 39196
rect 96676 39140 96680 39196
rect 96616 39136 96680 39140
rect 19576 38652 19640 38656
rect 19576 38596 19580 38652
rect 19580 38596 19636 38652
rect 19636 38596 19640 38652
rect 19576 38592 19640 38596
rect 19656 38652 19720 38656
rect 19656 38596 19660 38652
rect 19660 38596 19716 38652
rect 19716 38596 19720 38652
rect 19656 38592 19720 38596
rect 19736 38652 19800 38656
rect 19736 38596 19740 38652
rect 19740 38596 19796 38652
rect 19796 38596 19800 38652
rect 19736 38592 19800 38596
rect 19816 38652 19880 38656
rect 19816 38596 19820 38652
rect 19820 38596 19876 38652
rect 19876 38596 19880 38652
rect 19816 38592 19880 38596
rect 50296 38652 50360 38656
rect 50296 38596 50300 38652
rect 50300 38596 50356 38652
rect 50356 38596 50360 38652
rect 50296 38592 50360 38596
rect 50376 38652 50440 38656
rect 50376 38596 50380 38652
rect 50380 38596 50436 38652
rect 50436 38596 50440 38652
rect 50376 38592 50440 38596
rect 50456 38652 50520 38656
rect 50456 38596 50460 38652
rect 50460 38596 50516 38652
rect 50516 38596 50520 38652
rect 50456 38592 50520 38596
rect 50536 38652 50600 38656
rect 50536 38596 50540 38652
rect 50540 38596 50596 38652
rect 50596 38596 50600 38652
rect 50536 38592 50600 38596
rect 81016 38652 81080 38656
rect 81016 38596 81020 38652
rect 81020 38596 81076 38652
rect 81076 38596 81080 38652
rect 81016 38592 81080 38596
rect 81096 38652 81160 38656
rect 81096 38596 81100 38652
rect 81100 38596 81156 38652
rect 81156 38596 81160 38652
rect 81096 38592 81160 38596
rect 81176 38652 81240 38656
rect 81176 38596 81180 38652
rect 81180 38596 81236 38652
rect 81236 38596 81240 38652
rect 81176 38592 81240 38596
rect 81256 38652 81320 38656
rect 81256 38596 81260 38652
rect 81260 38596 81316 38652
rect 81316 38596 81320 38652
rect 81256 38592 81320 38596
rect 4216 38108 4280 38112
rect 4216 38052 4220 38108
rect 4220 38052 4276 38108
rect 4276 38052 4280 38108
rect 4216 38048 4280 38052
rect 4296 38108 4360 38112
rect 4296 38052 4300 38108
rect 4300 38052 4356 38108
rect 4356 38052 4360 38108
rect 4296 38048 4360 38052
rect 4376 38108 4440 38112
rect 4376 38052 4380 38108
rect 4380 38052 4436 38108
rect 4436 38052 4440 38108
rect 4376 38048 4440 38052
rect 4456 38108 4520 38112
rect 4456 38052 4460 38108
rect 4460 38052 4516 38108
rect 4516 38052 4520 38108
rect 4456 38048 4520 38052
rect 34936 38108 35000 38112
rect 34936 38052 34940 38108
rect 34940 38052 34996 38108
rect 34996 38052 35000 38108
rect 34936 38048 35000 38052
rect 35016 38108 35080 38112
rect 35016 38052 35020 38108
rect 35020 38052 35076 38108
rect 35076 38052 35080 38108
rect 35016 38048 35080 38052
rect 35096 38108 35160 38112
rect 35096 38052 35100 38108
rect 35100 38052 35156 38108
rect 35156 38052 35160 38108
rect 35096 38048 35160 38052
rect 35176 38108 35240 38112
rect 35176 38052 35180 38108
rect 35180 38052 35236 38108
rect 35236 38052 35240 38108
rect 35176 38048 35240 38052
rect 65656 38108 65720 38112
rect 65656 38052 65660 38108
rect 65660 38052 65716 38108
rect 65716 38052 65720 38108
rect 65656 38048 65720 38052
rect 65736 38108 65800 38112
rect 65736 38052 65740 38108
rect 65740 38052 65796 38108
rect 65796 38052 65800 38108
rect 65736 38048 65800 38052
rect 65816 38108 65880 38112
rect 65816 38052 65820 38108
rect 65820 38052 65876 38108
rect 65876 38052 65880 38108
rect 65816 38048 65880 38052
rect 65896 38108 65960 38112
rect 65896 38052 65900 38108
rect 65900 38052 65956 38108
rect 65956 38052 65960 38108
rect 65896 38048 65960 38052
rect 96376 38108 96440 38112
rect 96376 38052 96380 38108
rect 96380 38052 96436 38108
rect 96436 38052 96440 38108
rect 96376 38048 96440 38052
rect 96456 38108 96520 38112
rect 96456 38052 96460 38108
rect 96460 38052 96516 38108
rect 96516 38052 96520 38108
rect 96456 38048 96520 38052
rect 96536 38108 96600 38112
rect 96536 38052 96540 38108
rect 96540 38052 96596 38108
rect 96596 38052 96600 38108
rect 96536 38048 96600 38052
rect 96616 38108 96680 38112
rect 96616 38052 96620 38108
rect 96620 38052 96676 38108
rect 96676 38052 96680 38108
rect 96616 38048 96680 38052
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 50296 37564 50360 37568
rect 50296 37508 50300 37564
rect 50300 37508 50356 37564
rect 50356 37508 50360 37564
rect 50296 37504 50360 37508
rect 50376 37564 50440 37568
rect 50376 37508 50380 37564
rect 50380 37508 50436 37564
rect 50436 37508 50440 37564
rect 50376 37504 50440 37508
rect 50456 37564 50520 37568
rect 50456 37508 50460 37564
rect 50460 37508 50516 37564
rect 50516 37508 50520 37564
rect 50456 37504 50520 37508
rect 50536 37564 50600 37568
rect 50536 37508 50540 37564
rect 50540 37508 50596 37564
rect 50596 37508 50600 37564
rect 50536 37504 50600 37508
rect 81016 37564 81080 37568
rect 81016 37508 81020 37564
rect 81020 37508 81076 37564
rect 81076 37508 81080 37564
rect 81016 37504 81080 37508
rect 81096 37564 81160 37568
rect 81096 37508 81100 37564
rect 81100 37508 81156 37564
rect 81156 37508 81160 37564
rect 81096 37504 81160 37508
rect 81176 37564 81240 37568
rect 81176 37508 81180 37564
rect 81180 37508 81236 37564
rect 81236 37508 81240 37564
rect 81176 37504 81240 37508
rect 81256 37564 81320 37568
rect 81256 37508 81260 37564
rect 81260 37508 81316 37564
rect 81316 37508 81320 37564
rect 81256 37504 81320 37508
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 65656 37020 65720 37024
rect 65656 36964 65660 37020
rect 65660 36964 65716 37020
rect 65716 36964 65720 37020
rect 65656 36960 65720 36964
rect 65736 37020 65800 37024
rect 65736 36964 65740 37020
rect 65740 36964 65796 37020
rect 65796 36964 65800 37020
rect 65736 36960 65800 36964
rect 65816 37020 65880 37024
rect 65816 36964 65820 37020
rect 65820 36964 65876 37020
rect 65876 36964 65880 37020
rect 65816 36960 65880 36964
rect 65896 37020 65960 37024
rect 65896 36964 65900 37020
rect 65900 36964 65956 37020
rect 65956 36964 65960 37020
rect 65896 36960 65960 36964
rect 96376 37020 96440 37024
rect 96376 36964 96380 37020
rect 96380 36964 96436 37020
rect 96436 36964 96440 37020
rect 96376 36960 96440 36964
rect 96456 37020 96520 37024
rect 96456 36964 96460 37020
rect 96460 36964 96516 37020
rect 96516 36964 96520 37020
rect 96456 36960 96520 36964
rect 96536 37020 96600 37024
rect 96536 36964 96540 37020
rect 96540 36964 96596 37020
rect 96596 36964 96600 37020
rect 96536 36960 96600 36964
rect 96616 37020 96680 37024
rect 96616 36964 96620 37020
rect 96620 36964 96676 37020
rect 96676 36964 96680 37020
rect 96616 36960 96680 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 50296 36476 50360 36480
rect 50296 36420 50300 36476
rect 50300 36420 50356 36476
rect 50356 36420 50360 36476
rect 50296 36416 50360 36420
rect 50376 36476 50440 36480
rect 50376 36420 50380 36476
rect 50380 36420 50436 36476
rect 50436 36420 50440 36476
rect 50376 36416 50440 36420
rect 50456 36476 50520 36480
rect 50456 36420 50460 36476
rect 50460 36420 50516 36476
rect 50516 36420 50520 36476
rect 50456 36416 50520 36420
rect 50536 36476 50600 36480
rect 50536 36420 50540 36476
rect 50540 36420 50596 36476
rect 50596 36420 50600 36476
rect 50536 36416 50600 36420
rect 81016 36476 81080 36480
rect 81016 36420 81020 36476
rect 81020 36420 81076 36476
rect 81076 36420 81080 36476
rect 81016 36416 81080 36420
rect 81096 36476 81160 36480
rect 81096 36420 81100 36476
rect 81100 36420 81156 36476
rect 81156 36420 81160 36476
rect 81096 36416 81160 36420
rect 81176 36476 81240 36480
rect 81176 36420 81180 36476
rect 81180 36420 81236 36476
rect 81236 36420 81240 36476
rect 81176 36416 81240 36420
rect 81256 36476 81320 36480
rect 81256 36420 81260 36476
rect 81260 36420 81316 36476
rect 81316 36420 81320 36476
rect 81256 36416 81320 36420
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 65656 35932 65720 35936
rect 65656 35876 65660 35932
rect 65660 35876 65716 35932
rect 65716 35876 65720 35932
rect 65656 35872 65720 35876
rect 65736 35932 65800 35936
rect 65736 35876 65740 35932
rect 65740 35876 65796 35932
rect 65796 35876 65800 35932
rect 65736 35872 65800 35876
rect 65816 35932 65880 35936
rect 65816 35876 65820 35932
rect 65820 35876 65876 35932
rect 65876 35876 65880 35932
rect 65816 35872 65880 35876
rect 65896 35932 65960 35936
rect 65896 35876 65900 35932
rect 65900 35876 65956 35932
rect 65956 35876 65960 35932
rect 65896 35872 65960 35876
rect 96376 35932 96440 35936
rect 96376 35876 96380 35932
rect 96380 35876 96436 35932
rect 96436 35876 96440 35932
rect 96376 35872 96440 35876
rect 96456 35932 96520 35936
rect 96456 35876 96460 35932
rect 96460 35876 96516 35932
rect 96516 35876 96520 35932
rect 96456 35872 96520 35876
rect 96536 35932 96600 35936
rect 96536 35876 96540 35932
rect 96540 35876 96596 35932
rect 96596 35876 96600 35932
rect 96536 35872 96600 35876
rect 96616 35932 96680 35936
rect 96616 35876 96620 35932
rect 96620 35876 96676 35932
rect 96676 35876 96680 35932
rect 96616 35872 96680 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 50296 35388 50360 35392
rect 50296 35332 50300 35388
rect 50300 35332 50356 35388
rect 50356 35332 50360 35388
rect 50296 35328 50360 35332
rect 50376 35388 50440 35392
rect 50376 35332 50380 35388
rect 50380 35332 50436 35388
rect 50436 35332 50440 35388
rect 50376 35328 50440 35332
rect 50456 35388 50520 35392
rect 50456 35332 50460 35388
rect 50460 35332 50516 35388
rect 50516 35332 50520 35388
rect 50456 35328 50520 35332
rect 50536 35388 50600 35392
rect 50536 35332 50540 35388
rect 50540 35332 50596 35388
rect 50596 35332 50600 35388
rect 50536 35328 50600 35332
rect 81016 35388 81080 35392
rect 81016 35332 81020 35388
rect 81020 35332 81076 35388
rect 81076 35332 81080 35388
rect 81016 35328 81080 35332
rect 81096 35388 81160 35392
rect 81096 35332 81100 35388
rect 81100 35332 81156 35388
rect 81156 35332 81160 35388
rect 81096 35328 81160 35332
rect 81176 35388 81240 35392
rect 81176 35332 81180 35388
rect 81180 35332 81236 35388
rect 81236 35332 81240 35388
rect 81176 35328 81240 35332
rect 81256 35388 81320 35392
rect 81256 35332 81260 35388
rect 81260 35332 81316 35388
rect 81316 35332 81320 35388
rect 81256 35328 81320 35332
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 65656 34844 65720 34848
rect 65656 34788 65660 34844
rect 65660 34788 65716 34844
rect 65716 34788 65720 34844
rect 65656 34784 65720 34788
rect 65736 34844 65800 34848
rect 65736 34788 65740 34844
rect 65740 34788 65796 34844
rect 65796 34788 65800 34844
rect 65736 34784 65800 34788
rect 65816 34844 65880 34848
rect 65816 34788 65820 34844
rect 65820 34788 65876 34844
rect 65876 34788 65880 34844
rect 65816 34784 65880 34788
rect 65896 34844 65960 34848
rect 65896 34788 65900 34844
rect 65900 34788 65956 34844
rect 65956 34788 65960 34844
rect 65896 34784 65960 34788
rect 96376 34844 96440 34848
rect 96376 34788 96380 34844
rect 96380 34788 96436 34844
rect 96436 34788 96440 34844
rect 96376 34784 96440 34788
rect 96456 34844 96520 34848
rect 96456 34788 96460 34844
rect 96460 34788 96516 34844
rect 96516 34788 96520 34844
rect 96456 34784 96520 34788
rect 96536 34844 96600 34848
rect 96536 34788 96540 34844
rect 96540 34788 96596 34844
rect 96596 34788 96600 34844
rect 96536 34784 96600 34788
rect 96616 34844 96680 34848
rect 96616 34788 96620 34844
rect 96620 34788 96676 34844
rect 96676 34788 96680 34844
rect 96616 34784 96680 34788
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 50296 34300 50360 34304
rect 50296 34244 50300 34300
rect 50300 34244 50356 34300
rect 50356 34244 50360 34300
rect 50296 34240 50360 34244
rect 50376 34300 50440 34304
rect 50376 34244 50380 34300
rect 50380 34244 50436 34300
rect 50436 34244 50440 34300
rect 50376 34240 50440 34244
rect 50456 34300 50520 34304
rect 50456 34244 50460 34300
rect 50460 34244 50516 34300
rect 50516 34244 50520 34300
rect 50456 34240 50520 34244
rect 50536 34300 50600 34304
rect 50536 34244 50540 34300
rect 50540 34244 50596 34300
rect 50596 34244 50600 34300
rect 50536 34240 50600 34244
rect 81016 34300 81080 34304
rect 81016 34244 81020 34300
rect 81020 34244 81076 34300
rect 81076 34244 81080 34300
rect 81016 34240 81080 34244
rect 81096 34300 81160 34304
rect 81096 34244 81100 34300
rect 81100 34244 81156 34300
rect 81156 34244 81160 34300
rect 81096 34240 81160 34244
rect 81176 34300 81240 34304
rect 81176 34244 81180 34300
rect 81180 34244 81236 34300
rect 81236 34244 81240 34300
rect 81176 34240 81240 34244
rect 81256 34300 81320 34304
rect 81256 34244 81260 34300
rect 81260 34244 81316 34300
rect 81316 34244 81320 34300
rect 81256 34240 81320 34244
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 29500 31452 29564 31516
rect 102732 31452 102796 31516
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 51580 29412 51644 29476
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 79180 28052 79244 28116
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 52316 26692 52380 26756
rect 79548 26692 79612 26756
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 7604 26148 7668 26212
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 52316 25468 52380 25532
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 51948 24108 52012 24172
rect 79732 24108 79796 24172
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 12756 23428 12820 23492
rect 26372 23428 26436 23492
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 102732 23156 102796 23220
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 9812 22748 9876 22812
rect 52316 22808 52380 22812
rect 52316 22752 52366 22808
rect 52366 22752 52380 22808
rect 52316 22748 52380 22752
rect 78628 22748 78692 22812
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 21404 22068 21468 22132
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 78812 20028 78876 20092
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 9260 18668 9324 18732
rect 78260 18668 78324 18732
rect 79548 18668 79612 18732
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 9444 18048 9508 18052
rect 9444 17992 9494 18048
rect 9494 17992 9508 18048
rect 9444 17988 9508 17992
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 78628 17716 78692 17780
rect 79180 17716 79244 17780
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 20116 17308 20180 17372
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 18644 16628 18708 16692
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 16436 16008 16500 16012
rect 16436 15952 16450 16008
rect 16450 15952 16500 16008
rect 16436 15948 16500 15952
rect 79916 15948 79980 16012
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 21956 15328 22020 15332
rect 21956 15272 21970 15328
rect 21970 15272 22020 15328
rect 21956 15268 22020 15272
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 13676 14588 13740 14652
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
<< metal4 >>
rect 4208 43552 4528 44112
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 43014 4528 43488
rect 4208 42778 4250 43014
rect 4486 42778 4528 43014
rect 4208 42694 4528 42778
rect 4208 42464 4250 42694
rect 4486 42464 4528 42694
rect 4208 42400 4216 42464
rect 4280 42400 4296 42458
rect 4360 42400 4376 42458
rect 4440 42400 4456 42458
rect 4520 42400 4528 42464
rect 4208 41376 4528 42400
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 40288 4528 41312
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 39200 4528 40224
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 38112 4528 39136
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 37024 4528 38048
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 35936 4528 36960
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 19568 44096 19888 44112
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 43008 19888 44032
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 41920 19888 42944
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 40832 19888 41856
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 39744 19888 40768
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 38656 19888 39680
rect 34928 43552 35248 44112
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 43014 35248 43488
rect 34928 42778 34970 43014
rect 35206 42778 35248 43014
rect 34928 42694 35248 42778
rect 34928 42464 34970 42694
rect 35206 42464 35248 42694
rect 34928 42400 34936 42464
rect 35000 42400 35016 42458
rect 35080 42400 35096 42458
rect 35160 42400 35176 42458
rect 35240 42400 35248 42464
rect 34928 41376 35248 42400
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 40288 35248 41312
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 28947 39676 29013 39677
rect 28947 39612 28948 39676
rect 29012 39612 29013 39676
rect 28947 39611 29013 39612
rect 28950 39405 29010 39611
rect 28947 39404 29013 39405
rect 28947 39340 28948 39404
rect 29012 39340 29013 39404
rect 28947 39339 29013 39340
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 37568 19888 38592
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 34928 39200 35248 40224
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 38112 35248 39136
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 37024 35248 38048
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 35936 35248 36960
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33880 35248 34784
rect 50288 44096 50608 44112
rect 50288 44032 50296 44096
rect 50360 44032 50376 44096
rect 50440 44032 50456 44096
rect 50520 44032 50536 44096
rect 50600 44032 50608 44096
rect 50288 43008 50608 44032
rect 50288 42944 50296 43008
rect 50360 42944 50376 43008
rect 50440 42944 50456 43008
rect 50520 42944 50536 43008
rect 50600 42944 50608 43008
rect 50288 41920 50608 42944
rect 50288 41856 50296 41920
rect 50360 41856 50376 41920
rect 50440 41856 50456 41920
rect 50520 41856 50536 41920
rect 50600 41856 50608 41920
rect 50288 40832 50608 41856
rect 50288 40768 50296 40832
rect 50360 40768 50376 40832
rect 50440 40768 50456 40832
rect 50520 40768 50536 40832
rect 50600 40768 50608 40832
rect 50288 39744 50608 40768
rect 50288 39680 50296 39744
rect 50360 39680 50376 39744
rect 50440 39680 50456 39744
rect 50520 39680 50536 39744
rect 50600 39680 50608 39744
rect 50288 38656 50608 39680
rect 50288 38592 50296 38656
rect 50360 38592 50376 38656
rect 50440 38592 50456 38656
rect 50520 38592 50536 38656
rect 50600 38592 50608 38656
rect 50288 37568 50608 38592
rect 50288 37504 50296 37568
rect 50360 37504 50376 37568
rect 50440 37504 50456 37568
rect 50520 37504 50536 37568
rect 50600 37504 50608 37568
rect 50288 36480 50608 37504
rect 50288 36416 50296 36480
rect 50360 36416 50376 36480
rect 50440 36416 50456 36480
rect 50520 36416 50536 36480
rect 50600 36416 50608 36480
rect 50288 35392 50608 36416
rect 50288 35328 50296 35392
rect 50360 35328 50376 35392
rect 50440 35328 50456 35392
rect 50520 35328 50536 35392
rect 50600 35328 50608 35392
rect 50288 34304 50608 35328
rect 50288 34240 50296 34304
rect 50360 34240 50376 34304
rect 50440 34240 50456 34304
rect 50520 34240 50536 34304
rect 50600 34240 50608 34304
rect 50288 33880 50608 34240
rect 65648 43552 65968 44112
rect 65648 43488 65656 43552
rect 65720 43488 65736 43552
rect 65800 43488 65816 43552
rect 65880 43488 65896 43552
rect 65960 43488 65968 43552
rect 65648 43014 65968 43488
rect 65648 42778 65690 43014
rect 65926 42778 65968 43014
rect 65648 42694 65968 42778
rect 65648 42464 65690 42694
rect 65926 42464 65968 42694
rect 65648 42400 65656 42464
rect 65720 42400 65736 42458
rect 65800 42400 65816 42458
rect 65880 42400 65896 42458
rect 65960 42400 65968 42464
rect 65648 41376 65968 42400
rect 65648 41312 65656 41376
rect 65720 41312 65736 41376
rect 65800 41312 65816 41376
rect 65880 41312 65896 41376
rect 65960 41312 65968 41376
rect 65648 40288 65968 41312
rect 65648 40224 65656 40288
rect 65720 40224 65736 40288
rect 65800 40224 65816 40288
rect 65880 40224 65896 40288
rect 65960 40224 65968 40288
rect 65648 39200 65968 40224
rect 65648 39136 65656 39200
rect 65720 39136 65736 39200
rect 65800 39136 65816 39200
rect 65880 39136 65896 39200
rect 65960 39136 65968 39200
rect 65648 38112 65968 39136
rect 65648 38048 65656 38112
rect 65720 38048 65736 38112
rect 65800 38048 65816 38112
rect 65880 38048 65896 38112
rect 65960 38048 65968 38112
rect 65648 37024 65968 38048
rect 65648 36960 65656 37024
rect 65720 36960 65736 37024
rect 65800 36960 65816 37024
rect 65880 36960 65896 37024
rect 65960 36960 65968 37024
rect 65648 35936 65968 36960
rect 65648 35872 65656 35936
rect 65720 35872 65736 35936
rect 65800 35872 65816 35936
rect 65880 35872 65896 35936
rect 65960 35872 65968 35936
rect 65648 34848 65968 35872
rect 65648 34784 65656 34848
rect 65720 34784 65736 34848
rect 65800 34784 65816 34848
rect 65880 34784 65896 34848
rect 65960 34784 65968 34848
rect 65648 33880 65968 34784
rect 81008 44096 81328 44112
rect 81008 44032 81016 44096
rect 81080 44032 81096 44096
rect 81160 44032 81176 44096
rect 81240 44032 81256 44096
rect 81320 44032 81328 44096
rect 81008 43008 81328 44032
rect 81008 42944 81016 43008
rect 81080 42944 81096 43008
rect 81160 42944 81176 43008
rect 81240 42944 81256 43008
rect 81320 42944 81328 43008
rect 81008 41920 81328 42944
rect 81008 41856 81016 41920
rect 81080 41856 81096 41920
rect 81160 41856 81176 41920
rect 81240 41856 81256 41920
rect 81320 41856 81328 41920
rect 81008 40832 81328 41856
rect 81008 40768 81016 40832
rect 81080 40768 81096 40832
rect 81160 40768 81176 40832
rect 81240 40768 81256 40832
rect 81320 40768 81328 40832
rect 81008 39744 81328 40768
rect 81008 39680 81016 39744
rect 81080 39680 81096 39744
rect 81160 39680 81176 39744
rect 81240 39680 81256 39744
rect 81320 39680 81328 39744
rect 81008 38656 81328 39680
rect 81008 38592 81016 38656
rect 81080 38592 81096 38656
rect 81160 38592 81176 38656
rect 81240 38592 81256 38656
rect 81320 38592 81328 38656
rect 81008 37568 81328 38592
rect 81008 37504 81016 37568
rect 81080 37504 81096 37568
rect 81160 37504 81176 37568
rect 81240 37504 81256 37568
rect 81320 37504 81328 37568
rect 81008 36480 81328 37504
rect 81008 36416 81016 36480
rect 81080 36416 81096 36480
rect 81160 36416 81176 36480
rect 81240 36416 81256 36480
rect 81320 36416 81328 36480
rect 81008 35392 81328 36416
rect 81008 35328 81016 35392
rect 81080 35328 81096 35392
rect 81160 35328 81176 35392
rect 81240 35328 81256 35392
rect 81320 35328 81328 35392
rect 81008 34304 81328 35328
rect 81008 34240 81016 34304
rect 81080 34240 81096 34304
rect 81160 34240 81176 34304
rect 81240 34240 81256 34304
rect 81320 34240 81328 34304
rect 81008 33880 81328 34240
rect 96368 43552 96688 44112
rect 96368 43488 96376 43552
rect 96440 43488 96456 43552
rect 96520 43488 96536 43552
rect 96600 43488 96616 43552
rect 96680 43488 96688 43552
rect 96368 43014 96688 43488
rect 96368 42778 96410 43014
rect 96646 42778 96688 43014
rect 96368 42694 96688 42778
rect 96368 42464 96410 42694
rect 96646 42464 96688 42694
rect 96368 42400 96376 42464
rect 96440 42400 96456 42458
rect 96520 42400 96536 42458
rect 96600 42400 96616 42458
rect 96680 42400 96688 42464
rect 96368 41376 96688 42400
rect 96368 41312 96376 41376
rect 96440 41312 96456 41376
rect 96520 41312 96536 41376
rect 96600 41312 96616 41376
rect 96680 41312 96688 41376
rect 96368 40288 96688 41312
rect 96368 40224 96376 40288
rect 96440 40224 96456 40288
rect 96520 40224 96536 40288
rect 96600 40224 96616 40288
rect 96680 40224 96688 40288
rect 96368 39200 96688 40224
rect 96368 39136 96376 39200
rect 96440 39136 96456 39200
rect 96520 39136 96536 39200
rect 96600 39136 96616 39200
rect 96680 39136 96688 39200
rect 96368 38112 96688 39136
rect 96368 38048 96376 38112
rect 96440 38048 96456 38112
rect 96520 38048 96536 38112
rect 96600 38048 96616 38112
rect 96680 38048 96688 38112
rect 96368 37024 96688 38048
rect 96368 36960 96376 37024
rect 96440 36960 96456 37024
rect 96520 36960 96536 37024
rect 96600 36960 96616 37024
rect 96680 36960 96688 37024
rect 96368 35936 96688 36960
rect 96368 35872 96376 35936
rect 96440 35872 96456 35936
rect 96520 35872 96536 35936
rect 96600 35872 96616 35936
rect 96680 35872 96688 35936
rect 96368 34848 96688 35872
rect 96368 34784 96376 34848
rect 96440 34784 96456 34848
rect 96520 34784 96536 34848
rect 96600 34784 96616 34848
rect 96680 34784 96688 34848
rect 96368 33880 96688 34784
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 29499 31516 29565 31517
rect 29499 31452 29500 31516
rect 29564 31452 29565 31516
rect 29499 31451 29565 31452
rect 102731 31516 102797 31517
rect 102731 31452 102732 31516
rect 102796 31452 102797 31516
rect 102731 31451 102797 31452
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25014 19888 25536
rect 19568 24778 19610 25014
rect 19846 24778 19888 25014
rect 19568 24694 19888 24778
rect 19568 24512 19610 24694
rect 19846 24512 19888 24694
rect 19568 24448 19576 24512
rect 19640 24448 19656 24458
rect 19720 24448 19736 24458
rect 19800 24448 19816 24458
rect 19880 24448 19888 24512
rect 19568 23424 19888 24448
rect 26371 23492 26437 23493
rect 26371 23428 26372 23492
rect 26436 23428 26437 23492
rect 26371 23427 26437 23428
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 26374 21538 26434 23427
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20160 19888 21184
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 29502 14738 29562 31451
rect 51579 29476 51645 29477
rect 51579 29412 51580 29476
rect 51644 29412 51645 29476
rect 51579 29411 51645 29412
rect 51582 22898 51642 29411
rect 79179 28116 79245 28117
rect 79179 28052 79180 28116
rect 79244 28052 79245 28116
rect 79179 28051 79245 28052
rect 52315 26756 52381 26757
rect 52315 26692 52316 26756
rect 52380 26692 52381 26756
rect 52315 26691 52381 26692
rect 52318 26298 52378 26691
rect 52315 25532 52381 25533
rect 52315 25468 52316 25532
rect 52380 25468 52381 25532
rect 52315 25467 52381 25468
rect 51947 24172 52013 24173
rect 51947 24108 51948 24172
rect 52012 24108 52013 24172
rect 51947 24107 52013 24108
rect 51950 21538 52010 24107
rect 52318 23578 52378 25467
rect 52315 22812 52381 22813
rect 52315 22748 52316 22812
rect 52380 22748 52381 22812
rect 52315 22747 52381 22748
rect 78627 22812 78693 22813
rect 78627 22748 78628 22812
rect 78692 22748 78693 22812
rect 78627 22747 78693 22748
rect 52318 22218 52378 22747
rect 78630 17781 78690 22747
rect 78811 20092 78877 20093
rect 78811 20028 78812 20092
rect 78876 20028 78877 20092
rect 78811 20027 78877 20028
rect 78627 17780 78693 17781
rect 78627 17716 78628 17780
rect 78692 17716 78693 17780
rect 78627 17715 78693 17716
rect 78814 16778 78874 20027
rect 79182 18138 79242 28051
rect 79547 26756 79613 26757
rect 79547 26692 79548 26756
rect 79612 26692 79613 26756
rect 79547 26691 79613 26692
rect 79550 18733 79610 26691
rect 79731 24172 79797 24173
rect 79731 24108 79732 24172
rect 79796 24108 79797 24172
rect 79731 24107 79797 24108
rect 79547 18732 79613 18733
rect 79547 18668 79548 18732
rect 79612 18668 79613 18732
rect 79547 18667 79613 18668
rect 79734 18050 79794 24107
rect 102734 23221 102794 31451
rect 102731 23220 102797 23221
rect 102731 23156 102732 23220
rect 102796 23156 102797 23220
rect 102731 23155 102797 23156
rect 79550 17990 79794 18050
rect 79179 17780 79245 17781
rect 79179 17716 79180 17780
rect 79244 17716 79245 17780
rect 79179 17715 79245 17716
rect 79182 17458 79242 17715
rect 79550 15418 79610 17990
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7014 4528 7584
rect 4208 6778 4250 7014
rect 4486 6778 4528 7014
rect 4208 6694 4528 6778
rect 4208 6560 4250 6694
rect 4486 6560 4528 6694
rect 4208 6496 4216 6560
rect 4520 6496 4528 6560
rect 4208 6458 4250 6496
rect 4486 6458 4528 6496
rect 4208 5472 4528 6458
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 4384 4528 5408
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2128 19888 2688
<< via4 >>
rect 4250 42778 4486 43014
rect 4250 42464 4486 42694
rect 4250 42458 4280 42464
rect 4280 42458 4296 42464
rect 4296 42458 4360 42464
rect 4360 42458 4376 42464
rect 4376 42458 4440 42464
rect 4440 42458 4456 42464
rect 4456 42458 4486 42464
rect 34970 42778 35206 43014
rect 34970 42464 35206 42694
rect 34970 42458 35000 42464
rect 35000 42458 35016 42464
rect 35016 42458 35080 42464
rect 35080 42458 35096 42464
rect 35096 42458 35160 42464
rect 35160 42458 35176 42464
rect 35176 42458 35206 42464
rect 65690 42778 65926 43014
rect 65690 42464 65926 42694
rect 65690 42458 65720 42464
rect 65720 42458 65736 42464
rect 65736 42458 65800 42464
rect 65800 42458 65816 42464
rect 65816 42458 65880 42464
rect 65880 42458 65896 42464
rect 65896 42458 65926 42464
rect 96410 42778 96646 43014
rect 96410 42464 96646 42694
rect 96410 42458 96440 42464
rect 96440 42458 96456 42464
rect 96456 42458 96520 42464
rect 96520 42458 96536 42464
rect 96536 42458 96600 42464
rect 96600 42458 96616 42464
rect 96616 42458 96646 42464
rect 7518 26212 7754 26298
rect 7518 26148 7604 26212
rect 7604 26148 7668 26212
rect 7668 26148 7754 26212
rect 7518 26062 7754 26148
rect 19610 24778 19846 25014
rect 19610 24512 19846 24694
rect 19610 24458 19640 24512
rect 19640 24458 19656 24512
rect 19656 24458 19720 24512
rect 19720 24458 19736 24512
rect 19736 24458 19800 24512
rect 19800 24458 19816 24512
rect 19816 24458 19846 24512
rect 12670 23492 12906 23578
rect 12670 23428 12756 23492
rect 12756 23428 12820 23492
rect 12820 23428 12906 23492
rect 12670 23342 12906 23428
rect 9726 22812 9962 22898
rect 9726 22748 9812 22812
rect 9812 22748 9876 22812
rect 9876 22748 9962 22812
rect 9726 22662 9962 22748
rect 21318 22132 21554 22218
rect 21318 22068 21404 22132
rect 21404 22068 21468 22132
rect 21468 22068 21554 22132
rect 21318 21982 21554 22068
rect 26286 21302 26522 21538
rect 9174 18732 9410 18818
rect 9174 18668 9260 18732
rect 9260 18668 9324 18732
rect 9324 18668 9410 18732
rect 9174 18582 9410 18668
rect 9358 18052 9594 18138
rect 9358 17988 9444 18052
rect 9444 17988 9508 18052
rect 9508 17988 9594 18052
rect 9358 17902 9594 17988
rect 20030 17372 20266 17458
rect 20030 17308 20116 17372
rect 20116 17308 20180 17372
rect 20180 17308 20266 17372
rect 20030 17222 20266 17308
rect 18558 16692 18794 16778
rect 18558 16628 18644 16692
rect 18644 16628 18708 16692
rect 18708 16628 18794 16692
rect 18558 16542 18794 16628
rect 16350 16012 16586 16098
rect 16350 15948 16436 16012
rect 16436 15948 16500 16012
rect 16500 15948 16586 16012
rect 16350 15862 16586 15948
rect 13590 14652 13826 14738
rect 13590 14588 13676 14652
rect 13676 14588 13740 14652
rect 13740 14588 13826 14652
rect 13590 14502 13826 14588
rect 21870 15332 22106 15418
rect 21870 15268 21956 15332
rect 21956 15268 22020 15332
rect 22020 15268 22106 15332
rect 21870 15182 22106 15268
rect 52230 26062 52466 26298
rect 51494 22662 51730 22898
rect 52230 23342 52466 23578
rect 52230 21982 52466 22218
rect 51862 21302 52098 21538
rect 78174 18732 78410 18818
rect 78174 18668 78260 18732
rect 78260 18668 78324 18732
rect 78324 18668 78410 18732
rect 78174 18582 78410 18668
rect 79094 17902 79330 18138
rect 79094 17222 79330 17458
rect 78726 16542 78962 16778
rect 79830 16012 80066 16098
rect 79830 15948 79916 16012
rect 79916 15948 79980 16012
rect 79980 15948 80066 16012
rect 79830 15862 80066 15948
rect 79462 15182 79698 15418
rect 4250 6778 4486 7014
rect 4250 6560 4486 6694
rect 4250 6496 4280 6560
rect 4280 6496 4296 6560
rect 4296 6496 4360 6560
rect 4360 6496 4376 6560
rect 4376 6496 4440 6560
rect 4440 6496 4456 6560
rect 4456 6496 4486 6560
rect 4250 6458 4486 6496
rect 29414 14502 29650 14738
<< metal5 >>
rect 4208 43036 4528 43038
rect 34928 43036 35248 43038
rect 65648 43036 65968 43038
rect 96368 43036 96688 43038
rect 1104 43014 105616 43036
rect 1104 42778 4250 43014
rect 4486 42778 34970 43014
rect 35206 42778 65690 43014
rect 65926 42778 96410 43014
rect 96646 42778 105616 43014
rect 1104 42694 105616 42778
rect 1104 42458 4250 42694
rect 4486 42458 34970 42694
rect 35206 42458 65690 42694
rect 65926 42458 96410 42694
rect 96646 42458 105616 42694
rect 1104 42436 105616 42458
rect 4208 42434 4528 42436
rect 34928 42434 35248 42436
rect 65648 42434 65968 42436
rect 96368 42434 96688 42436
rect 7476 26298 52508 26340
rect 7476 26062 7518 26298
rect 7754 26062 52230 26298
rect 52466 26062 52508 26298
rect 7476 26020 52508 26062
rect 19568 25036 19888 25038
rect 1104 25014 105616 25036
rect 1104 24778 19610 25014
rect 19846 24778 105616 25014
rect 1104 24694 105616 24778
rect 1104 24458 19610 24694
rect 19846 24458 105616 24694
rect 1104 24436 105616 24458
rect 19568 24434 19888 24436
rect 12628 23578 52508 23620
rect 12628 23342 12670 23578
rect 12906 23342 52230 23578
rect 52466 23342 52508 23578
rect 12628 23300 52508 23342
rect 9684 22898 51772 22940
rect 9684 22662 9726 22898
rect 9962 22662 51494 22898
rect 51730 22662 51772 22898
rect 9684 22620 51772 22662
rect 21276 22218 52508 22260
rect 21276 21982 21318 22218
rect 21554 21982 52230 22218
rect 52466 21982 52508 22218
rect 21276 21940 52508 21982
rect 26244 21538 36132 21580
rect 26244 21302 26286 21538
rect 26522 21302 36132 21538
rect 26244 21260 36132 21302
rect 35812 20220 36132 21260
rect 45196 21538 52140 21580
rect 45196 21302 51862 21538
rect 52098 21302 52140 21538
rect 45196 21260 52140 21302
rect 45196 20220 45516 21260
rect 35812 19900 45516 20220
rect 9132 18818 78452 18860
rect 9132 18582 9174 18818
rect 9410 18582 78174 18818
rect 78410 18582 78452 18818
rect 9132 18540 78452 18582
rect 9316 18138 79372 18180
rect 9316 17902 9358 18138
rect 9594 17902 79094 18138
rect 79330 17902 79372 18138
rect 9316 17860 79372 17902
rect 19988 17458 79372 17500
rect 19988 17222 20030 17458
rect 20266 17222 79094 17458
rect 79330 17222 79372 17458
rect 19988 17180 79372 17222
rect 18516 16778 79004 16820
rect 18516 16542 18558 16778
rect 18794 16542 78726 16778
rect 78962 16542 79004 16778
rect 18516 16500 79004 16542
rect 16308 16098 80108 16140
rect 16308 15862 16350 16098
rect 16586 15862 79830 16098
rect 80066 15862 80108 16098
rect 16308 15820 80108 15862
rect 21828 15418 79740 15460
rect 21828 15182 21870 15418
rect 22106 15182 79462 15418
rect 79698 15182 79740 15418
rect 21828 15140 79740 15182
rect 13548 14738 29692 14780
rect 13548 14502 13590 14738
rect 13826 14502 29414 14738
rect 29650 14502 29692 14738
rect 13548 14460 29692 14502
rect 4208 7036 4528 7038
rect 1104 7014 105616 7036
rect 1104 6778 4250 7014
rect 4486 6778 105616 7014
rect 1104 6694 105616 6778
rect 1104 6458 4250 6694
rect 4486 6458 105616 6694
rect 1104 6436 105616 6458
rect 4208 6434 4528 6436
use sky130_fd_sc_hd__decap_8  FILLER_1_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 2484 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1607194113
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1607194113
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_152 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1607194113
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1607194113
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1483_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 3220 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_1_58
timestamp 1607194113
transform 1 0 6440 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_46
timestamp 1607194113
transform 1 0 5336 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1607194113
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__CLK $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 5152 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__D
timestamp 1607194113
transform 1 0 4968 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_74
timestamp 1607194113
transform 1 0 7912 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1607194113
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1607194113
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1607194113
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_740
timestamp 1607194113
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1607194113
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1607194113
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1607194113
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1607194113
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1484_
timestamp 1607194113
transform 1 0 8648 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_1_115
timestamp 1607194113
transform 1 0 11684 0 1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_103
timestamp 1607194113
transform 1 0 10580 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1607194113
transform 1 0 11960 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1607194113
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1484__CLK
timestamp 1607194113
transform 1 0 10396 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1607194113
transform 1 0 13524 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1607194113
transform 1 0 12420 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 12236 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_137
timestamp 1607194113
transform 1 0 13708 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1607194113
transform 1 0 12604 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_741
timestamp 1607194113
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1607194113
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1607194113
transform 1 0 14628 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1607194113
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_149
timestamp 1607194113
transform 1 0 14812 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1607194113
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1607194113
transform 1 0 16836 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1607194113
transform 1 0 15732 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1607194113
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1607194113
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1607194113
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1607194113
transform 1 0 18308 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1607194113
transform 1 0 17664 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_742
timestamp 1607194113
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1607194113
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1607194113
transform 1 0 20240 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1607194113
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1607194113
transform 1 0 20516 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1607194113
transform 1 0 19412 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1607194113
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_232
timestamp 1607194113
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_220
timestamp 1607194113
transform 1 0 21344 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1607194113
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1607194113
transform 1 0 23368 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_743
timestamp 1607194113
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1607194113
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1607194113
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1607194113
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1607194113
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1607194113
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1607194113
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1607194113
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1607194113
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1607194113
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1607194113
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1607194113
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1607194113
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_117
timestamp 1607194113
transform 1 0 11868 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1607194113
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_129
timestamp 1607194113
transform 1 0 12972 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1607194113
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_141
timestamp 1607194113
transform 1 0 14076 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1607194113
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1607194113
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1607194113
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1607194113
transform 1 0 18584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1607194113
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1607194113
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1607194113
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1607194113
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1607194113
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1607194113
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1607194113
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1485_
timestamp 1607194113
transform 1 0 2484 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_3_36
timestamp 1607194113
transform 1 0 4416 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1485__CLK
timestamp 1607194113
transform 1 0 4232 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_48
timestamp 1607194113
transform 1 0 5520 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_71
timestamp 1607194113
transform 1 0 7636 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_60
timestamp 1607194113
transform 1 0 6624 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1607194113
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:5.inst.g_clkdly15_2.dly $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 6808 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_3_91
timestamp 1607194113
transform 1 0 9476 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_83
timestamp 1607194113
transform 1 0 8740 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1341_
timestamp 1607194113
transform 1 0 9568 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_3_113
timestamp 1607194113
transform 1 0 11500 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1341__CLK
timestamp 1607194113
transform 1 0 11316 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1607194113
transform 1 0 13524 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1607194113
transform 1 0 12420 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1607194113
transform 1 0 12236 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1607194113
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1607194113
transform 1 0 14628 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1607194113
transform 1 0 16836 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1607194113
transform 1 0 15732 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1607194113
transform 1 0 19136 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1607194113
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1607194113
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1607194113
transform 1 0 20240 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1607194113
transform 1 0 22448 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1607194113
transform 1 0 21344 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1607194113
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1607194113
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1607194113
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1607194113
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1607194113
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1607194113
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1607194113
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_44
timestamp 1607194113
transform 1 0 5152 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1342_
timestamp 1607194113
transform 1 0 5520 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_4_69
timestamp 1607194113
transform 1 0 7452 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1342__CLK
timestamp 1607194113
transform 1 0 7268 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1607194113
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_89
timestamp 1607194113
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_81
timestamp 1607194113
transform 1 0 8556 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1607194113
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1333_
timestamp 1607194113
transform 1 0 10764 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_4_126
timestamp 1607194113
transform 1 0 12696 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1333__CLK
timestamp 1607194113
transform 1 0 12512 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:4.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 13248 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1607194113
transform 1 0 14076 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1607194113
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1340_
timestamp 1607194113
transform 1 0 15272 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_4_175
timestamp 1607194113
transform 1 0 17204 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1340__CLK
timestamp 1607194113
transform 1 0 17020 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_187
timestamp 1607194113
transform 1 0 18308 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1607194113
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_211
timestamp 1607194113
transform 1 0 20516 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_199
timestamp 1607194113
transform 1 0 19412 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1607194113
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1607194113
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1607194113
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1607194113
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1607194113
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1486_
timestamp 1607194113
transform 1 0 2484 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_5_36
timestamp 1607194113
transform 1 0 4416 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1486__CLK
timestamp 1607194113
transform 1 0 4232 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1607194113
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:6.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 4968 0 1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_5_62
timestamp 1607194113
transform 1 0 6808 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1607194113
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1334_
timestamp 1607194113
transform 1 0 6900 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_5_96
timestamp 1607194113
transform 1 0 9936 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_84
timestamp 1607194113
transform 1 0 8832 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1334__CLK
timestamp 1607194113
transform 1 0 8648 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_108
timestamp 1607194113
transform 1 0 11040 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1607194113
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1607194113
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1607194113
transform 1 0 12144 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1607194113
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_153
timestamp 1607194113
transform 1 0 15180 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_147
timestamp 1607194113
transform 1 0 14628 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1332__CLK
timestamp 1607194113
transform 1 0 15272 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1332_
timestamp 1607194113
transform 1 0 15456 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_5_175
timestamp 1607194113
transform 1 0 17204 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_5_196
timestamp 1607194113
transform 1 0 19136 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1607194113
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1607194113
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1339_
timestamp 1607194113
transform 1 0 19504 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_5_233
timestamp 1607194113
transform 1 0 22540 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_221
timestamp 1607194113
transform 1 0 21436 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1339__CLK
timestamp 1607194113
transform 1 0 21252 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_241
timestamp 1607194113
transform 1 0 23276 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1607194113
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1607194113
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1607194113
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1607194113
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1607194113
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1607194113
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1487_
timestamp 1607194113
transform 1 0 2484 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_7_38
timestamp 1607194113
transform 1 0 4600 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1607194113
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1487__CLK
timestamp 1607194113
transform 1 0 4416 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1487__D
timestamp 1607194113
transform 1 0 4232 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1607194113
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1343_
timestamp 1607194113
transform 1 0 4048 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_7_58
timestamp 1607194113
transform 1 0 6440 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_50
timestamp 1607194113
transform 1 0 5704 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1607194113
transform 1 0 5980 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1343__CLK
timestamp 1607194113
transform 1 0 5796 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_70
timestamp 1607194113
transform 1 0 7544 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_62
timestamp 1607194113
transform 1 0 6808 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_77
timestamp 1607194113
transform 1 0 8188 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1607194113
transform 1 0 7084 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1607194113
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1164_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 7820 0 1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_7_99
timestamp 1607194113
transform 1 0 10212 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_87
timestamp 1607194113
transform 1 0 9108 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1607194113
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_89
timestamp 1607194113
transform 1 0 9292 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1607194113
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_119
timestamp 1607194113
transform 1 0 12052 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_111
timestamp 1607194113
transform 1 0 11316 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_105
timestamp 1607194113
transform 1 0 10764 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _1165_
timestamp 1607194113
transform 1 0 11500 0 -1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1607194113
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1607194113
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_127
timestamp 1607194113
transform 1 0 12788 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1607194113
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_147
timestamp 1607194113
transform 1 0 14628 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_139
timestamp 1607194113
transform 1 0 13892 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1445__CLK
timestamp 1607194113
transform 1 0 14996 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1607194113
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1445_
timestamp 1607194113
transform 1 0 15272 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__o22a_4  _1166_
timestamp 1607194113
transform 1 0 14904 0 1 5984
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_7_176
timestamp 1607194113
transform 1 0 17296 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_164
timestamp 1607194113
transform 1 0 16192 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_173
timestamp 1607194113
transform 1 0 17020 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_196
timestamp 1607194113
transform 1 0 19136 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1607194113
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1607194113
transform 1 0 17848 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp 1607194113
transform 1 0 18860 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_6_185
timestamp 1607194113
transform 1 0 18124 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1607194113
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:3.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 19136 0 -1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_7_204
timestamp 1607194113
transform 1 0 19872 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_215
timestamp 1607194113
transform 1 0 20884 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_213
timestamp 1607194113
transform 1 0 20700 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_205
timestamp 1607194113
transform 1 0 19964 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1331__CLK
timestamp 1607194113
transform 1 0 20056 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1607194113
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1331_
timestamp 1607194113
transform 1 0 20240 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_7_227
timestamp 1607194113
transform 1 0 21988 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_221
timestamp 1607194113
transform 1 0 21436 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__CLK
timestamp 1607194113
transform 1 0 21528 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1346__D
timestamp 1607194113
transform 1 0 21712 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1346_
timestamp 1607194113
transform 1 0 21896 0 -1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_7_243
timestamp 1607194113
transform 1 0 23460 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_239
timestamp 1607194113
transform 1 0 23092 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1607194113
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1607194113
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1607194113
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1607194113
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1607194113
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1607194113
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1607194113
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_44
timestamp 1607194113
transform 1 0 5152 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1335_
timestamp 1607194113
transform 1 0 5428 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1607194113
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1335__CLK
timestamp 1607194113
transform 1 0 7176 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1607194113
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1607194113
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1607194113
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_105
timestamp 1607194113
transform 1 0 10764 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1446_
timestamp 1607194113
transform 1 0 11132 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_8_130
timestamp 1607194113
transform 1 0 13064 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1446__CLK
timestamp 1607194113
transform 1 0 12880 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0983_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 13800 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_8_145
timestamp 1607194113
transform 1 0 14444 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__B2
timestamp 1607194113
transform 1 0 14996 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1607194113
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1167_
timestamp 1607194113
transform 1 0 15272 0 -1 7072
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_8_168
timestamp 1607194113
transform 1 0 16560 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_196
timestamp 1607194113
transform 1 0 19136 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_192
timestamp 1607194113
transform 1 0 18768 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_180
timestamp 1607194113
transform 1 0 17664 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:2.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 19228 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_8_206
timestamp 1607194113
transform 1 0 20056 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1338__CLK
timestamp 1607194113
transform 1 0 20608 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_181
timestamp 1607194113
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1338_
timestamp 1607194113
transform 1 0 20884 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_8_234
timestamp 1607194113
transform 1 0 22632 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1607194113
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1607194113
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1488_
timestamp 1607194113
transform 1 0 2484 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_9_36
timestamp 1607194113
transform 1 0 4416 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1488__CLK
timestamp 1607194113
transform 1 0 4232 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_48
timestamp 1607194113
transform 1 0 5520 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_62
timestamp 1607194113
transform 1 0 6808 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1607194113
transform 1 0 6624 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_182
timestamp 1607194113
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1447_
timestamp 1607194113
transform 1 0 6992 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_9_97
timestamp 1607194113
transform 1 0 10028 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_85
timestamp 1607194113
transform 1 0 8924 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1447__CLK
timestamp 1607194113
transform 1 0 8740 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_109
timestamp 1607194113
transform 1 0 11132 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_135
timestamp 1607194113
transform 1 0 13524 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1607194113
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_121
timestamp 1607194113
transform 1 0 12236 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_183
timestamp 1607194113
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1444_
timestamp 1607194113
transform 1 0 13708 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_9_158
timestamp 1607194113
transform 1 0 15640 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1444__CLK
timestamp 1607194113
transform 1 0 15456 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_170
timestamp 1607194113
transform 1 0 16744 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_196
timestamp 1607194113
transform 1 0 19136 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1607194113
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1607194113
transform 1 0 17848 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_184
timestamp 1607194113
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:1.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 19320 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_9_207
timestamp 1607194113
transform 1 0 20148 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1330__CLK
timestamp 1607194113
transform 1 0 20700 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1330_
timestamp 1607194113
transform 1 0 20884 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_9_234
timestamp 1607194113
transform 1 0 22632 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_242
timestamp 1607194113
transform 1 0 23368 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_185
timestamp 1607194113
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1607194113
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1607194113
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1607194113
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1607194113
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1607194113
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_186
timestamp 1607194113
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1607194113
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1607194113
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _1162_
timestamp 1607194113
transform 1 0 7360 0 -1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_10_84
timestamp 1607194113
transform 1 0 8832 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__A2
timestamp 1607194113
transform 1 0 8648 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_187
timestamp 1607194113
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0969_
timestamp 1607194113
transform 1 0 9660 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_10_112
timestamp 1607194113
transform 1 0 11408 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_100
timestamp 1607194113
transform 1 0 10304 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _0976_
timestamp 1607194113
transform 1 0 11776 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_10_123
timestamp 1607194113
transform 1 0 12420 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A
timestamp 1607194113
transform 1 0 12972 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0982_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 13156 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_10_150
timestamp 1607194113
transform 1 0 14904 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_142
timestamp 1607194113
transform 1 0 14168 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__C
timestamp 1607194113
transform 1 0 13984 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A
timestamp 1607194113
transform 1 0 14996 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_188
timestamp 1607194113
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0990_
timestamp 1607194113
transform 1 0 15272 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_10_175
timestamp 1607194113
transform 1 0 17204 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_163
timestamp 1607194113
transform 1 0 16100 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_187
timestamp 1607194113
transform 1 0 18308 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1607194113
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_211
timestamp 1607194113
transform 1 0 20516 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_199
timestamp 1607194113
transform 1 0 19412 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_189
timestamp 1607194113
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1607194113
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1607194113
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1607194113
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1607194113
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1489_
timestamp 1607194113
transform 1 0 2484 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_11_36
timestamp 1607194113
transform 1 0 4416 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1489__CLK
timestamp 1607194113
transform 1 0 4232 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_48
timestamp 1607194113
transform 1 0 5520 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1607194113
transform 1 0 6624 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_190
timestamp 1607194113
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1448_
timestamp 1607194113
transform 1 0 6808 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_11_99
timestamp 1607194113
transform 1 0 10212 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_91
timestamp 1607194113
transform 1 0 9476 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_83
timestamp 1607194113
transform 1 0 8740 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1448__CLK
timestamp 1607194113
transform 1 0 8556 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__A
timestamp 1607194113
transform 1 0 10028 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1163_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 9660 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_119
timestamp 1607194113
transform 1 0 12052 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_111
timestamp 1607194113
transform 1 0 11316 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1607194113
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_191
timestamp 1607194113
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1168_
timestamp 1607194113
transform 1 0 13524 0 1 8160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_11_149
timestamp 1607194113
transform 1 0 14812 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1161_
timestamp 1607194113
transform 1 0 15548 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_173
timestamp 1607194113
transform 1 0 17020 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_161
timestamp 1607194113
transform 1 0 15916 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_190
timestamp 1607194113
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_184
timestamp 1607194113
transform 1 0 18032 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1607194113
transform 1 0 17756 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_192
timestamp 1607194113
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1337_
timestamp 1607194113
transform 1 0 18676 0 1 8160
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_11_212
timestamp 1607194113
transform 1 0 20608 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1337__CLK
timestamp 1607194113
transform 1 0 20424 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_236
timestamp 1607194113
transform 1 0 22816 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_224
timestamp 1607194113
transform 1 0 21712 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_193
timestamp 1607194113
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1607194113
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1607194113
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1607194113
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1607194113
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1607194113
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_194
timestamp 1607194113
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_56
timestamp 1607194113
transform 1 0 6256 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1607194113
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _0996_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 6348 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_12_64
timestamp 1607194113
transform 1 0 6992 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _0975_
timestamp 1607194113
transform 1 0 7728 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 1607194113
transform 1 0 9476 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_83
timestamp 1607194113
transform 1 0 8740 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__C
timestamp 1607194113
transform 1 0 8556 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_195
timestamp 1607194113
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0960_
timestamp 1607194113
transform 1 0 9660 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_12_112
timestamp 1607194113
transform 1 0 11408 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_100
timestamp 1607194113
transform 1 0 10304 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_124
timestamp 1607194113
transform 1 0 12512 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1443_
timestamp 1607194113
transform 1 0 12696 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_12_147
timestamp 1607194113
transform 1 0 14628 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1443__CLK
timestamp 1607194113
transform 1 0 14444 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__A
timestamp 1607194113
transform 1 0 15548 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_196
timestamp 1607194113
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1160_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 15272 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_171
timestamp 1607194113
transform 1 0 16836 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_159
timestamp 1607194113
transform 1 0 15732 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_189
timestamp 1607194113
transform 1 0 18492 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_183
timestamp 1607194113
transform 1 0 17940 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__clkdlybuf4s15_2  inst_core.g_test.i_minitdc.gen_delay:0.inst.g_clkdly15_2.dly
timestamp 1607194113
transform 1 0 18584 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_12_215
timestamp 1607194113
transform 1 0 20884 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_213
timestamp 1607194113
transform 1 0 20700 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_201
timestamp 1607194113
transform 1 0 19596 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_core.g_test.i_minitdc.gen_delay:0.inst.g_clkdly15_2.dly_A
timestamp 1607194113
transform 1 0 19412 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_197
timestamp 1607194113
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_219
timestamp 1607194113
transform 1 0 21252 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1347__CLK
timestamp 1607194113
transform 1 0 21344 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1347_
timestamp 1607194113
transform 1 0 21528 0 -1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_12_241
timestamp 1607194113
transform 1 0 23276 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1607194113
transform 1 0 2484 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1607194113
transform 1 0 1380 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1607194113
transform 1 0 1380 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1607194113
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1607194113
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1490_
timestamp 1607194113
transform 1 0 2484 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1607194113
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1607194113
transform 1 0 3588 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_36
timestamp 1607194113
transform 1 0 4416 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1490__CLK
timestamp 1607194113
transform 1 0 4232 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_202
timestamp 1607194113
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_56
timestamp 1607194113
transform 1 0 6256 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1607194113
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_48
timestamp 1607194113
transform 1 0 5520 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0940_
timestamp 1607194113
transform 1 0 6532 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_78
timestamp 1607194113
transform 1 0 8280 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_65
timestamp 1607194113
transform 1 0 7084 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_13_70
timestamp 1607194113
transform 1 0 7544 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_62
timestamp 1607194113
transform 1 0 6808 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_60
timestamp 1607194113
transform 1 0 6624 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A
timestamp 1607194113
transform 1 0 6900 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_198
timestamp 1607194113
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _0968_
timestamp 1607194113
transform 1 0 7728 0 1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _0956_
timestamp 1607194113
transform 1 0 7636 0 -1 10336
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1607194113
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 1607194113
transform 1 0 9384 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_96
timestamp 1607194113
transform 1 0 9936 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_83
timestamp 1607194113
transform 1 0 8740 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__C
timestamp 1607194113
transform 1 0 8556 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_203
timestamp 1607194113
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1002_
timestamp 1607194113
transform 1 0 9292 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_14_117
timestamp 1607194113
transform 1 0 11868 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1607194113
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_108
timestamp 1607194113
transform 1 0 11040 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_127
timestamp 1607194113
transform 1 0 12788 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_123
timestamp 1607194113
transform 1 0 12420 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_120
timestamp 1607194113
transform 1 0 12144 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_199
timestamp 1607194113
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1442_
timestamp 1607194113
transform 1 0 12236 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__o22a_4  _1169_
timestamp 1607194113
transform 1 0 12880 0 1 9248
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_14_157
timestamp 1607194113
transform 1 0 15548 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_150
timestamp 1607194113
transform 1 0 14904 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_142
timestamp 1607194113
transform 1 0 14168 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_156
timestamp 1607194113
transform 1 0 15456 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_144
timestamp 1607194113
transform 1 0 14352 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1442__CLK
timestamp 1607194113
transform 1 0 13984 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__B1
timestamp 1607194113
transform 1 0 14168 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204
timestamp 1607194113
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1607194113
transform 1 0 15272 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_169
timestamp 1607194113
transform 1 0 16652 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_168
timestamp 1607194113
transform 1 0 16560 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_193
timestamp 1607194113
transform 1 0 18860 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_181
timestamp 1607194113
transform 1 0 17756 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_192
timestamp 1607194113
transform 1 0 18768 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_184
timestamp 1607194113
transform 1 0 18032 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_180
timestamp 1607194113
transform 1 0 17664 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_200
timestamp 1607194113
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1329_
timestamp 1607194113
transform 1 0 18952 0 1 9248
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_14_213
timestamp 1607194113
transform 1 0 20700 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_205
timestamp 1607194113
transform 1 0 19964 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_215
timestamp 1607194113
transform 1 0 20884 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1348__CLK
timestamp 1607194113
transform 1 0 20884 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1329__CLK
timestamp 1607194113
transform 1 0 20700 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1607194113
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1348_
timestamp 1607194113
transform 1 0 21068 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_14_236
timestamp 1607194113
transform 1 0 22816 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_227
timestamp 1607194113
transform 1 0 21988 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_243
timestamp 1607194113
transform 1 0 23460 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_239
timestamp 1607194113
transform 1 0 23092 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_201
timestamp 1607194113
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1607194113
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1607194113
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1491_
timestamp 1607194113
transform 1 0 2484 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_15_36
timestamp 1607194113
transform 1 0 4416 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1491__CLK
timestamp 1607194113
transform 1 0 4232 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_56
timestamp 1607194113
transform 1 0 6256 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_48
timestamp 1607194113
transform 1 0 5520 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1297__B1
timestamp 1607194113
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_78
timestamp 1607194113
transform 1 0 8280 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1607194113
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1297_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 6808 0 1 10336
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_15_90
timestamp 1607194113
transform 1 0 9384 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_114
timestamp 1607194113
transform 1 0 11592 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_102
timestamp 1607194113
transform 1 0 10488 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1607194113
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1441_
timestamp 1607194113
transform 1 0 12420 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_15_156
timestamp 1607194113
transform 1 0 15456 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_144
timestamp 1607194113
transform 1 0 14352 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1441__CLK
timestamp 1607194113
transform 1 0 14168 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_168
timestamp 1607194113
transform 1 0 16560 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_180
timestamp 1607194113
transform 1 0 17664 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1328__CLK
timestamp 1607194113
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1607194113
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1328_
timestamp 1607194113
transform 1 0 18032 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_15_203
timestamp 1607194113
transform 1 0 19780 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1349__CLK
timestamp 1607194113
transform 1 0 20332 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1349_
timestamp 1607194113
transform 1 0 20516 0 1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_15_230
timestamp 1607194113
transform 1 0 22264 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_242
timestamp 1607194113
transform 1 0 23368 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1607194113
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1607194113
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1607194113
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1607194113
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1607194113
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1607194113
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1607194113
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_56
timestamp 1607194113
transform 1 0 6256 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1607194113
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_64
timestamp 1607194113
transform 1 0 6992 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1362_
timestamp 1607194113
transform 1 0 7084 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1607194113
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_86
timestamp 1607194113
transform 1 0 9016 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1362__CLK
timestamp 1607194113
transform 1 0 8832 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1607194113
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_117
timestamp 1607194113
transform 1 0 11868 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1607194113
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _1170_
timestamp 1607194113
transform 1 0 12604 0 -1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_16_154
timestamp 1607194113
transform 1 0 15272 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1607194113
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__B1
timestamp 1607194113
transform 1 0 13892 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1607194113
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_167
timestamp 1607194113
transform 1 0 16468 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_162
timestamp 1607194113
transform 1 0 16008 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 16192 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1336_
timestamp 1607194113
transform 1 0 17204 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_16_198
timestamp 1607194113
transform 1 0 19320 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__CLK
timestamp 1607194113
transform 1 0 19136 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1336__D
timestamp 1607194113
transform 1 0 18952 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1607194113
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_213
timestamp 1607194113
transform 1 0 20700 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_205
timestamp 1607194113
transform 1 0 19964 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_clk_i
timestamp 1607194113
transform 1 0 19688 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1607194113
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_227
timestamp 1607194113
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1607194113
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1607194113
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1607194113
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1492_
timestamp 1607194113
transform 1 0 2484 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_17_38
timestamp 1607194113
transform 1 0 4600 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1492__CLK
timestamp 1607194113
transform 1 0 4416 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1492__D
timestamp 1607194113
transform 1 0 4232 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_58
timestamp 1607194113
transform 1 0 6440 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_50
timestamp 1607194113
transform 1 0 5704 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_62
timestamp 1607194113
transform 1 0 6808 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1607194113
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1361_
timestamp 1607194113
transform 1 0 6992 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_17_97
timestamp 1607194113
transform 1 0 10028 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_85
timestamp 1607194113
transform 1 0 8924 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1361__CLK
timestamp 1607194113
transform 1 0 8740 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_109
timestamp 1607194113
transform 1 0 11132 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1607194113
transform 1 0 13524 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1607194113
transform 1 0 12420 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1607194113
transform 1 0 12236 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1607194113
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_147
timestamp 1607194113
transform 1 0 14628 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_172
timestamp 1607194113
transform 1 0 16928 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_159
timestamp 1607194113
transform 1 0 15732 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1286__A
timestamp 1607194113
transform 1 0 16744 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1286_
timestamp 1607194113
transform 1 0 16468 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_196
timestamp 1607194113
transform 1 0 19136 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1607194113
transform 1 0 18032 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_180
timestamp 1607194113
transform 1 0 17664 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1607194113
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1449_
timestamp 1607194113
transform 1 0 19504 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_17_232
timestamp 1607194113
transform 1 0 22448 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_221
timestamp 1607194113
transform 1 0 21436 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1449__CLK
timestamp 1607194113
transform 1 0 21252 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1304_
timestamp 1607194113
transform 1 0 22172 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1607194113
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1607194113
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1607194113
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1607194113
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_32
timestamp 1607194113
transform 1 0 4048 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1607194113
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1607194113
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_45
timestamp 1607194113
transform 1 0 5244 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_40
timestamp 1607194113
transform 1 0 4784 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1299__B1
timestamp 1607194113
transform 1 0 5796 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1299_
timestamp 1607194113
transform 1 0 5980 0 -1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _1296_
timestamp 1607194113
transform 1 0 4876 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_69
timestamp 1607194113
transform 1 0 7452 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1295_
timestamp 1607194113
transform 1 0 8188 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1607194113
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 1607194113
transform 1 0 9384 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_82
timestamp 1607194113
transform 1 0 8648 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1295__A
timestamp 1607194113
transform 1 0 8464 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1607194113
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1607194113
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1607194113
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_129
timestamp 1607194113
transform 1 0 12972 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_154
timestamp 1607194113
transform 1 0 15272 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1607194113
transform 1 0 14076 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1607194113
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1366_
timestamp 1607194113
transform 1 0 15640 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1366__CLK
timestamp 1607194113
transform 1 0 17388 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_188
timestamp 1607194113
transform 1 0 18400 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_179
timestamp 1607194113
transform 1 0 17572 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_clk_i
timestamp 1607194113
transform 1 0 18124 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_215
timestamp 1607194113
transform 1 0 20884 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1607194113
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_200
timestamp 1607194113
transform 1 0 19504 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1607194113
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1358__CLK
timestamp 1607194113
transform 1 0 21252 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1358_
timestamp 1607194113
transform 1 0 21436 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_18_240
timestamp 1607194113
transform 1 0 23184 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1607194113
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1607194113
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1607194113
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1607194113
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1607194113
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1607194113
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_36
timestamp 1607194113
transform 1 0 4416 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_32
timestamp 1607194113
transform 1 0 4048 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1607194113
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_27
timestamp 1607194113
transform 1 0 3588 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1301__B1
timestamp 1607194113
transform 1 0 4324 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1607194113
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1360_
timestamp 1607194113
transform 1 0 4508 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _1301_
timestamp 1607194113
transform 1 0 4508 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_20_58
timestamp 1607194113
transform 1 0 6440 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_53
timestamp 1607194113
transform 1 0 5980 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1360__CLK
timestamp 1607194113
transform 1 0 6256 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_75
timestamp 1607194113
transform 1 0 8004 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_62
timestamp 1607194113
transform 1 0 6808 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1298__A
timestamp 1607194113
transform 1 0 7820 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1303__B1
timestamp 1607194113
transform 1 0 7176 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1607194113
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1303_
timestamp 1607194113
transform 1 0 7360 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1298_
timestamp 1607194113
transform 1 0 7544 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1607194113
transform 1 0 10028 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_84
timestamp 1607194113
transform 1 0 8832 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_99
timestamp 1607194113
transform 1 0 10212 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_87
timestamp 1607194113
transform 1 0 9108 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1607194113
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1283_
timestamp 1607194113
transform 1 0 9660 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_109
timestamp 1607194113
transform 1 0 11132 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_116
timestamp 1607194113
transform 1 0 11776 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_104
timestamp 1607194113
transform 1 0 10672 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1285__B1
timestamp 1607194113
transform 1 0 11316 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1285_
timestamp 1607194113
transform 1 0 11500 0 -1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _1284_
timestamp 1607194113
transform 1 0 10304 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_129
timestamp 1607194113
transform 1 0 12972 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1607194113
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1367_
timestamp 1607194113
transform 1 0 12420 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1281_
timestamp 1607194113
transform 1 0 13708 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_142
timestamp 1607194113
transform 1 0 14168 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_148
timestamp 1607194113
transform 1 0 14720 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_144
timestamp 1607194113
transform 1 0 14352 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1367__CLK
timestamp 1607194113
transform 1 0 14168 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1281__A
timestamp 1607194113
transform 1 0 13984 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_clk_i
timestamp 1607194113
transform 1 0 14720 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_151
timestamp 1607194113
transform 1 0 14996 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1287__B1
timestamp 1607194113
transform 1 0 14812 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1607194113
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1607194113
transform 1 0 15272 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _1287_
timestamp 1607194113
transform 1 0 14996 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_19_167
timestamp 1607194113
transform 1 0 16468 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1365__CLK
timestamp 1607194113
transform 1 0 16376 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1365_
timestamp 1607194113
transform 1 0 16560 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_20_187
timestamp 1607194113
transform 1 0 18308 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1607194113
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1607194113
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_179
timestamp 1607194113
transform 1 0 17572 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1607194113
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_215
timestamp 1607194113
transform 1 0 20884 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_211
timestamp 1607194113
transform 1 0 20516 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_199
timestamp 1607194113
transform 1 0 19412 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_208
timestamp 1607194113
transform 1 0 20240 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1305__B1
timestamp 1607194113
transform 1 0 20424 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1607194113
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1305_
timestamp 1607194113
transform 1 0 20608 0 1 12512
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_20_223
timestamp 1607194113
transform 1 0 21620 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_228
timestamp 1607194113
transform 1 0 22080 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1357__CLK
timestamp 1607194113
transform 1 0 21712 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1357_
timestamp 1607194113
transform 1 0 21896 0 -1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_19_240
timestamp 1607194113
transform 1 0 23184 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1607194113
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1607194113
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1607194113
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1493_
timestamp 1607194113
transform 1 0 2484 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_21_38
timestamp 1607194113
transform 1 0 4600 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1493__CLK
timestamp 1607194113
transform 1 0 4416 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1493__D
timestamp 1607194113
transform 1 0 4232 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_55
timestamp 1607194113
transform 1 0 6164 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1300__A
timestamp 1607194113
transform 1 0 5980 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1300_
timestamp 1607194113
transform 1 0 5704 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_74
timestamp 1607194113
transform 1 0 7912 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1607194113
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1607194113
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1359_
timestamp 1607194113
transform 1 0 8004 0 1 13600
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_21_96
timestamp 1607194113
transform 1 0 9936 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1359__CLK
timestamp 1607194113
transform 1 0 9752 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_118
timestamp 1607194113
transform 1 0 11960 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_106
timestamp 1607194113
transform 1 0 10856 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1289_
timestamp 1607194113
transform 1 0 10488 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1607194113
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1607194113
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1607194113
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_147
timestamp 1607194113
transform 1 0 14628 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1290__B1
timestamp 1607194113
transform 1 0 14904 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_clk_i
timestamp 1607194113
transform 1 0 15088 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1290_
timestamp 1607194113
transform 1 0 15364 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_21_171
timestamp 1607194113
transform 1 0 16836 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_197
timestamp 1607194113
transform 1 0 19228 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_189
timestamp 1607194113
transform 1 0 18492 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1288__A
timestamp 1607194113
transform 1 0 18308 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1607194113
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1288_
timestamp 1607194113
transform 1 0 18032 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_205
timestamp 1607194113
transform 1 0 19964 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__A
timestamp 1607194113
transform 1 0 19412 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1307__B1
timestamp 1607194113
transform 1 0 20700 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1307_
timestamp 1607194113
transform 1 0 20884 0 1 13600
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _1159_
timestamp 1607194113
transform 1 0 19596 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_231
timestamp 1607194113
transform 1 0 22356 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_243
timestamp 1607194113
transform 1 0 23460 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1607194113
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1607194113
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1607194113
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1607194113
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1607194113
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1607194113
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1607194113
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_50
timestamp 1607194113
transform 1 0 5704 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_44
timestamp 1607194113
transform 1 0 5152 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__A
timestamp 1607194113
transform 1 0 5244 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0677_
timestamp 1607194113
transform 1 0 5428 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_74
timestamp 1607194113
transform 1 0 7912 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_62
timestamp 1607194113
transform 1 0 6808 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_93
timestamp 1607194113
transform 1 0 9660 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_22_86
timestamp 1607194113
transform 1 0 9016 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_80
timestamp 1607194113
transform 1 0 8464 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1302__A
timestamp 1607194113
transform 1 0 8832 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__A
timestamp 1607194113
transform 1 0 10212 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1607194113
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1302_
timestamp 1607194113
transform 1 0 8556 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_110
timestamp 1607194113
transform 1 0 11224 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _1011_
timestamp 1607194113
transform 1 0 10396 0 -1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_22_130
timestamp 1607194113
transform 1 0 13064 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_122
timestamp 1607194113
transform 1 0 12328 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1005_
timestamp 1607194113
transform 1 0 12420 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_22_154
timestamp 1607194113
transform 1 0 15272 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_147
timestamp 1607194113
transform 1 0 14628 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1363__CLK
timestamp 1607194113
transform 1 0 15640 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1293__A
timestamp 1607194113
transform 1 0 14444 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1607194113
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1293_
timestamp 1607194113
transform 1 0 14168 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1363_
timestamp 1607194113
transform 1 0 15824 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_22_187
timestamp 1607194113
transform 1 0 18308 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_179
timestamp 1607194113
transform 1 0 17572 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1292__B1
timestamp 1607194113
transform 1 0 18400 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1292_
timestamp 1607194113
transform 1 0 18584 0 -1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1607194113
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_206
timestamp 1607194113
transform 1 0 20056 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1607194113
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_238
timestamp 1607194113
transform 1 0 23000 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_227
timestamp 1607194113
transform 1 0 21988 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1306_
timestamp 1607194113
transform 1 0 22724 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1607194113
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1607194113
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1494_
timestamp 1607194113
transform 1 0 2484 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_23_38
timestamp 1607194113
transform 1 0 4600 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1494__CLK
timestamp 1607194113
transform 1 0 4416 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1494__D
timestamp 1607194113
transform 1 0 4232 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_48
timestamp 1607194113
transform 1 0 5520 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__A
timestamp 1607194113
transform 1 0 4968 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0680_
timestamp 1607194113
transform 1 0 5152 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_70
timestamp 1607194113
transform 1 0 7544 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_62
timestamp 1607194113
transform 1 0 6808 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_60
timestamp 1607194113
transform 1 0 6624 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__A
timestamp 1607194113
transform 1 0 7728 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1607194113
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1022_
timestamp 1607194113
transform 1 0 7912 0 1 14688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_23_95
timestamp 1607194113
transform 1 0 9844 0 1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_83
timestamp 1607194113
transform 1 0 8740 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1607194113
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__A
timestamp 1607194113
transform 1 0 11040 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1004_
timestamp 1607194113
transform 1 0 10396 0 1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_23_131
timestamp 1607194113
transform 1 0 13156 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_123
timestamp 1607194113
transform 1 0 12420 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_clk_i
timestamp 1607194113
transform 1 0 13248 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1607194113
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0958_
timestamp 1607194113
transform 1 0 13524 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_147
timestamp 1607194113
transform 1 0 14628 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_139
timestamp 1607194113
transform 1 0 13892 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1294__B1
timestamp 1607194113
transform 1 0 14720 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1294_
timestamp 1607194113
transform 1 0 14904 0 1 14688
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_23_178
timestamp 1607194113
transform 1 0 17480 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_166
timestamp 1607194113
transform 1 0 16376 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_196
timestamp 1607194113
transform 1 0 19136 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1607194113
transform 1 0 18032 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1607194113
transform 1 0 17848 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1607194113
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_204
timestamp 1607194113
transform 1 0 19872 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1364__CLK
timestamp 1607194113
transform 1 0 20148 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1364_
timestamp 1607194113
transform 1 0 20332 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_23_228
timestamp 1607194113
transform 1 0 22080 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_240
timestamp 1607194113
transform 1 0 23184 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1607194113
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1607194113
transform 1 0 2484 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1607194113
transform 1 0 1380 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1607194113
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_27
timestamp 1607194113
transform 1 0 3588 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1496__D
timestamp 1607194113
transform 1 0 3772 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1607194113
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1496_
timestamp 1607194113
transform 1 0 4048 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_24_53
timestamp 1607194113
transform 1 0 5980 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1496__CLK
timestamp 1607194113
transform 1 0 5796 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A
timestamp 1607194113
transform 1 0 6348 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0939_
timestamp 1607194113
transform 1 0 6532 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_71
timestamp 1607194113
transform 1 0 7636 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_63
timestamp 1607194113
transform 1 0 6900 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1012_
timestamp 1607194113
transform 1 0 7912 0 -1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_24_99
timestamp 1607194113
transform 1 0 10212 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_93
timestamp 1607194113
transform 1 0 9660 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1607194113
transform 1 0 9476 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_83
timestamp 1607194113
transform 1 0 8740 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__A
timestamp 1607194113
transform 1 0 8556 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1607194113
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1019_
timestamp 1607194113
transform 1 0 9936 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_4  _1020_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 10948 0 -1 15776
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_24_121
timestamp 1607194113
transform 1 0 12236 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__B
timestamp 1607194113
transform 1 0 13800 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1010_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 12972 0 -1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_24_154
timestamp 1607194113
transform 1 0 15272 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_148
timestamp 1607194113
transform 1 0 14720 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_140
timestamp 1607194113
transform 1 0 13984 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A1
timestamp 1607194113
transform 1 0 14996 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1607194113
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0955_
timestamp 1607194113
transform 1 0 15364 0 -1 15776
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_24_171
timestamp 1607194113
transform 1 0 16836 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A2
timestamp 1607194113
transform 1 0 16652 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_198
timestamp 1607194113
transform 1 0 19320 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_186
timestamp 1607194113
transform 1 0 18216 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp 1607194113
transform 1 0 17940 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_215
timestamp 1607194113
transform 1 0 20884 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_213
timestamp 1607194113
transform 1 0 20700 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_205
timestamp 1607194113
transform 1 0 19964 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1291__A
timestamp 1607194113
transform 1 0 19780 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1607194113
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1291_
timestamp 1607194113
transform 1 0 19504 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_223
timestamp 1607194113
transform 1 0 21620 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1408__CLK
timestamp 1607194113
transform 1 0 21712 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1408_
timestamp 1607194113
transform 1 0 21896 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1607194113
transform 1 0 1380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1607194113
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1495_
timestamp 1607194113
transform 1 0 2484 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_25_38
timestamp 1607194113
transform 1 0 4600 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__CLK
timestamp 1607194113
transform 1 0 4416 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__D
timestamp 1607194113
transform 1 0 4232 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_58
timestamp 1607194113
transform 1 0 6440 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_46
timestamp 1607194113
transform 1 0 5336 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0667__A
timestamp 1607194113
transform 1 0 4784 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0667_
timestamp 1607194113
transform 1 0 4968 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_73
timestamp 1607194113
transform 1 0 7820 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_62
timestamp 1607194113
transform 1 0 6808 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1607194113
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1003_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 6992 0 1 15776
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_25_91
timestamp 1607194113
transform 1 0 9476 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_85
timestamp 1607194113
transform 1 0 8924 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1009_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 9568 0 1 15776
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_25_119
timestamp 1607194113
transform 1 0 12052 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_107
timestamp 1607194113
transform 1 0 10948 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A2
timestamp 1607194113
transform 1 0 10764 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_132
timestamp 1607194113
transform 1 0 13248 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A
timestamp 1607194113
transform 1 0 13064 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1607194113
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _1007_
timestamp 1607194113
transform 1 0 12420 0 1 15776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_25_156
timestamp 1607194113
transform 1 0 15456 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_144
timestamp 1607194113
transform 1 0 14352 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_168
timestamp 1607194113
transform 1 0 16560 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_180
timestamp 1607194113
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1607194113
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_4  _0981_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 18032 0 1 15776
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_25_211
timestamp 1607194113
transform 1 0 20516 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_203
timestamp 1607194113
transform 1 0 19780 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__A1
timestamp 1607194113
transform 1 0 19596 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__B1
timestamp 1607194113
transform 1 0 20700 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1222_
timestamp 1607194113
transform 1 0 20884 0 1 15776
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_25_231
timestamp 1607194113
transform 1 0 22356 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_243
timestamp 1607194113
transform 1 0 23460 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1607194113
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_15
timestamp 1607194113
transform 1 0 2484 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1607194113
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_15
timestamp 1607194113
transform 1 0 2484 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1607194113
transform 1 0 1380 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__A
timestamp 1607194113
transform 1 0 2760 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A
timestamp 1607194113
transform 1 0 2668 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1607194113
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1607194113
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1607194113
transform 1 0 2852 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_22
timestamp 1607194113
transform 1 0 3128 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_23
timestamp 1607194113
transform 1 0 3220 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0668_
timestamp 1607194113
transform 1 0 2944 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_34
timestamp 1607194113
transform 1 0 4232 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_36
timestamp 1607194113
transform 1 0 4416 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_32
timestamp 1607194113
transform 1 0 4048 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__C
timestamp 1607194113
transform 1 0 4508 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1607194113
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0906_
timestamp 1607194113
transform 1 0 3864 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A
timestamp 1607194113
transform 1 0 4692 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1607194113
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1607194113
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_26_50
timestamp 1607194113
transform 1 0 5704 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__B
timestamp 1607194113
transform 1 0 4784 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _0948_
timestamp 1607194113
transform 1 0 6440 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _0866_
timestamp 1607194113
transform 1 0 4876 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _0669_
timestamp 1607194113
transform 1 0 4968 0 1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_27_79
timestamp 1607194113
transform 1 0 8372 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_79
timestamp 1607194113
transform 1 0 8372 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_67
timestamp 1607194113
transform 1 0 7268 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__A
timestamp 1607194113
transform 1 0 7820 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1607194113
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _0942_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 6808 0 1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _0679_
timestamp 1607194113
transform 1 0 8004 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_91
timestamp 1607194113
transform 1 0 9476 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_93
timestamp 1607194113
transform 1 0 9660 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1607194113
transform 1 0 9476 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__A
timestamp 1607194113
transform 1 0 10028 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1607194113
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1018_
timestamp 1607194113
transform 1 0 10212 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0908_
timestamp 1607194113
transform 1 0 9108 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_114
timestamp 1607194113
transform 1 0 11592 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_103
timestamp 1607194113
transform 1 0 10580 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_110
timestamp 1607194113
transform 1 0 11224 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_102
timestamp 1607194113
transform 1 0 10488 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__A
timestamp 1607194113
transform 1 0 10764 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1021_
timestamp 1607194113
transform 1 0 11408 0 -1 16864
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _1017_
timestamp 1607194113
transform 1 0 10948 0 1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_27_135
timestamp 1607194113
transform 1 0 13524 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1607194113
transform 1 0 12420 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_136
timestamp 1607194113
transform 1 0 13616 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_121
timestamp 1607194113
transform 1 0 12236 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1607194113
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0957_
timestamp 1607194113
transform 1 0 12972 0 -1 16864
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_27_141
timestamp 1607194113
transform 1 0 14076 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1607194113
transform 1 0 15272 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1607194113
transform 1 0 15088 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_148
timestamp 1607194113
transform 1 0 14720 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1607194113
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_4  _0989_
timestamp 1607194113
transform 1 0 14168 0 1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_8  FILLER_27_175
timestamp 1607194113
transform 1 0 17204 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_169
timestamp 1607194113
transform 1 0 16652 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_161
timestamp 1607194113
transform 1 0 15916 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_166
timestamp 1607194113
transform 1 0 16376 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A1
timestamp 1607194113
transform 1 0 15732 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0980_
timestamp 1607194113
transform 1 0 16928 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_4  _0967_
timestamp 1607194113
transform 1 0 16652 0 -1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_26_198
timestamp 1607194113
transform 1 0 19320 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_190
timestamp 1607194113
transform 1 0 18584 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A1
timestamp 1607194113
transform 1 0 18400 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A2
timestamp 1607194113
transform 1 0 18216 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1607194113
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_4  _0974_
timestamp 1607194113
transform 1 0 18032 0 1 16864
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _0943_
timestamp 1607194113
transform 1 0 18952 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1607194113
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1607194113
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A1
timestamp 1607194113
transform 1 0 19780 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__B2
timestamp 1607194113
transform 1 0 19964 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__A2
timestamp 1607194113
transform 1 0 20148 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A2
timestamp 1607194113
transform 1 0 19596 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1607194113
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0953_
timestamp 1607194113
transform 1 0 20332 0 1 16864
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_27_235
timestamp 1607194113
transform 1 0 22724 0 1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_223
timestamp 1607194113
transform 1 0 21620 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_238
timestamp 1607194113
transform 1 0 23000 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_227
timestamp 1607194113
transform 1 0 21988 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__A
timestamp 1607194113
transform 1 0 22816 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0947_
timestamp 1607194113
transform 1 0 22540 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_clk_i
timestamp 1607194113
transform 1 0 23276 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1607194113
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1607194113
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1607194113
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1607194113
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_39
timestamp 1607194113
transform 1 0 4692 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_32
timestamp 1607194113
transform 1 0 4048 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1607194113
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1607194113
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0905_
timestamp 1607194113
transform 1 0 4324 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_51
timestamp 1607194113
transform 1 0 5796 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0907_
timestamp 1607194113
transform 1 0 6532 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0678_
timestamp 1607194113
transform 1 0 5428 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_68
timestamp 1607194113
transform 1 0 7360 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _0941_
timestamp 1607194113
transform 1 0 8096 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1607194113
transform 1 0 9660 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1607194113
transform 1 0 9476 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_83
timestamp 1607194113
transform 1 0 8740 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1607194113
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1607194113
transform 1 0 11868 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1607194113
transform 1 0 10764 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_133
timestamp 1607194113
transform 1 0 13340 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_129
timestamp 1607194113
transform 1 0 12972 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0988_
timestamp 1607194113
transform 1 0 13064 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1607194113
transform 1 0 15272 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_145
timestamp 1607194113
transform 1 0 14444 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1607194113
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_178
timestamp 1607194113
transform 1 0 17480 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1607194113
transform 1 0 16376 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_194
timestamp 1607194113
transform 1 0 18952 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_184
timestamp 1607194113
transform 1 0 18032 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__A
timestamp 1607194113
transform 1 0 18768 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0977_
timestamp 1607194113
transform 1 0 18124 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1607194113
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_211
timestamp 1607194113
transform 1 0 20516 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_203
timestamp 1607194113
transform 1 0 19780 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1607194113
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp 1607194113
transform 1 0 19504 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_227
timestamp 1607194113
transform 1 0 21988 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__A
timestamp 1607194113
transform 1 0 23000 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1607194113
transform 1 0 22724 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_240
timestamp 1607194113
transform 1 0 23184 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1607194113
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1607194113
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1497_
timestamp 1607194113
transform 1 0 2484 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_29_38
timestamp 1607194113
transform 1 0 4600 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1497__CLK
timestamp 1607194113
transform 1 0 4416 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1497__D
timestamp 1607194113
transform 1 0 4232 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_53
timestamp 1607194113
transform 1 0 5980 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_46
timestamp 1607194113
transform 1 0 5336 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0681_
timestamp 1607194113
transform 1 0 5612 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_68
timestamp 1607194113
transform 1 0 7360 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_62
timestamp 1607194113
transform 1 0 6808 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1607194113
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a2111o_4  _1001_
timestamp 1607194113
transform 1 0 7452 0 1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_29_90
timestamp 1607194113
transform 1 0 9384 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__A1
timestamp 1607194113
transform 1 0 9200 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__A2
timestamp 1607194113
transform 1 0 9016 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_109
timestamp 1607194113
transform 1 0 11132 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_102
timestamp 1607194113
transform 1 0 10488 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0949_
timestamp 1607194113
transform 1 0 10764 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_131
timestamp 1607194113
transform 1 0 13156 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_123
timestamp 1607194113
transform 1 0 12420 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_121
timestamp 1607194113
transform 1 0 12236 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1607194113
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _1000_
timestamp 1607194113
transform 1 0 13248 0 1 17952
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_29_151
timestamp 1607194113
transform 1 0 14996 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__B1
timestamp 1607194113
transform 1 0 14812 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_173
timestamp 1607194113
transform 1 0 17020 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_163
timestamp 1607194113
transform 1 0 16100 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A
timestamp 1607194113
transform 1 0 16192 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0962_
timestamp 1607194113
transform 1 0 16376 0 1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_29_184
timestamp 1607194113
transform 1 0 18032 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1607194113
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A2
timestamp 1607194113
transform 1 0 18584 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__B2
timestamp 1607194113
transform 1 0 18768 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1607194113
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0965_
timestamp 1607194113
transform 1 0 18952 0 1 17952
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_29_208
timestamp 1607194113
transform 1 0 20240 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__B1
timestamp 1607194113
transform 1 0 20792 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1223_
timestamp 1607194113
transform 1 0 20976 0 1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1607194113
transform 1 0 22448 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1607194113
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1607194113
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1607194113
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1607194113
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1607194113
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1607194113
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1607194113
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_59
timestamp 1607194113
transform 1 0 6532 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_30_44
timestamp 1607194113
transform 1 0 5152 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__and4_4  _1282_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 5704 0 -1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_4  _0995_
timestamp 1607194113
transform 1 0 7268 0 -1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1607194113
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_88
timestamp 1607194113
transform 1 0 9200 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A1
timestamp 1607194113
transform 1 0 9016 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A2
timestamp 1607194113
transform 1 0 8832 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1607194113
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_117
timestamp 1607194113
transform 1 0 11868 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1607194113
transform 1 0 10764 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_125
timestamp 1607194113
transform 1 0 12604 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_4  _0994_
timestamp 1607194113
transform 1 0 12880 0 -1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_6  FILLER_30_147
timestamp 1607194113
transform 1 0 14628 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__A3
timestamp 1607194113
transform 1 0 14444 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1607194113
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0984_
timestamp 1607194113
transform 1 0 15272 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_30_175
timestamp 1607194113
transform 1 0 17204 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_163
timestamp 1607194113
transform 1 0 16100 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A
timestamp 1607194113
transform 1 0 15916 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_192
timestamp 1607194113
transform 1 0 18768 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__A
timestamp 1607194113
transform 1 0 18584 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0970_
timestamp 1607194113
transform 1 0 17940 0 -1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_30_215
timestamp 1607194113
transform 1 0 20884 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_212
timestamp 1607194113
transform 1 0 20608 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_204
timestamp 1607194113
transform 1 0 19872 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1607194113
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_223
timestamp 1607194113
transform 1 0 21620 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1407__CLK
timestamp 1607194113
transform 1 0 21712 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1407_
timestamp 1607194113
transform 1 0 21896 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1607194113
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1607194113
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1607194113
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1607194113
transform 1 0 4692 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1607194113
transform 1 0 3588 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1607194113
transform 1 0 6532 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1607194113
transform 1 0 5796 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_73
timestamp 1607194113
transform 1 0 7820 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_62
timestamp 1607194113
transform 1 0 6808 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1607194113
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _0993_
timestamp 1607194113
transform 1 0 6992 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_31_92
timestamp 1607194113
transform 1 0 9568 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__D
timestamp 1607194113
transform 1 0 9384 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _1158_
timestamp 1607194113
transform 1 0 10120 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _0999_
timestamp 1607194113
transform 1 0 8556 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_31_119
timestamp 1607194113
transform 1 0 12052 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_107
timestamp 1607194113
transform 1 0 10948 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_129
timestamp 1607194113
transform 1 0 12972 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__A
timestamp 1607194113
transform 1 0 12788 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__A2
timestamp 1607194113
transform 1 0 13156 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__A3
timestamp 1607194113
transform 1 0 13340 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1607194113
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _1272_
timestamp 1607194113
transform 1 0 13524 0 1 19040
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _0950_
timestamp 1607194113
transform 1 0 12420 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_154
timestamp 1607194113
transform 1 0 15272 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__A
timestamp 1607194113
transform 1 0 15640 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1272__B1
timestamp 1607194113
transform 1 0 15088 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_167
timestamp 1607194113
transform 1 0 16468 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _0946_
timestamp 1607194113
transform 1 0 15824 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_31_187
timestamp 1607194113
transform 1 0 18308 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_179
timestamp 1607194113
transform 1 0 17572 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1607194113
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1607194113
transform 1 0 18032 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_203
timestamp 1607194113
transform 1 0 19780 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_199
timestamp 1607194113
transform 1 0 19412 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__A2_N
timestamp 1607194113
transform 1 0 19872 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__B2
timestamp 1607194113
transform 1 0 20056 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__B1
timestamp 1607194113
transform 1 0 20240 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1209_
timestamp 1607194113
transform 1 0 20424 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_31_238
timestamp 1607194113
transform 1 0 23000 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_226
timestamp 1607194113
transform 1 0 21896 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1607194113
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1607194113
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1607194113
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1607194113
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1607194113
transform 1 0 4048 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1607194113
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1607194113
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_56
timestamp 1607194113
transform 1 0 6256 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_44
timestamp 1607194113
transform 1 0 5152 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__D
timestamp 1607194113
transform 1 0 6072 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _1219_
timestamp 1607194113
transform 1 0 5244 0 -1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_32_79
timestamp 1607194113
transform 1 0 8372 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__A2
timestamp 1607194113
transform 1 0 8188 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__B1
timestamp 1607194113
transform 1 0 8004 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _0992_
timestamp 1607194113
transform 1 0 6808 0 -1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1607194113
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_91
timestamp 1607194113
transform 1 0 9476 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1607194113
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_117
timestamp 1607194113
transform 1 0 11868 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1607194113
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_123
timestamp 1607194113
transform 1 0 12420 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__A2
timestamp 1607194113
transform 1 0 12512 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__A3
timestamp 1607194113
transform 1 0 12696 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _1271_
timestamp 1607194113
transform 1 0 12880 0 -1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_32_158
timestamp 1607194113
transform 1 0 15640 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_147
timestamp 1607194113
transform 1 0 14628 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1271__B1
timestamp 1607194113
transform 1 0 14444 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1607194113
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0961_
timestamp 1607194113
transform 1 0 15272 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_170
timestamp 1607194113
transform 1 0 16744 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_194
timestamp 1607194113
transform 1 0 18952 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_182
timestamp 1607194113
transform 1 0 17848 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_215
timestamp 1607194113
transform 1 0 20884 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_206
timestamp 1607194113
transform 1 0 20056 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1417__CLK
timestamp 1607194113
transform 1 0 20608 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1607194113
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1417_
timestamp 1607194113
transform 1 0 20976 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_32_235
timestamp 1607194113
transform 1 0 22724 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1607194113
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1607194113
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1607194113
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1607194113
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1607194113
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1498_
timestamp 1607194113
transform 1 0 2484 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1607194113
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1607194113
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_36
timestamp 1607194113
transform 1 0 4416 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1498__CLK
timestamp 1607194113
transform 1 0 4232 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1607194113
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_56
timestamp 1607194113
transform 1 0 6256 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1607194113
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_48
timestamp 1607194113
transform 1 0 5520 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_62
timestamp 1607194113
transform 1 0 6808 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_62
timestamp 1607194113
transform 1 0 6808 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_60
timestamp 1607194113
transform 1 0 6624 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__D
timestamp 1607194113
transform 1 0 6900 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1607194113
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _0682_
timestamp 1607194113
transform 1 0 7084 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A2
timestamp 1607194113
transform 1 0 8280 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__B1
timestamp 1607194113
transform 1 0 8096 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_74
timestamp 1607194113
transform 1 0 7912 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_4  _0998_
timestamp 1607194113
transform 1 0 6900 0 1 20128
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1607194113
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_86
timestamp 1607194113
transform 1 0 9016 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_92
timestamp 1607194113
transform 1 0 9568 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_80
timestamp 1607194113
transform 1 0 8464 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1607194113
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_117
timestamp 1607194113
transform 1 0 11868 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1607194113
transform 1 0 10764 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_116
timestamp 1607194113
transform 1 0 11776 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_104
timestamp 1607194113
transform 1 0 10672 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_123
timestamp 1607194113
transform 1 0 12420 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_135
timestamp 1607194113
transform 1 0 13524 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1607194113
transform 1 0 12420 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1376__CLK
timestamp 1607194113
transform 1 0 12512 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1375__CLK
timestamp 1607194113
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1607194113
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1376_
timestamp 1607194113
transform 1 0 12696 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1375_
timestamp 1607194113
transform 1 0 13800 0 1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_34_158
timestamp 1607194113
transform 1 0 15640 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_145
timestamp 1607194113
transform 1 0 14444 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_157
timestamp 1607194113
transform 1 0 15548 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1607194113
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0945_
timestamp 1607194113
transform 1 0 15272 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_170
timestamp 1607194113
transform 1 0 16744 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1607194113
transform 1 0 16652 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_194
timestamp 1607194113
transform 1 0 18952 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_182
timestamp 1607194113
transform 1 0 17848 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_196
timestamp 1607194113
transform 1 0 19136 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1607194113
transform 1 0 18032 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_181
timestamp 1607194113
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1607194113
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_215
timestamp 1607194113
transform 1 0 20884 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_206
timestamp 1607194113
transform 1 0 20056 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_200
timestamp 1607194113
transform 1 0 19504 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__A2_N
timestamp 1607194113
transform 1 0 19596 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__B2
timestamp 1607194113
transform 1 0 19780 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__B1
timestamp 1607194113
transform 1 0 19964 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1607194113
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1208_
timestamp 1607194113
transform 1 0 20148 0 1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_33_236
timestamp 1607194113
transform 1 0 22816 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_223
timestamp 1607194113
transform 1 0 21620 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1416__CLK
timestamp 1607194113
transform 1 0 21436 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A
timestamp 1607194113
transform 1 0 22632 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1416_
timestamp 1607194113
transform 1 0 21620 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0951_
timestamp 1607194113
transform 1 0 22356 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_242
timestamp 1607194113
transform 1 0 23368 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1607194113
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1607194113
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1607194113
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1499_
timestamp 1607194113
transform 1 0 2484 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_35_38
timestamp 1607194113
transform 1 0 4600 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1499__CLK
timestamp 1607194113
transform 1 0 4416 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1499__D
timestamp 1607194113
transform 1 0 4232 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_35_58
timestamp 1607194113
transform 1 0 6440 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_50
timestamp 1607194113
transform 1 0 5704 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_79
timestamp 1607194113
transform 1 0 8372 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_74
timestamp 1607194113
transform 1 0 7912 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_66
timestamp 1607194113
transform 1 0 7176 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1607194113
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1025_
timestamp 1607194113
transform 1 0 8004 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0670_
timestamp 1607194113
transform 1 0 6808 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_91
timestamp 1607194113
transform 1 0 9476 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1220_
timestamp 1607194113
transform 1 0 9108 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_119
timestamp 1607194113
transform 1 0 12052 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_115
timestamp 1607194113
transform 1 0 11684 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_103
timestamp 1607194113
transform 1 0 10580 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1372__CLK
timestamp 1607194113
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1607194113
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1372_
timestamp 1607194113
transform 1 0 12420 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_35_154
timestamp 1607194113
transform 1 0 15272 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_142
timestamp 1607194113
transform 1 0 14168 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_178
timestamp 1607194113
transform 1 0 17480 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_166
timestamp 1607194113
transform 1 0 16376 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_184
timestamp 1607194113
transform 1 0 18032 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_182
timestamp 1607194113
transform 1 0 17848 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__B1
timestamp 1607194113
transform 1 0 18216 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1607194113
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1225_
timestamp 1607194113
transform 1 0 18400 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_35_216
timestamp 1607194113
transform 1 0 20976 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_204
timestamp 1607194113
transform 1 0 19872 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_234
timestamp 1607194113
transform 1 0 22632 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_228
timestamp 1607194113
transform 1 0 22080 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__A
timestamp 1607194113
transform 1 0 22448 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1607194113
transform 1 0 22172 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_242
timestamp 1607194113
transform 1 0 23368 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1607194113
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1607194113
transform 1 0 2484 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1607194113
transform 1 0 1380 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1607194113
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1607194113
transform 1 0 3588 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1607194113
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1500_
timestamp 1607194113
transform 1 0 4048 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_36_53
timestamp 1607194113
transform 1 0 5980 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1500__CLK
timestamp 1607194113
transform 1 0 5796 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1231__B1
timestamp 1607194113
transform 1 0 6532 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_77
timestamp 1607194113
transform 1 0 8188 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__a2bb2o_4  _1231_
timestamp 1607194113
transform 1 0 6716 0 -1 22304
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_36_97
timestamp 1607194113
transform 1 0 10028 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_89
timestamp 1607194113
transform 1 0 9292 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1607194113
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1224_
timestamp 1607194113
transform 1 0 9660 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_116
timestamp 1607194113
transform 1 0 11776 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_109
timestamp 1607194113
transform 1 0 11132 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1016_
timestamp 1607194113
transform 1 0 11500 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__A2
timestamp 1607194113
transform 1 0 12144 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__A3
timestamp 1607194113
transform 1 0 12328 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _1275_
timestamp 1607194113
transform 1 0 12512 0 -1 22304
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_12  FILLER_36_154
timestamp 1607194113
transform 1 0 15272 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_151
timestamp 1607194113
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_143
timestamp 1607194113
transform 1 0 14260 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1275__B1
timestamp 1607194113
transform 1 0 14076 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1607194113
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_174
timestamp 1607194113
transform 1 0 17112 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_166
timestamp 1607194113
transform 1 0 16376 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1221_
timestamp 1607194113
transform 1 0 17296 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_180
timestamp 1607194113
transform 1 0 17664 0 -1 22304
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A2
timestamp 1607194113
transform 1 0 18216 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__B2
timestamp 1607194113
transform 1 0 18400 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0972_
timestamp 1607194113
transform 1 0 18584 0 -1 22304
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_36_206
timestamp 1607194113
transform 1 0 20056 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__A
timestamp 1607194113
transform 1 0 21160 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A1
timestamp 1607194113
transform 1 0 19872 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1607194113
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1607194113
transform 1 0 20884 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_232
timestamp 1607194113
transform 1 0 22448 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_220
timestamp 1607194113
transform 1 0 21344 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_244
timestamp 1607194113
transform 1 0 23552 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1607194113
transform 1 0 1380 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1607194113
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1482_
timestamp 1607194113
transform 1 0 2484 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_37_38
timestamp 1607194113
transform 1 0 4600 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1482__CLK
timestamp 1607194113
transform 1 0 4416 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1482__D
timestamp 1607194113
transform 1 0 4232 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_58
timestamp 1607194113
transform 1 0 6440 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_50
timestamp 1607194113
transform 1 0 5704 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_66
timestamp 1607194113
transform 1 0 7176 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_62
timestamp 1607194113
transform 1 0 6808 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1607194113
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1401_
timestamp 1607194113
transform 1 0 7268 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_37_97
timestamp 1607194113
transform 1 0 10028 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_88
timestamp 1607194113
transform 1 0 9200 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1401__CLK
timestamp 1607194113
transform 1 0 9016 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A
timestamp 1607194113
transform 1 0 9568 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp 1607194113
transform 1 0 9752 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_117
timestamp 1607194113
transform 1 0 11868 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_109
timestamp 1607194113
transform 1 0 11132 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__A2
timestamp 1607194113
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__B1
timestamp 1607194113
transform 1 0 13708 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1607194113
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _1015_
timestamp 1607194113
transform 1 0 12420 0 1 22304
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_37_151
timestamp 1607194113
transform 1 0 14996 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_139
timestamp 1607194113
transform 1 0 13892 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_175
timestamp 1607194113
transform 1 0 17204 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_163
timestamp 1607194113
transform 1 0 16100 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_37_196
timestamp 1607194113
transform 1 0 19136 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1607194113
transform 1 0 18032 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1607194113
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1406__CLK
timestamp 1607194113
transform 1 0 19412 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1406_
timestamp 1607194113
transform 1 0 19596 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_37_232
timestamp 1607194113
transform 1 0 22448 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_220
timestamp 1607194113
transform 1 0 21344 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1607194113
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1607194113
transform 1 0 2484 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1607194113
transform 1 0 1380 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1607194113
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1607194113
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1607194113
transform 1 0 3588 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1607194113
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_44
timestamp 1607194113
transform 1 0 5152 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1230__B1
timestamp 1607194113
transform 1 0 5244 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1230_
timestamp 1607194113
transform 1 0 5428 0 -1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_38_75
timestamp 1607194113
transform 1 0 8004 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_63
timestamp 1607194113
transform 1 0 6900 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1228_
timestamp 1607194113
transform 1 0 7636 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_96
timestamp 1607194113
transform 1 0 9936 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_91
timestamp 1607194113
transform 1 0 9476 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_87
timestamp 1607194113
transform 1 0 9108 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1607194113
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1024_
timestamp 1607194113
transform 1 0 9660 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_108
timestamp 1607194113
transform 1 0 11040 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__B2
timestamp 1607194113
transform 1 0 11592 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0987_
timestamp 1607194113
transform 1 0 11776 0 -1 23392
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_38_130
timestamp 1607194113
transform 1 0 13064 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_154
timestamp 1607194113
transform 1 0 15272 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_150
timestamp 1607194113
transform 1 0 14904 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_142
timestamp 1607194113
transform 1 0 14168 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1607194113
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_178
timestamp 1607194113
transform 1 0 17480 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_38_166
timestamp 1607194113
transform 1 0 16376 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1405_
timestamp 1607194113
transform 1 0 18032 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_38_215
timestamp 1607194113
transform 1 0 20884 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_213
timestamp 1607194113
transform 1 0 20700 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_205
timestamp 1607194113
transform 1 0 19964 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1405__CLK
timestamp 1607194113
transform 1 0 19780 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1607194113
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_223
timestamp 1607194113
transform 1 0 21620 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1356__CLK
timestamp 1607194113
transform 1 0 21712 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1356_
timestamp 1607194113
transform 1 0 21896 0 -1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1607194113
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1607194113
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1607194113
transform 1 0 1380 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1607194113
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1607194113
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1501_
timestamp 1607194113
transform 1 0 2484 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_40_32
timestamp 1607194113
transform 1 0 4048 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1607194113
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_36
timestamp 1607194113
transform 1 0 4416 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1501__CLK
timestamp 1607194113
transform 1 0 4232 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1607194113
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_40
timestamp 1607194113
transform 1 0 4784 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_48
timestamp 1607194113
transform 1 0 5520 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1229__B1
timestamp 1607194113
transform 1 0 5060 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1229_
timestamp 1607194113
transform 1 0 5244 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_40_61
timestamp 1607194113
transform 1 0 6716 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_66
timestamp 1607194113
transform 1 0 7176 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_62
timestamp 1607194113
transform 1 0 6808 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_60
timestamp 1607194113
transform 1 0 6624 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A
timestamp 1607194113
transform 1 0 7268 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1607194113
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0997_
timestamp 1607194113
transform 1 0 7268 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1607194113
transform 1 0 7452 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__A
timestamp 1607194113
transform 1 0 7544 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_72
timestamp 1607194113
transform 1 0 7728 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_72
timestamp 1607194113
transform 1 0 7728 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_93
timestamp 1607194113
transform 1 0 9660 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_84
timestamp 1607194113
transform 1 0 8832 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_84
timestamp 1607194113
transform 1 0 8832 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__B1
timestamp 1607194113
transform 1 0 9936 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1607194113
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1227_
timestamp 1607194113
transform 1 0 10120 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_40_105
timestamp 1607194113
transform 1 0 10764 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_114
timestamp 1607194113
transform 1 0 11592 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1404_
timestamp 1607194113
transform 1 0 10856 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_40_127
timestamp 1607194113
transform 1 0 12788 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_127
timestamp 1607194113
transform 1 0 12788 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1404__CLK
timestamp 1607194113
transform 1 0 12604 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1232__B1
timestamp 1607194113
transform 1 0 13524 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1607194113
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1232_
timestamp 1607194113
transform 1 0 13708 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _0952_
timestamp 1607194113
transform 1 0 12420 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_139
timestamp 1607194113
transform 1 0 13892 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_153
timestamp 1607194113
transform 1 0 15180 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1400__CLK
timestamp 1607194113
transform 1 0 14996 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1607194113
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1400_
timestamp 1607194113
transform 1 0 15272 0 -1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_40_173
timestamp 1607194113
transform 1 0 17020 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_177
timestamp 1607194113
transform 1 0 17388 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_165
timestamp 1607194113
transform 1 0 16284 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A2
timestamp 1607194113
transform 1 0 17756 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__B2
timestamp 1607194113
transform 1 0 17940 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__B1
timestamp 1607194113
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1607194113
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1226_
timestamp 1607194113
transform 1 0 18032 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__o22a_4  _0979_
timestamp 1607194113
transform 1 0 18124 0 -1 24480
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_39_200
timestamp 1607194113
transform 1 0 19504 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A
timestamp 1607194113
transform 1 0 20056 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A1
timestamp 1607194113
transform 1 0 19412 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1607194113
transform 1 0 20240 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_218
timestamp 1607194113
transform 1 0 21160 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_213
timestamp 1607194113
transform 1 0 20700 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_39_217
timestamp 1607194113
transform 1 0 21068 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_211
timestamp 1607194113
transform 1 0 20516 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1311__B1
timestamp 1607194113
transform 1 0 21160 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1607194113
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1314_
timestamp 1607194113
transform 1 0 20884 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_201
timestamp 1607194113
transform 1 0 19596 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_229
timestamp 1607194113
transform 1 0 22172 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_39_236
timestamp 1607194113
transform 1 0 22816 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_clk_i
timestamp 1607194113
transform 1 0 22908 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1312_
timestamp 1607194113
transform 1 0 21896 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1311_
timestamp 1607194113
transform 1 0 21344 0 1 23392
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_40_240
timestamp 1607194113
transform 1 0 23184 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1607194113
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1308_
timestamp 1607194113
transform 1 0 23368 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1607194113
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1607194113
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1502_
timestamp 1607194113
transform 1 0 2484 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_41_38
timestamp 1607194113
transform 1 0 4600 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1502__CLK
timestamp 1607194113
transform 1 0 4416 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1502__D
timestamp 1607194113
transform 1 0 4232 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_58
timestamp 1607194113
transform 1 0 6440 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_50
timestamp 1607194113
transform 1 0 5704 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1607194113
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1402_
timestamp 1607194113
transform 1 0 6808 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_41_95
timestamp 1607194113
transform 1 0 9844 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_83
timestamp 1607194113
transform 1 0 8740 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1402__CLK
timestamp 1607194113
transform 1 0 8556 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_113
timestamp 1607194113
transform 1 0 11500 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_107
timestamp 1607194113
transform 1 0 10948 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_clk_i
timestamp 1607194113
transform 1 0 11224 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_41_132
timestamp 1607194113
transform 1 0 13248 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_128
timestamp 1607194113
transform 1 0 12880 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_121
timestamp 1607194113
transform 1 0 12236 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A
timestamp 1607194113
transform 1 0 12696 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1315__A
timestamp 1607194113
transform 1 0 13340 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1607194113
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1315_
timestamp 1607194113
transform 1 0 13524 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1607194113
transform 1 0 12420 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_41_151
timestamp 1607194113
transform 1 0 14996 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_139
timestamp 1607194113
transform 1 0 13892 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__A
timestamp 1607194113
transform 1 0 15548 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1014_
timestamp 1607194113
transform 1 0 15272 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_171
timestamp 1607194113
transform 1 0 16836 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_159
timestamp 1607194113
transform 1 0 15732 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1607194113
transform 1 0 18032 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1309__A
timestamp 1607194113
transform 1 0 19136 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1607194113
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1309_
timestamp 1607194113
transform 1 0 19320 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_214
timestamp 1607194113
transform 1 0 20792 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_202
timestamp 1607194113
transform 1 0 19688 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1355__CLK
timestamp 1607194113
transform 1 0 20884 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1355_
timestamp 1607194113
transform 1 0 21068 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_41_236
timestamp 1607194113
transform 1 0 22816 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1607194113
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1607194113
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1607194113
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1607194113
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1607194113
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1607194113
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1607194113
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_44
timestamp 1607194113
transform 1 0 5152 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _1403_
timestamp 1607194113
transform 1 0 5704 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_42_71
timestamp 1607194113
transform 1 0 7636 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1403__CLK
timestamp 1607194113
transform 1 0 7452 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_93
timestamp 1607194113
transform 1 0 9660 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_91
timestamp 1607194113
transform 1 0 9476 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_83
timestamp 1607194113
transform 1 0 8740 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1607194113
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_111
timestamp 1607194113
transform 1 0 11316 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_105
timestamp 1607194113
transform 1 0 10764 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_4  _1171_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 11408 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_42_136
timestamp 1607194113
transform 1 0 13616 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_123
timestamp 1607194113
transform 1 0 12420 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__A
timestamp 1607194113
transform 1 0 12236 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1233__A
timestamp 1607194113
transform 1 0 12788 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1233_
timestamp 1607194113
transform 1 0 12972 0 -1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_42_154
timestamp 1607194113
transform 1 0 15272 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_147
timestamp 1607194113
transform 1 0 14628 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_clk_i
timestamp 1607194113
transform 1 0 14352 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1607194113
transform 1 0 15180 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_178
timestamp 1607194113
transform 1 0 17480 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_42_166
timestamp 1607194113
transform 1 0 16376 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_184
timestamp 1607194113
transform 1 0 18032 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1316__B1
timestamp 1607194113
transform 1 0 18124 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1316_
timestamp 1607194113
transform 1 0 18308 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_42_211
timestamp 1607194113
transform 1 0 20516 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_203
timestamp 1607194113
transform 1 0 19780 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1313__B1
timestamp 1607194113
transform 1 0 20608 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1607194113
transform 1 0 20792 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1313_
timestamp 1607194113
transform 1 0 20884 0 -1 25568
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_42_231
timestamp 1607194113
transform 1 0 22356 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_243
timestamp 1607194113
transform 1 0 23460 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1607194113
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1607194113
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1503_
timestamp 1607194113
transform 1 0 2484 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_43_36
timestamp 1607194113
transform 1 0 4416 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1503__CLK
timestamp 1607194113
transform 1 0 4232 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_48
timestamp 1607194113
transform 1 0 5520 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_70
timestamp 1607194113
transform 1 0 7544 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_62
timestamp 1607194113
transform 1 0 6808 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_60
timestamp 1607194113
transform 1 0 6624 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1607194113
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0683_
timestamp 1607194113
transform 1 0 7636 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_43_94
timestamp 1607194113
transform 1 0 9752 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_82
timestamp 1607194113
transform 1 0 8648 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A
timestamp 1607194113
transform 1 0 8464 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_118
timestamp 1607194113
transform 1 0 11960 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_106
timestamp 1607194113
transform 1 0 10856 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_127
timestamp 1607194113
transform 1 0 12788 0 1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1353__CLK
timestamp 1607194113
transform 1 0 13340 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1607194113
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1353_
timestamp 1607194113
transform 1 0 13524 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _0671_
timestamp 1607194113
transform 1 0 12420 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_154
timestamp 1607194113
transform 1 0 15272 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_178
timestamp 1607194113
transform 1 0 17480 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_166
timestamp 1607194113
transform 1 0 16376 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_196
timestamp 1607194113
transform 1 0 19136 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_184
timestamp 1607194113
transform 1 0 18032 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_182
timestamp 1607194113
transform 1 0 17848 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1607194113
transform 1 0 17940 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1354__CLK
timestamp 1607194113
transform 1 0 19412 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1354_
timestamp 1607194113
transform 1 0 19596 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_43_232
timestamp 1607194113
transform 1 0 22448 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_220
timestamp 1607194113
transform 1 0 21344 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1607194113
transform 1 0 23552 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1607194113
transform 1 0 2484 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1607194113
transform 1 0 1380 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1607194113
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_32
timestamp 1607194113
transform 1 0 4048 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_27
timestamp 1607194113
transform 1 0 3588 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1607194113
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_56
timestamp 1607194113
transform 1 0 6256 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_44
timestamp 1607194113
transform 1 0 5152 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1517_
timestamp 1607194113
transform 1 0 6440 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_44_79
timestamp 1607194113
transform 1 0 8372 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1517__CLK
timestamp 1607194113
transform 1 0 8188 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_93
timestamp 1607194113
transform 1 0 9660 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_91
timestamp 1607194113
transform 1 0 9476 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1607194113
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_118
timestamp 1607194113
transform 1 0 11960 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_44_107
timestamp 1607194113
transform 1 0 10948 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A
timestamp 1607194113
transform 1 0 10396 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_clk_i
timestamp 1607194113
transform 1 0 11684 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0867_
timestamp 1607194113
transform 1 0 10580 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_126
timestamp 1607194113
transform 1 0 12696 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1318__B1
timestamp 1607194113
transform 1 0 12788 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1318_
timestamp 1607194113
transform 1 0 12972 0 -1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_44_157
timestamp 1607194113
transform 1 0 15548 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_145
timestamp 1607194113
transform 1 0 14444 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1607194113
transform 1 0 15180 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1317_
timestamp 1607194113
transform 1 0 15272 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_177
timestamp 1607194113
transform 1 0 17388 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_169
timestamp 1607194113
transform 1 0 16652 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1352__CLK
timestamp 1607194113
transform 1 0 19320 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1352_
timestamp 1607194113
transform 1 0 17572 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_44_212
timestamp 1607194113
transform 1 0 20608 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_200
timestamp 1607194113
transform 1 0 19504 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1607194113
transform 1 0 20792 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1310_
timestamp 1607194113
transform 1 0 20884 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_231
timestamp 1607194113
transform 1 0 22356 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_219
timestamp 1607194113
transform 1 0 21252 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_243
timestamp 1607194113
transform 1 0 23460 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_239
timestamp 1607194113
transform 1 0 23092 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0730_
timestamp 1607194113
transform 1 0 23184 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1607194113
transform 1 0 1380 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1607194113
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1504_
timestamp 1607194113
transform 1 0 2484 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_45_36
timestamp 1607194113
transform 1 0 4416 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1504__CLK
timestamp 1607194113
transform 1 0 4232 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_53
timestamp 1607194113
transform 1 0 5980 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_48
timestamp 1607194113
transform 1 0 5520 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0685_
timestamp 1607194113
transform 1 0 5704 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1607194113
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1412_
timestamp 1607194113
transform 1 0 6808 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_45_95
timestamp 1607194113
transform 1 0 9844 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_83
timestamp 1607194113
transform 1 0 8740 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1412__CLK
timestamp 1607194113
transform 1 0 8556 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_45_119
timestamp 1607194113
transform 1 0 12052 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_107
timestamp 1607194113
transform 1 0 10948 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__B1
timestamp 1607194113
transform 1 0 12144 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1607194113
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1214_
timestamp 1607194113
transform 1 0 12420 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_45_151
timestamp 1607194113
transform 1 0 14996 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_139
timestamp 1607194113
transform 1 0 13892 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_175
timestamp 1607194113
transform 1 0 17204 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_163
timestamp 1607194113
transform 1 0 16100 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_189
timestamp 1607194113
transform 1 0 18492 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_184
timestamp 1607194113
transform 1 0 18032 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1607194113
transform 1 0 17940 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1319_
timestamp 1607194113
transform 1 0 18216 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_45_201
timestamp 1607194113
transform 1 0 19596 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__B1
timestamp 1607194113
transform 1 0 19688 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1212_
timestamp 1607194113
transform 1 0 19872 0 1 26656
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_45_234
timestamp 1607194113
transform 1 0 22632 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_222
timestamp 1607194113
transform 1 0 21528 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__A1_N
timestamp 1607194113
transform 1 0 21344 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_242
timestamp 1607194113
transform 1 0 23368 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1607194113
transform 1 0 23552 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1607194113
transform 1 0 1380 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1607194113
transform 1 0 2484 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1607194113
transform 1 0 1380 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1607194113
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1607194113
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1505_
timestamp 1607194113
transform 1 0 2484 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_47_36
timestamp 1607194113
transform 1 0 4416 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_32
timestamp 1607194113
transform 1 0 4048 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_27
timestamp 1607194113
transform 1 0 3588 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1505__CLK
timestamp 1607194113
transform 1 0 4232 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1607194113
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_48
timestamp 1607194113
transform 1 0 5520 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_56
timestamp 1607194113
transform 1 0 6256 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_44
timestamp 1607194113
transform 1 0 5152 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_66
timestamp 1607194113
transform 1 0 7176 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_62
timestamp 1607194113
transform 1 0 6808 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_60
timestamp 1607194113
transform 1 0 6624 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_46_60
timestamp 1607194113
transform 1 0 6624 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__A1_N
timestamp 1607194113
transform 1 0 8372 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__B1
timestamp 1607194113
transform 1 0 6716 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1607194113
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1215_
timestamp 1607194113
transform 1 0 6900 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__a211o_4  _0684_
timestamp 1607194113
transform 1 0 7268 0 1 27744
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_47_93
timestamp 1607194113
transform 1 0 9660 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_81
timestamp 1607194113
transform 1 0 8556 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_96
timestamp 1607194113
transform 1 0 9936 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_89
timestamp 1607194113
transform 1 0 9292 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_81
timestamp 1607194113
transform 1 0 8556 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1607194113
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0735_
timestamp 1607194113
transform 1 0 9660 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_114
timestamp 1607194113
transform 1 0 11592 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_109
timestamp 1607194113
transform 1 0 11132 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_105
timestamp 1607194113
transform 1 0 10764 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_108
timestamp 1607194113
transform 1 0 11040 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1213_
timestamp 1607194113
transform 1 0 11224 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_123
timestamp 1607194113
transform 1 0 12420 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_120
timestamp 1607194113
transform 1 0 12144 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1413__CLK
timestamp 1607194113
transform 1 0 12512 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1607194113
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1413_
timestamp 1607194113
transform 1 0 12696 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1371_
timestamp 1607194113
transform 1 0 13524 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_47_156
timestamp 1607194113
transform 1 0 15456 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_145
timestamp 1607194113
transform 1 0 14444 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1371__CLK
timestamp 1607194113
transform 1 0 15272 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A
timestamp 1607194113
transform 1 0 15548 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1607194113
transform 1 0 15180 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1607194113
transform 1 0 15272 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_168
timestamp 1607194113
transform 1 0 16560 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_159
timestamp 1607194113
transform 1 0 15732 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1320__B1
timestamp 1607194113
transform 1 0 16284 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1320_
timestamp 1607194113
transform 1 0 16468 0 -1 27744
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_47_195
timestamp 1607194113
transform 1 0 19044 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_184
timestamp 1607194113
transform 1 0 18032 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_180
timestamp 1607194113
transform 1 0 17664 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_195
timestamp 1607194113
transform 1 0 19044 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_183
timestamp 1607194113
transform 1 0 17940 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_clk_i
timestamp 1607194113
transform 1 0 18768 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1607194113
transform 1 0 17940 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_47_207
timestamp 1607194113
transform 1 0 20148 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_215
timestamp 1607194113
transform 1 0 20884 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_213
timestamp 1607194113
transform 1 0 20700 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_207
timestamp 1607194113
transform 1 0 20148 0 -1 27744
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1351__CLK
timestamp 1607194113
transform 1 0 20240 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1607194113
transform 1 0 20792 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1351_
timestamp 1607194113
transform 1 0 20424 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_47_229
timestamp 1607194113
transform 1 0 22172 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1414__CLK
timestamp 1607194113
transform 1 0 21436 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1414_
timestamp 1607194113
transform 1 0 21620 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_47_241
timestamp 1607194113
transform 1 0 23276 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_46_242
timestamp 1607194113
transform 1 0 23368 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1607194113
transform 1 0 23552 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1607194113
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1607194113
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1607194113
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_27
timestamp 1607194113
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1607194113
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0921_
timestamp 1607194113
transform 1 0 4048 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_48_55
timestamp 1607194113
transform 1 0 6164 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_43
timestamp 1607194113
transform 1 0 5060 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__B
timestamp 1607194113
transform 1 0 4876 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_79
timestamp 1607194113
transform 1 0 8372 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_67
timestamp 1607194113
transform 1 0 7268 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_93
timestamp 1607194113
transform 1 0 9660 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_91
timestamp 1607194113
transform 1 0 9476 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1607194113
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_117
timestamp 1607194113
transform 1 0 11868 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_105
timestamp 1607194113
transform 1 0 10764 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_134
timestamp 1607194113
transform 1 0 13432 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_48_125
timestamp 1607194113
transform 1 0 12604 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1013_
timestamp 1607194113
transform 1 0 12788 0 -1 28832
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_48_157
timestamp 1607194113
transform 1 0 15548 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_145
timestamp 1607194113
transform 1 0 14444 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0944__A
timestamp 1607194113
transform 1 0 13984 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1607194113
transform 1 0 15180 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0944_
timestamp 1607194113
transform 1 0 14168 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0822_
timestamp 1607194113
transform 1 0 15272 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_169
timestamp 1607194113
transform 1 0 16652 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_165
timestamp 1607194113
transform 1 0 16284 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_clk_i
timestamp 1607194113
transform 1 0 16376 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_48_187
timestamp 1607194113
transform 1 0 18308 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_181
timestamp 1607194113
transform 1 0 17756 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1324__B1
timestamp 1607194113
transform 1 0 18400 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1324_
timestamp 1607194113
transform 1 0 18584 0 -1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_48_215
timestamp 1607194113
transform 1 0 20884 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_206
timestamp 1607194113
transform 1 0 20056 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1350__CLK
timestamp 1607194113
transform 1 0 20608 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1607194113
transform 1 0 20792 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1350_
timestamp 1607194113
transform 1 0 20976 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_48_235
timestamp 1607194113
transform 1 0 22724 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1607194113
transform 1 0 1380 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1607194113
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1506_
timestamp 1607194113
transform 1 0 2484 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_49_36
timestamp 1607194113
transform 1 0 4416 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1506__CLK
timestamp 1607194113
transform 1 0 4232 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_48
timestamp 1607194113
transform 1 0 5520 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_74
timestamp 1607194113
transform 1 0 7912 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_62
timestamp 1607194113
transform 1 0 6808 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_60
timestamp 1607194113
transform 1 0 6624 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1607194113
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1411_
timestamp 1607194113
transform 1 0 8188 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_49_98
timestamp 1607194113
transform 1 0 10120 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1411__CLK
timestamp 1607194113
transform 1 0 9936 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_119
timestamp 1607194113
transform 1 0 12052 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_107
timestamp 1607194113
transform 1 0 10948 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0675_
timestamp 1607194113
transform 1 0 10672 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_131
timestamp 1607194113
transform 1 0 13156 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_123
timestamp 1607194113
transform 1 0 12420 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__B1
timestamp 1607194113
transform 1 0 13340 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1607194113
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1277_
timestamp 1607194113
transform 1 0 13524 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_49_153
timestamp 1607194113
transform 1 0 15180 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1277__A1_N
timestamp 1607194113
transform 1 0 14996 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_177
timestamp 1607194113
transform 1 0 17388 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_165
timestamp 1607194113
transform 1 0 16284 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_184
timestamp 1607194113
transform 1 0 18032 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1322__B1
timestamp 1607194113
transform 1 0 19136 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1607194113
transform 1 0 17940 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1322_
timestamp 1607194113
transform 1 0 19320 0 1 28832
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_49_214
timestamp 1607194113
transform 1 0 20792 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_236
timestamp 1607194113
transform 1 0 22816 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_49_225
timestamp 1607194113
transform 1 0 21804 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1323_
timestamp 1607194113
transform 1 0 22540 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1321_
timestamp 1607194113
transform 1 0 21528 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1607194113
transform 1 0 23552 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_50_11
timestamp 1607194113
transform 1 0 2116 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_3
timestamp 1607194113
transform 1 0 1380 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1607194113
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0901_
timestamp 1607194113
transform 1 0 2392 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_50_25
timestamp 1607194113
transform 1 0 3404 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__B
timestamp 1607194113
transform 1 0 3220 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1607194113
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1507_
timestamp 1607194113
transform 1 0 4048 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1607194113
transform 1 0 5980 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1507__CLK
timestamp 1607194113
transform 1 0 5796 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_65
timestamp 1607194113
transform 1 0 7084 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__B1
timestamp 1607194113
transform 1 0 7176 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1216_
timestamp 1607194113
transform 1 0 7360 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_50_93
timestamp 1607194113
transform 1 0 9660 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_86
timestamp 1607194113
transform 1 0 9016 0 -1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__A1_N
timestamp 1607194113
transform 1 0 8832 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1607194113
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1518_
timestamp 1607194113
transform 1 0 9844 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_50_116
timestamp 1607194113
transform 1 0 11776 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1518__CLK
timestamp 1607194113
transform 1 0 11592 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_128
timestamp 1607194113
transform 1 0 12880 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_140
timestamp 1607194113
transform 1 0 13984 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__A2_N
timestamp 1607194113
transform 1 0 14996 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_clk_i
timestamp 1607194113
transform 1 0 14720 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1607194113
transform 1 0 15180 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1006_
timestamp 1607194113
transform 1 0 15272 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_50_172
timestamp 1607194113
transform 1 0 16928 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__A1_N
timestamp 1607194113
transform 1 0 16744 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_196
timestamp 1607194113
transform 1 0 19136 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_184
timestamp 1607194113
transform 1 0 18032 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_208
timestamp 1607194113
transform 1 0 20240 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__B1
timestamp 1607194113
transform 1 0 20608 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1607194113
transform 1 0 20792 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1274_
timestamp 1607194113
transform 1 0 20884 0 -1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_50_233
timestamp 1607194113
transform 1 0 22540 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1274__A1_N
timestamp 1607194113
transform 1 0 22356 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_15
timestamp 1607194113
transform 1 0 2484 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1607194113
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1607194113
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_51_37
timestamp 1607194113
transform 1 0 4508 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_51_23
timestamp 1607194113
transform 1 0 3220 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__B
timestamp 1607194113
transform 1 0 4324 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0899_
timestamp 1607194113
transform 1 0 3496 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_51_54
timestamp 1607194113
transform 1 0 6072 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__B
timestamp 1607194113
transform 1 0 5888 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0914_
timestamp 1607194113
transform 1 0 5060 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_51_74
timestamp 1607194113
transform 1 0 7912 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_62
timestamp 1607194113
transform 1 0 6808 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_60
timestamp 1607194113
transform 1 0 6624 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1607194113
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_93
timestamp 1607194113
transform 1 0 9660 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_86
timestamp 1607194113
transform 1 0 9016 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A
timestamp 1607194113
transform 1 0 9476 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0781_
timestamp 1607194113
transform 1 0 9200 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_51_116
timestamp 1607194113
transform 1 0 11776 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__B
timestamp 1607194113
transform 1 0 11592 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _0674_
timestamp 1607194113
transform 1 0 10764 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_51_128
timestamp 1607194113
transform 1 0 12880 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__A
timestamp 1607194113
transform 1 0 12696 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1607194113
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0672_
timestamp 1607194113
transform 1 0 12420 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_140
timestamp 1607194113
transform 1 0 13984 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1278__B1
timestamp 1607194113
transform 1 0 15088 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1278_
timestamp 1607194113
transform 1 0 15272 0 1 29920
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_51_172
timestamp 1607194113
transform 1 0 16928 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1278__A1_N
timestamp 1607194113
transform 1 0 16744 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_196
timestamp 1607194113
transform 1 0 19136 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_184
timestamp 1607194113
transform 1 0 18032 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_180
timestamp 1607194113
transform 1 0 17664 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1607194113
transform 1 0 17940 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_202
timestamp 1607194113
transform 1 0 19688 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1373__CLK
timestamp 1607194113
transform 1 0 19780 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1373_
timestamp 1607194113
transform 1 0 19964 0 1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_51_235
timestamp 1607194113
transform 1 0 22724 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_224
timestamp 1607194113
transform 1 0 21712 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__A
timestamp 1607194113
transform 1 0 22264 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0820_
timestamp 1607194113
transform 1 0 22448 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_51_243
timestamp 1607194113
transform 1 0 23460 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1607194113
transform 1 0 23552 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_18
timestamp 1607194113
transform 1 0 2760 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_11
timestamp 1607194113
transform 1 0 2116 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_3
timestamp 1607194113
transform 1 0 1380 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1607194113
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1607194113
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1607194113
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1607194113
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0895_
timestamp 1607194113
transform 1 0 2392 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_53_37
timestamp 1607194113
transform 1 0 4508 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_27
timestamp 1607194113
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__B
timestamp 1607194113
transform 1 0 4324 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1607194113
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0928_
timestamp 1607194113
transform 1 0 3496 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _0912_
timestamp 1607194113
transform 1 0 4048 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_53_54
timestamp 1607194113
transform 1 0 6072 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_55
timestamp 1607194113
transform 1 0 6164 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_43
timestamp 1607194113
transform 1 0 5060 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__B
timestamp 1607194113
transform 1 0 5888 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__B
timestamp 1607194113
transform 1 0 4876 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0936_
timestamp 1607194113
transform 1 0 5060 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_53_74
timestamp 1607194113
transform 1 0 7912 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_62
timestamp 1607194113
transform 1 0 6808 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_60
timestamp 1607194113
transform 1 0 6624 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_79
timestamp 1607194113
transform 1 0 8372 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_67
timestamp 1607194113
transform 1 0 7268 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1607194113
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_98
timestamp 1607194113
transform 1 0 10120 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_91
timestamp 1607194113
transform 1 0 9476 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1519__CLK
timestamp 1607194113
transform 1 0 10212 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__A
timestamp 1607194113
transform 1 0 9936 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1607194113
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1519_
timestamp 1607194113
transform 1 0 8464 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0666_
timestamp 1607194113
transform 1 0 9660 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_116
timestamp 1607194113
transform 1 0 11776 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_53_101
timestamp 1607194113
transform 1 0 10396 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__A2
timestamp 1607194113
transform 1 0 11960 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A
timestamp 1607194113
transform 1 0 11592 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1023_
timestamp 1607194113
transform 1 0 10948 0 1 31008
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_4  _0673_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 10856 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_135
timestamp 1607194113
transform 1 0 13524 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_123
timestamp 1607194113
transform 1 0 12420 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_132
timestamp 1607194113
transform 1 0 13248 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_120
timestamp 1607194113
transform 1 0 12144 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1607194113
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_143
timestamp 1607194113
transform 1 0 14260 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_154
timestamp 1607194113
transform 1 0 15272 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_52_145
timestamp 1607194113
transform 1 0 14444 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_140
timestamp 1607194113
transform 1 0 13984 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1607194113
transform 1 0 15180 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1369_
timestamp 1607194113
transform 1 0 14352 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1234_
timestamp 1607194113
transform 1 0 14168 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_174
timestamp 1607194113
transform 1 0 17112 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_53_165
timestamp 1607194113
transform 1 0 16284 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1370__CLK
timestamp 1607194113
transform 1 0 16008 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1369__CLK
timestamp 1607194113
transform 1 0 16100 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1370_
timestamp 1607194113
transform 1 0 16192 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0798_
timestamp 1607194113
transform 1 0 16836 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_53_196
timestamp 1607194113
transform 1 0 19136 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_184
timestamp 1607194113
transform 1 0 18032 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_182
timestamp 1607194113
transform 1 0 17848 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_195
timestamp 1607194113
transform 1 0 19044 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_183
timestamp 1607194113
transform 1 0 17940 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1607194113
transform 1 0 17940 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_202
timestamp 1607194113
transform 1 0 19688 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_215
timestamp 1607194113
transform 1 0 20884 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_52_213
timestamp 1607194113
transform 1 0 20700 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_207
timestamp 1607194113
transform 1 0 20148 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__B1
timestamp 1607194113
transform 1 0 19780 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__B1
timestamp 1607194113
transform 1 0 20976 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1607194113
transform 1 0 20792 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1273_
timestamp 1607194113
transform 1 0 21160 0 -1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _1211_
timestamp 1607194113
transform 1 0 19964 0 1 31008
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_53_238
timestamp 1607194113
transform 1 0 23000 0 1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_231
timestamp 1607194113
transform 1 0 22356 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_223
timestamp 1607194113
transform 1 0 21620 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_236
timestamp 1607194113
transform 1 0 22816 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A
timestamp 1607194113
transform 1 0 22816 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1273__A1_N
timestamp 1607194113
transform 1 0 22632 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__A1_N
timestamp 1607194113
transform 1 0 21436 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0824_
timestamp 1607194113
transform 1 0 22540 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1607194113
transform 1 0 23552 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_54_11
timestamp 1607194113
transform 1 0 2116 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_3
timestamp 1607194113
transform 1 0 1380 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1607194113
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0932_
timestamp 1607194113
transform 1 0 2392 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_54_25
timestamp 1607194113
transform 1 0 3404 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__B
timestamp 1607194113
transform 1 0 3220 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1607194113
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0926_
timestamp 1607194113
transform 1 0 4048 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_54_53
timestamp 1607194113
transform 1 0 5980 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_43
timestamp 1607194113
transform 1 0 5060 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__B
timestamp 1607194113
transform 1 0 4876 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0922_
timestamp 1607194113
transform 1 0 5612 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_77
timestamp 1607194113
transform 1 0 8188 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_65
timestamp 1607194113
transform 1 0 7084 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_84
timestamp 1607194113
transform 1 0 8832 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1607194113
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1327_
timestamp 1607194113
transform 1 0 8556 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _1325_
timestamp 1607194113
transform 1 0 9660 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_119
timestamp 1607194113
transform 1 0 12052 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_107
timestamp 1607194113
transform 1 0 10948 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1325__A2
timestamp 1607194113
transform 1 0 10764 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_131
timestamp 1607194113
transform 1 0 13156 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1210_
timestamp 1607194113
transform 1 0 13524 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_154
timestamp 1607194113
transform 1 0 15272 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1607194113
transform 1 0 14076 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__A
timestamp 1607194113
transform 1 0 13892 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1607194113
transform 1 0 15180 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1240_
timestamp 1607194113
transform 1 0 15456 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_172
timestamp 1607194113
transform 1 0 16928 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_54_160
timestamp 1607194113
transform 1 0 15824 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1276__A
timestamp 1607194113
transform 1 0 16376 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1276_
timestamp 1607194113
transform 1 0 16560 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1607194113
transform 1 0 19228 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_185
timestamp 1607194113
transform 1 0 18124 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__A
timestamp 1607194113
transform 1 0 17940 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0853_
timestamp 1607194113
transform 1 0 17664 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_215
timestamp 1607194113
transform 1 0 20884 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_213
timestamp 1607194113
transform 1 0 20700 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_209
timestamp 1607194113
transform 1 0 20332 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1607194113
transform 1 0 20792 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_54_223
timestamp 1607194113
transform 1 0 21620 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1374__CLK
timestamp 1607194113
transform 1 0 21712 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1374_
timestamp 1607194113
transform 1 0 21896 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_55_15
timestamp 1607194113
transform 1 0 2484 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1607194113
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1607194113
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1508_
timestamp 1607194113
transform 1 0 2668 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_55_38
timestamp 1607194113
transform 1 0 4600 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1508__CLK
timestamp 1607194113
transform 1 0 4416 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_55_55
timestamp 1607194113
transform 1 0 6164 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__B
timestamp 1607194113
transform 1 0 5980 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0934_
timestamp 1607194113
transform 1 0 5152 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_55_74
timestamp 1607194113
transform 1 0 7912 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_62
timestamp 1607194113
transform 1 0 6808 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1607194113
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_92
timestamp 1607194113
transform 1 0 9568 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_86
timestamp 1607194113
transform 1 0 9016 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__or3_4  _1326_
timestamp 1607194113
transform 1 0 9660 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_55_116
timestamp 1607194113
transform 1 0 11776 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_104
timestamp 1607194113
transform 1 0 10672 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1326__B
timestamp 1607194113
transform 1 0 10488 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_127
timestamp 1607194113
transform 1 0 12788 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1607194113
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1172_
timestamp 1607194113
transform 1 0 12420 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_139
timestamp 1607194113
transform 1 0 13892 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__A1_N
timestamp 1607194113
transform 1 0 15640 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1279__B1
timestamp 1607194113
transform 1 0 13984 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1279_
timestamp 1607194113
transform 1 0 14168 0 1 32096
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_55_172
timestamp 1607194113
transform 1 0 16928 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_160
timestamp 1607194113
transform 1 0 15824 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_184
timestamp 1607194113
transform 1 0 18032 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_180
timestamp 1607194113
transform 1 0 17664 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1607194113
transform 1 0 17940 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1410_
timestamp 1607194113
transform 1 0 18124 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_55_216
timestamp 1607194113
transform 1 0 20976 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_206
timestamp 1607194113
transform 1 0 20056 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1410__CLK
timestamp 1607194113
transform 1 0 19872 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1269__A
timestamp 1607194113
transform 1 0 20424 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1269_
timestamp 1607194113
transform 1 0 20608 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_236
timestamp 1607194113
transform 1 0 22816 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_232
timestamp 1607194113
transform 1 0 22448 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_228
timestamp 1607194113
transform 1 0 22080 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0739_
timestamp 1607194113
transform 1 0 22540 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1607194113
transform 1 0 23552 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1607194113
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1607194113
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1607194113
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_37
timestamp 1607194113
transform 1 0 4508 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_27
timestamp 1607194113
transform 1 0 3588 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A
timestamp 1607194113
transform 1 0 4324 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1607194113
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0860_
timestamp 1607194113
transform 1 0 4048 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_43
timestamp 1607194113
transform 1 0 5060 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1509_
timestamp 1607194113
transform 1 0 5152 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_56_77
timestamp 1607194113
transform 1 0 8188 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1607194113
transform 1 0 7084 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1509__CLK
timestamp 1607194113
transform 1 0 6900 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_93
timestamp 1607194113
transform 1 0 9660 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_89
timestamp 1607194113
transform 1 0 9292 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1607194113
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_56_111
timestamp 1607194113
transform 1 0 11316 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_105
timestamp 1607194113
transform 1 0 10764 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1280__B1
timestamp 1607194113
transform 1 0 11408 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1280_
timestamp 1607194113
transform 1 0 11592 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_56_130
timestamp 1607194113
transform 1 0 13064 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1181_
timestamp 1607194113
transform 1 0 13800 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_158
timestamp 1607194113
transform 1 0 15640 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_150
timestamp 1607194113
transform 1 0 14904 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_142
timestamp 1607194113
transform 1 0 14168 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1607194113
transform 1 0 15180 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1235_
timestamp 1607194113
transform 1 0 15272 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_56_170
timestamp 1607194113
transform 1 0 16744 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__B1
timestamp 1607194113
transform 1 0 17020 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1217_
timestamp 1607194113
transform 1 0 17204 0 -1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_56_193
timestamp 1607194113
transform 1 0 18860 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__A1_N
timestamp 1607194113
transform 1 0 18676 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_215
timestamp 1607194113
transform 1 0 20884 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_212
timestamp 1607194113
transform 1 0 20608 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_204
timestamp 1607194113
transform 1 0 19872 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1607194113
transform 1 0 20792 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0699_
timestamp 1607194113
transform 1 0 19596 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_56_223
timestamp 1607194113
transform 1 0 21620 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1415__CLK
timestamp 1607194113
transform 1 0 21712 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1415_
timestamp 1607194113
transform 1 0 21896 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1607194113
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1607194113
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1607194113
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_57_35
timestamp 1607194113
transform 1 0 4324 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_27
timestamp 1607194113
transform 1 0 3588 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _0861_
timestamp 1607194113
transform 1 0 4600 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_54
timestamp 1607194113
transform 1 0 6072 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_42
timestamp 1607194113
transform 1 0 4968 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_74
timestamp 1607194113
transform 1 0 7912 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_62
timestamp 1607194113
transform 1 0 6808 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_60
timestamp 1607194113
transform 1 0 6624 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1607194113
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_98
timestamp 1607194113
transform 1 0 10120 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_57_86
timestamp 1607194113
transform 1 0 9016 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_114
timestamp 1607194113
transform 1 0 11592 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_57_106
timestamp 1607194113
transform 1 0 10856 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__A
timestamp 1607194113
transform 1 0 11408 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0665_
timestamp 1607194113
transform 1 0 11040 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1368__CLK
timestamp 1607194113
transform 1 0 12144 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1607194113
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1368_
timestamp 1607194113
transform 1 0 12420 0 1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_57_154
timestamp 1607194113
transform 1 0 15272 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_142
timestamp 1607194113
transform 1 0 14168 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_178
timestamp 1607194113
transform 1 0 17480 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_166
timestamp 1607194113
transform 1 0 16376 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_196
timestamp 1607194113
transform 1 0 19136 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_184
timestamp 1607194113
transform 1 0 18032 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_182
timestamp 1607194113
transform 1 0 17848 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1607194113
transform 1 0 17940 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__B1
timestamp 1607194113
transform 1 0 20240 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1270_
timestamp 1607194113
transform 1 0 20424 0 1 33184
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_57_230
timestamp 1607194113
transform 1 0 22264 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__A2_N
timestamp 1607194113
transform 1 0 22080 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1270__A1_N
timestamp 1607194113
transform 1 0 21896 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_242
timestamp 1607194113
transform 1 0 23368 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1607194113
transform 1 0 23552 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1607194113
transform 1 0 2484 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1607194113
transform 1 0 1380 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1607194113
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_32
timestamp 1607194113
transform 1 0 4048 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_27
timestamp 1607194113
transform 1 0 3588 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1607194113
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_45
timestamp 1607194113
transform 1 0 5244 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_40
timestamp 1607194113
transform 1 0 4784 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0884_
timestamp 1607194113
transform 1 0 5980 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _0880_
timestamp 1607194113
transform 1 0 4876 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_74
timestamp 1607194113
transform 1 0 7912 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_62
timestamp 1607194113
transform 1 0 6808 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_93
timestamp 1607194113
transform 1 0 9660 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_86
timestamp 1607194113
transform 1 0 9016 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A
timestamp 1607194113
transform 1 0 9844 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1607194113
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0800_
timestamp 1607194113
transform 1 0 10028 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_58_115
timestamp 1607194113
transform 1 0 11684 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_58_108
timestamp 1607194113
transform 1 0 11040 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_100
timestamp 1607194113
transform 1 0 10304 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1176_
timestamp 1607194113
transform 1 0 11316 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__B1
timestamp 1607194113
transform 1 0 12236 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1218_
timestamp 1607194113
transform 1 0 12420 0 -1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_58_157
timestamp 1607194113
transform 1 0 15548 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1607194113
transform 1 0 14076 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__A1_N
timestamp 1607194113
transform 1 0 13892 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1607194113
transform 1 0 15180 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0704_
timestamp 1607194113
transform 1 0 15272 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_169
timestamp 1607194113
transform 1 0 16652 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_193
timestamp 1607194113
transform 1 0 18860 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_58_181
timestamp 1607194113
transform 1 0 17756 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_215
timestamp 1607194113
transform 1 0 20884 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_206
timestamp 1607194113
transform 1 0 20056 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_199
timestamp 1607194113
transform 1 0 19412 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__A
timestamp 1607194113
transform 1 0 19504 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1607194113
transform 1 0 20792 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1377_
timestamp 1607194113
transform 1 0 21068 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1206_
timestamp 1607194113
transform 1 0 19688 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_238
timestamp 1607194113
transform 1 0 23000 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1377__CLK
timestamp 1607194113
transform 1 0 22816 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1607194113
transform 1 0 2484 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1607194113
transform 1 0 1380 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1607194113
transform 1 0 1380 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1607194113
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1607194113
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1510_
timestamp 1607194113
transform 1 0 2484 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_60_32
timestamp 1607194113
transform 1 0 4048 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_27
timestamp 1607194113
transform 1 0 3588 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_36
timestamp 1607194113
transform 1 0 4416 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1510__CLK
timestamp 1607194113
transform 1 0 4232 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1607194113
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_59
timestamp 1607194113
transform 1 0 6532 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_60_44
timestamp 1607194113
transform 1 0 5152 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_53
timestamp 1607194113
transform 1 0 5980 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _0888_
timestamp 1607194113
transform 1 0 5152 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _0886_
timestamp 1607194113
transform 1 0 5704 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_60_76
timestamp 1607194113
transform 1 0 8096 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_71
timestamp 1607194113
transform 1 0 7636 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1607194113
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0938_
timestamp 1607194113
transform 1 0 7268 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_4  _0892_
timestamp 1607194113
transform 1 0 6808 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_60_93
timestamp 1607194113
transform 1 0 9660 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_88
timestamp 1607194113
transform 1 0 9200 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_95
timestamp 1607194113
transform 1 0 9844 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_83
timestamp 1607194113
transform 1 0 8740 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1607194113
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_117
timestamp 1607194113
transform 1 0 11868 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_105
timestamp 1607194113
transform 1 0 10764 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_114
timestamp 1607194113
transform 1 0 11592 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_107
timestamp 1607194113
transform 1 0 10948 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0803_
timestamp 1607194113
transform 1 0 11316 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_125
timestamp 1607194113
transform 1 0 12604 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_59_129
timestamp 1607194113
transform 1 0 12972 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_59_123
timestamp 1607194113
transform 1 0 12420 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1607194113
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1409_
timestamp 1607194113
transform 1 0 13064 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__o22a_4  _0706_
timestamp 1607194113
transform 1 0 12880 0 -1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_60_154
timestamp 1607194113
transform 1 0 15272 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_152
timestamp 1607194113
transform 1 0 15088 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_148
timestamp 1607194113
transform 1 0 14720 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_151
timestamp 1607194113
transform 1 0 14996 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1409__CLK
timestamp 1607194113
transform 1 0 14812 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__A2
timestamp 1607194113
transform 1 0 14536 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__B2
timestamp 1607194113
transform 1 0 14352 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__B1
timestamp 1607194113
transform 1 0 14168 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1607194113
transform 1 0 15180 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_178
timestamp 1607194113
transform 1 0 17480 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_60_166
timestamp 1607194113
transform 1 0 16376 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_175
timestamp 1607194113
transform 1 0 17204 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_163
timestamp 1607194113
transform 1 0 16100 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_194
timestamp 1607194113
transform 1 0 18952 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_184
timestamp 1607194113
transform 1 0 18032 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__B1
timestamp 1607194113
transform 1 0 18032 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1607194113
transform 1 0 17940 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1258_
timestamp 1607194113
transform 1 0 18216 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _1173_
timestamp 1607194113
transform 1 0 18584 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_215
timestamp 1607194113
transform 1 0 20884 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_212
timestamp 1607194113
transform 1 0 20608 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_204
timestamp 1607194113
transform 1 0 19872 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_206
timestamp 1607194113
transform 1 0 20056 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__B2
timestamp 1607194113
transform 1 0 20148 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1258__A1_N
timestamp 1607194113
transform 1 0 19688 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__B1
timestamp 1607194113
transform 1 0 20332 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1607194113
transform 1 0 20792 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1207_
timestamp 1607194113
transform 1 0 20516 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_60_223
timestamp 1607194113
transform 1 0 21620 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_231
timestamp 1607194113
transform 1 0 22356 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__A2_N
timestamp 1607194113
transform 1 0 22172 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__A1_N
timestamp 1607194113
transform 1 0 21988 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1418_
timestamp 1607194113
transform 1 0 21804 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_59_243
timestamp 1607194113
transform 1 0 23460 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1418__CLK
timestamp 1607194113
transform 1 0 23552 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1607194113
transform 1 0 23552 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1607194113
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1607194113
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1511_
timestamp 1607194113
transform 1 0 2484 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_61_36
timestamp 1607194113
transform 1 0 4416 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1511__CLK
timestamp 1607194113
transform 1 0 4232 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_53
timestamp 1607194113
transform 1 0 5980 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _0894_
timestamp 1607194113
transform 1 0 5152 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_61_78
timestamp 1607194113
transform 1 0 8280 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_62
timestamp 1607194113
transform 1 0 6808 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1607194113
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _0917_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 7084 0 1 35360
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_61_95
timestamp 1607194113
transform 1 0 9844 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A
timestamp 1607194113
transform 1 0 9660 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0915_
timestamp 1607194113
transform 1 0 9016 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_61_119
timestamp 1607194113
transform 1 0 12052 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_111
timestamp 1607194113
transform 1 0 11316 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_103
timestamp 1607194113
transform 1 0 10580 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A
timestamp 1607194113
transform 1 0 10764 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0868_
timestamp 1607194113
transform 1 0 10948 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_123
timestamp 1607194113
transform 1 0 12420 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__B2
timestamp 1607194113
transform 1 0 13800 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1607194113
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0804_
timestamp 1607194113
transform 1 0 12512 0 1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_61_142
timestamp 1607194113
transform 1 0 14168 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__A2
timestamp 1607194113
transform 1 0 13984 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0937_
timestamp 1607194113
transform 1 0 14536 0 1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_61_176
timestamp 1607194113
transform 1 0 17296 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_164
timestamp 1607194113
transform 1 0 16192 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__B1
timestamp 1607194113
transform 1 0 16008 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__A1
timestamp 1607194113
transform 1 0 15824 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_182
timestamp 1607194113
transform 1 0 17848 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1607194113
transform 1 0 17940 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1426_
timestamp 1607194113
transform 1 0 18032 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_61_215
timestamp 1607194113
transform 1 0 20884 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_211
timestamp 1607194113
transform 1 0 20516 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_205
timestamp 1607194113
transform 1 0 19964 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1426__CLK
timestamp 1607194113
transform 1 0 19780 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0829_
timestamp 1607194113
transform 1 0 20608 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_227
timestamp 1607194113
transform 1 0 21988 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_243
timestamp 1607194113
transform 1 0 23460 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_239
timestamp 1607194113
transform 1 0 23092 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1607194113
transform 1 0 23552 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1607194113
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1607194113
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1607194113
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_32
timestamp 1607194113
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_27
timestamp 1607194113
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1607194113
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_56
timestamp 1607194113
transform 1 0 6256 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_44
timestamp 1607194113
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_68
timestamp 1607194113
transform 1 0 7360 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _0916_
timestamp 1607194113
transform 1 0 7728 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_93
timestamp 1607194113
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_88
timestamp 1607194113
transform 1 0 9200 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__B1
timestamp 1607194113
transform 1 0 9016 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__A1
timestamp 1607194113
transform 1 0 8832 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1607194113
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_117
timestamp 1607194113
transform 1 0 11868 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_105
timestamp 1607194113
transform 1 0 10764 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1236__A
timestamp 1607194113
transform 1 0 11684 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1236_
timestamp 1607194113
transform 1 0 11316 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_132
timestamp 1607194113
transform 1 0 13248 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A
timestamp 1607194113
transform 1 0 13800 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0707_
timestamp 1607194113
transform 1 0 12420 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_62_154
timestamp 1607194113
transform 1 0 15272 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_152
timestamp 1607194113
transform 1 0 15088 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_144
timestamp 1607194113
transform 1 0 14352 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1607194113
transform 1 0 15180 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0863_
timestamp 1607194113
transform 1 0 13984 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_166
timestamp 1607194113
transform 1 0 16376 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__B1
timestamp 1607194113
transform 1 0 17480 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_198
timestamp 1607194113
transform 1 0 19320 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__A1_N
timestamp 1607194113
transform 1 0 19136 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1195_
timestamp 1607194113
transform 1 0 17664 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_62_218
timestamp 1607194113
transform 1 0 21160 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_210
timestamp 1607194113
transform 1 0 20424 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1607194113
transform 1 0 20792 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0747_
timestamp 1607194113
transform 1 0 20884 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_230
timestamp 1607194113
transform 1 0 22264 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_242
timestamp 1607194113
transform 1 0 23368 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1607194113
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1607194113
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1344_
timestamp 1607194113
transform 1 0 2484 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_63_38
timestamp 1607194113
transform 1 0 4600 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__CLK
timestamp 1607194113
transform 1 0 4416 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1344__D
timestamp 1607194113
transform 1 0 4232 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_58
timestamp 1607194113
transform 1 0 6440 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_50
timestamp 1607194113
transform 1 0 5704 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_63_76
timestamp 1607194113
transform 1 0 8096 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_62
timestamp 1607194113
transform 1 0 6808 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1607194113
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _0910_
timestamp 1607194113
transform 1 0 6900 0 1 36448
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__B1
timestamp 1607194113
transform 1 0 10120 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A1
timestamp 1607194113
transform 1 0 9936 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _0909_
timestamp 1607194113
transform 1 0 8832 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_112
timestamp 1607194113
transform 1 0 11408 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_100
timestamp 1607194113
transform 1 0 10304 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_132
timestamp 1607194113
transform 1 0 13248 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_120
timestamp 1607194113
transform 1 0 12144 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1607194113
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0805_
timestamp 1607194113
transform 1 0 12420 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_63_158
timestamp 1607194113
transform 1 0 15640 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_146
timestamp 1607194113
transform 1 0 14536 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__A
timestamp 1607194113
transform 1 0 14352 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1182_
timestamp 1607194113
transform 1 0 13984 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_175
timestamp 1607194113
transform 1 0 17204 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_166
timestamp 1607194113
transform 1 0 16376 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__A
timestamp 1607194113
transform 1 0 16652 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1192_
timestamp 1607194113
transform 1 0 16836 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_192
timestamp 1607194113
transform 1 0 18768 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_184
timestamp 1607194113
transform 1 0 18032 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1607194113
transform 1 0 17940 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1385_
timestamp 1607194113
transform 1 0 19044 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_63_216
timestamp 1607194113
transform 1 0 20976 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1385__CLK
timestamp 1607194113
transform 1 0 20792 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_236
timestamp 1607194113
transform 1 0 22816 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_228
timestamp 1607194113
transform 1 0 22080 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1262__A
timestamp 1607194113
transform 1 0 22264 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1262_
timestamp 1607194113
transform 1 0 22448 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1607194113
transform 1 0 23552 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1607194113
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1607194113
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1607194113
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_27
timestamp 1607194113
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1607194113
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1513_
timestamp 1607194113
transform 1 0 4048 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1607194113
transform 1 0 5980 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1513__CLK
timestamp 1607194113
transform 1 0 5796 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_65
timestamp 1607194113
transform 1 0 7084 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _0903_
timestamp 1607194113
transform 1 0 8188 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_64_93
timestamp 1607194113
transform 1 0 9660 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_86
timestamp 1607194113
transform 1 0 9016 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__A
timestamp 1607194113
transform 1 0 8832 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1607194113
transform 1 0 9568 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_117
timestamp 1607194113
transform 1 0 11868 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_105
timestamp 1607194113
transform 1 0 10764 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_132
timestamp 1607194113
transform 1 0 13248 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__B
timestamp 1607194113
transform 1 0 13064 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0802_
timestamp 1607194113
transform 1 0 13800 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0703_
timestamp 1607194113
transform 1 0 12420 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_64_154
timestamp 1607194113
transform 1 0 15272 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_147
timestamp 1607194113
transform 1 0 14628 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__B
timestamp 1607194113
transform 1 0 14444 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1607194113
transform 1 0 15180 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_178
timestamp 1607194113
transform 1 0 17480 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_166
timestamp 1607194113
transform 1 0 16376 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__B1
timestamp 1607194113
transform 1 0 18032 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1194_
timestamp 1607194113
transform 1 0 18216 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_64_204
timestamp 1607194113
transform 1 0 19872 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__A1_N
timestamp 1607194113
transform 1 0 19688 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__B1
timestamp 1607194113
transform 1 0 20608 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1607194113
transform 1 0 20792 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1257_
timestamp 1607194113
transform 1 0 20884 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_64_237
timestamp 1607194113
transform 1 0 22908 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_233
timestamp 1607194113
transform 1 0 22540 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__A
timestamp 1607194113
transform 1 0 23000 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1257__A1_N
timestamp 1607194113
transform 1 0 22356 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_244
timestamp 1607194113
transform 1 0 23552 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1189_
timestamp 1607194113
transform 1 0 23184 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1607194113
transform 1 0 1380 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1607194113
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1512_
timestamp 1607194113
transform 1 0 2484 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_65_36
timestamp 1607194113
transform 1 0 4416 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1512__CLK
timestamp 1607194113
transform 1 0 4232 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_65_58
timestamp 1607194113
transform 1 0 6440 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_46
timestamp 1607194113
transform 1 0 5336 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0862_
timestamp 1607194113
transform 1 0 4968 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_62
timestamp 1607194113
transform 1 0 6808 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1607194113
transform 1 0 6716 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0883_
timestamp 1607194113
transform 1 0 7544 0 1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_65_96
timestamp 1607194113
transform 1 0 9936 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_84
timestamp 1607194113
transform 1 0 8832 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_108
timestamp 1607194113
transform 1 0 11040 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_120
timestamp 1607194113
transform 1 0 12144 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1607194113
transform 1 0 12328 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1435_
timestamp 1607194113
transform 1 0 12420 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_65_156
timestamp 1607194113
transform 1 0 15456 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_144
timestamp 1607194113
transform 1 0 14352 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1435__CLK
timestamp 1607194113
transform 1 0 14168 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_168
timestamp 1607194113
transform 1 0 16560 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_191
timestamp 1607194113
transform 1 0 18676 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_184
timestamp 1607194113
transform 1 0 18032 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_180
timestamp 1607194113
transform 1 0 17664 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1255__A
timestamp 1607194113
transform 1 0 18492 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1607194113
transform 1 0 17940 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1386_
timestamp 1607194113
transform 1 0 19228 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _1255_
timestamp 1607194113
transform 1 0 18124 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_218
timestamp 1607194113
transform 1 0 21160 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1386__CLK
timestamp 1607194113
transform 1 0 20976 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_227
timestamp 1607194113
transform 1 0 21988 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0806_
timestamp 1607194113
transform 1 0 21712 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_65_243
timestamp 1607194113
transform 1 0 23460 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_239
timestamp 1607194113
transform 1 0 23092 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1607194113
transform 1 0 23552 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_3
timestamp 1607194113
transform 1 0 1380 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_15
timestamp 1607194113
transform 1 0 2484 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_3
timestamp 1607194113
transform 1 0 1380 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1607194113
transform 1 0 1104 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1607194113
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1514_
timestamp 1607194113
transform 1 0 2484 0 1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_67_36
timestamp 1607194113
transform 1 0 4416 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_27
timestamp 1607194113
transform 1 0 3588 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1514__CLK
timestamp 1607194113
transform 1 0 4232 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1607194113
transform 1 0 3956 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0875_
timestamp 1607194113
transform 1 0 4048 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_67_48
timestamp 1607194113
transform 1 0 5520 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_55
timestamp 1607194113
transform 1 0 6164 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_43
timestamp 1607194113
transform 1 0 5060 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__B
timestamp 1607194113
transform 1 0 4876 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_62
timestamp 1607194113
transform 1 0 6808 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_60
timestamp 1607194113
transform 1 0 6624 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_72
timestamp 1607194113
transform 1 0 7728 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_67
timestamp 1607194113
transform 1 0 7268 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1607194113
transform 1 0 6716 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0885_
timestamp 1607194113
transform 1 0 7544 0 1 38624
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _0882_
timestamp 1607194113
transform 1 0 7360 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_88
timestamp 1607194113
transform 1 0 9200 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_93
timestamp 1607194113
transform 1 0 9660 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_84
timestamp 1607194113
transform 1 0 8832 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__B1
timestamp 1607194113
transform 1 0 9016 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__A1
timestamp 1607194113
transform 1 0 8832 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1246__B1
timestamp 1607194113
transform 1 0 9936 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1607194113
transform 1 0 9568 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1246_
timestamp 1607194113
transform 1 0 10120 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _0881_
timestamp 1607194113
transform 1 0 8464 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_114
timestamp 1607194113
transform 1 0 11592 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_105
timestamp 1607194113
transform 1 0 10764 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__B1
timestamp 1607194113
transform 1 0 11040 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1183_
timestamp 1607194113
transform 1 0 11224 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_67_123
timestamp 1607194113
transform 1 0 12420 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_126
timestamp 1607194113
transform 1 0 12696 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A
timestamp 1607194113
transform 1 0 13708 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1607194113
transform 1 0 12328 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1394_
timestamp 1607194113
transform 1 0 12696 0 1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0702_
timestamp 1607194113
transform 1 0 13432 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_156
timestamp 1607194113
transform 1 0 15456 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_147
timestamp 1607194113
transform 1 0 14628 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_154
timestamp 1607194113
transform 1 0 15272 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_151
timestamp 1607194113
transform 1 0 14996 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_139
timestamp 1607194113
transform 1 0 13892 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1394__CLK
timestamp 1607194113
transform 1 0 14444 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__A
timestamp 1607194113
transform 1 0 14996 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1607194113
transform 1 0 15180 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0801_
timestamp 1607194113
transform 1 0 15180 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_168
timestamp 1607194113
transform 1 0 16560 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_178
timestamp 1607194113
transform 1 0 17480 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_166
timestamp 1607194113
transform 1 0 16376 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_184
timestamp 1607194113
transform 1 0 18032 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_180
timestamp 1607194113
transform 1 0 17664 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_186
timestamp 1607194113
transform 1 0 18216 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__B1
timestamp 1607194113
transform 1 0 18400 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1607194113
transform 1 0 17940 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1427_
timestamp 1607194113
transform 1 0 19136 0 1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _1193_
timestamp 1607194113
transform 1 0 18584 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1607194113
transform 1 0 21068 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_208
timestamp 1607194113
transform 1 0 20240 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1427__CLK
timestamp 1607194113
transform 1 0 20884 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__A1_N
timestamp 1607194113
transform 1 0 20424 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__A1_N
timestamp 1607194113
transform 1 0 20056 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1256__B1
timestamp 1607194113
transform 1 0 20608 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1607194113
transform 1 0 20792 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1256_
timestamp 1607194113
transform 1 0 20884 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_67_238
timestamp 1607194113
transform 1 0 23000 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_226
timestamp 1607194113
transform 1 0 21896 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_231
timestamp 1607194113
transform 1 0 22356 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0902_
timestamp 1607194113
transform 1 0 21620 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_243
timestamp 1607194113
transform 1 0 23460 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1607194113
transform 1 0 23552 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_11
timestamp 1607194113
transform 1 0 2116 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_3
timestamp 1607194113
transform 1 0 1380 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1607194113
transform 1 0 1104 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_4  _0873_
timestamp 1607194113
transform 1 0 2392 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_68_25
timestamp 1607194113
transform 1 0 3404 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__B
timestamp 1607194113
transform 1 0 3220 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1607194113
transform 1 0 3956 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0871_
timestamp 1607194113
transform 1 0 4048 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_68_55
timestamp 1607194113
transform 1 0 6164 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_43
timestamp 1607194113
transform 1 0 5060 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__B
timestamp 1607194113
transform 1 0 4876 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__B1
timestamp 1607194113
transform 1 0 6256 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__A1
timestamp 1607194113
transform 1 0 6440 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_74
timestamp 1607194113
transform 1 0 7912 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _0893_
timestamp 1607194113
transform 1 0 6624 0 -1 39712
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_68_98
timestamp 1607194113
transform 1 0 10120 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_86
timestamp 1607194113
transform 1 0 9016 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__A
timestamp 1607194113
transform 1 0 9936 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1607194113
transform 1 0 9568 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0676_
timestamp 1607194113
transform 1 0 9660 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_68_110
timestamp 1607194113
transform 1 0 11224 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1248_
timestamp 1607194113
transform 1 0 11776 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_122
timestamp 1607194113
transform 1 0 12328 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1248__A
timestamp 1607194113
transform 1 0 12144 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__B1
timestamp 1607194113
transform 1 0 12696 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1184_
timestamp 1607194113
transform 1 0 12880 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_68_158
timestamp 1607194113
transform 1 0 15640 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_152
timestamp 1607194113
transform 1 0 15088 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_146
timestamp 1607194113
transform 1 0 14536 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__A1_N
timestamp 1607194113
transform 1 0 14352 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1607194113
transform 1 0 15180 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0864_
timestamp 1607194113
transform 1 0 15272 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_170
timestamp 1607194113
transform 1 0 16744 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_194
timestamp 1607194113
transform 1 0 18952 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_182
timestamp 1607194113
transform 1 0 17848 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_218
timestamp 1607194113
transform 1 0 21160 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_208
timestamp 1607194113
transform 1 0 20240 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_202
timestamp 1607194113
transform 1 0 19688 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__A
timestamp 1607194113
transform 1 0 20056 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1607194113
transform 1 0 20792 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0904_
timestamp 1607194113
transform 1 0 19780 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0710_
timestamp 1607194113
transform 1 0 20884 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_230
timestamp 1607194113
transform 1 0 22264 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_242
timestamp 1607194113
transform 1 0 23368 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1607194113
transform 1 0 1380 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__B1
timestamp 1607194113
transform 1 0 2484 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1607194113
transform 1 0 1104 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1251_
timestamp 1607194113
transform 1 0 2668 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_69_35
timestamp 1607194113
transform 1 0 4324 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1251__A1_N
timestamp 1607194113
transform 1 0 4140 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_69_58
timestamp 1607194113
transform 1 0 6440 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_50
timestamp 1607194113
transform 1 0 5704 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_4  _0879_
timestamp 1607194113
transform 1 0 4876 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_69_70
timestamp 1607194113
transform 1 0 7544 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_62
timestamp 1607194113
transform 1 0 6808 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1607194113
transform 1 0 6716 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0887_
timestamp 1607194113
transform 1 0 7728 0 1 39712
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_69_90
timestamp 1607194113
transform 1 0 9384 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__B1
timestamp 1607194113
transform 1 0 9200 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__A1
timestamp 1607194113
transform 1 0 9016 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_114
timestamp 1607194113
transform 1 0 11592 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_102
timestamp 1607194113
transform 1 0 10488 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_123
timestamp 1607194113
transform 1 0 12420 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__B1
timestamp 1607194113
transform 1 0 12788 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1607194113
transform 1 0 12328 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1247_
timestamp 1607194113
transform 1 0 12972 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_69_157
timestamp 1607194113
transform 1 0 15548 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_147
timestamp 1607194113
transform 1 0 14628 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1247__A1_N
timestamp 1607194113
transform 1 0 14444 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0869_
timestamp 1607194113
transform 1 0 15180 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1607194113
transform 1 0 16652 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_196
timestamp 1607194113
transform 1 0 19136 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_184
timestamp 1607194113
transform 1 0 18032 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_181
timestamp 1607194113
transform 1 0 17756 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1607194113
transform 1 0 17940 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_204
timestamp 1607194113
transform 1 0 19872 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1387_
timestamp 1607194113
transform 1 0 19964 0 1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_69_238
timestamp 1607194113
transform 1 0 23000 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_226
timestamp 1607194113
transform 1 0 21896 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1387__CLK
timestamp 1607194113
transform 1 0 21712 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1607194113
transform 1 0 23552 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1607194113
transform 1 0 2484 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1607194113
transform 1 0 1380 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1607194113
transform 1 0 1104 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_70_27
timestamp 1607194113
transform 1 0 3588 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_593
timestamp 1607194113
transform 1 0 3956 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _0877_
timestamp 1607194113
transform 1 0 4048 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_70_52
timestamp 1607194113
transform 1 0 5888 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_43
timestamp 1607194113
transform 1 0 5060 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__B
timestamp 1607194113
transform 1 0 4876 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0808_
timestamp 1607194113
transform 1 0 5612 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_79
timestamp 1607194113
transform 1 0 8372 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_64
timestamp 1607194113
transform 1 0 6992 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0891_
timestamp 1607194113
transform 1 0 7084 0 -1 40800
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_70_93
timestamp 1607194113
transform 1 0 9660 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_91
timestamp 1607194113
transform 1 0 9476 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_594
timestamp 1607194113
transform 1 0 9568 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_105
timestamp 1607194113
transform 1 0 10764 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__B1
timestamp 1607194113
transform 1 0 11132 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1249_
timestamp 1607194113
transform 1 0 11316 0 -1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_70_129
timestamp 1607194113
transform 1 0 12972 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1249__A1_N
timestamp 1607194113
transform 1 0 12788 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1245_
timestamp 1607194113
transform 1 0 13524 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_154
timestamp 1607194113
transform 1 0 15272 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_70_151
timestamp 1607194113
transform 1 0 14996 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_139
timestamp 1607194113
transform 1 0 13892 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_595
timestamp 1607194113
transform 1 0 15180 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_171
timestamp 1607194113
transform 1 0 16836 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_162
timestamp 1607194113
transform 1 0 16008 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1241__A
timestamp 1607194113
transform 1 0 16284 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1241_
timestamp 1607194113
transform 1 0 16468 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_195
timestamp 1607194113
transform 1 0 19044 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_183
timestamp 1607194113
transform 1 0 17940 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_211
timestamp 1607194113
transform 1 0 20516 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_207
timestamp 1607194113
transform 1 0 20148 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A2
timestamp 1607194113
transform 1 0 20608 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_596
timestamp 1607194113
transform 1 0 20792 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0876_
timestamp 1607194113
transform 1 0 20884 0 -1 40800
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_70_233
timestamp 1607194113
transform 1 0 22540 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__B1
timestamp 1607194113
transform 1 0 22356 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A1
timestamp 1607194113
transform 1 0 22172 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_71_15
timestamp 1607194113
transform 1 0 2484 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1607194113
transform 1 0 1380 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1607194113
transform 1 0 1104 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1390_
timestamp 1607194113
transform 1 0 2760 0 1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_71_39
timestamp 1607194113
transform 1 0 4692 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1390__CLK
timestamp 1607194113
transform 1 0 4508 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_59
timestamp 1607194113
transform 1 0 6532 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_51
timestamp 1607194113
transform 1 0 5796 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_78
timestamp 1607194113
transform 1 0 8280 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_74
timestamp 1607194113
transform 1 0 7912 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_62
timestamp 1607194113
transform 1 0 6808 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_612
timestamp 1607194113
transform 1 0 6716 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1607194113
transform 1 0 8372 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_96
timestamp 1607194113
transform 1 0 9936 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_84
timestamp 1607194113
transform 1 0 8832 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__A
timestamp 1607194113
transform 1 0 8648 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_108
timestamp 1607194113
transform 1 0 11040 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_71_123
timestamp 1607194113
transform 1 0 12420 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_120
timestamp 1607194113
transform 1 0 12144 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_613
timestamp 1607194113
transform 1 0 12328 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1392_
timestamp 1607194113
transform 1 0 12696 0 1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_71_157
timestamp 1607194113
transform 1 0 15548 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_147
timestamp 1607194113
transform 1 0 14628 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1392__CLK
timestamp 1607194113
transform 1 0 14444 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1237_
timestamp 1607194113
transform 1 0 15180 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1607194113
transform 1 0 16652 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_196
timestamp 1607194113
transform 1 0 19136 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_184
timestamp 1607194113
transform 1 0 18032 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_181
timestamp 1607194113
transform 1 0 17756 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_614
timestamp 1607194113
transform 1 0 17940 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1428_
timestamp 1607194113
transform 1 0 19688 0 1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_71_233
timestamp 1607194113
transform 1 0 22540 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_229
timestamp 1607194113
transform 1 0 22172 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_223
timestamp 1607194113
transform 1 0 21620 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1428__CLK
timestamp 1607194113
transform 1 0 21436 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0810_
timestamp 1607194113
transform 1 0 22264 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_71_241
timestamp 1607194113
transform 1 0 23276 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_615
timestamp 1607194113
transform 1 0 23552 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_73_15
timestamp 1607194113
transform 1 0 2484 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1607194113
transform 1 0 1380 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1607194113
transform 1 0 2484 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1607194113
transform 1 0 1380 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1607194113
transform 1 0 1104 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1607194113
transform 1 0 1104 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1431_
timestamp 1607194113
transform 1 0 2760 0 1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_73_39
timestamp 1607194113
transform 1 0 4692 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_32
timestamp 1607194113
transform 1 0 4048 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_27
timestamp 1607194113
transform 1 0 3588 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1431__CLK
timestamp 1607194113
transform 1 0 4508 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_630
timestamp 1607194113
transform 1 0 3956 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_59
timestamp 1607194113
transform 1 0 6532 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_51
timestamp 1607194113
transform 1 0 5796 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_56
timestamp 1607194113
transform 1 0 6256 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_44
timestamp 1607194113
transform 1 0 5152 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_74
timestamp 1607194113
transform 1 0 7912 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_62
timestamp 1607194113
transform 1 0 6808 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_78
timestamp 1607194113
transform 1 0 8280 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1250__B1
timestamp 1607194113
transform 1 0 6624 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_649
timestamp 1607194113
transform 1 0 6716 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1250_
timestamp 1607194113
transform 1 0 6808 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_73_80
timestamp 1607194113
transform 1 0 8464 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_72_97
timestamp 1607194113
transform 1 0 10028 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_93
timestamp 1607194113
transform 1 0 9660 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_90
timestamp 1607194113
transform 1 0 9384 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__B1
timestamp 1607194113
transform 1 0 10120 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_631
timestamp 1607194113
transform 1 0 9568 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1432_
timestamp 1607194113
transform 1 0 8556 0 1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_73_114
timestamp 1607194113
transform 1 0 11592 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_73_102
timestamp 1607194113
transform 1 0 10488 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_72_118
timestamp 1607194113
transform 1 0 11960 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1432__CLK
timestamp 1607194113
transform 1 0 10304 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__A
timestamp 1607194113
transform 1 0 11408 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__A1_N
timestamp 1607194113
transform 1 0 11776 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1186_
timestamp 1607194113
transform 1 0 10304 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _1185_
timestamp 1607194113
transform 1 0 11040 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_135
timestamp 1607194113
transform 1 0 13524 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_123
timestamp 1607194113
transform 1 0 12420 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_130
timestamp 1607194113
transform 1 0 13064 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_650
timestamp 1607194113
transform 1 0 12328 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_147
timestamp 1607194113
transform 1 0 14628 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_154
timestamp 1607194113
transform 1 0 15272 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_145
timestamp 1607194113
transform 1 0 14444 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__B1
timestamp 1607194113
transform 1 0 15364 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_632
timestamp 1607194113
transform 1 0 15180 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1180_
timestamp 1607194113
transform 1 0 15548 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__o22a_4  _0878_
timestamp 1607194113
transform 1 0 15364 0 -1 41888
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _0831_
timestamp 1607194113
transform 1 0 14168 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_175
timestamp 1607194113
transform 1 0 17204 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_175
timestamp 1607194113
transform 1 0 17204 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A2
timestamp 1607194113
transform 1 0 17020 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__B1
timestamp 1607194113
transform 1 0 16836 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A1
timestamp 1607194113
transform 1 0 16652 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__A1_N
timestamp 1607194113
transform 1 0 17020 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_190
timestamp 1607194113
transform 1 0 18584 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_73_184
timestamp 1607194113
transform 1 0 18032 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_187
timestamp 1607194113
transform 1 0 18308 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_651
timestamp 1607194113
transform 1 0 17940 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0812_
timestamp 1607194113
transform 1 0 18308 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_202
timestamp 1607194113
transform 1 0 19688 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_72_211
timestamp 1607194113
transform 1 0 20516 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_199
timestamp 1607194113
transform 1 0 19412 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__B1
timestamp 1607194113
transform 1 0 19872 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_633
timestamp 1607194113
transform 1 0 20792 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1396_
timestamp 1607194113
transform 1 0 20884 0 -1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _1243_
timestamp 1607194113
transform 1 0 20056 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_73_236
timestamp 1607194113
transform 1 0 22816 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_232
timestamp 1607194113
transform 1 0 22448 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_224
timestamp 1607194113
transform 1 0 21712 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_236
timestamp 1607194113
transform 1 0 22816 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1396__CLK
timestamp 1607194113
transform 1 0 22632 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1243__A1_N
timestamp 1607194113
transform 1 0 21528 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0715_
timestamp 1607194113
transform 1 0 22540 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_652
timestamp 1607194113
transform 1 0 23552 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_3
timestamp 1607194113
transform 1 0 1380 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__B1
timestamp 1607194113
transform 1 0 1564 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1607194113
transform 1 0 1104 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _1188_
timestamp 1607194113
transform 1 0 1748 0 -1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_74_36
timestamp 1607194113
transform 1 0 4416 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_32
timestamp 1607194113
transform 1 0 4048 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_25
timestamp 1607194113
transform 1 0 3404 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__A1_N
timestamp 1607194113
transform 1 0 3220 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_667
timestamp 1607194113
transform 1 0 3956 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0712_
timestamp 1607194113
transform 1 0 4140 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_48
timestamp 1607194113
transform 1 0 5520 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_60
timestamp 1607194113
transform 1 0 6624 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__B1
timestamp 1607194113
transform 1 0 7176 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1187_
timestamp 1607194113
transform 1 0 7360 0 -1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_74_98
timestamp 1607194113
transform 1 0 10120 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_74_84
timestamp 1607194113
transform 1 0 8832 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__A
timestamp 1607194113
transform 1 0 9936 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_668
timestamp 1607194113
transform 1 0 9568 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0889_
timestamp 1607194113
transform 1 0 9660 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_74_104
timestamp 1607194113
transform 1 0 10672 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1433_
timestamp 1607194113
transform 1 0 10764 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_74_138
timestamp 1607194113
transform 1 0 13800 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_126
timestamp 1607194113
transform 1 0 12696 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1433__CLK
timestamp 1607194113
transform 1 0 12512 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_154
timestamp 1607194113
transform 1 0 15272 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_150
timestamp 1607194113
transform 1 0 14904 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_669
timestamp 1607194113
transform 1 0 15180 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_166
timestamp 1607194113
transform 1 0 16376 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1395_
timestamp 1607194113
transform 1 0 16744 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_74_191
timestamp 1607194113
transform 1 0 18676 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1395__CLK
timestamp 1607194113
transform 1 0 18492 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_215
timestamp 1607194113
transform 1 0 20884 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_74_211
timestamp 1607194113
transform 1 0 20516 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_74_203
timestamp 1607194113
transform 1 0 19780 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_670
timestamp 1607194113
transform 1 0 20792 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1437__CLK
timestamp 1607194113
transform 1 0 23000 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1437_
timestamp 1607194113
transform 1 0 21252 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_74_240
timestamp 1607194113
transform 1 0 23184 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_75_11
timestamp 1607194113
transform 1 0 2116 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_3
timestamp 1607194113
transform 1 0 1380 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__D
timestamp 1607194113
transform 1 0 2300 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1607194113
transform 1 0 1104 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1345_
timestamp 1607194113
transform 1 0 2484 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_36
timestamp 1607194113
transform 1 0 4416 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1345__CLK
timestamp 1607194113
transform 1 0 4232 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_48
timestamp 1607194113
transform 1 0 5520 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_62
timestamp 1607194113
transform 1 0 6808 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_60
timestamp 1607194113
transform 1 0 6624 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_686
timestamp 1607194113
transform 1 0 6716 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1391_
timestamp 1607194113
transform 1 0 7544 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_91
timestamp 1607194113
transform 1 0 9476 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1391__CLK
timestamp 1607194113
transform 1 0 9292 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_115
timestamp 1607194113
transform 1 0 11684 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_103
timestamp 1607194113
transform 1 0 10580 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_138
timestamp 1607194113
transform 1 0 13800 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_126
timestamp 1607194113
transform 1 0 12696 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_121
timestamp 1607194113
transform 1 0 12236 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_687
timestamp 1607194113
transform 1 0 12328 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0752_
timestamp 1607194113
transform 1 0 12420 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_75_150
timestamp 1607194113
transform 1 0 14904 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _1436_
timestamp 1607194113
transform 1 0 15456 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_75_177
timestamp 1607194113
transform 1 0 17388 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1436__CLK
timestamp 1607194113
transform 1 0 17204 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_187
timestamp 1607194113
transform 1 0 18308 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_688
timestamp 1607194113
transform 1 0 17940 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0717_
timestamp 1607194113
transform 1 0 18032 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_75_207
timestamp 1607194113
transform 1 0 20148 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_199
timestamp 1607194113
transform 1 0 19412 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__B1
timestamp 1607194113
transform 1 0 20240 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1179_
timestamp 1607194113
transform 1 0 20424 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_75_228
timestamp 1607194113
transform 1 0 22080 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__A1_N
timestamp 1607194113
transform 1 0 21896 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_240
timestamp 1607194113
transform 1 0 23184 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_689
timestamp 1607194113
transform 1 0 23552 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1607194113
transform 1 0 2484 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1607194113
transform 1 0 1380 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1607194113
transform 1 0 1104 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_32
timestamp 1607194113
transform 1 0 4048 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_27
timestamp 1607194113
transform 1 0 3588 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_704
timestamp 1607194113
transform 1 0 3956 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_56
timestamp 1607194113
transform 1 0 6256 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_44
timestamp 1607194113
transform 1 0 5152 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_75
timestamp 1607194113
transform 1 0 8004 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_63
timestamp 1607194113
transform 1 0 6900 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_705
timestamp 1607194113
transform 1 0 6808 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_94
timestamp 1607194113
transform 1 0 9752 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_87
timestamp 1607194113
transform 1 0 9108 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_706
timestamp 1607194113
transform 1 0 9660 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_118
timestamp 1607194113
transform 1 0 11960 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_106
timestamp 1607194113
transform 1 0 10856 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_137
timestamp 1607194113
transform 1 0 13708 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_125
timestamp 1607194113
transform 1 0 12604 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_707
timestamp 1607194113
transform 1 0 12512 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_76_156
timestamp 1607194113
transform 1 0 15456 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_149
timestamp 1607194113
transform 1 0 14812 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__B1
timestamp 1607194113
transform 1 0 15548 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_708
timestamp 1607194113
transform 1 0 15364 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_177
timestamp 1607194113
transform 1 0 17388 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1244__A1_N
timestamp 1607194113
transform 1 0 17204 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1244_
timestamp 1607194113
transform 1 0 15732 0 -1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_76_187
timestamp 1607194113
transform 1 0 18308 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_185
timestamp 1607194113
transform 1 0 18124 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_709
timestamp 1607194113
transform 1 0 18216 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_218
timestamp 1607194113
transform 1 0 21160 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_211
timestamp 1607194113
transform 1 0 20516 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_199
timestamp 1607194113
transform 1 0 19412 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_710
timestamp 1607194113
transform 1 0 21068 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_230
timestamp 1607194113
transform 1 0 22264 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_242
timestamp 1607194113
transform 1 0 23368 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_245
timestamp 1607194113
transform 1 0 23644 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_249
timestamp 1607194113
transform 1 0 24012 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1607194113
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1607194113
transform -1 0 24656 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1607194113
transform -1 0 24656 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_251
timestamp 1607194113
transform 1 0 24196 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1607194113
transform -1 0 24656 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_251
timestamp 1607194113
transform 1 0 24196 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_245
timestamp 1607194113
transform 1 0 23644 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1607194113
transform -1 0 24656 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1607194113
transform -1 0 24656 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_252
timestamp 1607194113
transform 1 0 24288 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_246
timestamp 1607194113
transform 1 0 23736 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_7_245
timestamp 1607194113
transform 1 0 23644 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_245
timestamp 1607194113
transform 1 0 23644 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_5_245
timestamp 1607194113
transform 1 0 23644 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1607194113
transform -1 0 24656 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1607194113
transform -1 0 24656 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1607194113
transform -1 0 24656 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1607194113
transform -1 0 24656 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_245
timestamp 1607194113
transform 1 0 23644 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_245
timestamp 1607194113
transform 1 0 23644 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_251
timestamp 1607194113
transform 1 0 24196 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_245
timestamp 1607194113
transform 1 0 23644 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1607194113
transform -1 0 24656 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1607194113
transform -1 0 24656 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1607194113
transform -1 0 24656 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1607194113
transform -1 0 24656 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1607194113
transform -1 0 24656 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_245
timestamp 1607194113
transform 1 0 23644 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_251
timestamp 1607194113
transform 1 0 24196 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_245
timestamp 1607194113
transform 1 0 23644 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_252
timestamp 1607194113
transform 1 0 24288 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1607194113
transform 1 0 23920 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1607194113
transform -1 0 24656 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1607194113
transform -1 0 24656 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1607194113
transform -1 0 24656 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1607194113
transform -1 0 24656 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_245
timestamp 1607194113
transform 1 0 23644 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_252
timestamp 1607194113
transform 1 0 24288 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1607194113
transform -1 0 24656 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1607194113
transform -1 0 24656 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_245
timestamp 1607194113
transform 1 0 23644 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1607194113
transform -1 0 24656 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_250
timestamp 1607194113
transform 1 0 24104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_245
timestamp 1607194113
transform 1 0 23644 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1607194113
transform -1 0 24656 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1607194113
transform -1 0 24656 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_250
timestamp 1607194113
transform 1 0 24104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_245
timestamp 1607194113
transform 1 0 23644 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_24_245
timestamp 1607194113
transform 1 0 23644 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_245
timestamp 1607194113
transform 1 0 23644 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1607194113
transform -1 0 24656 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1607194113
transform -1 0 24656 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1607194113
transform -1 0 24656 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1607194113
transform -1 0 24656 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_252
timestamp 1607194113
transform 1 0 24288 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_245
timestamp 1607194113
transform 1 0 23644 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1607194113
transform -1 0 24656 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1607194113
transform -1 0 24656 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_245
timestamp 1607194113
transform 1 0 23644 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1607194113
transform -1 0 24656 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_245
timestamp 1607194113
transform 1 0 23644 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_30_245
timestamp 1607194113
transform 1 0 23644 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1607194113
transform -1 0 24656 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1607194113
transform -1 0 24656 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_35_245
timestamp 1607194113
transform 1 0 23644 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_250
timestamp 1607194113
transform 1 0 24104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_245
timestamp 1607194113
transform 1 0 23644 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_32_247
timestamp 1607194113
transform 1 0 23828 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1607194113
transform -1 0 24656 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1607194113
transform -1 0 24656 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1607194113
transform -1 0 24656 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1607194113
transform -1 0 24656 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_245
timestamp 1607194113
transform 1 0 23644 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_37_245
timestamp 1607194113
transform 1 0 23644 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_clk_i_A
timestamp 1607194113
transform 1 0 23920 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_clk_i
timestamp 1607194113
transform 1 0 24104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1607194113
transform -1 0 24656 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1607194113
transform -1 0 24656 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1607194113
transform -1 0 24656 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_39_245
timestamp 1607194113
transform 1 0 23644 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1607194113
transform -1 0 24656 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_245
timestamp 1607194113
transform 1 0 23644 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1607194113
transform -1 0 24656 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_251
timestamp 1607194113
transform 1 0 24196 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_41_245
timestamp 1607194113
transform 1 0 23644 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1607194113
transform -1 0 24656 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1607194113
transform -1 0 24656 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_245
timestamp 1607194113
transform 1 0 23644 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1607194113
transform -1 0 24656 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_251
timestamp 1607194113
transform 1 0 24196 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1607194113
transform -1 0 24656 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_245
timestamp 1607194113
transform 1 0 23644 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1607194113
transform -1 0 24656 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_46_250
timestamp 1607194113
transform 1 0 24104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1607194113
transform -1 0 24656 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_48_247
timestamp 1607194113
transform 1 0 23828 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_245
timestamp 1607194113
transform 1 0 23644 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1607194113
transform -1 0 24656 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1607194113
transform -1 0 24656 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_49_245
timestamp 1607194113
transform 1 0 23644 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1607194113
transform -1 0 24656 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_245
timestamp 1607194113
transform 1 0 23644 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1607194113
transform -1 0 24656 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_245
timestamp 1607194113
transform 1 0 23644 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1607194113
transform -1 0 24656 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_52_252
timestamp 1607194113
transform 1 0 24288 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_248
timestamp 1607194113
transform 1 0 23920 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1607194113
transform -1 0 24656 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_245
timestamp 1607194113
transform 1 0 23644 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1607194113
transform -1 0 24656 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_55_245
timestamp 1607194113
transform 1 0 23644 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_245
timestamp 1607194113
transform 1 0 23644 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1607194113
transform -1 0 24656 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1607194113
transform -1 0 24656 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_245
timestamp 1607194113
transform 1 0 23644 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1607194113
transform -1 0 24656 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_245
timestamp 1607194113
transform 1 0 23644 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1607194113
transform -1 0 24656 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_58_250
timestamp 1607194113
transform 1 0 24104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1607194113
transform -1 0 24656 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_260
timestamp 1607194113
transform 1 0 25024 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_251
timestamp 1607194113
transform 1 0 24196 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1266__A
timestamp 1607194113
transform 1 0 24012 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1266_
timestamp 1607194113
transform 1 0 23644 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0728_
timestamp 1607194113
transform 1 0 24748 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_279
timestamp 1607194113
transform 1 0 26772 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_272
timestamp 1607194113
transform 1 0 26128 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__A
timestamp 1607194113
transform 1 0 26220 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1203_
timestamp 1607194113
transform 1 0 26404 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_303
timestamp 1607194113
transform 1 0 28980 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_291
timestamp 1607194113
transform 1 0 27876 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_318
timestamp 1607194113
transform 1 0 30360 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_306
timestamp 1607194113
transform 1 0 29256 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__A1_N
timestamp 1607194113
transform 1 0 30728 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1607194113
transform 1 0 29164 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__A2_N
timestamp 1607194113
transform 1 0 32568 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__B2
timestamp 1607194113
transform 1 0 32384 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0783_
timestamp 1607194113
transform 1 0 30912 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_59_356
timestamp 1607194113
transform 1 0 33856 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_344
timestamp 1607194113
transform 1 0 32752 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_381
timestamp 1607194113
transform 1 0 36156 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_367
timestamp 1607194113
transform 1 0 34868 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_364
timestamp 1607194113
transform 1 0 34592 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__A
timestamp 1607194113
transform 1 0 35604 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1607194113
transform 1 0 34776 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0923_
timestamp 1607194113
transform 1 0 35788 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_393
timestamp 1607194113
transform 1 0 37260 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__A1_N
timestamp 1607194113
transform 1 0 37444 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__B1
timestamp 1607194113
transform 1 0 37628 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0701_
timestamp 1607194113
transform 1 0 37812 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_59_419
timestamp 1607194113
transform 1 0 39652 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__A2_N
timestamp 1607194113
transform 1 0 39468 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__B2
timestamp 1607194113
transform 1 0 39284 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_428
timestamp 1607194113
transform 1 0 40480 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__A2_N
timestamp 1607194113
transform 1 0 41216 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__B2
timestamp 1607194113
transform 1 0 41400 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__B1
timestamp 1607194113
transform 1 0 41584 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1607194113
transform 1 0 40388 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1205_
timestamp 1607194113
transform 1 0 41768 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_59_458
timestamp 1607194113
transform 1 0 43240 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_482
timestamp 1607194113
transform 1 0 45448 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_470
timestamp 1607194113
transform 1 0 44344 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1607194113
transform 1 0 46000 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_255
timestamp 1607194113
transform 1 0 24564 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_60_246
timestamp 1607194113
transform 1 0 23736 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__A
timestamp 1607194113
transform 1 0 25116 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0897_
timestamp 1607194113
transform 1 0 25300 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0819_
timestamp 1607194113
transform 1 0 24288 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_276
timestamp 1607194113
transform 1 0 26496 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_267
timestamp 1607194113
transform 1 0 25668 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1607194113
transform 1 0 26404 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_297
timestamp 1607194113
transform 1 0 28428 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_60_288
timestamp 1607194113
transform 1 0 27600 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1259__A
timestamp 1607194113
transform 1 0 27876 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1261__B1
timestamp 1607194113
transform 1 0 28980 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1259_
timestamp 1607194113
transform 1 0 28060 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_321
timestamp 1607194113
transform 1 0 30636 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _1261_
timestamp 1607194113
transform 1 0 29164 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_60_335
timestamp 1607194113
transform 1 0 31924 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_329
timestamp 1607194113
transform 1 0 31372 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__B1
timestamp 1607194113
transform 1 0 31740 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A1_N
timestamp 1607194113
transform 1 0 31556 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1607194113
transform 1 0 32016 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0854_
timestamp 1607194113
transform 1 0 32108 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_60_357
timestamp 1607194113
transform 1 0 33948 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A2_N
timestamp 1607194113
transform 1 0 33764 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A
timestamp 1607194113
transform 1 0 34316 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__B2
timestamp 1607194113
transform 1 0 33580 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0924_
timestamp 1607194113
transform 1 0 34500 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_367
timestamp 1607194113
transform 1 0 34868 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__B2
timestamp 1607194113
transform 1 0 35420 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0925_
timestamp 1607194113
transform 1 0 35604 0 -1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_60_398
timestamp 1607194113
transform 1 0 37720 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_391
timestamp 1607194113
transform 1 0 37076 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A2
timestamp 1607194113
transform 1 0 36892 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__A1_N
timestamp 1607194113
transform 1 0 37260 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__B1
timestamp 1607194113
transform 1 0 37444 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1607194113
transform 1 0 37628 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0799_
timestamp 1607194113
transform 1 0 37812 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_60_419
timestamp 1607194113
transform 1 0 39652 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__A2_N
timestamp 1607194113
transform 1 0 39468 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__B2
timestamp 1607194113
transform 1 0 39284 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_427
timestamp 1607194113
transform 1 0 40388 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__A2_N
timestamp 1607194113
transform 1 0 40480 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__B2
timestamp 1607194113
transform 1 0 40664 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1268__B1
timestamp 1607194113
transform 1 0 40848 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1268_
timestamp 1607194113
transform 1 0 41032 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_60_457
timestamp 1607194113
transform 1 0 43148 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_60_450
timestamp 1607194113
transform 1 0 42504 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__B2
timestamp 1607194113
transform 1 0 42964 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__A2
timestamp 1607194113
transform 1 0 42780 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1607194113
transform 1 0 43240 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0935_
timestamp 1607194113
transform 1 0 43332 0 -1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_60_473
timestamp 1607194113
transform 1 0 44620 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_485
timestamp 1607194113
transform 1 0 45724 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_61_264
timestamp 1607194113
transform 1 0 25392 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_257
timestamp 1607194113
transform 1 0 24748 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_245
timestamp 1607194113
transform 1 0 23644 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__B1
timestamp 1607194113
transform 1 0 23920 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A1
timestamp 1607194113
transform 1 0 24104 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A
timestamp 1607194113
transform 1 0 24840 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0913_
timestamp 1607194113
transform 1 0 24288 0 -1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__buf_2  _0896_
timestamp 1607194113
transform 1 0 25024 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_62_276
timestamp 1607194113
transform 1 0 26496 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_62_274
timestamp 1607194113
transform 1 0 26312 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_266
timestamp 1607194113
transform 1 0 25576 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__A
timestamp 1607194113
transform 1 0 26772 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1607194113
transform 1 0 26404 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1196_
timestamp 1607194113
transform 1 0 26956 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_4  _0920_
timestamp 1607194113
transform 1 0 26128 0 1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_62_297
timestamp 1607194113
transform 1 0 28428 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_285
timestamp 1607194113
transform 1 0 27324 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_298
timestamp 1607194113
transform 1 0 28520 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_286
timestamp 1607194113
transform 1 0 27416 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__B1
timestamp 1607194113
transform 1 0 28612 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1198_
timestamp 1607194113
transform 1 0 28796 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_62_317
timestamp 1607194113
transform 1 0 30268 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_314
timestamp 1607194113
transform 1 0 29992 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_306
timestamp 1607194113
transform 1 0 29256 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_304
timestamp 1607194113
transform 1 0 29072 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1607194113
transform 1 0 29164 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1424_
timestamp 1607194113
transform 1 0 30268 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_62_340
timestamp 1607194113
transform 1 0 32384 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_328
timestamp 1607194113
transform 1 0 31280 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_338
timestamp 1607194113
transform 1 0 32200 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1424__CLK
timestamp 1607194113
transform 1 0 32016 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1607194113
transform 1 0 32016 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0919_
timestamp 1607194113
transform 1 0 32108 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0918_
timestamp 1607194113
transform 1 0 31004 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_352
timestamp 1607194113
transform 1 0 33488 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_362
timestamp 1607194113
transform 1 0 34408 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_350
timestamp 1607194113
transform 1 0 33304 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_370
timestamp 1607194113
transform 1 0 35144 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_364
timestamp 1607194113
transform 1 0 34592 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_61_367
timestamp 1607194113
transform 1 0 34868 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__B1
timestamp 1607194113
transform 1 0 35236 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__B1
timestamp 1607194113
transform 1 0 35144 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1607194113
transform 1 0 34776 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1260_
timestamp 1607194113
transform 1 0 35328 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _1197_
timestamp 1607194113
transform 1 0 35420 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_62_398
timestamp 1607194113
transform 1 0 37720 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_391
timestamp 1607194113
transform 1 0 37076 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_402
timestamp 1607194113
transform 1 0 38088 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_390
timestamp 1607194113
transform 1 0 36984 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1260__A1_N
timestamp 1607194113
transform 1 0 36800 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__A1_N
timestamp 1607194113
transform 1 0 36892 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1607194113
transform 1 0 37628 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_415
timestamp 1607194113
transform 1 0 39284 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_410
timestamp 1607194113
transform 1 0 38824 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_414
timestamp 1607194113
transform 1 0 39192 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0796_
timestamp 1607194113
transform 1 0 39008 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_439
timestamp 1607194113
transform 1 0 41492 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_427
timestamp 1607194113
transform 1 0 40388 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_440
timestamp 1607194113
transform 1 0 41584 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_428
timestamp 1607194113
transform 1 0 40480 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_426
timestamp 1607194113
transform 1 0 40296 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1607194113
transform 1 0 40388 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_455
timestamp 1607194113
transform 1 0 42964 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_451
timestamp 1607194113
transform 1 0 42596 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1419__CLK
timestamp 1607194113
transform 1 0 43056 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1378__CLK
timestamp 1607194113
transform 1 0 42688 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1607194113
transform 1 0 43240 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1419_
timestamp 1607194113
transform 1 0 43332 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1378_
timestamp 1607194113
transform 1 0 42872 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_62_478
timestamp 1607194113
transform 1 0 45080 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1607194113
transform 1 0 44620 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_485
timestamp 1607194113
transform 1 0 45724 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1607194113
transform 1 0 46000 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_245
timestamp 1607194113
transform 1 0 23644 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__B1
timestamp 1607194113
transform 1 0 24012 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A1
timestamp 1607194113
transform 1 0 24196 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0911_
timestamp 1607194113
transform 1 0 24380 0 1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_63_267
timestamp 1607194113
transform 1 0 25668 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _0898_
timestamp 1607194113
transform 1 0 26404 0 1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1607194113
transform 1 0 28060 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__B1
timestamp 1607194113
transform 1 0 27876 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A1
timestamp 1607194113
transform 1 0 27692 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_314
timestamp 1607194113
transform 1 0 29992 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_306
timestamp 1607194113
transform 1 0 29256 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1607194113
transform 1 0 29164 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1383_
timestamp 1607194113
transform 1 0 30268 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_63_338
timestamp 1607194113
transform 1 0 32200 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1383__CLK
timestamp 1607194113
transform 1 0 32016 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_359
timestamp 1607194113
transform 1 0 34132 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_347
timestamp 1607194113
transform 1 0 33028 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_clk_i
timestamp 1607194113
transform 1 0 32752 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_367
timestamp 1607194113
transform 1 0 34868 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_365
timestamp 1607194113
transform 1 0 34684 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__B2
timestamp 1607194113
transform 1 0 35420 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__B1
timestamp 1607194113
transform 1 0 35604 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1607194113
transform 1 0 34776 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1200_
timestamp 1607194113
transform 1 0 35788 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1607194113
transform 1 0 37260 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_418
timestamp 1607194113
transform 1 0 39560 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_413
timestamp 1607194113
transform 1 0 39100 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_405
timestamp 1607194113
transform 1 0 38364 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0697_
timestamp 1607194113
transform 1 0 39284 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_440
timestamp 1607194113
transform 1 0 41584 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_428
timestamp 1607194113
transform 1 0 40480 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_426
timestamp 1607194113
transform 1 0 40296 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1607194113
transform 1 0 40388 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_452
timestamp 1607194113
transform 1 0 42688 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_482
timestamp 1607194113
transform 1 0 45448 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_470
timestamp 1607194113
transform 1 0 44344 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_464
timestamp 1607194113
transform 1 0 43792 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0846_
timestamp 1607194113
transform 1 0 44068 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1607194113
transform 1 0 46000 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_252
timestamp 1607194113
transform 1 0 24288 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0900_
timestamp 1607194113
transform 1 0 24380 0 -1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_64_276
timestamp 1607194113
transform 1 0 26496 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_271
timestamp 1607194113
transform 1 0 26036 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__B1
timestamp 1607194113
transform 1 0 25852 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A1
timestamp 1607194113
transform 1 0 25668 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1607194113
transform 1 0 26404 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_284
timestamp 1607194113
transform 1 0 27232 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__A1_N
timestamp 1607194113
transform 1 0 28980 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1253__B1
timestamp 1607194113
transform 1 0 27324 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1253_
timestamp 1607194113
transform 1 0 27508 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_64_317
timestamp 1607194113
transform 1 0 30268 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_305
timestamp 1607194113
transform 1 0 29164 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_337
timestamp 1607194113
transform 1 0 32108 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_335
timestamp 1607194113
transform 1 0 31924 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_329
timestamp 1607194113
transform 1 0 31372 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__A
timestamp 1607194113
transform 1 0 32476 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1607194113
transform 1 0 32016 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1199_
timestamp 1607194113
transform 1 0 32660 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_64_359
timestamp 1607194113
transform 1 0 34132 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_347
timestamp 1607194113
transform 1 0 33028 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_clk_i
timestamp 1607194113
transform 1 0 34408 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_365
timestamp 1607194113
transform 1 0 34684 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__B2
timestamp 1607194113
transform 1 0 35052 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1263__B1
timestamp 1607194113
transform 1 0 35236 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1263_
timestamp 1607194113
transform 1 0 35420 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_64_389
timestamp 1607194113
transform 1 0 36892 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1382__CLK
timestamp 1607194113
transform 1 0 37444 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1607194113
transform 1 0 37628 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1382_
timestamp 1607194113
transform 1 0 37720 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_64_417
timestamp 1607194113
transform 1 0 39468 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_64_434
timestamp 1607194113
transform 1 0 41032 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__C
timestamp 1607194113
transform 1 0 40020 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0815_
timestamp 1607194113
transform 1 0 40204 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_64_459
timestamp 1607194113
transform 1 0 43332 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_446
timestamp 1607194113
transform 1 0 42136 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1607194113
transform 1 0 43240 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_467
timestamp 1607194113
transform 1 0 44068 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_463
timestamp 1607194113
transform 1 0 43700 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1384__CLK
timestamp 1607194113
transform 1 0 44620 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1384_
timestamp 1607194113
transform 1 0 44804 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0770_
timestamp 1607194113
transform 1 0 43792 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_65_257
timestamp 1607194113
transform 1 0 24748 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_245
timestamp 1607194113
transform 1 0 23644 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__B1
timestamp 1607194113
transform 1 0 25300 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_283
timestamp 1607194113
transform 1 0 27140 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__A1_N
timestamp 1607194113
transform 1 0 26956 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1191_
timestamp 1607194113
transform 1 0 25484 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_65_303
timestamp 1607194113
transform 1 0 28980 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_295
timestamp 1607194113
transform 1 0 28244 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_318
timestamp 1607194113
transform 1 0 30360 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_306
timestamp 1607194113
transform 1 0 29256 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1607194113
transform 1 0 29164 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1430__CLK
timestamp 1607194113
transform 1 0 31464 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_clk_i
timestamp 1607194113
transform 1 0 31648 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1430_
timestamp 1607194113
transform 1 0 31924 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_65_354
timestamp 1607194113
transform 1 0 33672 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_379
timestamp 1607194113
transform 1 0 35972 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_367
timestamp 1607194113
transform 1 0 34868 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1607194113
transform 1 0 34776 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_391
timestamp 1607194113
transform 1 0 37076 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1423__CLK
timestamp 1607194113
transform 1 0 37628 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1423_
timestamp 1607194113
transform 1 0 37812 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_65_418
timestamp 1607194113
transform 1 0 39560 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_437
timestamp 1607194113
transform 1 0 41308 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_424
timestamp 1607194113
transform 1 0 40112 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__C
timestamp 1607194113
transform 1 0 40204 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1607194113
transform 1 0 40388 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0720_
timestamp 1607194113
transform 1 0 40480 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_65_461
timestamp 1607194113
transform 1 0 43516 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1607194113
transform 1 0 42412 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__B2
timestamp 1607194113
transform 1 0 45448 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A2_N
timestamp 1607194113
transform 1 0 45264 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0828_
timestamp 1607194113
transform 1 0 43792 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_65_484
timestamp 1607194113
transform 1 0 45632 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1607194113
transform 1 0 46000 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_255
timestamp 1607194113
transform 1 0 24564 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_276
timestamp 1607194113
transform 1 0 26496 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_66_267
timestamp 1607194113
transform 1 0 25668 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1607194113
transform 1 0 26404 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_66_284
timestamp 1607194113
transform 1 0 27232 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__B1
timestamp 1607194113
transform 1 0 27508 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1190_
timestamp 1607194113
transform 1 0 27692 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_319
timestamp 1607194113
transform 1 0 30452 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_307
timestamp 1607194113
transform 1 0 29348 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__A1_N
timestamp 1607194113
transform 1 0 29164 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_337
timestamp 1607194113
transform 1 0 32108 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_335
timestamp 1607194113
transform 1 0 31924 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_331
timestamp 1607194113
transform 1 0 31556 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1607194113
transform 1 0 32016 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_354
timestamp 1607194113
transform 1 0 33672 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _0856_
timestamp 1607194113
transform 1 0 32844 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_66_378
timestamp 1607194113
transform 1 0 35880 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_366
timestamp 1607194113
transform 1 0 34776 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_398
timestamp 1607194113
transform 1 0 37720 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_396
timestamp 1607194113
transform 1 0 37536 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_390
timestamp 1607194113
transform 1 0 36984 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1607194113
transform 1 0 37628 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0797_
timestamp 1607194113
transform 1 0 38824 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_442
timestamp 1607194113
transform 1 0 41768 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_430
timestamp 1607194113
transform 1 0 40664 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__B2
timestamp 1607194113
transform 1 0 40480 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__A2_N
timestamp 1607194113
transform 1 0 40296 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_459
timestamp 1607194113
transform 1 0 43332 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_66_454
timestamp 1607194113
transform 1 0 42872 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1607194113
transform 1 0 43240 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_66_467
timestamp 1607194113
transform 1 0 44068 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0746_
timestamp 1607194113
transform 1 0 44252 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__B2
timestamp 1607194113
transform 1 0 45908 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A2_N
timestamp 1607194113
transform 1 0 45724 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_254
timestamp 1607194113
transform 1 0 24472 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_257
timestamp 1607194113
transform 1 0 24748 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_245
timestamp 1607194113
transform 1 0 23644 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_276
timestamp 1607194113
transform 1 0 26496 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_274
timestamp 1607194113
transform 1 0 26312 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_266
timestamp 1607194113
transform 1 0 25576 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_67_269
timestamp 1607194113
transform 1 0 25852 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1607194113
transform 1 0 26404 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1429_
timestamp 1607194113
transform 1 0 26128 0 1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_68_292
timestamp 1607194113
transform 1 0 27968 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_284
timestamp 1607194113
transform 1 0 27232 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1607194113
transform 1 0 28060 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1429__CLK
timestamp 1607194113
transform 1 0 27876 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1252__A
timestamp 1607194113
transform 1 0 27416 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1252_
timestamp 1607194113
transform 1 0 27600 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_316
timestamp 1607194113
transform 1 0 30176 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_304
timestamp 1607194113
transform 1 0 29072 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_321
timestamp 1607194113
transform 1 0 30636 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_309
timestamp 1607194113
transform 1 0 29532 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1607194113
transform 1 0 29164 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0768_
timestamp 1607194113
transform 1 0 29256 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_328
timestamp 1607194113
transform 1 0 31280 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_329
timestamp 1607194113
transform 1 0 31372 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__B1
timestamp 1607194113
transform 1 0 31556 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__B1
timestamp 1607194113
transform 1 0 31740 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__A1_N
timestamp 1607194113
transform 1 0 31556 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__A1_N
timestamp 1607194113
transform 1 0 31740 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_335
timestamp 1607194113
transform 1 0 31924 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1607194113
transform 1 0 32016 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0851_
timestamp 1607194113
transform 1 0 32108 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _0777_
timestamp 1607194113
transform 1 0 31924 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_68_357
timestamp 1607194113
transform 1 0 33948 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_363
timestamp 1607194113
transform 1 0 34500 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_355
timestamp 1607194113
transform 1 0 33764 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__A2_N
timestamp 1607194113
transform 1 0 33580 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__A2_N
timestamp 1607194113
transform 1 0 33764 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__B2
timestamp 1607194113
transform 1 0 33396 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__B2
timestamp 1607194113
transform 1 0 33580 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0785_
timestamp 1607194113
transform 1 0 34316 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_68_382
timestamp 1607194113
transform 1 0 36248 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_370
timestamp 1607194113
transform 1 0 35144 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_379
timestamp 1607194113
transform 1 0 35972 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_367
timestamp 1607194113
transform 1 0 34868 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1607194113
transform 1 0 34776 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_398
timestamp 1607194113
transform 1 0 37720 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_394
timestamp 1607194113
transform 1 0 37352 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_391
timestamp 1607194113
transform 1 0 37076 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1607194113
transform 1 0 37628 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_410
timestamp 1607194113
transform 1 0 38824 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_421
timestamp 1607194113
transform 1 0 39836 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_409
timestamp 1607194113
transform 1 0 38732 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_403
timestamp 1607194113
transform 1 0 38180 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__B
timestamp 1607194113
transform 1 0 39652 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0814_
timestamp 1607194113
transform 1 0 38824 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__a2bb2o_4  _0698_
timestamp 1607194113
transform 1 0 39192 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_68_434
timestamp 1607194113
transform 1 0 41032 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_440
timestamp 1607194113
transform 1 0 41584 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_428
timestamp 1607194113
transform 1 0 40480 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__B2
timestamp 1607194113
transform 1 0 40848 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__A2_N
timestamp 1607194113
transform 1 0 40664 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1607194113
transform 1 0 40388 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_459
timestamp 1607194113
transform 1 0 43332 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_446
timestamp 1607194113
transform 1 0 42136 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_452
timestamp 1607194113
transform 1 0 42688 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__A1_N
timestamp 1607194113
transform 1 0 43424 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__B1
timestamp 1607194113
transform 1 0 43608 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1607194113
transform 1 0 43240 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_463
timestamp 1607194113
transform 1 0 43700 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__A2_N
timestamp 1607194113
transform 1 0 45448 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__B2
timestamp 1607194113
transform 1 0 45264 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A1_N
timestamp 1607194113
transform 1 0 43792 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__B1
timestamp 1607194113
transform 1 0 43976 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0830_
timestamp 1607194113
transform 1 0 43792 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _0749_
timestamp 1607194113
transform 1 0 44160 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_68_488
timestamp 1607194113
transform 1 0 46000 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_484
timestamp 1607194113
transform 1 0 45632 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A2_N
timestamp 1607194113
transform 1 0 45816 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__B2
timestamp 1607194113
transform 1 0 45632 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1607194113
transform 1 0 46000 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_69_257
timestamp 1607194113
transform 1 0 24748 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_245
timestamp 1607194113
transform 1 0 23644 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__B1
timestamp 1607194113
transform 1 0 25024 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1254_
timestamp 1607194113
transform 1 0 25208 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_69_280
timestamp 1607194113
transform 1 0 26864 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1254__A1_N
timestamp 1607194113
transform 1 0 26680 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_301
timestamp 1607194113
transform 1 0 28796 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_289
timestamp 1607194113
transform 1 0 27692 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0844_
timestamp 1607194113
transform 1 0 27416 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_318
timestamp 1607194113
transform 1 0 30360 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_306
timestamp 1607194113
transform 1 0 29256 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1607194113
transform 1 0 29164 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_69_330
timestamp 1607194113
transform 1 0 31464 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A1_N
timestamp 1607194113
transform 1 0 31556 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0784_
timestamp 1607194113
transform 1 0 31740 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_69_353
timestamp 1607194113
transform 1 0 33580 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A2_N
timestamp 1607194113
transform 1 0 33396 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__B2
timestamp 1607194113
transform 1 0 33212 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_379
timestamp 1607194113
transform 1 0 35972 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_367
timestamp 1607194113
transform 1 0 34868 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_365
timestamp 1607194113
transform 1 0 34684 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1607194113
transform 1 0 34776 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__B1
timestamp 1607194113
transform 1 0 37076 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0711_
timestamp 1607194113
transform 1 0 37260 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_69_413
timestamp 1607194113
transform 1 0 39100 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__B2
timestamp 1607194113
transform 1 0 38916 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__A2_N
timestamp 1607194113
transform 1 0 38732 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_437
timestamp 1607194113
transform 1 0 41308 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_425
timestamp 1607194113
transform 1 0 40204 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1607194113
transform 1 0 40388 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0719_
timestamp 1607194113
transform 1 0 40480 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_69_460
timestamp 1607194113
transform 1 0 43424 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_452
timestamp 1607194113
transform 1 0 42688 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_445
timestamp 1607194113
transform 1 0 42044 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_clk_i_A
timestamp 1607194113
transform 1 0 42504 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_clk_i
timestamp 1607194113
transform 1 0 42228 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _0847_
timestamp 1607194113
transform 1 0 43516 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_69_479
timestamp 1607194113
transform 1 0 45172 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A2_N
timestamp 1607194113
transform 1 0 44988 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_487
timestamp 1607194113
transform 1 0 45908 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1607194113
transform 1 0 46000 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_257
timestamp 1607194113
transform 1 0 24748 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_245
timestamp 1607194113
transform 1 0 23644 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_269
timestamp 1607194113
transform 1 0 25852 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_597
timestamp 1607194113
transform 1 0 26404 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1388_
timestamp 1607194113
transform 1 0 26496 0 -1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_70_297
timestamp 1607194113
transform 1 0 28428 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1388__CLK
timestamp 1607194113
transform 1 0 28244 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_320
timestamp 1607194113
transform 1 0 30544 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_309
timestamp 1607194113
transform 1 0 29532 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_clk_i
timestamp 1607194113
transform 1 0 30268 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_70_332
timestamp 1607194113
transform 1 0 31648 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__B1
timestamp 1607194113
transform 1 0 31832 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_598
timestamp 1607194113
transform 1 0 32016 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0780_
timestamp 1607194113
transform 1 0 32108 0 -1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_70_357
timestamp 1607194113
transform 1 0 33948 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__B2
timestamp 1607194113
transform 1 0 33764 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A2_N
timestamp 1607194113
transform 1 0 33580 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_381
timestamp 1607194113
transform 1 0 36156 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_369
timestamp 1607194113
transform 1 0 35052 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_393
timestamp 1607194113
transform 1 0 37260 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__A1_N
timestamp 1607194113
transform 1 0 37444 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_599
timestamp 1607194113
transform 1 0 37628 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0716_
timestamp 1607194113
transform 1 0 37720 0 -1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_70_418
timestamp 1607194113
transform 1 0 39560 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__A2_N
timestamp 1607194113
transform 1 0 39376 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__B2
timestamp 1607194113
transform 1 0 39192 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_442
timestamp 1607194113
transform 1 0 41768 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_430
timestamp 1607194113
transform 1 0 40664 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__B1
timestamp 1607194113
transform 1 0 42872 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__A1_N
timestamp 1607194113
transform 1 0 43056 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_600
timestamp 1607194113
transform 1 0 43240 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0769_
timestamp 1607194113
transform 1 0 43332 0 -1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_70_479
timestamp 1607194113
transform 1 0 45172 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__A2_N
timestamp 1607194113
transform 1 0 44988 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__B2
timestamp 1607194113
transform 1 0 44804 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_257
timestamp 1607194113
transform 1 0 24748 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_245
timestamp 1607194113
transform 1 0 23644 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__A
timestamp 1607194113
transform 1 0 24932 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1177_
timestamp 1607194113
transform 1 0 25116 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_265
timestamp 1607194113
transform 1 0 25484 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A2
timestamp 1607194113
transform 1 0 26036 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0870_
timestamp 1607194113
transform 1 0 26220 0 1 40800
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_71_303
timestamp 1607194113
transform 1 0 28980 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_291
timestamp 1607194113
transform 1 0 27876 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__B1
timestamp 1607194113
transform 1 0 27692 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A1
timestamp 1607194113
transform 1 0 27508 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_318
timestamp 1607194113
transform 1 0 30360 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_306
timestamp 1607194113
transform 1 0 29256 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_616
timestamp 1607194113
transform 1 0 29164 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_71_326
timestamp 1607194113
transform 1 0 31096 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__A1_N
timestamp 1607194113
transform 1 0 31372 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__B1
timestamp 1607194113
transform 1 0 31556 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0852_
timestamp 1607194113
transform 1 0 31740 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_71_360
timestamp 1607194113
transform 1 0 34224 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_71_353
timestamp 1607194113
transform 1 0 33580 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__B2
timestamp 1607194113
transform 1 0 33396 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__A2_N
timestamp 1607194113
transform 1 0 33212 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_clk_i
timestamp 1607194113
transform 1 0 33948 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_379
timestamp 1607194113
transform 1 0 35972 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_367
timestamp 1607194113
transform 1 0 34868 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_617
timestamp 1607194113
transform 1 0 34776 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_387
timestamp 1607194113
transform 1 0 36708 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__B1
timestamp 1607194113
transform 1 0 36800 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0807_
timestamp 1607194113
transform 1 0 36984 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_71_422
timestamp 1607194113
transform 1 0 39928 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_410
timestamp 1607194113
transform 1 0 38824 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__B2
timestamp 1607194113
transform 1 0 38640 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__A2_N
timestamp 1607194113
transform 1 0 38456 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_440
timestamp 1607194113
transform 1 0 41584 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_428
timestamp 1607194113
transform 1 0 40480 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_426
timestamp 1607194113
transform 1 0 40296 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_618
timestamp 1607194113
transform 1 0 40388 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_452
timestamp 1607194113
transform 1 0 42688 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_482
timestamp 1607194113
transform 1 0 45448 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A2_N
timestamp 1607194113
transform 1 0 45264 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0772_
timestamp 1607194113
transform 1 0 43792 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_619
timestamp 1607194113
transform 1 0 46000 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_72_248
timestamp 1607194113
transform 1 0 23920 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A2
timestamp 1607194113
transform 1 0 24196 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0874_
timestamp 1607194113
transform 1 0 24380 0 -1 41888
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_72_271
timestamp 1607194113
transform 1 0 26036 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__A2
timestamp 1607194113
transform 1 0 26220 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__B1
timestamp 1607194113
transform 1 0 25852 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A1
timestamp 1607194113
transform 1 0 25668 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_634
timestamp 1607194113
transform 1 0 26404 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0872_
timestamp 1607194113
transform 1 0 26496 0 -1 41888
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_72_294
timestamp 1607194113
transform 1 0 28152 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__B1
timestamp 1607194113
transform 1 0 27968 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__A1
timestamp 1607194113
transform 1 0 27784 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_318
timestamp 1607194113
transform 1 0 30360 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_306
timestamp 1607194113
transform 1 0 29256 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_clk_i
timestamp 1607194113
transform 1 0 30728 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_72_335
timestamp 1607194113
transform 1 0 31924 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_325
timestamp 1607194113
transform 1 0 31004 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__B1
timestamp 1607194113
transform 1 0 31740 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A1_N
timestamp 1607194113
transform 1 0 31556 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_635
timestamp 1607194113
transform 1 0 32016 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0855_
timestamp 1607194113
transform 1 0 32108 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A2_N
timestamp 1607194113
transform 1 0 33764 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__A2_N
timestamp 1607194113
transform 1 0 34132 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__B2
timestamp 1607194113
transform 1 0 33948 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__B2
timestamp 1607194113
transform 1 0 33580 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1238_
timestamp 1607194113
transform 1 0 34316 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_72_379
timestamp 1607194113
transform 1 0 35972 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__A1_N
timestamp 1607194113
transform 1 0 35788 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_398
timestamp 1607194113
transform 1 0 37720 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_391
timestamp 1607194113
transform 1 0 37076 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A1_N
timestamp 1607194113
transform 1 0 37444 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_636
timestamp 1607194113
transform 1 0 37628 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0811_
timestamp 1607194113
transform 1 0 37812 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_72_419
timestamp 1607194113
transform 1 0 39652 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A2_N
timestamp 1607194113
transform 1 0 39468 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__B2
timestamp 1607194113
transform 1 0 39284 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_431
timestamp 1607194113
transform 1 0 40756 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_459
timestamp 1607194113
transform 1 0 43332 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_450
timestamp 1607194113
transform 1 0 42504 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_443
timestamp 1607194113
transform 1 0 41860 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A1_N
timestamp 1607194113
transform 1 0 43516 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_637
timestamp 1607194113
transform 1 0 43240 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0839_
timestamp 1607194113
transform 1 0 42228 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__B1
timestamp 1607194113
transform 1 0 43700 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A2_N
timestamp 1607194113
transform 1 0 45356 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0753_
timestamp 1607194113
transform 1 0 43884 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_72_485
timestamp 1607194113
transform 1 0 45724 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__B2
timestamp 1607194113
transform 1 0 45540 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_257
timestamp 1607194113
transform 1 0 24748 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_245
timestamp 1607194113
transform 1 0 23644 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_265
timestamp 1607194113
transform 1 0 25484 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__A2_N
timestamp 1607194113
transform 1 0 25576 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__B1
timestamp 1607194113
transform 1 0 25760 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1178_
timestamp 1607194113
transform 1 0 25944 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_73_300
timestamp 1607194113
transform 1 0 28704 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_288
timestamp 1607194113
transform 1 0 27600 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__A1_N
timestamp 1607194113
transform 1 0 27416 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_318
timestamp 1607194113
transform 1 0 30360 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_306
timestamp 1607194113
transform 1 0 29256 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_304
timestamp 1607194113
transform 1 0 29072 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_653
timestamp 1607194113
transform 1 0 29164 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_330
timestamp 1607194113
transform 1 0 31464 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__A2_N
timestamp 1607194113
transform 1 0 32016 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__B2
timestamp 1607194113
transform 1 0 32200 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__B1
timestamp 1607194113
transform 1 0 32384 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1174_
timestamp 1607194113
transform 1 0 32568 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_73_363
timestamp 1607194113
transform 1 0 34500 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_73_358
timestamp 1607194113
transform 1 0 34040 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__A1_N
timestamp 1607194113
transform 1 0 34316 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1238__B1
timestamp 1607194113
transform 1 0 34132 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_379
timestamp 1607194113
transform 1 0 35972 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_367
timestamp 1607194113
transform 1 0 34868 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_654
timestamp 1607194113
transform 1 0 34776 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_387
timestamp 1607194113
transform 1 0 36708 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__A1_N
timestamp 1607194113
transform 1 0 36800 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__B1
timestamp 1607194113
transform 1 0 36984 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0718_
timestamp 1607194113
transform 1 0 37168 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_73_419
timestamp 1607194113
transform 1 0 39652 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_73_412
timestamp 1607194113
transform 1 0 39008 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__A2_N
timestamp 1607194113
transform 1 0 38824 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__B2
timestamp 1607194113
transform 1 0 38640 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0848_
timestamp 1607194113
transform 1 0 39376 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_431
timestamp 1607194113
transform 1 0 40756 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_655
timestamp 1607194113
transform 1 0 40388 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0773_
timestamp 1607194113
transform 1 0 40480 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1440__CLK
timestamp 1607194113
transform 1 0 41860 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1440_
timestamp 1607194113
transform 1 0 42044 0 1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_73_475
timestamp 1607194113
transform 1 0 44804 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_464
timestamp 1607194113
transform 1 0 43792 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0762_
timestamp 1607194113
transform 1 0 44528 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_73_487
timestamp 1607194113
transform 1 0 45908 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_656
timestamp 1607194113
transform 1 0 46000 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_257
timestamp 1607194113
transform 1 0 24748 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_245
timestamp 1607194113
transform 1 0 23644 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_246
timestamp 1607194113
transform 1 0 23736 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__A2_N
timestamp 1607194113
transform 1 0 23828 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__B1
timestamp 1607194113
transform 1 0 24012 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1242_
timestamp 1607194113
transform 1 0 24196 0 -1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_75_277
timestamp 1607194113
transform 1 0 26588 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_269
timestamp 1607194113
transform 1 0 25852 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_276
timestamp 1607194113
transform 1 0 26496 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_74_269
timestamp 1607194113
transform 1 0 25852 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1242__A1_N
timestamp 1607194113
transform 1 0 25668 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_671
timestamp 1607194113
transform 1 0 26404 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1438_
timestamp 1607194113
transform 1 0 26680 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1397_
timestamp 1607194113
transform 1 0 26680 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_75_299
timestamp 1607194113
transform 1 0 28612 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_74_299
timestamp 1607194113
transform 1 0 28612 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1438__CLK
timestamp 1607194113
transform 1 0 28428 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1397__CLK
timestamp 1607194113
transform 1 0 28428 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_318
timestamp 1607194113
transform 1 0 30360 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_306
timestamp 1607194113
transform 1 0 29256 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_320
timestamp 1607194113
transform 1 0 30544 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_308
timestamp 1607194113
transform 1 0 29440 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_690
timestamp 1607194113
transform 1 0 29164 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0765_
timestamp 1607194113
transform 1 0 29164 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_75_330
timestamp 1607194113
transform 1 0 31464 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_332
timestamp 1607194113
transform 1 0 31648 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__A2_N
timestamp 1607194113
transform 1 0 32016 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__B2
timestamp 1607194113
transform 1 0 32200 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__A2_N
timestamp 1607194113
transform 1 0 32108 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__B2
timestamp 1607194113
transform 1 0 32292 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__B1
timestamp 1607194113
transform 1 0 32476 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__B1
timestamp 1607194113
transform 1 0 32384 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_672
timestamp 1607194113
transform 1 0 32016 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1239_
timestamp 1607194113
transform 1 0 32568 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _1175_
timestamp 1607194113
transform 1 0 32660 0 -1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_75_360
timestamp 1607194113
transform 1 0 34224 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_74_361
timestamp 1607194113
transform 1 0 34316 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1239__A1_N
timestamp 1607194113
transform 1 0 34040 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__A1_N
timestamp 1607194113
transform 1 0 34132 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_379
timestamp 1607194113
transform 1 0 35972 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_367
timestamp 1607194113
transform 1 0 34868 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_365
timestamp 1607194113
transform 1 0 34684 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1398__CLK
timestamp 1607194113
transform 1 0 34776 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_691
timestamp 1607194113
transform 1 0 34776 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1398_
timestamp 1607194113
transform 1 0 34960 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_75_387
timestamp 1607194113
transform 1 0 36708 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_387
timestamp 1607194113
transform 1 0 36708 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__A1_N
timestamp 1607194113
transform 1 0 36800 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__B1
timestamp 1607194113
transform 1 0 36984 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_398
timestamp 1607194113
transform 1 0 37720 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_395
timestamp 1607194113
transform 1 0 37444 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1439__CLK
timestamp 1607194113
transform 1 0 37812 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_673
timestamp 1607194113
transform 1 0 37628 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1439_
timestamp 1607194113
transform 1 0 37996 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__a2bb2o_4  _0813_
timestamp 1607194113
transform 1 0 37168 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_75_412
timestamp 1607194113
transform 1 0 39008 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_420
timestamp 1607194113
transform 1 0 39744 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__A2_N
timestamp 1607194113
transform 1 0 38824 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__B2
timestamp 1607194113
transform 1 0 38640 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_428
timestamp 1607194113
transform 1 0 40480 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_75_424
timestamp 1607194113
transform 1 0 40112 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_432
timestamp 1607194113
transform 1 0 40848 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1399__CLK
timestamp 1607194113
transform 1 0 40848 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_692
timestamp 1607194113
transform 1 0 40388 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1399_
timestamp 1607194113
transform 1 0 41032 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_75_453
timestamp 1607194113
transform 1 0 42780 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_459
timestamp 1607194113
transform 1 0 43332 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_456
timestamp 1607194113
transform 1 0 43056 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_444
timestamp 1607194113
transform 1 0 41952 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_674
timestamp 1607194113
transform 1 0 43240 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_477
timestamp 1607194113
transform 1 0 44988 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_465
timestamp 1607194113
transform 1 0 43884 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A1_N
timestamp 1607194113
transform 1 0 44436 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__B1
timestamp 1607194113
transform 1 0 44620 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0767_
timestamp 1607194113
transform 1 0 44804 0 -1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_75_485
timestamp 1607194113
transform 1 0 45724 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_693
timestamp 1607194113
transform 1 0 46000 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_261
timestamp 1607194113
transform 1 0 25116 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_249
timestamp 1607194113
transform 1 0 24012 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_711
timestamp 1607194113
transform 1 0 23920 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_280
timestamp 1607194113
transform 1 0 26864 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_273
timestamp 1607194113
transform 1 0 26220 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_712
timestamp 1607194113
transform 1 0 26772 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_298
timestamp 1607194113
transform 1 0 28520 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_292
timestamp 1607194113
transform 1 0 27968 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0842_
timestamp 1607194113
transform 1 0 28244 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_323
timestamp 1607194113
transform 1 0 30820 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_311
timestamp 1607194113
transform 1 0 29716 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_713
timestamp 1607194113
transform 1 0 29624 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_342
timestamp 1607194113
transform 1 0 32568 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_335
timestamp 1607194113
transform 1 0 31924 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_714
timestamp 1607194113
transform 1 0 32476 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_354
timestamp 1607194113
transform 1 0 33672 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_373
timestamp 1607194113
transform 1 0 35420 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_366
timestamp 1607194113
transform 1 0 34776 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_715
timestamp 1607194113
transform 1 0 35328 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_397
timestamp 1607194113
transform 1 0 37628 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_385
timestamp 1607194113
transform 1 0 36524 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_416
timestamp 1607194113
transform 1 0 39376 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_404
timestamp 1607194113
transform 1 0 38272 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_716
timestamp 1607194113
transform 1 0 38180 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_435
timestamp 1607194113
transform 1 0 41124 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_428
timestamp 1607194113
transform 1 0 40480 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_717
timestamp 1607194113
transform 1 0 41032 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_459
timestamp 1607194113
transform 1 0 43332 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_447
timestamp 1607194113
transform 1 0 42228 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_466
timestamp 1607194113
transform 1 0 43976 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__B1
timestamp 1607194113
transform 1 0 44068 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A1_N
timestamp 1607194113
transform 1 0 44252 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_718
timestamp 1607194113
transform 1 0 43884 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0774_
timestamp 1607194113
transform 1 0 44436 0 -1 44064
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__B2
timestamp 1607194113
transform 1 0 45908 0 -1 44064
box -38 -48 222 592
use delayline_9_ms  inst_tdelay_line
timestamp 1607276512
transform 1 0 26680 0 1 3761
box 800 801 23264 27367
use sky130_fd_sc_hd__decap_12  FILLER_59_501
timestamp 1607194113
transform 1 0 47196 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_489
timestamp 1607194113
transform 1 0 46092 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_513
timestamp 1607194113
transform 1 0 48300 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_i_A
timestamp 1607194113
transform 1 0 48392 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk_i $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 48576 0 1 34272
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_59_550
timestamp 1607194113
transform 1 0 51704 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_548
timestamp 1607194113
transform 1 0 51520 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_536
timestamp 1607194113
transform 1 0 50416 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1607194113
transform 1 0 51612 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_clk_i_A
timestamp 1607194113
transform 1 0 52256 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_clk_i
timestamp 1607194113
transform 1 0 52440 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1515_
timestamp 1607194113
transform 1 0 52716 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_59_592
timestamp 1607194113
transform 1 0 55568 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_inp_i
timestamp 1607194113
transform 1 0 54648 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[8]
timestamp 1607194113
transform 1 0 54464 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[7]
timestamp 1607194113
transform 1 0 54832 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[6]
timestamp 1607194113
transform 1 0 55384 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[4]
timestamp 1607194113
transform 1 0 55200 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[2]
timestamp 1607194113
transform 1 0 55016 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_59_609
timestamp 1607194113
transform 1 0 57132 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_604
timestamp 1607194113
transform 1 0 56672 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A1_N
timestamp 1607194113
transform 1 0 56948 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__B1
timestamp 1607194113
transform 1 0 56764 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1607194113
transform 1 0 57224 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0825_
timestamp 1607194113
transform 1 0 57316 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_59_631
timestamp 1607194113
transform 1 0 59156 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__B2
timestamp 1607194113
transform 1 0 58972 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A2_N
timestamp 1607194113
transform 1 0 58788 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_655
timestamp 1607194113
transform 1 0 61364 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_643
timestamp 1607194113
transform 1 0 60260 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__A1_N
timestamp 1607194113
transform 1 0 62468 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__B1
timestamp 1607194113
transform 1 0 62652 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1607194113
transform 1 0 62836 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0727_
timestamp 1607194113
transform 1 0 62928 0 1 34272
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_59_692
timestamp 1607194113
transform 1 0 64768 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__A2_N
timestamp 1607194113
transform 1 0 64584 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__B2
timestamp 1607194113
transform 1 0 64400 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_700
timestamp 1607194113
transform 1 0 65504 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1516__CLK
timestamp 1607194113
transform 1 0 65780 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1516_
timestamp 1607194113
transform 1 0 65964 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_59_724
timestamp 1607194113
transform 1 0 67712 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1607194113
transform 1 0 68448 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_493
timestamp 1607194113
transform 1 0 46460 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A1_N
timestamp 1607194113
transform 1 0 46552 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__B1
timestamp 1607194113
transform 1 0 46736 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0740_
timestamp 1607194113
transform 1 0 46920 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_60_520
timestamp 1607194113
transform 1 0 48944 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_518
timestamp 1607194113
transform 1 0 48760 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__B2
timestamp 1607194113
transform 1 0 48576 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A2_N
timestamp 1607194113
transform 1 0 48392 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__B1
timestamp 1607194113
transform 1 0 49680 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__A1_N
timestamp 1607194113
transform 1 0 49864 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1607194113
transform 1 0 48852 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__B2
timestamp 1607194113
transform 1 0 51704 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__A2_N
timestamp 1607194113
transform 1 0 51520 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0732_
timestamp 1607194113
transform 1 0 50048 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_60_570
timestamp 1607194113
transform 1 0 53544 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_60_564
timestamp 1607194113
transform 1 0 52992 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_552
timestamp 1607194113
transform 1 0 51888 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1607194113
transform 1 0 53268 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_587
timestamp 1607194113
transform 1 0 55108 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_579
timestamp 1607194113
transform 1 0 54372 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_574
timestamp 1607194113
transform 1 0 53912 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1515__CLK
timestamp 1607194113
transform 1 0 54924 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[5]
timestamp 1607194113
transform 1 0 54740 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[3]
timestamp 1607194113
transform 1 0 54556 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[1]
timestamp 1607194113
transform 1 0 54188 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_idelay_line_en_i[0]
timestamp 1607194113
transform 1 0 54004 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1607194113
transform 1 0 54464 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__B1
timestamp 1607194113
transform 1 0 56396 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__A1_N
timestamp 1607194113
transform 1 0 56580 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__B2
timestamp 1607194113
transform 1 0 56212 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0821_
timestamp 1607194113
transform 1 0 56764 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_60_625
timestamp 1607194113
transform 1 0 58604 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__B2
timestamp 1607194113
transform 1 0 58420 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__A2_N
timestamp 1607194113
transform 1 0 58236 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_654
timestamp 1607194113
transform 1 0 61272 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_642
timestamp 1607194113
transform 1 0 60168 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_637
timestamp 1607194113
transform 1 0 59708 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1607194113
transform 1 0 60076 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_60_658
timestamp 1607194113
transform 1 0 61640 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A1_N
timestamp 1607194113
transform 1 0 61732 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__B1
timestamp 1607194113
transform 1 0 61916 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0818_
timestamp 1607194113
transform 1 0 62100 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_60_694
timestamp 1607194113
transform 1 0 64952 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_60_683
timestamp 1607194113
transform 1 0 63940 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A2_N
timestamp 1607194113
transform 1 0 63756 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__B2
timestamp 1607194113
transform 1 0 63572 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0788_
timestamp 1607194113
transform 1 0 64676 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_60_703
timestamp 1607194113
transform 1 0 65780 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__A2_N
timestamp 1607194113
transform 1 0 65872 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__B2
timestamp 1607194113
transform 1 0 66056 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__B1
timestamp 1607194113
transform 1 0 66240 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1607194113
transform 1 0 65688 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1204_
timestamp 1607194113
transform 1 0 66424 0 -1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_60_726
timestamp 1607194113
transform 1 0 67896 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_502
timestamp 1607194113
transform 1 0 47288 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_490
timestamp 1607194113
transform 1 0 46184 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_501
timestamp 1607194113
transform 1 0 47196 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_489
timestamp 1607194113
transform 1 0 46092 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_518
timestamp 1607194113
transform 1 0 48760 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_514
timestamp 1607194113
transform 1 0 48392 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_517
timestamp 1607194113
transform 1 0 48668 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_513
timestamp 1607194113
transform 1 0 48300 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A1_N
timestamp 1607194113
transform 1 0 48760 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1607194113
transform 1 0 48852 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_62_520
timestamp 1607194113
transform 1 0 48944 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__B1
timestamp 1607194113
transform 1 0 49036 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__B1
timestamp 1607194113
transform 1 0 48944 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A1_N
timestamp 1607194113
transform 1 0 49220 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0759_
timestamp 1607194113
transform 1 0 49404 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _0736_
timestamp 1607194113
transform 1 0 49128 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_62_545
timestamp 1607194113
transform 1 0 51244 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_548
timestamp 1607194113
transform 1 0 51520 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_542
timestamp 1607194113
transform 1 0 50968 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__B2
timestamp 1607194113
transform 1 0 50784 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A2_N
timestamp 1607194113
transform 1 0 50600 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__B2
timestamp 1607194113
transform 1 0 51060 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A2_N
timestamp 1607194113
transform 1 0 50876 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1607194113
transform 1 0 51612 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0741_
timestamp 1607194113
transform 1 0 51704 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_62_569
timestamp 1607194113
transform 1 0 53452 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_557
timestamp 1607194113
transform 1 0 52348 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_571
timestamp 1607194113
transform 1 0 53636 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_559
timestamp 1607194113
transform 1 0 52532 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_581
timestamp 1607194113
transform 1 0 54556 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_577
timestamp 1607194113
transform 1 0 54188 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_579
timestamp 1607194113
transform 1 0 54372 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__B1
timestamp 1607194113
transform 1 0 54648 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A1_N
timestamp 1607194113
transform 1 0 54832 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1607194113
transform 1 0 54464 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0838_
timestamp 1607194113
transform 1 0 55016 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  FILLER_62_593
timestamp 1607194113
transform 1 0 55660 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__B1
timestamp 1607194113
transform 1 0 55936 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__B1
timestamp 1607194113
transform 1 0 56488 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A1_N
timestamp 1607194113
transform 1 0 56120 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_609
timestamp 1607194113
transform 1 0 57132 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_606
timestamp 1607194113
transform 1 0 56856 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A2_N
timestamp 1607194113
transform 1 0 56672 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A1_N
timestamp 1607194113
transform 1 0 56948 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1607194113
transform 1 0 57224 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0837_
timestamp 1607194113
transform 1 0 56304 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _0823_
timestamp 1607194113
transform 1 0 57316 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_62_633
timestamp 1607194113
transform 1 0 59340 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_620
timestamp 1607194113
transform 1 0 58144 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_631
timestamp 1607194113
transform 1 0 59156 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__B2
timestamp 1607194113
transform 1 0 58972 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A2_N
timestamp 1607194113
transform 1 0 58788 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__B2
timestamp 1607194113
transform 1 0 57960 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A2_N
timestamp 1607194113
transform 1 0 57776 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0826_
timestamp 1607194113
transform 1 0 58512 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_62_654
timestamp 1607194113
transform 1 0 61272 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_642
timestamp 1607194113
transform 1 0 60168 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_655
timestamp 1607194113
transform 1 0 61364 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_643
timestamp 1607194113
transform 1 0 60260 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1607194113
transform 1 0 60076 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_662
timestamp 1607194113
transform 1 0 62008 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_61_672
timestamp 1607194113
transform 1 0 62928 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_667
timestamp 1607194113
transform 1 0 62468 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__B2
timestamp 1607194113
transform 1 0 62284 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__B2
timestamp 1607194113
transform 1 0 63020 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A2
timestamp 1607194113
transform 1 0 62468 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A2
timestamp 1607194113
transform 1 0 63204 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1607194113
transform 1 0 62836 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0927_
timestamp 1607194113
transform 1 0 62652 0 -1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_62_695
timestamp 1607194113
transform 1 0 65044 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_683
timestamp 1607194113
transform 1 0 63940 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_691
timestamp 1607194113
transform 1 0 64676 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _0933_
timestamp 1607194113
transform 1 0 63388 0 1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_62_715
timestamp 1607194113
transform 1 0 66884 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_703
timestamp 1607194113
transform 1 0 65780 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_701
timestamp 1607194113
transform 1 0 65596 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_699
timestamp 1607194113
transform 1 0 65412 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__A2_N
timestamp 1607194113
transform 1 0 65688 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__B2
timestamp 1607194113
transform 1 0 65872 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1267__B1
timestamp 1607194113
transform 1 0 66056 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1607194113
transform 1 0 65688 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1267_
timestamp 1607194113
transform 1 0 66240 0 1 35360
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_62_727
timestamp 1607194113
transform 1 0 67988 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_724
timestamp 1607194113
transform 1 0 67712 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1607194113
transform 1 0 68448 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_489
timestamp 1607194113
transform 1 0 46092 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1425__CLK
timestamp 1607194113
transform 1 0 46828 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1425_
timestamp 1607194113
transform 1 0 47012 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__B1
timestamp 1607194113
transform 1 0 48760 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0760_
timestamp 1607194113
transform 1 0 48944 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_63_550
timestamp 1607194113
transform 1 0 51704 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A2_N
timestamp 1607194113
transform 1 0 51244 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__B2
timestamp 1607194113
transform 1 0 51428 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1607194113
transform 1 0 51612 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0764_
timestamp 1607194113
transform 1 0 50416 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_63_556
timestamp 1607194113
transform 1 0 52256 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__B1
timestamp 1607194113
transform 1 0 52348 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0836_
timestamp 1607194113
transform 1 0 52532 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_1  FILLER_63_583
timestamp 1607194113
transform 1 0 54740 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_579
timestamp 1607194113
transform 1 0 54372 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__B2
timestamp 1607194113
transform 1 0 54832 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__A2
timestamp 1607194113
transform 1 0 55016 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A2_N
timestamp 1607194113
transform 1 0 54188 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__B2
timestamp 1607194113
transform 1 0 54004 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0931_
timestamp 1607194113
transform 1 0 55200 0 1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_63_609
timestamp 1607194113
transform 1 0 57132 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_63_602
timestamp 1607194113
transform 1 0 56488 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__A2_N
timestamp 1607194113
transform 1 0 56764 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__B2
timestamp 1607194113
transform 1 0 56948 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1265__B1
timestamp 1607194113
transform 1 0 56580 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1607194113
transform 1 0 57224 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _1265_
timestamp 1607194113
transform 1 0 57316 0 1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_63_627
timestamp 1607194113
transform 1 0 58788 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_651
timestamp 1607194113
transform 1 0 60996 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_639
timestamp 1607194113
transform 1 0 59892 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_672
timestamp 1607194113
transform 1 0 62928 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_663
timestamp 1607194113
transform 1 0 62100 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1607194113
transform 1 0 62836 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_63_684
timestamp 1607194113
transform 1 0 64032 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1422__CLK
timestamp 1607194113
transform 1 0 64308 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1422_
timestamp 1607194113
transform 1 0 64492 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_63_708
timestamp 1607194113
transform 1 0 66240 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_720
timestamp 1607194113
transform 1 0 67344 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1607194113
transform 1 0 68448 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_506
timestamp 1607194113
transform 1 0 47656 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_494
timestamp 1607194113
transform 1 0 46552 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0833_
timestamp 1607194113
transform 1 0 47840 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_64_526
timestamp 1607194113
transform 1 0 49496 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_520
timestamp 1607194113
transform 1 0 48944 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_511
timestamp 1607194113
transform 1 0 48116 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A1_N
timestamp 1607194113
transform 1 0 49312 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1607194113
transform 1 0 48852 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0754_
timestamp 1607194113
transform 1 0 49036 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__B2
timestamp 1607194113
transform 1 0 51704 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__B1
timestamp 1607194113
transform 1 0 50048 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0758_
timestamp 1607194113
transform 1 0 50232 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_64_566
timestamp 1607194113
transform 1 0 53176 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_554
timestamp 1607194113
transform 1 0 52072 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A2_N
timestamp 1607194113
transform 1 0 51888 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_590
timestamp 1607194113
transform 1 0 55384 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_578
timestamp 1607194113
transform 1 0 54280 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1607194113
transform 1 0 54464 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0841_
timestamp 1607194113
transform 1 0 54556 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_64_598
timestamp 1607194113
transform 1 0 56120 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__A2_N
timestamp 1607194113
transform 1 0 56212 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__B2
timestamp 1607194113
transform 1 0 56396 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__B1
timestamp 1607194113
transform 1 0 56580 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1202_
timestamp 1607194113
transform 1 0 56764 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_64_633
timestamp 1607194113
transform 1 0 59340 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_621
timestamp 1607194113
transform 1 0 58236 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_654
timestamp 1607194113
transform 1 0 61272 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_642
timestamp 1607194113
transform 1 0 60168 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1607194113
transform 1 0 60076 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_662
timestamp 1607194113
transform 1 0 62008 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__A2_N
timestamp 1607194113
transform 1 0 62192 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__B2
timestamp 1607194113
transform 1 0 62376 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__B1
timestamp 1607194113
transform 1 0 62560 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1201_
timestamp 1607194113
transform 1 0 62744 0 -1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_64_686
timestamp 1607194113
transform 1 0 64216 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_715
timestamp 1607194113
transform 1 0 66884 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_703
timestamp 1607194113
transform 1 0 65780 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_698
timestamp 1607194113
transform 1 0 65320 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1607194113
transform 1 0 65688 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_727
timestamp 1607194113
transform 1 0 67988 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_501
timestamp 1607194113
transform 1 0 47196 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_489
timestamp 1607194113
transform 1 0 46092 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_525
timestamp 1607194113
transform 1 0 49404 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_513
timestamp 1607194113
transform 1 0 48300 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_548
timestamp 1607194113
transform 1 0 51520 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_65_543
timestamp 1607194113
transform 1 0 51060 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_537
timestamp 1607194113
transform 1 0 50508 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A1_N
timestamp 1607194113
transform 1 0 51336 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__B1
timestamp 1607194113
transform 1 0 51152 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1607194113
transform 1 0 51612 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0840_
timestamp 1607194113
transform 1 0 51704 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_65_568
timestamp 1607194113
transform 1 0 53360 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A2_N
timestamp 1607194113
transform 1 0 53176 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_65_592
timestamp 1607194113
transform 1 0 55568 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_580
timestamp 1607194113
transform 1 0 54464 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_611
timestamp 1607194113
transform 1 0 57316 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_602
timestamp 1607194113
transform 1 0 56488 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_598
timestamp 1607194113
transform 1 0 56120 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1380__CLK
timestamp 1607194113
transform 1 0 57408 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1607194113
transform 1 0 57224 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0929_
timestamp 1607194113
transform 1 0 56212 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_633
timestamp 1607194113
transform 1 0 59340 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1380_
timestamp 1607194113
transform 1 0 57592 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_65_650
timestamp 1607194113
transform 1 0 60904 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__D
timestamp 1607194113
transform 1 0 59708 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__B
timestamp 1607194113
transform 1 0 59892 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0787_
timestamp 1607194113
transform 1 0 60076 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_65_672
timestamp 1607194113
transform 1 0 62928 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_670
timestamp 1607194113
transform 1 0 62744 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_662
timestamp 1607194113
transform 1 0 62008 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1607194113
transform 1 0 62836 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_684
timestamp 1607194113
transform 1 0 64032 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1381__CLK
timestamp 1607194113
transform 1 0 64216 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1381_
timestamp 1607194113
transform 1 0 64400 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_65_707
timestamp 1607194113
transform 1 0 66148 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_731
timestamp 1607194113
transform 1 0 68356 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_719
timestamp 1607194113
transform 1 0 67252 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1607194113
transform 1 0 68448 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_501
timestamp 1607194113
transform 1 0 47196 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_489
timestamp 1607194113
transform 1 0 46092 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_528
timestamp 1607194113
transform 1 0 49680 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_520
timestamp 1607194113
transform 1 0 48944 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_66_513
timestamp 1607194113
transform 1 0 48300 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__A1_N
timestamp 1607194113
transform 1 0 49772 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1607194113
transform 1 0 48852 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__B1
timestamp 1607194113
transform 1 0 49956 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__A2_N
timestamp 1607194113
transform 1 0 51612 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0763_
timestamp 1607194113
transform 1 0 50140 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_551
timestamp 1607194113
transform 1 0 51796 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _0858_
timestamp 1607194113
transform 1 0 52900 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_66_581
timestamp 1607194113
transform 1 0 54556 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_574
timestamp 1607194113
transform 1 0 53912 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__A
timestamp 1607194113
transform 1 0 53728 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1607194113
transform 1 0 54464 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_606
timestamp 1607194113
transform 1 0 56856 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_601
timestamp 1607194113
transform 1 0 56396 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_593
timestamp 1607194113
transform 1 0 55660 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1421__CLK
timestamp 1607194113
transform 1 0 57408 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0930_
timestamp 1607194113
transform 1 0 56580 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_633
timestamp 1607194113
transform 1 0 59340 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1421_
timestamp 1607194113
transform 1 0 57592 0 -1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_66_654
timestamp 1607194113
transform 1 0 61272 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_642
timestamp 1607194113
transform 1 0 60168 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1607194113
transform 1 0 60076 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_662
timestamp 1607194113
transform 1 0 62008 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__A2_N
timestamp 1607194113
transform 1 0 62100 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__B2
timestamp 1607194113
transform 1 0 62284 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1264__B1
timestamp 1607194113
transform 1 0 62468 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _1264_
timestamp 1607194113
transform 1 0 62652 0 -1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_66_685
timestamp 1607194113
transform 1 0 64124 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_715
timestamp 1607194113
transform 1 0 66884 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_703
timestamp 1607194113
transform 1 0 65780 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_701
timestamp 1607194113
transform 1 0 65596 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_697
timestamp 1607194113
transform 1 0 65228 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1607194113
transform 1 0 65688 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1389__CLK
timestamp 1607194113
transform 1 0 67252 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1389__D
timestamp 1607194113
transform 1 0 67436 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1389_
timestamp 1607194113
transform 1 0 67620 0 -1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_68_501
timestamp 1607194113
transform 1 0 47196 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_498
timestamp 1607194113
transform 1 0 46920 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _0786_
timestamp 1607194113
transform 1 0 46092 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0756_
timestamp 1607194113
transform 1 0 46368 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_68_518
timestamp 1607194113
transform 1 0 48760 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_68_513
timestamp 1607194113
transform 1 0 48300 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_514
timestamp 1607194113
transform 1 0 48392 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_510
timestamp 1607194113
transform 1 0 48024 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A1_N
timestamp 1607194113
transform 1 0 48576 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__B1
timestamp 1607194113
transform 1 0 48392 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__B1
timestamp 1607194113
transform 1 0 48484 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1607194113
transform 1 0 48852 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0834_
timestamp 1607194113
transform 1 0 48944 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _0755_
timestamp 1607194113
transform 1 0 48668 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_67_539
timestamp 1607194113
transform 1 0 50692 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__B2
timestamp 1607194113
transform 1 0 50508 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__B2
timestamp 1607194113
transform 1 0 50600 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A2_N
timestamp 1607194113
transform 1 0 50324 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A2_N
timestamp 1607194113
transform 1 0 50416 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A1_N
timestamp 1607194113
transform 1 0 50140 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_544
timestamp 1607194113
transform 1 0 51152 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_540
timestamp 1607194113
transform 1 0 50784 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_clk_i_A
timestamp 1607194113
transform 1 0 51428 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__D
timestamp 1607194113
transform 1 0 51428 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A1_N
timestamp 1607194113
transform 1 0 51244 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_clk_i
timestamp 1607194113
transform 1 0 51612 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1607194113
transform 1 0 51612 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0857_
timestamp 1607194113
transform 1 0 51704 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_67_571
timestamp 1607194113
transform 1 0 53636 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_559
timestamp 1607194113
transform 1 0 52532 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A2_N
timestamp 1607194113
transform 1 0 53544 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__B2
timestamp 1607194113
transform 1 0 53360 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0809_
timestamp 1607194113
transform 1 0 51888 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_6  FILLER_68_572
timestamp 1607194113
transform 1 0 53728 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_591
timestamp 1607194113
transform 1 0 55476 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_579
timestamp 1607194113
transform 1 0 54372 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_575
timestamp 1607194113
transform 1 0 54004 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__CLK
timestamp 1607194113
transform 1 0 54556 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1434__D
timestamp 1607194113
transform 1 0 54280 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_clk_i
timestamp 1607194113
transform 1 0 54096 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1607194113
transform 1 0 54464 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1434_
timestamp 1607194113
transform 1 0 54740 0 -1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_68_602
timestamp 1607194113
transform 1 0 56488 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_611
timestamp 1607194113
transform 1 0 57316 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_67_609
timestamp 1607194113
transform 1 0 57132 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_67_603
timestamp 1607194113
transform 1 0 56580 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1607194113
transform 1 0 57224 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_614
timestamp 1607194113
transform 1 0 57592 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_619
timestamp 1607194113
transform 1 0 58052 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__B1
timestamp 1607194113
transform 1 0 58236 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__A2_N
timestamp 1607194113
transform 1 0 59340 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0817_
timestamp 1607194113
transform 1 0 57868 0 -1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _0724_
timestamp 1607194113
transform 1 0 58420 0 1 38624
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_68_637
timestamp 1607194113
transform 1 0 59708 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_641
timestamp 1607194113
transform 1 0 60076 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__B1
timestamp 1607194113
transform 1 0 59524 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__A2_N
timestamp 1607194113
transform 1 0 59892 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1607194113
transform 1 0 60076 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0827_
timestamp 1607194113
transform 1 0 60168 0 -1 39712
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_4  _0742_
timestamp 1607194113
transform 1 0 60628 0 1 38624
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_68_668
timestamp 1607194113
transform 1 0 62560 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_662
timestamp 1607194113
transform 1 0 62008 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_68_656
timestamp 1607194113
transform 1 0 61456 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_672
timestamp 1607194113
transform 1 0 62928 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_669
timestamp 1607194113
transform 1 0 62652 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_661
timestamp 1607194113
transform 1 0 61916 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_clk_i_A
timestamp 1607194113
transform 1 0 62100 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_clk_i
timestamp 1607194113
transform 1 0 62284 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1607194113
transform 1 0 62836 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_692
timestamp 1607194113
transform 1 0 64768 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_680
timestamp 1607194113
transform 1 0 63664 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_696
timestamp 1607194113
transform 1 0 65136 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_684
timestamp 1607194113
transform 1 0 64032 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_700
timestamp 1607194113
transform 1 0 65504 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_717
timestamp 1607194113
transform 1 0 67068 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_705
timestamp 1607194113
transform 1 0 65964 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1476__CLK
timestamp 1607194113
transform 1 0 65780 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__A
timestamp 1607194113
transform 1 0 65780 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1607194113
transform 1 0 65688 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1476_
timestamp 1607194113
transform 1 0 65964 0 -1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0776_
timestamp 1607194113
transform 1 0 65504 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_724
timestamp 1607194113
transform 1 0 67712 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_729
timestamp 1607194113
transform 1 0 68172 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1607194113
transform 1 0 68448 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_501
timestamp 1607194113
transform 1 0 47196 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_489
timestamp 1607194113
transform 1 0 46092 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_521
timestamp 1607194113
transform 1 0 49036 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_513
timestamp 1607194113
transform 1 0 48300 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__or4_4  _0835_
timestamp 1607194113
transform 1 0 49312 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_69_550
timestamp 1607194113
transform 1 0 51704 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_545
timestamp 1607194113
transform 1 0 51244 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_533
timestamp 1607194113
transform 1 0 50140 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__A1_N
timestamp 1607194113
transform 1 0 51428 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1607194113
transform 1 0 51612 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_571
timestamp 1607194113
transform 1 0 53636 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__A2_N
timestamp 1607194113
transform 1 0 53452 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__B2
timestamp 1607194113
transform 1 0 53268 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0714_
timestamp 1607194113
transform 1 0 51796 0 1 39712
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_69_591
timestamp 1607194113
transform 1 0 55476 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_579
timestamp 1607194113
transform 1 0 54372 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_575
timestamp 1607194113
transform 1 0 54004 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_clk_i
timestamp 1607194113
transform 1 0 54096 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_69_609
timestamp 1607194113
transform 1 0 57132 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_603
timestamp 1607194113
transform 1 0 56580 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__CLK
timestamp 1607194113
transform 1 0 56948 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1393__D
timestamp 1607194113
transform 1 0 56764 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1607194113
transform 1 0 57224 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1393_
timestamp 1607194113
transform 1 0 57316 0 1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_69_630
timestamp 1607194113
transform 1 0 59064 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_654
timestamp 1607194113
transform 1 0 61272 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_642
timestamp 1607194113
transform 1 0 60168 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_69_672
timestamp 1607194113
transform 1 0 62928 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_69_670
timestamp 1607194113
transform 1 0 62744 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_666
timestamp 1607194113
transform 1 0 62376 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1607194113
transform 1 0 62836 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0721_
timestamp 1607194113
transform 1 0 63204 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_69_678
timestamp 1607194113
transform 1 0 63480 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1475__CLK
timestamp 1607194113
transform 1 0 64032 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1475_
timestamp 1607194113
transform 1 0 64216 0 1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_69_705
timestamp 1607194113
transform 1 0 65964 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1075_
timestamp 1607194113
transform 1 0 66700 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_69_724
timestamp 1607194113
transform 1 0 67712 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__A
timestamp 1607194113
transform 1 0 67528 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1607194113
transform 1 0 68448 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_503
timestamp 1607194113
transform 1 0 47380 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_491
timestamp 1607194113
transform 1 0 46276 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_524
timestamp 1607194113
transform 1 0 49312 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_520
timestamp 1607194113
transform 1 0 48944 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_515
timestamp 1607194113
transform 1 0 48484 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_601
timestamp 1607194113
transform 1 0 48852 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0850_
timestamp 1607194113
transform 1 0 49404 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_70_546
timestamp 1607194113
transform 1 0 51336 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_534
timestamp 1607194113
transform 1 0 50232 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_570
timestamp 1607194113
transform 1 0 53544 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_558
timestamp 1607194113
transform 1 0 52440 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_589
timestamp 1607194113
transform 1 0 55292 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_581
timestamp 1607194113
transform 1 0 54556 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_578
timestamp 1607194113
transform 1 0 54280 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_602
timestamp 1607194113
transform 1 0 54464 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1054_
timestamp 1607194113
transform 1 0 54648 0 -1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_70_613
timestamp 1607194113
transform 1 0 57500 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_601
timestamp 1607194113
transform 1 0 56396 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_630
timestamp 1607194113
transform 1 0 59064 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_70_619
timestamp 1607194113
transform 1 0 58052 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0816_
timestamp 1607194113
transform 1 0 58788 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0723_
timestamp 1607194113
transform 1 0 57776 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_654
timestamp 1607194113
transform 1 0 61272 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_642
timestamp 1607194113
transform 1 0 60168 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_638
timestamp 1607194113
transform 1 0 59800 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_603
timestamp 1607194113
transform 1 0 60076 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_666
timestamp 1607194113
transform 1 0 62376 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _1077_
timestamp 1607194113
transform 1 0 62744 0 -1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_70_696
timestamp 1607194113
transform 1 0 65136 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_677
timestamp 1607194113
transform 1 0 63388 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__A
timestamp 1607194113
transform 1 0 64952 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1078_
timestamp 1607194113
transform 1 0 64124 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_70_712
timestamp 1607194113
transform 1 0 66608 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__A
timestamp 1607194113
transform 1 0 65504 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_604
timestamp 1607194113
transform 1 0 65688 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1074_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 65780 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_70_727
timestamp 1607194113
transform 1 0 67988 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__A
timestamp 1607194113
transform 1 0 67160 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1070_
timestamp 1607194113
transform 1 0 67344 0 -1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_71_501
timestamp 1607194113
transform 1 0 47196 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_489
timestamp 1607194113
transform 1 0 46092 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__A1_N
timestamp 1607194113
transform 1 0 47932 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__B1
timestamp 1607194113
transform 1 0 48116 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__A2_N
timestamp 1607194113
transform 1 0 49772 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0832_
timestamp 1607194113
transform 1 0 48300 0 1 40800
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_71_550
timestamp 1607194113
transform 1 0 51704 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_71_545
timestamp 1607194113
transform 1 0 51244 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_533
timestamp 1607194113
transform 1 0 50140 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__B2
timestamp 1607194113
transform 1 0 49956 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_620
timestamp 1607194113
transform 1 0 51612 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_563
timestamp 1607194113
transform 1 0 52900 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_558
timestamp 1607194113
transform 1 0 52440 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0771_
timestamp 1607194113
transform 1 0 52624 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_71_575
timestamp 1607194113
transform 1 0 54004 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1481__CLK
timestamp 1607194113
transform 1 0 54556 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1481_
timestamp 1607194113
transform 1 0 54740 0 1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_71_611
timestamp 1607194113
transform 1 0 57316 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_602
timestamp 1607194113
transform 1 0 56488 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_621
timestamp 1607194113
transform 1 0 57224 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_623
timestamp 1607194113
transform 1 0 58420 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_647
timestamp 1607194113
transform 1 0 60628 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_635
timestamp 1607194113
transform 1 0 59524 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_672
timestamp 1607194113
transform 1 0 62928 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_659
timestamp 1607194113
transform 1 0 61732 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_622
timestamp 1607194113
transform 1 0 62836 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_683
timestamp 1607194113
transform 1 0 63940 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1076_
timestamp 1607194113
transform 1 0 63664 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1068_
timestamp 1607194113
transform 1 0 64676 0 1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_71_713
timestamp 1607194113
transform 1 0 66700 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_698
timestamp 1607194113
transform 1 0 65320 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1069_
timestamp 1607194113
transform 1 0 66056 0 1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_71_731
timestamp 1607194113
transform 1 0 68356 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_725
timestamp 1607194113
transform 1 0 67804 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_623
timestamp 1607194113
transform 1 0 68448 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_498
timestamp 1607194113
transform 1 0 46920 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__or4_4  _0775_
timestamp 1607194113
transform 1 0 46092 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_72_518
timestamp 1607194113
transform 1 0 48760 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_510
timestamp 1607194113
transform 1 0 48024 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__B1
timestamp 1607194113
transform 1 0 48576 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A1_N
timestamp 1607194113
transform 1 0 48392 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_638
timestamp 1607194113
transform 1 0 48852 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0849_
timestamp 1607194113
transform 1 0 48944 0 -1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_72_550
timestamp 1607194113
transform 1 0 51704 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_538
timestamp 1607194113
transform 1 0 50600 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__B2
timestamp 1607194113
transform 1 0 50416 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_72_562
timestamp 1607194113
transform 1 0 52808 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1055_
timestamp 1607194113
transform 1 0 53084 0 -1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_72_581
timestamp 1607194113
transform 1 0 54556 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_72_572
timestamp 1607194113
transform 1 0 53728 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_639
timestamp 1607194113
transform 1 0 54464 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1056_
timestamp 1607194113
transform 1 0 54924 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_72_608
timestamp 1607194113
transform 1 0 57040 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_596
timestamp 1607194113
transform 1 0 55936 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A
timestamp 1607194113
transform 1 0 55752 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_631
timestamp 1607194113
transform 1 0 59156 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_72_620
timestamp 1607194113
transform 1 0 58144 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__A
timestamp 1607194113
transform 1 0 58696 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1607194113
transform 1 0 58880 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_647
timestamp 1607194113
transform 1 0 60628 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_639
timestamp 1607194113
transform 1 0 59892 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__A
timestamp 1607194113
transform 1 0 60444 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_640
timestamp 1607194113
transform 1 0 60076 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1607194113
transform 1 0 60168 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_72_675
timestamp 1607194113
transform 1 0 63204 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_671
timestamp 1607194113
transform 1 0 62836 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_659
timestamp 1607194113
transform 1 0 61732 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_694
timestamp 1607194113
transform 1 0 64952 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_72_681
timestamp 1607194113
transform 1 0 63756 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A
timestamp 1607194113
transform 1 0 63572 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1032_
timestamp 1607194113
transform 1 0 64308 0 -1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1031_
timestamp 1607194113
transform 1 0 63296 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_712
timestamp 1607194113
transform 1 0 66608 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__A
timestamp 1607194113
transform 1 0 65504 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_641
timestamp 1607194113
transform 1 0 65688 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1050_
timestamp 1607194113
transform 1 0 65780 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_72_724
timestamp 1607194113
transform 1 0 67712 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_501
timestamp 1607194113
transform 1 0 47196 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_489
timestamp 1607194113
transform 1 0 46092 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__B1
timestamp 1607194113
transform 1 0 47564 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__A1_N
timestamp 1607194113
transform 1 0 47748 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0845_
timestamp 1607194113
transform 1 0 47932 0 1 41888
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_12  FILLER_73_529
timestamp 1607194113
transform 1 0 49772 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__A2_N
timestamp 1607194113
transform 1 0 49588 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__B2
timestamp 1607194113
transform 1 0 49404 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_541
timestamp 1607194113
transform 1 0 50876 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_657
timestamp 1607194113
transform 1 0 51612 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0696_
timestamp 1607194113
transform 1 0 51704 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_565
timestamp 1607194113
transform 1 0 53084 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_553
timestamp 1607194113
transform 1 0 51980 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__A1
timestamp 1607194113
transform 1 0 53452 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1059_
timestamp 1607194113
transform 1 0 53636 0 1 41888
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_73_587
timestamp 1607194113
transform 1 0 55108 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__B1
timestamp 1607194113
transform 1 0 54924 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_611
timestamp 1607194113
transform 1 0 57316 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_608
timestamp 1607194113
transform 1 0 57040 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_596
timestamp 1607194113
transform 1 0 55936 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_658
timestamp 1607194113
transform 1 0 57224 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1053_
timestamp 1607194113
transform 1 0 55660 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_73_623
timestamp 1607194113
transform 1 0 58420 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_4  _1066_
timestamp 1607194113
transform 1 0 58972 0 1 41888
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_73_645
timestamp 1607194113
transform 1 0 60444 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__B1
timestamp 1607194113
transform 1 0 60260 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1064_
timestamp 1607194113
transform 1 0 60996 0 1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_73_672
timestamp 1607194113
transform 1 0 62928 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_670
timestamp 1607194113
transform 1 0 62744 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_658
timestamp 1607194113
transform 1 0 61640 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_659
timestamp 1607194113
transform 1 0 62836 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_680
timestamp 1607194113
transform 1 0 63664 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__B1
timestamp 1607194113
transform 1 0 65136 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1079_
timestamp 1607194113
transform 1 0 63848 0 1 41888
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_73_717
timestamp 1607194113
transform 1 0 67068 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_710
timestamp 1607194113
transform 1 0 66424 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_698
timestamp 1607194113
transform 1 0 65320 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A
timestamp 1607194113
transform 1 0 66884 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1030_
timestamp 1607194113
transform 1 0 66608 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_73_729
timestamp 1607194113
transform 1 0 68172 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_660
timestamp 1607194113
transform 1 0 68448 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_75_509
timestamp 1607194113
transform 1 0 47932 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_75_501
timestamp 1607194113
transform 1 0 47196 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_489
timestamp 1607194113
transform 1 0 46092 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_507
timestamp 1607194113
transform 1 0 47748 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_495
timestamp 1607194113
transform 1 0 46644 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A2_N
timestamp 1607194113
transform 1 0 46460 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__B2
timestamp 1607194113
transform 1 0 46276 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_520
timestamp 1607194113
transform 1 0 48944 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__A1_N
timestamp 1607194113
transform 1 0 48208 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__B1
timestamp 1607194113
transform 1 0 48392 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_675
timestamp 1607194113
transform 1 0 48852 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0843_
timestamp 1607194113
transform 1 0 48576 0 1 42976
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_75_550
timestamp 1607194113
transform 1 0 51704 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_75_546
timestamp 1607194113
transform 1 0 51336 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_534
timestamp 1607194113
transform 1 0 50232 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_532
timestamp 1607194113
transform 1 0 50048 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1480__CLK
timestamp 1607194113
transform 1 0 50784 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__A2_N
timestamp 1607194113
transform 1 0 50048 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_694
timestamp 1607194113
transform 1 0 51612 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1480_
timestamp 1607194113
transform 1 0 50968 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_75_558
timestamp 1607194113
transform 1 0 52440 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_554
timestamp 1607194113
transform 1 0 52072 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_561
timestamp 1607194113
transform 1 0 52716 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1479_
timestamp 1607194113
transform 1 0 53176 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1060_
timestamp 1607194113
transform 1 0 53452 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0664_
timestamp 1607194113
transform 1 0 52164 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_587
timestamp 1607194113
transform 1 0 55108 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_590
timestamp 1607194113
transform 1 0 55384 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_572
timestamp 1607194113
transform 1 0 53728 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1479__CLK
timestamp 1607194113
transform 1 0 54924 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A
timestamp 1607194113
transform 1 0 55200 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_676
timestamp 1607194113
transform 1 0 54464 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1052_
timestamp 1607194113
transform 1 0 54556 0 -1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_75_611
timestamp 1607194113
transform 1 0 57316 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_607
timestamp 1607194113
transform 1 0 56948 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_75_599
timestamp 1607194113
transform 1 0 56212 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_606
timestamp 1607194113
transform 1 0 56856 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_602
timestamp 1607194113
transform 1 0 56488 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__A
timestamp 1607194113
transform 1 0 56948 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_695
timestamp 1607194113
transform 1 0 57224 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1063_
timestamp 1607194113
transform 1 0 57132 0 -1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_75_623
timestamp 1607194113
transform 1 0 58420 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_633
timestamp 1607194113
transform 1 0 59340 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_74_616
timestamp 1607194113
transform 1 0 57776 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1478__CLK
timestamp 1607194113
transform 1 0 58604 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1478_
timestamp 1607194113
transform 1 0 58788 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__or3_4  _1051_
timestamp 1607194113
transform 1 0 58512 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_75_646
timestamp 1607194113
transform 1 0 60536 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_653
timestamp 1607194113
transform 1 0 61180 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__A
timestamp 1607194113
transform 1 0 60996 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_677
timestamp 1607194113
transform 1 0 60076 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1065_
timestamp 1607194113
transform 1 0 60168 0 -1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_75_672
timestamp 1607194113
transform 1 0 62928 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_670
timestamp 1607194113
transform 1 0 62744 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_658
timestamp 1607194113
transform 1 0 61640 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_670
timestamp 1607194113
transform 1 0 62744 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_662
timestamp 1607194113
transform 1 0 62008 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1474__CLK
timestamp 1607194113
transform 1 0 62928 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_696
timestamp 1607194113
transform 1 0 62836 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1474_
timestamp 1607194113
transform 1 0 63112 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1062_
timestamp 1607194113
transform 1 0 61732 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_695
timestamp 1607194113
transform 1 0 65044 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_683
timestamp 1607194113
transform 1 0 63940 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_693
timestamp 1607194113
transform 1 0 64860 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1080_
timestamp 1607194113
transform 1 0 63664 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_707
timestamp 1607194113
transform 1 0 66148 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_703
timestamp 1607194113
transform 1 0 65780 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_74_699
timestamp 1607194113
transform 1 0 65412 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1477__CLK
timestamp 1607194113
transform 1 0 65504 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_678
timestamp 1607194113
transform 1 0 65688 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1477_
timestamp 1607194113
transform 1 0 65872 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1073_
timestamp 1607194113
transform 1 0 66332 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_75_729
timestamp 1607194113
transform 1 0 68172 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_75_721
timestamp 1607194113
transform 1 0 67436 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_74_723
timestamp 1607194113
transform 1 0 67620 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_697
timestamp 1607194113
transform 1 0 68448 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1072_
timestamp 1607194113
transform 1 0 68356 0 -1 42976
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_76_509
timestamp 1607194113
transform 1 0 47932 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_497
timestamp 1607194113
transform 1 0 46828 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_495
timestamp 1607194113
transform 1 0 46644 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_489
timestamp 1607194113
transform 1 0 46092 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_719
timestamp 1607194113
transform 1 0 46736 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_528
timestamp 1607194113
transform 1 0 49680 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_521
timestamp 1607194113
transform 1 0 49036 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_720
timestamp 1607194113
transform 1 0 49588 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_540
timestamp 1607194113
transform 1 0 50784 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_559
timestamp 1607194113
transform 1 0 52532 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_552
timestamp 1607194113
transform 1 0 51888 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_721
timestamp 1607194113
transform 1 0 52440 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0766_
timestamp 1607194113
transform 1 0 53636 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_590
timestamp 1607194113
transform 1 0 55384 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_587
timestamp 1607194113
transform 1 0 55108 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_575
timestamp 1607194113
transform 1 0 54004 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_722
timestamp 1607194113
transform 1 0 55292 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_602
timestamp 1607194113
transform 1 0 56488 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_627
timestamp 1607194113
transform 1 0 58788 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_621
timestamp 1607194113
transform 1 0 58236 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_76_614
timestamp 1607194113
transform 1 0 57592 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_723
timestamp 1607194113
transform 1 0 58144 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1067_
timestamp 1607194113
transform 1 0 58512 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_652
timestamp 1607194113
transform 1 0 61088 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_650
timestamp 1607194113
transform 1 0 60904 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_642
timestamp 1607194113
transform 1 0 60168 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_724
timestamp 1607194113
transform 1 0 60996 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1061_
timestamp 1607194113
transform 1 0 59524 0 -1 44064
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_76_664
timestamp 1607194113
transform 1 0 62192 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_695
timestamp 1607194113
transform 1 0 65044 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_683
timestamp 1607194113
transform 1 0 63940 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_676
timestamp 1607194113
transform 1 0 63296 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_725
timestamp 1607194113
transform 1 0 63848 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_714
timestamp 1607194113
transform 1 0 66792 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_707
timestamp 1607194113
transform 1 0 66148 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_726
timestamp 1607194113
transform 1 0 66700 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_726
timestamp 1607194113
transform 1 0 67896 0 -1 44064
box -38 -48 1142 592
use delayline_9_ms  inst_idelay_line
timestamp 1607276512
transform 1 0 53176 0 1 3761
box 800 801 23264 27367
use sky130_fd_sc_hd__decap_12  FILLER_59_745
timestamp 1607194113
transform 1 0 69644 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_733
timestamp 1607194113
transform 1 0 68540 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_769
timestamp 1607194113
transform 1 0 71852 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_757
timestamp 1607194113
transform 1 0 70748 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_781
timestamp 1607194113
transform 1 0 72956 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_806
timestamp 1607194113
transform 1 0 75256 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_794
timestamp 1607194113
transform 1 0 74152 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1607194113
transform 1 0 74060 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1451__CLK
timestamp 1607194113
transform 1 0 75992 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1451_
timestamp 1607194113
transform 1 0 76176 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_59_848
timestamp 1607194113
transform 1 0 79120 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_59_835
timestamp 1607194113
transform 1 0 77924 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A
timestamp 1607194113
transform 1 0 78936 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0761_
timestamp 1607194113
transform 1 0 78660 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_866
timestamp 1607194113
transform 1 0 80776 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_858
timestamp 1607194113
transform 1 0 80040 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[7]
timestamp 1607194113
transform 1 0 80960 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[5]
timestamp 1607194113
transform 1 0 81144 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1607194113
transform 1 0 79672 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1044_
timestamp 1607194113
transform 1 0 79764 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1454__CLK
timestamp 1607194113
transform 1 0 82524 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[3]
timestamp 1607194113
transform 1 0 81328 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[2]
timestamp 1607194113
transform 1 0 81512 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[1]
timestamp 1607194113
transform 1 0 82340 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[0]
timestamp 1607194113
transform 1 0 82156 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_inp_i
timestamp 1607194113
transform 1 0 81972 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1454_
timestamp 1607194113
transform 1 0 82708 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _1148_
timestamp 1607194113
transform 1 0 81696 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_59_906
timestamp 1607194113
transform 1 0 84456 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_59_922
timestamp 1607194113
transform 1 0 85928 0 1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_914
timestamp 1607194113
transform 1 0 85192 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__A
timestamp 1607194113
transform 1 0 85744 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1607194113
transform 1 0 85284 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0738_
timestamp 1607194113
transform 1 0 85376 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0737_
timestamp 1607194113
transform 1 0 86480 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_949
timestamp 1607194113
transform 1 0 88412 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_943
timestamp 1607194113
transform 1 0 87860 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_931
timestamp 1607194113
transform 1 0 86756 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A
timestamp 1607194113
transform 1 0 88228 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0782_
timestamp 1607194113
transform 1 0 87952 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_59_962
timestamp 1607194113
transform 1 0 89608 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__B
timestamp 1607194113
transform 1 0 88780 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1043_
timestamp 1607194113
transform 1 0 88964 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_59_974
timestamp 1607194113
transform 1 0 90712 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1607194113
transform 1 0 90896 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_734
timestamp 1607194113
transform 1 0 68632 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1379_
timestamp 1607194113
transform 1 0 68816 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_60_764
timestamp 1607194113
transform 1 0 71392 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_757
timestamp 1607194113
transform 1 0 70748 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1379__CLK
timestamp 1607194113
transform 1 0 70564 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1607194113
transform 1 0 71300 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_776
timestamp 1607194113
transform 1 0 72496 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1450_
timestamp 1607194113
transform 1 0 72864 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_60_801
timestamp 1607194113
transform 1 0 74796 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1450__CLK
timestamp 1607194113
transform 1 0 74612 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__A
timestamp 1607194113
transform 1 0 75164 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1155_
timestamp 1607194113
transform 1 0 75348 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_60_829
timestamp 1607194113
transform 1 0 77372 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_816
timestamp 1607194113
transform 1 0 76176 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__B
timestamp 1607194113
transform 1 0 75992 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1607194113
transform 1 0 76912 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0700_
timestamp 1607194113
transform 1 0 77004 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_835
timestamp 1607194113
transform 1 0 77924 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1452__CLK
timestamp 1607194113
transform 1 0 78016 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1452_
timestamp 1607194113
transform 1 0 78200 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_60_869
timestamp 1607194113
transform 1 0 81052 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_857
timestamp 1607194113
transform 1 0 79948 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_886
timestamp 1607194113
transform 1 0 82616 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_60_883
timestamp 1607194113
transform 1 0 82340 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[8]
timestamp 1607194113
transform 1 0 82156 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[6]
timestamp 1607194113
transform 1 0 81972 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_inst_rdelay_line_en_i[4]
timestamp 1607194113
transform 1 0 81788 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1607194113
transform 1 0 82524 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_910
timestamp 1607194113
transform 1 0 84824 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__B1
timestamp 1607194113
transform 1 0 83168 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__A1
timestamp 1607194113
transform 1 0 84640 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1147_
timestamp 1607194113
transform 1 0 83352 0 -1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_60_925
timestamp 1607194113
transform 1 0 86204 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__A
timestamp 1607194113
transform 1 0 86020 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1137_
timestamp 1607194113
transform 1 0 85376 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_60_950
timestamp 1607194113
transform 1 0 88504 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_945
timestamp 1607194113
transform 1 0 88044 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_937
timestamp 1607194113
transform 1 0 87308 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1607194113
transform 1 0 88136 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1144_
timestamp 1607194113
transform 1 0 88228 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1456__CLK
timestamp 1607194113
transform 1 0 89056 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1456_
timestamp 1607194113
transform 1 0 89240 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_62_750
timestamp 1607194113
transform 1 0 70104 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_739
timestamp 1607194113
transform 1 0 69092 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_733
timestamp 1607194113
transform 1 0 68540 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1420_
timestamp 1607194113
transform 1 0 68816 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0689_
timestamp 1607194113
transform 1 0 69828 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_767
timestamp 1607194113
transform 1 0 71668 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_762
timestamp 1607194113
transform 1 0 71208 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_766
timestamp 1607194113
transform 1 0 71576 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_757
timestamp 1607194113
transform 1 0 70748 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1420__CLK
timestamp 1607194113
transform 1 0 70564 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1607194113
transform 1 0 71300 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0793_
timestamp 1607194113
transform 1 0 71392 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0692_
timestamp 1607194113
transform 1 0 71300 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_792
timestamp 1607194113
transform 1 0 73968 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_779
timestamp 1607194113
transform 1 0 72772 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_790
timestamp 1607194113
transform 1 0 73784 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_778
timestamp 1607194113
transform 1 0 72680 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__A
timestamp 1607194113
transform 1 0 73784 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__B
timestamp 1607194113
transform 1 0 73600 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _1157_
timestamp 1607194113
transform 1 0 72956 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_62_804
timestamp 1607194113
transform 1 0 75072 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_811
timestamp 1607194113
transform 1 0 75716 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_799
timestamp 1607194113
transform 1 0 74612 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__A
timestamp 1607194113
transform 1 0 74428 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1607194113
transform 1 0 74060 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0705_
timestamp 1607194113
transform 1 0 74152 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_825
timestamp 1607194113
transform 1 0 77004 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_62_816
timestamp 1607194113
transform 1 0 76176 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_61_825
timestamp 1607194113
transform 1 0 77004 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_815
timestamp 1607194113
transform 1 0 76084 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__A
timestamp 1607194113
transform 1 0 77556 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1607194113
transform 1 0 76912 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1156_
timestamp 1607194113
transform 1 0 76176 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1153_
timestamp 1607194113
transform 1 0 77556 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_62_842
timestamp 1607194113
transform 1 0 78568 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_61_844
timestamp 1607194113
transform 1 0 78752 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__C
timestamp 1607194113
transform 1 0 78568 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__A
timestamp 1607194113
transform 1 0 78384 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1154_
timestamp 1607194113
transform 1 0 79120 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _1046_
timestamp 1607194113
transform 1 0 77740 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_62_869
timestamp 1607194113
transform 1 0 81052 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_857
timestamp 1607194113
transform 1 0 79948 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_864
timestamp 1607194113
transform 1 0 80592 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_852
timestamp 1607194113
transform 1 0 79488 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__A
timestamp 1607194113
transform 1 0 80408 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1607194113
transform 1 0 79672 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1149_
timestamp 1607194113
transform 1 0 79764 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_62_886
timestamp 1607194113
transform 1 0 82616 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_881
timestamp 1607194113
transform 1 0 82156 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_888
timestamp 1607194113
transform 1 0 82800 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_876
timestamp 1607194113
transform 1 0 81696 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1607194113
transform 1 0 82524 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_898
timestamp 1607194113
transform 1 0 83720 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_61_904
timestamp 1607194113
transform 1 0 84272 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_896
timestamp 1607194113
transform 1 0 83536 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1457__CLK
timestamp 1607194113
transform 1 0 83996 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__A
timestamp 1607194113
transform 1 0 84088 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1457_
timestamp 1607194113
transform 1 0 84180 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_2  _0734_
timestamp 1607194113
transform 1 0 83720 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_922
timestamp 1607194113
transform 1 0 85928 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_929
timestamp 1607194113
transform 1 0 86572 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_912
timestamp 1607194113
transform 1 0 85008 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A
timestamp 1607194113
transform 1 0 86388 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__B
timestamp 1607194113
transform 1 0 86204 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1607194113
transform 1 0 85284 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1047_
timestamp 1607194113
transform 1 0 85376 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0733_
timestamp 1607194113
transform 1 0 86664 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_62_947
timestamp 1607194113
transform 1 0 88228 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_945
timestamp 1607194113
transform 1 0 88044 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_933
timestamp 1607194113
transform 1 0 86940 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_941
timestamp 1607194113
transform 1 0 87676 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1607194113
transform 1 0 88136 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1138_
timestamp 1607194113
transform 1 0 87952 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_62_964
timestamp 1607194113
transform 1 0 89792 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_61_968
timestamp 1607194113
transform 1 0 90160 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_951
timestamp 1607194113
transform 1 0 88596 0 1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__A
timestamp 1607194113
transform 1 0 88780 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__A
timestamp 1607194113
transform 1 0 89148 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1143_
timestamp 1607194113
transform 1 0 88964 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1142_
timestamp 1607194113
transform 1 0 89332 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_62_975
timestamp 1607194113
transform 1 0 90804 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__A
timestamp 1607194113
transform 1 0 90712 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1607194113
transform 1 0 90896 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1042_
timestamp 1607194113
transform 1 0 90528 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_744
timestamp 1607194113
transform 1 0 69552 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_63_733
timestamp 1607194113
transform 1 0 68540 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _0791_
timestamp 1607194113
transform 1 0 69276 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _0694_
timestamp 1607194113
transform 1 0 70288 0 1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_63_770
timestamp 1607194113
transform 1 0 71944 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__A2
timestamp 1607194113
transform 1 0 71760 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__B2
timestamp 1607194113
transform 1 0 71576 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_790
timestamp 1607194113
transform 1 0 73784 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_782
timestamp 1607194113
transform 1 0 73048 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_806
timestamp 1607194113
transform 1 0 75256 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_794
timestamp 1607194113
transform 1 0 74152 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1607194113
transform 1 0 74060 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_818
timestamp 1607194113
transform 1 0 76360 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _1152_
timestamp 1607194113
transform 1 0 76728 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_845
timestamp 1607194113
transform 1 0 78844 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_63_834
timestamp 1607194113
transform 1 0 77832 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__A
timestamp 1607194113
transform 1 0 78384 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1045_
timestamp 1607194113
transform 1 0 78568 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_864
timestamp 1607194113
transform 1 0 80592 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_853
timestamp 1607194113
transform 1 0 79580 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__A
timestamp 1607194113
transform 1 0 80408 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1607194113
transform 1 0 79672 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1150_
timestamp 1607194113
transform 1 0 79764 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_63_890
timestamp 1607194113
transform 1 0 82984 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_878
timestamp 1607194113
transform 1 0 81880 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_872
timestamp 1607194113
transform 1 0 81328 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _1117_
timestamp 1607194113
transform 1 0 81512 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_902
timestamp 1607194113
transform 1 0 84088 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__A1
timestamp 1607194113
transform 1 0 84824 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_929
timestamp 1607194113
transform 1 0 86572 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_914
timestamp 1607194113
transform 1 0 85192 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__B1
timestamp 1607194113
transform 1 0 85008 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1607194113
transform 1 0 85284 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1139_
timestamp 1607194113
transform 1 0 85376 0 1 36448
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_63_941
timestamp 1607194113
transform 1 0 87676 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_970
timestamp 1607194113
transform 1 0 90344 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_953
timestamp 1607194113
transform 1 0 88780 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__A
timestamp 1607194113
transform 1 0 90160 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1145_
timestamp 1607194113
transform 1 0 89516 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1607194113
transform 1 0 90896 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_739
timestamp 1607194113
transform 1 0 69092 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0792_
timestamp 1607194113
transform 1 0 69276 0 -1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_64_759
timestamp 1607194113
transform 1 0 70932 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__A2
timestamp 1607194113
transform 1 0 70748 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__B2
timestamp 1607194113
transform 1 0 70564 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1607194113
transform 1 0 71300 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0794_
timestamp 1607194113
transform 1 0 71392 0 -1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_64_782
timestamp 1607194113
transform 1 0 73048 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__A2
timestamp 1607194113
transform 1 0 72864 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__B2
timestamp 1607194113
transform 1 0 72680 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_809
timestamp 1607194113
transform 1 0 75532 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_802
timestamp 1607194113
transform 1 0 74888 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_794
timestamp 1607194113
transform 1 0 74152 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1027_
timestamp 1607194113
transform 1 0 75164 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_821
timestamp 1607194113
transform 1 0 76636 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1453__CLK
timestamp 1607194113
transform 1 0 76728 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1607194113
transform 1 0 76912 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1453_
timestamp 1607194113
transform 1 0 77004 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_64_844
timestamp 1607194113
transform 1 0 78752 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_868
timestamp 1607194113
transform 1 0 80960 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_856
timestamp 1607194113
transform 1 0 79856 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_886
timestamp 1607194113
transform 1 0 82616 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_884
timestamp 1607194113
transform 1 0 82432 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_880
timestamp 1607194113
transform 1 0 82064 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__A
timestamp 1607194113
transform 1 0 82708 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1607194113
transform 1 0 82524 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1114_
timestamp 1607194113
transform 1 0 82892 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_64_896
timestamp 1607194113
transform 1 0 83536 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__A1
timestamp 1607194113
transform 1 0 84272 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1140_
timestamp 1607194113
transform 1 0 84456 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_930
timestamp 1607194113
transform 1 0 86664 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_918
timestamp 1607194113
transform 1 0 85560 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_947
timestamp 1607194113
transform 1 0 88228 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_942
timestamp 1607194113
transform 1 0 87768 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1607194113
transform 1 0 88136 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_959
timestamp 1607194113
transform 1 0 89332 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__A
timestamp 1607194113
transform 1 0 90252 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _1108_
timestamp 1607194113
transform 1 0 89424 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_64_971
timestamp 1607194113
transform 1 0 90436 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_65_743
timestamp 1607194113
transform 1 0 69460 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_733
timestamp 1607194113
transform 1 0 68540 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _0695_
timestamp 1607194113
transform 1 0 68632 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_4  _0691_
timestamp 1607194113
transform 1 0 70196 0 1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_65_769
timestamp 1607194113
transform 1 0 71852 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__A2
timestamp 1607194113
transform 1 0 71668 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__B2
timestamp 1607194113
transform 1 0 71484 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_65_790
timestamp 1607194113
transform 1 0 73784 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_782
timestamp 1607194113
transform 1 0 73048 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0795_
timestamp 1607194113
transform 1 0 72220 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_65_806
timestamp 1607194113
transform 1 0 75256 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_794
timestamp 1607194113
transform 1 0 74152 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1607194113
transform 1 0 74060 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_818
timestamp 1607194113
transform 1 0 76360 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__B1
timestamp 1607194113
transform 1 0 76636 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _1151_
timestamp 1607194113
transform 1 0 76820 0 1 37536
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_65_848
timestamp 1607194113
transform 1 0 79120 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_65_836
timestamp 1607194113
transform 1 0 78016 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_867
timestamp 1607194113
transform 1 0 80868 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_855
timestamp 1607194113
transform 1 0 79764 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1463__CLK
timestamp 1607194113
transform 1 0 81144 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1607194113
transform 1 0 79672 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_891
timestamp 1607194113
transform 1 0 83076 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _1463_
timestamp 1607194113
transform 1 0 81328 0 1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_65_906
timestamp 1607194113
transform 1 0 84456 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__A
timestamp 1607194113
transform 1 0 83628 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1119_
timestamp 1607194113
transform 1 0 83812 0 1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_65_923
timestamp 1607194113
transform 1 0 86020 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_65_916
timestamp 1607194113
transform 1 0 85376 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_65_914
timestamp 1607194113
transform 1 0 85192 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1607194113
transform 1 0 85284 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0744_
timestamp 1607194113
transform 1 0 85652 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_947
timestamp 1607194113
transform 1 0 88228 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_935
timestamp 1607194113
transform 1 0 87124 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_970
timestamp 1607194113
transform 1 0 90344 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_65_955
timestamp 1607194113
transform 1 0 88964 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__A
timestamp 1607194113
transform 1 0 89148 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__B
timestamp 1607194113
transform 1 0 90160 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _1109_
timestamp 1607194113
transform 1 0 89332 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1607194113
transform 1 0 90896 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_742
timestamp 1607194113
transform 1 0 69368 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__A
timestamp 1607194113
transform 1 0 70104 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _0686_
timestamp 1607194113
transform 1 0 70288 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_66_762
timestamp 1607194113
transform 1 0 71208 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_66_755
timestamp 1607194113
transform 1 0 70564 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__A1
timestamp 1607194113
transform 1 0 71024 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__B1
timestamp 1607194113
transform 1 0 70840 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1607194113
transform 1 0 71300 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0688_
timestamp 1607194113
transform 1 0 71392 0 -1 38624
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_66_790
timestamp 1607194113
transform 1 0 73784 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_778
timestamp 1607194113
transform 1 0 72680 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_809
timestamp 1607194113
transform 1 0 75532 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_797
timestamp 1607194113
transform 1 0 74428 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_clk_i
timestamp 1607194113
transform 1 0 74152 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_825
timestamp 1607194113
transform 1 0 77004 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_66_821
timestamp 1607194113
transform 1 0 76636 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1607194113
transform 1 0 76912 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0745_
timestamp 1607194113
transform 1 0 77372 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_846
timestamp 1607194113
transform 1 0 78936 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_834
timestamp 1607194113
transform 1 0 77832 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__A
timestamp 1607194113
transform 1 0 77648 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_870
timestamp 1607194113
transform 1 0 81144 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_858
timestamp 1607194113
transform 1 0 80040 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_879
timestamp 1607194113
transform 1 0 81972 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A
timestamp 1607194113
transform 1 0 81788 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__A
timestamp 1607194113
transform 1 0 82340 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1607194113
transform 1 0 82524 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1120_
timestamp 1607194113
transform 1 0 82616 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0690_
timestamp 1607194113
transform 1 0 81512 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_907
timestamp 1607194113
transform 1 0 84548 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_895
timestamp 1607194113
transform 1 0 83444 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__B
timestamp 1607194113
transform 1 0 84732 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A
timestamp 1607194113
transform 1 0 84916 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_924
timestamp 1607194113
transform 1 0 86112 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__D
timestamp 1607194113
transform 1 0 85928 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1041_
timestamp 1607194113
transform 1 0 85100 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_66_947
timestamp 1607194113
transform 1 0 88228 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_944
timestamp 1607194113
transform 1 0 87952 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_936
timestamp 1607194113
transform 1 0 87216 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1607194113
transform 1 0 88136 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1040_
timestamp 1607194113
transform 1 0 88412 0 -1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_66_964
timestamp 1607194113
transform 1 0 89792 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__B1
timestamp 1607194113
transform 1 0 90068 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__A1
timestamp 1607194113
transform 1 0 90252 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__A
timestamp 1607194113
transform 1 0 89608 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__C
timestamp 1607194113
transform 1 0 89424 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__D
timestamp 1607194113
transform 1 0 89240 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1128_
timestamp 1607194113
transform 1 0 90436 0 -1 38624
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_68_748
timestamp 1607194113
transform 1 0 69920 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_736
timestamp 1607194113
transform 1 0 68816 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_748
timestamp 1607194113
transform 1 0 69920 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_733
timestamp 1607194113
transform 1 0 68540 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0789_
timestamp 1607194113
transform 1 0 69644 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_768
timestamp 1607194113
transform 1 0 71760 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_764
timestamp 1607194113
transform 1 0 71392 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_760
timestamp 1607194113
transform 1 0 71024 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_67_770
timestamp 1607194113
transform 1 0 71944 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__B1
timestamp 1607194113
transform 1 0 70472 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1607194113
transform 1 0 71300 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1094_
timestamp 1607194113
transform 1 0 71484 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _0790_
timestamp 1607194113
transform 1 0 70656 0 1 38624
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_68_779
timestamp 1607194113
transform 1 0 72772 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_781
timestamp 1607194113
transform 1 0 72956 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_clk_i_A
timestamp 1607194113
transform 1 0 72496 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_clk_i
timestamp 1607194113
transform 1 0 72680 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1471_
timestamp 1607194113
transform 1 0 73508 0 -1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__inv_2  _0687_
timestamp 1607194113
transform 1 0 72496 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_808
timestamp 1607194113
transform 1 0 75440 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_801
timestamp 1607194113
transform 1 0 74796 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1471__CLK
timestamp 1607194113
transform 1 0 75256 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1607194113
transform 1 0 74060 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1091_
timestamp 1607194113
transform 1 0 74152 0 1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_68_825
timestamp 1607194113
transform 1 0 77004 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_820
timestamp 1607194113
transform 1 0 76544 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_821
timestamp 1607194113
transform 1 0 76636 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_813
timestamp 1607194113
transform 1 0 75900 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1466__CLK
timestamp 1607194113
transform 1 0 77188 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1464__CLK
timestamp 1607194113
transform 1 0 76820 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1607194113
transform 1 0 76912 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1466_
timestamp 1607194113
transform 1 0 77372 0 -1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1464_
timestamp 1607194113
transform 1 0 77004 0 1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_68_848
timestamp 1607194113
transform 1 0 79120 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_67_844
timestamp 1607194113
transform 1 0 78752 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_68_859
timestamp 1607194113
transform 1 0 80132 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_867
timestamp 1607194113
transform 1 0 80868 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_855
timestamp 1607194113
transform 1 0 79764 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_852
timestamp 1607194113
transform 1 0 79488 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1607194113
transform 1 0 79672 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1107_
timestamp 1607194113
transform 1 0 79856 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1102_
timestamp 1607194113
transform 1 0 81236 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_68_890
timestamp 1607194113
transform 1 0 82984 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_886
timestamp 1607194113
transform 1 0 82616 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_882
timestamp 1607194113
transform 1 0 82248 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_874
timestamp 1607194113
transform 1 0 81512 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_890
timestamp 1607194113
transform 1 0 82984 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__A
timestamp 1607194113
transform 1 0 81972 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1607194113
transform 1 0 82524 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1118_
timestamp 1607194113
transform 1 0 82708 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _1115_
timestamp 1607194113
transform 1 0 82156 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_67_909
timestamp 1607194113
transform 1 0 84732 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__B1
timestamp 1607194113
transform 1 0 83536 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__B
timestamp 1607194113
transform 1 0 83352 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__C
timestamp 1607194113
transform 1 0 84548 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__A
timestamp 1607194113
transform 1 0 83536 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1121_
timestamp 1607194113
transform 1 0 83720 0 -1 39712
box -38 -48 1326 592
use sky130_fd_sc_hd__or4_4  _1110_
timestamp 1607194113
transform 1 0 83720 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_68_926
timestamp 1607194113
transform 1 0 86296 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_68_914
timestamp 1607194113
transform 1 0 85192 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_67_925
timestamp 1607194113
transform 1 0 86204 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__A
timestamp 1607194113
transform 1 0 86020 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__A1
timestamp 1607194113
transform 1 0 85008 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__A
timestamp 1607194113
transform 1 0 86112 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1607194113
transform 1 0 85284 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1113_
timestamp 1607194113
transform 1 0 85376 0 1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0709_
timestamp 1607194113
transform 1 0 85744 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_947
timestamp 1607194113
transform 1 0 88228 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_945
timestamp 1607194113
transform 1 0 88044 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_937
timestamp 1607194113
transform 1 0 87308 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_941
timestamp 1607194113
transform 1 0 87676 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_931
timestamp 1607194113
transform 1 0 86756 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__A
timestamp 1607194113
transform 1 0 87124 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1607194113
transform 1 0 88136 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1048_
timestamp 1607194113
transform 1 0 86848 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0743_
timestamp 1607194113
transform 1 0 86848 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_968
timestamp 1607194113
transform 1 0 90160 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_963
timestamp 1607194113
transform 1 0 89700 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_955
timestamp 1607194113
transform 1 0 88964 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_951
timestamp 1607194113
transform 1 0 88596 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_965
timestamp 1607194113
transform 1 0 89884 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_953
timestamp 1607194113
transform 1 0 88780 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1122_
timestamp 1607194113
transform 1 0 88688 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0713_
timestamp 1607194113
transform 1 0 89884 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_68_976
timestamp 1607194113
transform 1 0 90896 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_973
timestamp 1607194113
transform 1 0 90620 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1607194113
transform 1 0 90896 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_745
timestamp 1607194113
transform 1 0 69644 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_733
timestamp 1607194113
transform 1 0 68540 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_753
timestamp 1607194113
transform 1 0 70380 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1470__CLK
timestamp 1607194113
transform 1 0 70564 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1470_
timestamp 1607194113
transform 1 0 70748 0 1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_69_788
timestamp 1607194113
transform 1 0 73600 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_776
timestamp 1607194113
transform 1 0 72496 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_clk_i
timestamp 1607194113
transform 1 0 73784 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_803
timestamp 1607194113
transform 1 0 74980 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1607194113
transform 1 0 74060 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1092_
timestamp 1607194113
transform 1 0 74152 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_69_827
timestamp 1607194113
transform 1 0 77188 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_815
timestamp 1607194113
transform 1 0 76084 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0757_
timestamp 1607194113
transform 1 0 77464 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_847
timestamp 1607194113
transform 1 0 79028 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_835
timestamp 1607194113
transform 1 0 77924 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__A
timestamp 1607194113
transform 1 0 77740 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__B1
timestamp 1607194113
transform 1 0 79396 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__A1
timestamp 1607194113
transform 1 0 79212 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_871
timestamp 1607194113
transform 1 0 81236 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_853
timestamp 1607194113
transform 1 0 79580 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__A2
timestamp 1607194113
transform 1 0 81052 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1607194113
transform 1 0 79672 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1106_
timestamp 1607194113
transform 1 0 79764 0 1 39712
box -38 -48 1326 592
use sky130_fd_sc_hd__and3_4  _1116_
timestamp 1607194113
transform 1 0 82340 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_69_909
timestamp 1607194113
transform 1 0 84732 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_69_900
timestamp 1607194113
transform 1 0 83904 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_892
timestamp 1607194113
transform 1 0 83168 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__A
timestamp 1607194113
transform 1 0 84548 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0722_
timestamp 1607194113
transform 1 0 84180 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__B1
timestamp 1607194113
transform 1 0 85100 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__A1
timestamp 1607194113
transform 1 0 86572 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1607194113
transform 1 0 85284 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1111_
timestamp 1607194113
transform 1 0 85376 0 1 39712
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_1  FILLER_69_949
timestamp 1607194113
transform 1 0 88412 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_69_943
timestamp 1607194113
transform 1 0 87860 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_931
timestamp 1607194113
transform 1 0 86756 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0708_
timestamp 1607194113
transform 1 0 88504 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_965
timestamp 1607194113
transform 1 0 89884 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_69_953
timestamp 1607194113
transform 1 0 88780 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_973
timestamp 1607194113
transform 1 0 90620 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1460__CLK
timestamp 1607194113
transform 1 0 90712 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1607194113
transform 1 0 90896 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_751
timestamp 1607194113
transform 1 0 70196 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_739
timestamp 1607194113
transform 1 0 69092 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_767
timestamp 1607194113
transform 1 0 71668 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_605
timestamp 1607194113
transform 1 0 71300 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1090_
timestamp 1607194113
transform 1 0 71392 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_791
timestamp 1607194113
transform 1 0 73876 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__B1
timestamp 1607194113
transform 1 0 73692 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _1093_
timestamp 1607194113
transform 1 0 72404 0 -1 40800
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_70_809
timestamp 1607194113
transform 1 0 75532 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_799
timestamp 1607194113
transform 1 0 74612 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A
timestamp 1607194113
transform 1 0 75348 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1081_
timestamp 1607194113
transform 1 0 74704 0 -1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_70_825
timestamp 1607194113
transform 1 0 77004 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_821
timestamp 1607194113
transform 1 0 76636 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_606
timestamp 1607194113
transform 1 0 76912 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_849
timestamp 1607194113
transform 1 0 79212 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_837
timestamp 1607194113
transform 1 0 78108 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_861
timestamp 1607194113
transform 1 0 80316 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__A
timestamp 1607194113
transform 1 0 80592 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1095_
timestamp 1607194113
transform 1 0 80776 0 -1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_70_883
timestamp 1607194113
transform 1 0 82340 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_875
timestamp 1607194113
transform 1 0 81604 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__B
timestamp 1607194113
transform 1 0 81420 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_607
timestamp 1607194113
transform 1 0 82524 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1103_
timestamp 1607194113
transform 1 0 82616 0 -1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_70_907
timestamp 1607194113
transform 1 0 84548 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_895
timestamp 1607194113
transform 1 0 83444 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__A
timestamp 1607194113
transform 1 0 83260 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1112_
timestamp 1607194113
transform 1 0 85652 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_947
timestamp 1607194113
transform 1 0 88228 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_945
timestamp 1607194113
transform 1 0 88044 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_933
timestamp 1607194113
transform 1 0 86940 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__A1
timestamp 1607194113
transform 1 0 86756 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_608
timestamp 1607194113
transform 1 0 88136 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1462__CLK
timestamp 1607194113
transform 1 0 88964 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1462_
timestamp 1607194113
transform 1 0 89148 0 -1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_70_976
timestamp 1607194113
transform 1 0 90896 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_745
timestamp 1607194113
transform 1 0 69644 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_733
timestamp 1607194113
transform 1 0 68540 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_772
timestamp 1607194113
transform 1 0 72128 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_71_765
timestamp 1607194113
transform 1 0 71484 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_757
timestamp 1607194113
transform 1 0 70748 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__A
timestamp 1607194113
transform 1 0 71944 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1036_
timestamp 1607194113
transform 1 0 71668 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_71_785
timestamp 1607194113
transform 1 0 73324 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1082_
timestamp 1607194113
transform 1 0 72680 0 1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_71_807
timestamp 1607194113
transform 1 0 75348 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_794
timestamp 1607194113
transform 1 0 74152 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__C
timestamp 1607194113
transform 1 0 75164 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_624
timestamp 1607194113
transform 1 0 74060 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _1049_
timestamp 1607194113
transform 1 0 74336 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_71_831
timestamp 1607194113
transform 1 0 77556 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_819
timestamp 1607194113
transform 1 0 76452 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_844
timestamp 1607194113
transform 1 0 78752 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_839
timestamp 1607194113
transform 1 0 78292 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1105_
timestamp 1607194113
transform 1 0 78384 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_859
timestamp 1607194113
transform 1 0 80132 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_855
timestamp 1607194113
transform 1 0 79764 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_71_852
timestamp 1607194113
transform 1 0 79488 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__D
timestamp 1607194113
transform 1 0 80224 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A
timestamp 1607194113
transform 1 0 80408 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_625
timestamp 1607194113
transform 1 0 79672 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1035_
timestamp 1607194113
transform 1 0 80592 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_71_890
timestamp 1607194113
transform 1 0 82984 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_885
timestamp 1607194113
transform 1 0 82524 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_873
timestamp 1607194113
transform 1 0 81420 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _0748_
timestamp 1607194113
transform 1 0 82616 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_902
timestamp 1607194113
transform 1 0 84088 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_928
timestamp 1607194113
transform 1 0 86480 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_71_916
timestamp 1607194113
transform 1 0 85376 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_914
timestamp 1607194113
transform 1 0 85192 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_626
timestamp 1607194113
transform 1 0 85284 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_934
timestamp 1607194113
transform 1 0 87032 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1465__CLK
timestamp 1607194113
transform 1 0 87124 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1465_
timestamp 1607194113
transform 1 0 87308 0 1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_71_968
timestamp 1607194113
transform 1 0 90160 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_71_956
timestamp 1607194113
transform 1 0 89056 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_627
timestamp 1607194113
transform 1 0 90896 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_748
timestamp 1607194113
transform 1 0 69920 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_736
timestamp 1607194113
transform 1 0 68816 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_771
timestamp 1607194113
transform 1 0 72036 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_764
timestamp 1607194113
transform 1 0 71392 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_72_760
timestamp 1607194113
transform 1 0 71024 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_642
timestamp 1607194113
transform 1 0 71300 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _0750_
timestamp 1607194113
transform 1 0 71760 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_72_789
timestamp 1607194113
transform 1 0 73692 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_777
timestamp 1607194113
transform 1 0 72588 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__D
timestamp 1607194113
transform 1 0 72680 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1038_
timestamp 1607194113
transform 1 0 72864 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_72_804
timestamp 1607194113
transform 1 0 75072 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _1083_
timestamp 1607194113
transform 1 0 74428 0 -1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_72_825
timestamp 1607194113
transform 1 0 77004 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_72_816
timestamp 1607194113
transform 1 0 76176 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_643
timestamp 1607194113
transform 1 0 76912 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_841
timestamp 1607194113
transform 1 0 78476 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_833
timestamp 1607194113
transform 1 0 77740 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__A
timestamp 1607194113
transform 1 0 78292 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0779_
timestamp 1607194113
transform 1 0 77924 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_869
timestamp 1607194113
transform 1 0 81052 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_865
timestamp 1607194113
transform 1 0 80684 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_853
timestamp 1607194113
transform 1 0 79580 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _1096_
timestamp 1607194113
transform 1 0 81144 0 -1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_72_877
timestamp 1607194113
transform 1 0 81788 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_644
timestamp 1607194113
transform 1 0 82524 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__and3_4  _1104_
timestamp 1607194113
transform 1 0 82616 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_72_906
timestamp 1607194113
transform 1 0 84456 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_72_895
timestamp 1607194113
transform 1 0 83444 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1607194113
transform 1 0 84180 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_930
timestamp 1607194113
transform 1 0 86664 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_918
timestamp 1607194113
transform 1 0 85560 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_947
timestamp 1607194113
transform 1 0 88228 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_942
timestamp 1607194113
transform 1 0 87768 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_645
timestamp 1607194113
transform 1 0 88136 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_959
timestamp 1607194113
transform 1 0 89332 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_971
timestamp 1607194113
transform 1 0 90436 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_749
timestamp 1607194113
transform 1 0 70012 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_741
timestamp 1607194113
transform 1 0 69276 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_733
timestamp 1607194113
transform 1 0 68540 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A
timestamp 1607194113
transform 1 0 69828 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0751_
timestamp 1607194113
transform 1 0 69460 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_73_767
timestamp 1607194113
transform 1 0 71668 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__A1
timestamp 1607194113
transform 1 0 70380 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1086_
timestamp 1607194113
transform 1 0 70564 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_785
timestamp 1607194113
transform 1 0 73324 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_775
timestamp 1607194113
transform 1 0 72404 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1084_
timestamp 1607194113
transform 1 0 72680 0 1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_73_803
timestamp 1607194113
transform 1 0 74980 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_661
timestamp 1607194113
transform 1 0 74060 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _1088_
timestamp 1607194113
transform 1 0 74152 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_73_824
timestamp 1607194113
transform 1 0 76912 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_819
timestamp 1607194113
transform 1 0 76452 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_815
timestamp 1607194113
transform 1 0 76084 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1058_
timestamp 1607194113
transform 1 0 76544 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_73_848
timestamp 1607194113
transform 1 0 79120 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_73_836
timestamp 1607194113
transform 1 0 78016 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _1071_
timestamp 1607194113
transform 1 0 77648 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_871
timestamp 1607194113
transform 1 0 81236 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_859
timestamp 1607194113
transform 1 0 80132 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_855
timestamp 1607194113
transform 1 0 79764 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_662
timestamp 1607194113
transform 1 0 79672 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _1087_
timestamp 1607194113
transform 1 0 80868 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0778_
timestamp 1607194113
transform 1 0 79856 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_73_883
timestamp 1607194113
transform 1 0 82340 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1467__CLK
timestamp 1607194113
transform 1 0 82616 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1467_
timestamp 1607194113
transform 1 0 82800 0 1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_73_907
timestamp 1607194113
transform 1 0 84548 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_928
timestamp 1607194113
transform 1 0 86480 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_916
timestamp 1607194113
transform 1 0 85376 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_663
timestamp 1607194113
transform 1 0 85284 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_940
timestamp 1607194113
transform 1 0 87584 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_964
timestamp 1607194113
transform 1 0 89792 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_952
timestamp 1607194113
transform 1 0 88688 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_664
timestamp 1607194113
transform 1 0 90896 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_75_751
timestamp 1607194113
transform 1 0 70196 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_75_745
timestamp 1607194113
transform 1 0 69644 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_733
timestamp 1607194113
transform 1 0 68540 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_746
timestamp 1607194113
transform 1 0 69736 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__B1
timestamp 1607194113
transform 1 0 69552 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1473_
timestamp 1607194113
transform 1 0 70288 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_74_758
timestamp 1607194113
transform 1 0 70840 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1473__CLK
timestamp 1607194113
transform 1 0 72036 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__A1
timestamp 1607194113
transform 1 0 71116 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_679
timestamp 1607194113
transform 1 0 71300 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1085_
timestamp 1607194113
transform 1 0 71392 0 -1 42976
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_75_785
timestamp 1607194113
transform 1 0 73324 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_773
timestamp 1607194113
transform 1 0 72220 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_779
timestamp 1607194113
transform 1 0 72772 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1472__CLK
timestamp 1607194113
transform 1 0 73876 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__B1
timestamp 1607194113
transform 1 0 72588 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_803
timestamp 1607194113
transform 1 0 74980 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A
timestamp 1607194113
transform 1 0 75532 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_698
timestamp 1607194113
transform 1 0 74060 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1472_
timestamp 1607194113
transform 1 0 74060 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__and3_4  _1089_
timestamp 1607194113
transform 1 0 74152 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _1026_
timestamp 1607194113
transform 1 0 75716 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_75_827
timestamp 1607194113
transform 1 0 77188 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_815
timestamp 1607194113
transform 1 0 76084 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_830
timestamp 1607194113
transform 1 0 77464 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_74_812
timestamp 1607194113
transform 1 0 75808 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__A
timestamp 1607194113
transform 1 0 77280 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_680
timestamp 1607194113
transform 1 0 76912 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1057_
timestamp 1607194113
transform 1 0 77004 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_75_848
timestamp 1607194113
transform 1 0 79120 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_833
timestamp 1607194113
transform 1 0 77740 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_838
timestamp 1607194113
transform 1 0 78200 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1469__CLK
timestamp 1607194113
transform 1 0 78384 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__A1
timestamp 1607194113
transform 1 0 78936 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1469_
timestamp 1607194113
transform 1 0 78568 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _1099_
timestamp 1607194113
transform 1 0 77832 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_867
timestamp 1607194113
transform 1 0 80868 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_855
timestamp 1607194113
transform 1 0 79764 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_869
timestamp 1607194113
transform 1 0 81052 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_861
timestamp 1607194113
transform 1 0 80316 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_699
timestamp 1607194113
transform 1 0 79672 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1097_
timestamp 1607194113
transform 1 0 81144 0 -1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_75_888
timestamp 1607194113
transform 1 0 82800 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_886
timestamp 1607194113
transform 1 0 82616 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_877
timestamp 1607194113
transform 1 0 81788 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1468__CLK
timestamp 1607194113
transform 1 0 82340 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_681
timestamp 1607194113
transform 1 0 82524 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1468_
timestamp 1607194113
transform 1 0 82708 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2_4  _1100_
timestamp 1607194113
transform 1 0 81972 0 1 42976
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_75_901
timestamp 1607194113
transform 1 0 83996 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_906
timestamp 1607194113
transform 1 0 84456 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__A
timestamp 1607194113
transform 1 0 83812 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp 1607194113
transform 1 0 83536 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_928
timestamp 1607194113
transform 1 0 86480 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_916
timestamp 1607194113
transform 1 0 85376 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_913
timestamp 1607194113
transform 1 0 85100 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_930
timestamp 1607194113
transform 1 0 86664 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_918
timestamp 1607194113
transform 1 0 85560 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_700
timestamp 1607194113
transform 1 0 85284 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_940
timestamp 1607194113
transform 1 0 87584 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_947
timestamp 1607194113
transform 1 0 88228 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_942
timestamp 1607194113
transform 1 0 87768 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_682
timestamp 1607194113
transform 1 0 88136 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_964
timestamp 1607194113
transform 1 0 89792 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_952
timestamp 1607194113
transform 1 0 88688 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_959
timestamp 1607194113
transform 1 0 89332 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_971
timestamp 1607194113
transform 1 0 90436 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_701
timestamp 1607194113
transform 1 0 90896 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_745
timestamp 1607194113
transform 1 0 69644 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_738
timestamp 1607194113
transform 1 0 69000 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_727
timestamp 1607194113
transform 1 0 69552 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_769
timestamp 1607194113
transform 1 0 71852 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_757
timestamp 1607194113
transform 1 0 70748 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_788
timestamp 1607194113
transform 1 0 73600 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_776
timestamp 1607194113
transform 1 0 72496 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_728
timestamp 1607194113
transform 1 0 72404 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1607194113
transform 1 0 73784 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_807
timestamp 1607194113
transform 1 0 75348 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_803
timestamp 1607194113
transform 1 0 74980 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_76_795
timestamp 1607194113
transform 1 0 74244 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A
timestamp 1607194113
transform 1 0 74060 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_729
timestamp 1607194113
transform 1 0 75256 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_831
timestamp 1607194113
transform 1 0 77556 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_819
timestamp 1607194113
transform 1 0 76452 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_838
timestamp 1607194113
transform 1 0 78200 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__B1
timestamp 1607194113
transform 1 0 78384 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__A1
timestamp 1607194113
transform 1 0 78568 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_730
timestamp 1607194113
transform 1 0 78108 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__a21oi_4  _1098_
timestamp 1607194113
transform 1 0 78752 0 -1 44064
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_76_869
timestamp 1607194113
transform 1 0 81052 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_865
timestamp 1607194113
transform 1 0 80684 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_76_857
timestamp 1607194113
transform 1 0 79948 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_731
timestamp 1607194113
transform 1 0 80960 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_889
timestamp 1607194113
transform 1 0 82892 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_76_877
timestamp 1607194113
transform 1 0 81788 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _1101_
timestamp 1607194113
transform 1 0 82064 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_76_900
timestamp 1607194113
transform 1 0 83904 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_897
timestamp 1607194113
transform 1 0 83628 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_732
timestamp 1607194113
transform 1 0 83812 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_924
timestamp 1607194113
transform 1 0 86112 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_912
timestamp 1607194113
transform 1 0 85008 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_733
timestamp 1607194113
transform 1 0 86664 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_943
timestamp 1607194113
transform 1 0 87860 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_931
timestamp 1607194113
transform 1 0 86756 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_962
timestamp 1607194113
transform 1 0 89608 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_955
timestamp 1607194113
transform 1 0 88964 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_734
timestamp 1607194113
transform 1 0 89516 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_974
timestamp 1607194113
transform 1 0 90712 0 -1 44064
box -38 -48 1142 592
use delayline_9_ms  inst_rdelay_line
timestamp 1607276512
transform 1 0 80960 0 1 3761
box 800 801 23264 27367
use sky130_fd_sc_hd__decap_12  FILLER_60_989
timestamp 1607194113
transform 1 0 92092 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_977
timestamp 1607194113
transform 1 0 90988 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_59_996
timestamp 1607194113
transform 1 0 92736 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_984
timestamp 1607194113
transform 1 0 91632 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _1141_
timestamp 1607194113
transform 1 0 90988 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _0731_
timestamp 1607194113
transform 1 0 91724 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_1001
timestamp 1607194113
transform 1 0 93196 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1008
timestamp 1607194113
transform 1 0 93840 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1455__CLK
timestamp 1607194113
transform 1 0 93564 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1607194113
transform 1 0 93748 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1455_
timestamp 1607194113
transform 1 0 93840 0 -1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1027
timestamp 1607194113
transform 1 0 95588 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_1036
timestamp 1607194113
transform 1 0 96416 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_1032
timestamp 1607194113
transform 1 0 96048 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1020
timestamp 1607194113
transform 1 0 94944 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1051
timestamp 1607194113
transform 1 0 97796 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1039
timestamp 1607194113
transform 1 0 96692 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1050
timestamp 1607194113
transform 1 0 97704 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1038
timestamp 1607194113
transform 1 0 96600 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1607194113
transform 1 0 96508 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1069
timestamp 1607194113
transform 1 0 99452 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_1067
timestamp 1607194113
transform 1 0 99268 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_1063
timestamp 1607194113
transform 1 0 98900 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1074
timestamp 1607194113
transform 1 0 99912 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1062
timestamp 1607194113
transform 1 0 98808 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1607194113
transform 1 0 99360 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1093
timestamp 1607194113
transform 1 0 101660 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1081
timestamp 1607194113
transform 1 0 100556 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1086
timestamp 1607194113
transform 1 0 101016 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1105
timestamp 1607194113
transform 1 0 102764 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1111
timestamp 1607194113
transform 1 0 103316 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_1099
timestamp 1607194113
transform 1 0 102212 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1607194113
transform 1 0 102120 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_60_1130
timestamp 1607194113
transform 1 0 105064 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_1117
timestamp 1607194113
transform 1 0 103868 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_1131
timestamp 1607194113
transform 1 0 105156 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_1123
timestamp 1607194113
transform 1 0 104420 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1607194113
transform 1 0 104972 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1607194113
transform -1 0 105616 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1607194113
transform -1 0 105616 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_62_995
timestamp 1607194113
transform 1 0 92644 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_987
timestamp 1607194113
transform 1 0 91908 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_986
timestamp 1607194113
transform 1 0 91816 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _1146_
timestamp 1607194113
transform 1 0 90988 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1136_
timestamp 1607194113
transform 1 0 92736 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_61_1012
timestamp 1607194113
transform 1 0 94208 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_998
timestamp 1607194113
transform 1 0 92920 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__A
timestamp 1607194113
transform 1 0 94576 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__A
timestamp 1607194113
transform 1 0 94024 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _0726_
timestamp 1607194113
transform 1 0 93656 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_1008
timestamp 1607194113
transform 1 0 93840 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_62_999
timestamp 1607194113
transform 1 0 93012 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1458__CLK
timestamp 1607194113
transform 1 0 94392 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1607194113
transform 1 0 93748 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1458_
timestamp 1607194113
transform 1 0 94576 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_62_1035
timestamp 1607194113
transform 1 0 96324 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1025
timestamp 1607194113
transform 1 0 95404 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _1130_
timestamp 1607194113
transform 1 0 94760 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1047
timestamp 1607194113
transform 1 0 97428 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1053
timestamp 1607194113
transform 1 0 97980 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1041
timestamp 1607194113
transform 1 0 96876 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1607194113
transform 1 0 96508 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _0729_
timestamp 1607194113
transform 1 0 97060 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0725_
timestamp 1607194113
transform 1 0 96600 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1069
timestamp 1607194113
transform 1 0 99452 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_1067
timestamp 1607194113
transform 1 0 99268 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_1059
timestamp 1607194113
transform 1 0 98532 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1065
timestamp 1607194113
transform 1 0 99084 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1607194113
transform 1 0 99360 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1093
timestamp 1607194113
transform 1 0 101660 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1081
timestamp 1607194113
transform 1 0 100556 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_1089
timestamp 1607194113
transform 1 0 101292 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1077
timestamp 1607194113
transform 1 0 100188 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1105
timestamp 1607194113
transform 1 0 102764 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1111
timestamp 1607194113
transform 1 0 103316 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_1099
timestamp 1607194113
transform 1 0 102212 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_1097
timestamp 1607194113
transform 1 0 102028 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1607194113
transform 1 0 102120 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_1130
timestamp 1607194113
transform 1 0 105064 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_1117
timestamp 1607194113
transform 1 0 103868 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_1131
timestamp 1607194113
transform 1 0 105156 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_1123
timestamp 1607194113
transform 1 0 104420 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1607194113
transform 1 0 104972 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1607194113
transform -1 0 105616 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1607194113
transform -1 0 105616 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_989
timestamp 1607194113
transform 1 0 92092 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_979
timestamp 1607194113
transform 1 0 91172 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_994
timestamp 1607194113
transform 1 0 92552 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_982
timestamp 1607194113
transform 1 0 91448 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A
timestamp 1607194113
transform 1 0 91264 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__A
timestamp 1607194113
transform 1 0 91264 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1126_
timestamp 1607194113
transform 1 0 91448 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _0693_
timestamp 1607194113
transform 1 0 90988 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_986
timestamp 1607194113
transform 1 0 91816 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__A
timestamp 1607194113
transform 1 0 91632 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1123_
timestamp 1607194113
transform 1 0 90988 0 1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_64_1008
timestamp 1607194113
transform 1 0 93840 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_64_1001
timestamp 1607194113
transform 1 0 93196 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_1001
timestamp 1607194113
transform 1 0 93196 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__B1
timestamp 1607194113
transform 1 0 93564 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__A1
timestamp 1607194113
transform 1 0 93748 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1607194113
transform 1 0 93748 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _1135_
timestamp 1607194113
transform 1 0 93932 0 1 36448
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_4  _1133_
timestamp 1607194113
transform 1 0 94024 0 -1 37536
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1131_
timestamp 1607194113
transform 1 0 92920 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_65_1011
timestamp 1607194113
transform 1 0 94116 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_65_998
timestamp 1607194113
transform 1 0 92920 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__A
timestamp 1607194113
transform 1 0 93104 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1127_
timestamp 1607194113
transform 1 0 93288 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_65_1029
timestamp 1607194113
transform 1 0 95772 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_1017
timestamp 1607194113
transform 1 0 94668 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_1017
timestamp 1607194113
transform 1 0 94668 0 -1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1035
timestamp 1607194113
transform 1 0 96324 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1023
timestamp 1607194113
transform 1 0 95220 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1459__CLK
timestamp 1607194113
transform 1 0 95220 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__A
timestamp 1607194113
transform 1 0 94760 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1459_
timestamp 1607194113
transform 1 0 95404 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__and3_4  _1134_
timestamp 1607194113
transform 1 0 94944 0 1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1056
timestamp 1607194113
transform 1 0 98256 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1044
timestamp 1607194113
transform 1 0 97152 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1047
timestamp 1607194113
transform 1 0 97428 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__A
timestamp 1607194113
transform 1 0 97244 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1607194113
transform 1 0 96508 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _1132_
timestamp 1607194113
transform 1 0 96600 0 1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1053
timestamp 1607194113
transform 1 0 97980 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1041
timestamp 1607194113
transform 1 0 96876 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1607194113
transform 1 0 96508 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1607194113
transform 1 0 96600 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1065
timestamp 1607194113
transform 1 0 99084 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1069
timestamp 1607194113
transform 1 0 99452 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1071
timestamp 1607194113
transform 1 0 99636 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1059
timestamp 1607194113
transform 1 0 98532 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1607194113
transform 1 0 99360 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_1089
timestamp 1607194113
transform 1 0 101292 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1077
timestamp 1607194113
transform 1 0 100188 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1093
timestamp 1607194113
transform 1 0 101660 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1081
timestamp 1607194113
transform 1 0 100556 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_1095
timestamp 1607194113
transform 1 0 101844 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1083
timestamp 1607194113
transform 1 0 100740 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1111
timestamp 1607194113
transform 1 0 103316 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_1099
timestamp 1607194113
transform 1 0 102212 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_1097
timestamp 1607194113
transform 1 0 102028 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1105
timestamp 1607194113
transform 1 0 102764 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1111
timestamp 1607194113
transform 1 0 103316 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_1099
timestamp 1607194113
transform 1 0 102212 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1607194113
transform 1 0 102120 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1607194113
transform 1 0 102120 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_1130
timestamp 1607194113
transform 1 0 105064 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_1117
timestamp 1607194113
transform 1 0 103868 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_1131
timestamp 1607194113
transform 1 0 105156 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_1123
timestamp 1607194113
transform 1 0 104420 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1607194113
transform 1 0 104972 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1607194113
transform -1 0 105616 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1607194113
transform -1 0 105616 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_1131
timestamp 1607194113
transform 1 0 105156 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_1123
timestamp 1607194113
transform 1 0 104420 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1607194113
transform -1 0 105616 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_992
timestamp 1607194113
transform 1 0 92368 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_980
timestamp 1607194113
transform 1 0 91264 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_994
timestamp 1607194113
transform 1 0 92552 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_986
timestamp 1607194113
transform 1 0 91816 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_67_977
timestamp 1607194113
transform 1 0 90988 0 1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_985
timestamp 1607194113
transform 1 0 91724 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1129_
timestamp 1607194113
transform 1 0 90988 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _1125_
timestamp 1607194113
transform 1 0 92644 0 1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1124_
timestamp 1607194113
transform 1 0 91540 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_66_1008
timestamp 1607194113
transform 1 0 93840 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_1005
timestamp 1607194113
transform 1 0 93564 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_997
timestamp 1607194113
transform 1 0 92828 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1461__CLK
timestamp 1607194113
transform 1 0 94116 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1607194113
transform 1 0 93748 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1461_
timestamp 1607194113
transform 1 0 94300 0 -1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1008
timestamp 1607194113
transform 1 0 93840 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_1004
timestamp 1607194113
transform 1 0 93472 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1016
timestamp 1607194113
transform 1 0 94576 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1004
timestamp 1607194113
transform 1 0 93472 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__A
timestamp 1607194113
transform 1 0 93288 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1607194113
transform 1 0 93748 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1032
timestamp 1607194113
transform 1 0 96048 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1020
timestamp 1607194113
transform 1 0 94944 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_1036
timestamp 1607194113
transform 1 0 96416 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_1028
timestamp 1607194113
transform 1 0 95680 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1032
timestamp 1607194113
transform 1 0 96048 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1056
timestamp 1607194113
transform 1 0 98256 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1044
timestamp 1607194113
transform 1 0 97152 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1050
timestamp 1607194113
transform 1 0 97704 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1038
timestamp 1607194113
transform 1 0 96600 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1056
timestamp 1607194113
transform 1 0 98256 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1044
timestamp 1607194113
transform 1 0 97152 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1607194113
transform 1 0 96508 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1069
timestamp 1607194113
transform 1 0 99452 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1074
timestamp 1607194113
transform 1 0 99912 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1062
timestamp 1607194113
transform 1 0 98808 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1069
timestamp 1607194113
transform 1 0 99452 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1607194113
transform 1 0 99360 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1607194113
transform 1 0 99360 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1093
timestamp 1607194113
transform 1 0 101660 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1081
timestamp 1607194113
transform 1 0 100556 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1086
timestamp 1607194113
transform 1 0 101016 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1093
timestamp 1607194113
transform 1 0 101660 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1081
timestamp 1607194113
transform 1 0 100556 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1105
timestamp 1607194113
transform 1 0 102764 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1111
timestamp 1607194113
transform 1 0 103316 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_1099
timestamp 1607194113
transform 1 0 102212 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1105
timestamp 1607194113
transform 1 0 102764 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1607194113
transform 1 0 102120 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_66_1130
timestamp 1607194113
transform 1 0 105064 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_1117
timestamp 1607194113
transform 1 0 103868 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1607194113
transform 1 0 104972 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1607194113
transform -1 0 105616 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_68_1130
timestamp 1607194113
transform 1 0 105064 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_1117
timestamp 1607194113
transform 1 0 103868 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_1131
timestamp 1607194113
transform 1 0 105156 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_1123
timestamp 1607194113
transform 1 0 104420 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1607194113
transform 1 0 104972 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1607194113
transform -1 0 105616 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1607194113
transform -1 0 105616 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_989
timestamp 1607194113
transform 1 0 92092 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_977
timestamp 1607194113
transform 1 0 90988 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_988
timestamp 1607194113
transform 1 0 92000 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_996
timestamp 1607194113
transform 1 0 92736 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1460_
timestamp 1607194113
transform 1 0 90988 0 1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1013
timestamp 1607194113
transform 1 0 94300 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1001
timestamp 1607194113
transform 1 0 93196 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1008
timestamp 1607194113
transform 1 0 93840 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_1006
timestamp 1607194113
transform 1 0 93656 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_1000
timestamp 1607194113
transform 1 0 93104 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1008
timestamp 1607194113
transform 1 0 93840 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_609
timestamp 1607194113
transform 1 0 93748 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1025
timestamp 1607194113
transform 1 0 95404 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1032
timestamp 1607194113
transform 1 0 96048 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1020
timestamp 1607194113
transform 1 0 94944 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_1036
timestamp 1607194113
transform 1 0 96416 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_1032
timestamp 1607194113
transform 1 0 96048 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1020
timestamp 1607194113
transform 1 0 94944 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1050
timestamp 1607194113
transform 1 0 97704 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1038
timestamp 1607194113
transform 1 0 96600 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1056
timestamp 1607194113
transform 1 0 98256 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1044
timestamp 1607194113
transform 1 0 97152 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1050
timestamp 1607194113
transform 1 0 97704 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1038
timestamp 1607194113
transform 1 0 96600 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_628
timestamp 1607194113
transform 1 0 96508 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_591
timestamp 1607194113
transform 1 0 96508 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1074
timestamp 1607194113
transform 1 0 99912 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1062
timestamp 1607194113
transform 1 0 98808 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1069
timestamp 1607194113
transform 1 0 99452 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1074
timestamp 1607194113
transform 1 0 99912 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1062
timestamp 1607194113
transform 1 0 98808 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_610
timestamp 1607194113
transform 1 0 99360 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1086
timestamp 1607194113
transform 1 0 101016 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1093
timestamp 1607194113
transform 1 0 101660 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1081
timestamp 1607194113
transform 1 0 100556 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1086
timestamp 1607194113
transform 1 0 101016 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1111
timestamp 1607194113
transform 1 0 103316 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_1099
timestamp 1607194113
transform 1 0 102212 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1105
timestamp 1607194113
transform 1 0 102764 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1111
timestamp 1607194113
transform 1 0 103316 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_1099
timestamp 1607194113
transform 1 0 102212 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_629
timestamp 1607194113
transform 1 0 102120 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_592
timestamp 1607194113
transform 1 0 102120 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_1131
timestamp 1607194113
transform 1 0 105156 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_1123
timestamp 1607194113
transform 1 0 104420 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1607194113
transform -1 0 105616 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_70_1130
timestamp 1607194113
transform 1 0 105064 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_1117
timestamp 1607194113
transform 1 0 103868 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_611
timestamp 1607194113
transform 1 0 104972 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1607194113
transform -1 0 105616 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_1131
timestamp 1607194113
transform 1 0 105156 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_1123
timestamp 1607194113
transform 1 0 104420 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1607194113
transform -1 0 105616 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_995
timestamp 1607194113
transform 1 0 92644 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_983
timestamp 1607194113
transform 1 0 91540 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_989
timestamp 1607194113
transform 1 0 92092 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_977
timestamp 1607194113
transform 1 0 90988 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_995
timestamp 1607194113
transform 1 0 92644 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_983
timestamp 1607194113
transform 1 0 91540 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1008
timestamp 1607194113
transform 1 0 93840 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1013
timestamp 1607194113
transform 1 0 94300 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1001
timestamp 1607194113
transform 1 0 93196 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1008
timestamp 1607194113
transform 1 0 93840 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_683
timestamp 1607194113
transform 1 0 93748 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_646
timestamp 1607194113
transform 1 0 93748 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1032
timestamp 1607194113
transform 1 0 96048 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1020
timestamp 1607194113
transform 1 0 94944 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1025
timestamp 1607194113
transform 1 0 95404 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1032
timestamp 1607194113
transform 1 0 96048 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1020
timestamp 1607194113
transform 1 0 94944 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1056
timestamp 1607194113
transform 1 0 98256 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1044
timestamp 1607194113
transform 1 0 97152 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1050
timestamp 1607194113
transform 1 0 97704 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1038
timestamp 1607194113
transform 1 0 96600 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1056
timestamp 1607194113
transform 1 0 98256 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1044
timestamp 1607194113
transform 1 0 97152 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_665
timestamp 1607194113
transform 1 0 96508 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1069
timestamp 1607194113
transform 1 0 99452 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1074
timestamp 1607194113
transform 1 0 99912 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1062
timestamp 1607194113
transform 1 0 98808 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1069
timestamp 1607194113
transform 1 0 99452 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_684
timestamp 1607194113
transform 1 0 99360 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_647
timestamp 1607194113
transform 1 0 99360 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1093
timestamp 1607194113
transform 1 0 101660 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1081
timestamp 1607194113
transform 1 0 100556 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1086
timestamp 1607194113
transform 1 0 101016 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1093
timestamp 1607194113
transform 1 0 101660 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1081
timestamp 1607194113
transform 1 0 100556 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1105
timestamp 1607194113
transform 1 0 102764 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1111
timestamp 1607194113
transform 1 0 103316 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_1099
timestamp 1607194113
transform 1 0 102212 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1105
timestamp 1607194113
transform 1 0 102764 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_666
timestamp 1607194113
transform 1 0 102120 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_72_1130
timestamp 1607194113
transform 1 0 105064 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_1117
timestamp 1607194113
transform 1 0 103868 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_648
timestamp 1607194113
transform 1 0 104972 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1607194113
transform -1 0 105616 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_1131
timestamp 1607194113
transform 1 0 105156 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_1123
timestamp 1607194113
transform 1 0 104420 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1607194113
transform -1 0 105616 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_74_1130
timestamp 1607194113
transform 1 0 105064 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_1117
timestamp 1607194113
transform 1 0 103868 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_685
timestamp 1607194113
transform 1 0 104972 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1607194113
transform -1 0 105616 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_993
timestamp 1607194113
transform 1 0 92460 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_986
timestamp 1607194113
transform 1 0 91816 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_989
timestamp 1607194113
transform 1 0 92092 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_977
timestamp 1607194113
transform 1 0 90988 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_735
timestamp 1607194113
transform 1 0 92368 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1005
timestamp 1607194113
transform 1 0 93564 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1013
timestamp 1607194113
transform 1 0 94300 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1001
timestamp 1607194113
transform 1 0 93196 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1036
timestamp 1607194113
transform 1 0 96416 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1024
timestamp 1607194113
transform 1 0 95312 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_1017
timestamp 1607194113
transform 1 0 94668 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1025
timestamp 1607194113
transform 1 0 95404 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_736
timestamp 1607194113
transform 1 0 95220 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1055
timestamp 1607194113
transform 1 0 98164 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_1048
timestamp 1607194113
transform 1 0 97520 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1050
timestamp 1607194113
transform 1 0 97704 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1038
timestamp 1607194113
transform 1 0 96600 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_737
timestamp 1607194113
transform 1 0 98072 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_702
timestamp 1607194113
transform 1 0 96508 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1067
timestamp 1607194113
transform 1 0 99268 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1074
timestamp 1607194113
transform 1 0 99912 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1062
timestamp 1607194113
transform 1 0 98808 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1086
timestamp 1607194113
transform 1 0 101016 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_1079
timestamp 1607194113
transform 1 0 100372 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1086
timestamp 1607194113
transform 1 0 101016 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_738
timestamp 1607194113
transform 1 0 100924 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_1110
timestamp 1607194113
transform 1 0 103224 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1098
timestamp 1607194113
transform 1 0 102120 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1111
timestamp 1607194113
transform 1 0 103316 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_1099
timestamp 1607194113
transform 1 0 102212 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_703
timestamp 1607194113
transform 1 0 102120 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_1129
timestamp 1607194113
transform 1 0 104972 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_1117
timestamp 1607194113
transform 1 0 103868 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_1131
timestamp 1607194113
transform 1 0 105156 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_1123
timestamp 1607194113
transform 1 0 104420 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_739
timestamp 1607194113
transform 1 0 103776 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1607194113
transform -1 0 105616 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1607194113
transform -1 0 105616 0 1 42976
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 280 800 400 6 bus_in[0]
port 0 nsew default input
rlabel metal3 s 0 12112 800 12232 6 bus_in[10]
port 1 nsew default input
rlabel metal3 s 0 13200 800 13320 6 bus_in[11]
port 2 nsew default input
rlabel metal3 s 0 14424 800 14544 6 bus_in[12]
port 3 nsew default input
rlabel metal3 s 0 15648 800 15768 6 bus_in[13]
port 4 nsew default input
rlabel metal3 s 0 16872 800 16992 6 bus_in[14]
port 5 nsew default input
rlabel metal3 s 0 17960 800 18080 6 bus_in[15]
port 6 nsew default input
rlabel metal3 s 0 19184 800 19304 6 bus_in[16]
port 7 nsew default input
rlabel metal3 s 0 20408 800 20528 6 bus_in[17]
port 8 nsew default input
rlabel metal3 s 0 21496 800 21616 6 bus_in[18]
port 9 nsew default input
rlabel metal3 s 0 22720 800 22840 6 bus_in[19]
port 10 nsew default input
rlabel metal3 s 0 1368 800 1488 6 bus_in[1]
port 11 nsew default input
rlabel metal3 s 0 23944 800 24064 6 bus_in[20]
port 12 nsew default input
rlabel metal3 s 0 25168 800 25288 6 bus_in[21]
port 13 nsew default input
rlabel metal3 s 0 26256 800 26376 6 bus_in[22]
port 14 nsew default input
rlabel metal3 s 0 27480 800 27600 6 bus_in[23]
port 15 nsew default input
rlabel metal3 s 0 28704 800 28824 6 bus_in[24]
port 16 nsew default input
rlabel metal3 s 0 29792 800 29912 6 bus_in[25]
port 17 nsew default input
rlabel metal3 s 0 31016 800 31136 6 bus_in[26]
port 18 nsew default input
rlabel metal3 s 0 32240 800 32360 6 bus_in[27]
port 19 nsew default input
rlabel metal3 s 0 33464 800 33584 6 bus_in[28]
port 20 nsew default input
rlabel metal3 s 0 34552 800 34672 6 bus_in[29]
port 21 nsew default input
rlabel metal3 s 0 2592 800 2712 6 bus_in[2]
port 22 nsew default input
rlabel metal3 s 0 35776 800 35896 6 bus_in[30]
port 23 nsew default input
rlabel metal3 s 0 37000 800 37120 6 bus_in[31]
port 24 nsew default input
rlabel metal3 s 0 38088 800 38208 6 bus_in[32]
port 25 nsew default input
rlabel metal3 s 0 39312 800 39432 6 bus_in[33]
port 26 nsew default input
rlabel metal3 s 0 40536 800 40656 6 bus_in[34]
port 27 nsew default input
rlabel metal3 s 0 41760 800 41880 6 bus_in[35]
port 28 nsew default input
rlabel metal3 s 0 42304 800 42424 6 bus_in[36]
port 29 nsew default input
rlabel metal3 s 0 42848 800 42968 6 bus_in[37]
port 30 nsew default input
rlabel metal3 s 0 43528 800 43648 6 bus_in[38]
port 31 nsew default input
rlabel metal3 s 0 44072 800 44192 6 bus_in[39]
port 32 nsew default input
rlabel metal3 s 0 3816 800 3936 6 bus_in[3]
port 33 nsew default input
rlabel metal3 s 0 44616 800 44736 6 bus_in[40]
port 34 nsew default input
rlabel metal3 s 0 45296 800 45416 6 bus_in[41]
port 35 nsew default input
rlabel metal3 s 0 4904 800 5024 6 bus_in[4]
port 36 nsew default input
rlabel metal3 s 0 6128 800 6248 6 bus_in[5]
port 37 nsew default input
rlabel metal3 s 0 7352 800 7472 6 bus_in[6]
port 38 nsew default input
rlabel metal3 s 0 8576 800 8696 6 bus_in[7]
port 39 nsew default input
rlabel metal3 s 0 9664 800 9784 6 bus_in[8]
port 40 nsew default input
rlabel metal3 s 0 10888 800 11008 6 bus_in[9]
port 41 nsew default input
rlabel metal3 s 0 824 800 944 6 bus_out[0]
port 42 nsew default tristate
rlabel metal3 s 0 12656 800 12776 6 bus_out[10]
port 43 nsew default tristate
rlabel metal3 s 0 13880 800 14000 6 bus_out[11]
port 44 nsew default tristate
rlabel metal3 s 0 14968 800 15088 6 bus_out[12]
port 45 nsew default tristate
rlabel metal3 s 0 16192 800 16312 6 bus_out[13]
port 46 nsew default tristate
rlabel metal3 s 0 17416 800 17536 6 bus_out[14]
port 47 nsew default tristate
rlabel metal3 s 0 18640 800 18760 6 bus_out[15]
port 48 nsew default tristate
rlabel metal3 s 0 19728 800 19848 6 bus_out[16]
port 49 nsew default tristate
rlabel metal3 s 0 20952 800 21072 6 bus_out[17]
port 50 nsew default tristate
rlabel metal3 s 0 22176 800 22296 6 bus_out[18]
port 51 nsew default tristate
rlabel metal3 s 0 23400 800 23520 6 bus_out[19]
port 52 nsew default tristate
rlabel metal3 s 0 2048 800 2168 6 bus_out[1]
port 53 nsew default tristate
rlabel metal3 s 0 24488 800 24608 6 bus_out[20]
port 54 nsew default tristate
rlabel metal3 s 0 25712 800 25832 6 bus_out[21]
port 55 nsew default tristate
rlabel metal3 s 0 26936 800 27056 6 bus_out[22]
port 56 nsew default tristate
rlabel metal3 s 0 28024 800 28144 6 bus_out[23]
port 57 nsew default tristate
rlabel metal3 s 0 29248 800 29368 6 bus_out[24]
port 58 nsew default tristate
rlabel metal3 s 0 30472 800 30592 6 bus_out[25]
port 59 nsew default tristate
rlabel metal3 s 0 31696 800 31816 6 bus_out[26]
port 60 nsew default tristate
rlabel metal3 s 0 32784 800 32904 6 bus_out[27]
port 61 nsew default tristate
rlabel metal3 s 0 34008 800 34128 6 bus_out[28]
port 62 nsew default tristate
rlabel metal3 s 0 35232 800 35352 6 bus_out[29]
port 63 nsew default tristate
rlabel metal3 s 0 3136 800 3256 6 bus_out[2]
port 64 nsew default tristate
rlabel metal3 s 0 36320 800 36440 6 bus_out[30]
port 65 nsew default tristate
rlabel metal3 s 0 37544 800 37664 6 bus_out[31]
port 66 nsew default tristate
rlabel metal3 s 0 38768 800 38888 6 bus_out[32]
port 67 nsew default tristate
rlabel metal3 s 0 39992 800 40112 6 bus_out[33]
port 68 nsew default tristate
rlabel metal3 s 0 41080 800 41200 6 bus_out[34]
port 69 nsew default tristate
rlabel metal3 s 0 4360 800 4480 6 bus_out[3]
port 70 nsew default tristate
rlabel metal3 s 0 5584 800 5704 6 bus_out[4]
port 71 nsew default tristate
rlabel metal3 s 0 6672 800 6792 6 bus_out[5]
port 72 nsew default tristate
rlabel metal3 s 0 7896 800 8016 6 bus_out[6]
port 73 nsew default tristate
rlabel metal3 s 0 9120 800 9240 6 bus_out[7]
port 74 nsew default tristate
rlabel metal3 s 0 10344 800 10464 6 bus_out[8]
port 75 nsew default tristate
rlabel metal3 s 0 11432 800 11552 6 bus_out[9]
port 76 nsew default tristate
rlabel metal2 s 53378 0 53434 800 6 clk_i
port 77 nsew default input
rlabel metal3 s 0 45840 800 45960 6 out1_o
port 78 nsew default tristate
rlabel metal3 s 105920 23128 106720 23248 6 out2_o
port 79 nsew default tristate
rlabel metal2 s 53378 45440 53434 46240 6 rst_n_i
port 80 nsew default input
rlabel metal5 s 1104 6436 105616 7036 6 VPWR
port 81 nsew default input
rlabel metal5 s 1104 24436 105616 25036 6 VGND
port 82 nsew default input
<< properties >>
string FIXED_BBOX 0 0 106720 46240
<< end >>
