magic
tech sky130A
magscale 1 2
timestamp 1608318970
<< metal1 >>
rect 287698 700544 287704 700596
rect 287756 700584 287762 700596
rect 332502 700584 332508 700596
rect 287756 700556 332508 700584
rect 287756 700544 287762 700556
rect 332502 700544 332508 700556
rect 332560 700544 332566 700596
rect 305638 700476 305644 700528
rect 305696 700516 305702 700528
rect 397454 700516 397460 700528
rect 305696 700488 397460 700516
rect 305696 700476 305702 700488
rect 397454 700476 397460 700488
rect 397512 700476 397518 700528
rect 313918 700408 313924 700460
rect 313976 700448 313982 700460
rect 413646 700448 413652 700460
rect 313976 700420 413652 700448
rect 313976 700408 313982 700420
rect 413646 700408 413652 700420
rect 413704 700408 413710 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 138658 700340 138664 700392
rect 138716 700380 138722 700392
rect 154114 700380 154120 700392
rect 138716 700352 154120 700380
rect 138716 700340 138722 700352
rect 154114 700340 154120 700352
rect 154172 700340 154178 700392
rect 308398 700340 308404 700392
rect 308456 700380 308462 700392
rect 462314 700380 462320 700392
rect 308456 700352 462320 700380
rect 308456 700340 308462 700352
rect 462314 700340 462320 700352
rect 462372 700340 462378 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 8938 700312 8944 700324
rect 8168 700284 8944 700312
rect 8168 700272 8174 700284
rect 8938 700272 8944 700284
rect 8996 700272 9002 700324
rect 89162 700272 89168 700324
rect 89220 700312 89226 700324
rect 138750 700312 138756 700324
rect 89220 700284 138756 700312
rect 89220 700272 89226 700284
rect 138750 700272 138756 700284
rect 138808 700272 138814 700324
rect 202782 700272 202788 700324
rect 202840 700312 202846 700324
rect 250898 700312 250904 700324
rect 202840 700284 250904 700312
rect 202840 700272 202846 700284
rect 250898 700272 250904 700284
rect 250956 700272 250962 700324
rect 267642 700272 267648 700324
rect 267700 700312 267706 700324
rect 282270 700312 282276 700324
rect 267700 700284 282276 700312
rect 267700 700272 267706 700284
rect 282270 700272 282276 700284
rect 282328 700272 282334 700324
rect 309778 700272 309784 700324
rect 309836 700312 309842 700324
rect 527174 700312 527180 700324
rect 309836 700284 527180 700312
rect 309836 700272 309842 700284
rect 527174 700272 527180 700284
rect 527232 700272 527238 700324
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 250898 699116 250904 699168
rect 250956 699156 250962 699168
rect 253198 699156 253204 699168
rect 250956 699128 253204 699156
rect 250956 699116 250962 699128
rect 253198 699116 253204 699128
rect 253256 699116 253262 699168
rect 283282 698232 283288 698284
rect 283340 698272 283346 698284
rect 283926 698272 283932 698284
rect 283340 698244 283932 698272
rect 283340 698232 283346 698244
rect 283926 698232 283932 698244
rect 283984 698232 283990 698284
rect 576118 696940 576124 696992
rect 576176 696980 576182 696992
rect 580166 696980 580172 696992
rect 576176 696952 580172 696980
rect 576176 696940 576182 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 133138 696872 133144 696924
rect 133196 696912 133202 696924
rect 137830 696912 137836 696924
rect 133196 696884 137836 696912
rect 133196 696872 133202 696884
rect 137830 696872 137836 696884
rect 137888 696872 137894 696924
rect 253198 696872 253204 696924
rect 253256 696912 253262 696924
rect 260006 696912 260012 696924
rect 253256 696884 260012 696912
rect 253256 696872 253262 696884
rect 260006 696872 260012 696884
rect 260064 696872 260070 696924
rect 260006 694764 260012 694816
rect 260064 694804 260070 694816
rect 266998 694804 267004 694816
rect 260064 694776 267004 694804
rect 260064 694764 260070 694776
rect 266998 694764 267004 694776
rect 267056 694764 267062 694816
rect 218974 694152 218980 694204
rect 219032 694192 219038 694204
rect 219158 694192 219164 694204
rect 219032 694164 219164 694192
rect 219032 694152 219038 694164
rect 219158 694152 219164 694164
rect 219216 694152 219222 694204
rect 283098 694084 283104 694136
rect 283156 694124 283162 694136
rect 283282 694124 283288 694136
rect 283156 694096 283288 694124
rect 283156 694084 283162 694096
rect 283282 694084 283288 694096
rect 283340 694084 283346 694136
rect 219158 688684 219164 688696
rect 219084 688656 219164 688684
rect 219084 688628 219112 688656
rect 219158 688644 219164 688656
rect 219216 688644 219222 688696
rect 219066 688576 219072 688628
rect 219124 688576 219130 688628
rect 283006 684496 283012 684548
rect 283064 684536 283070 684548
rect 283098 684536 283104 684548
rect 283064 684508 283104 684536
rect 283064 684496 283070 684508
rect 283098 684496 283104 684508
rect 283156 684496 283162 684548
rect 3510 681708 3516 681760
rect 3568 681748 3574 681760
rect 453298 681748 453304 681760
rect 3568 681720 453304 681748
rect 3568 681708 3574 681720
rect 453298 681708 453304 681720
rect 453356 681708 453362 681760
rect 218790 676132 218796 676184
rect 218848 676172 218854 676184
rect 218974 676172 218980 676184
rect 218848 676144 218980 676172
rect 218848 676132 218854 676144
rect 218974 676132 218980 676144
rect 219032 676132 219038 676184
rect 122098 675452 122104 675504
rect 122156 675492 122162 675504
rect 133138 675492 133144 675504
rect 122156 675464 133144 675492
rect 122156 675452 122162 675464
rect 133138 675452 133144 675464
rect 133196 675452 133202 675504
rect 266998 670624 267004 670676
rect 267056 670664 267062 670676
rect 268378 670664 268384 670676
rect 267056 670636 268384 670664
rect 267056 670624 267062 670636
rect 268378 670624 268384 670636
rect 268436 670624 268442 670676
rect 218790 666544 218796 666596
rect 218848 666584 218854 666596
rect 219066 666584 219072 666596
rect 218848 666556 219072 666584
rect 218848 666544 218854 666556
rect 219066 666544 219072 666556
rect 219124 666544 219130 666596
rect 283098 666544 283104 666596
rect 283156 666584 283162 666596
rect 283374 666584 283380 666596
rect 283156 666556 283380 666584
rect 283156 666544 283162 666556
rect 283374 666544 283380 666556
rect 283432 666544 283438 666596
rect 283098 661716 283104 661768
rect 283156 661756 283162 661768
rect 283374 661756 283380 661768
rect 283156 661728 283380 661756
rect 283156 661716 283162 661728
rect 283374 661716 283380 661728
rect 283432 661716 283438 661768
rect 268378 661172 268384 661224
rect 268436 661212 268442 661224
rect 270402 661212 270408 661224
rect 268436 661184 270408 661212
rect 268436 661172 268442 661184
rect 270402 661172 270408 661184
rect 270460 661172 270466 661224
rect 219158 659608 219164 659660
rect 219216 659648 219222 659660
rect 219342 659648 219348 659660
rect 219216 659620 219348 659648
rect 219216 659608 219222 659620
rect 219342 659608 219348 659620
rect 219400 659608 219406 659660
rect 116578 658520 116584 658572
rect 116636 658560 116642 658572
rect 122098 658560 122104 658572
rect 116636 658532 122104 658560
rect 116636 658520 116642 658532
rect 122098 658520 122104 658532
rect 122156 658520 122162 658572
rect 270402 656888 270408 656940
rect 270460 656928 270466 656940
rect 270460 656900 270540 656928
rect 270460 656888 270466 656900
rect 219066 656820 219072 656872
rect 219124 656860 219130 656872
rect 219342 656860 219348 656872
rect 219124 656832 219348 656860
rect 219124 656820 219130 656832
rect 219342 656820 219348 656832
rect 219400 656820 219406 656872
rect 270512 656860 270540 656900
rect 283098 656888 283104 656940
rect 283156 656928 283162 656940
rect 283190 656928 283196 656940
rect 283156 656900 283196 656928
rect 283156 656888 283162 656900
rect 283190 656888 283196 656900
rect 283248 656888 283254 656940
rect 273254 656860 273260 656872
rect 270512 656832 273260 656860
rect 273254 656820 273260 656832
rect 273312 656820 273318 656872
rect 273254 654100 273260 654152
rect 273312 654140 273318 654152
rect 273312 654112 274680 654140
rect 273312 654100 273318 654112
rect 274652 654072 274680 654112
rect 276658 654072 276664 654084
rect 274652 654044 276664 654072
rect 276658 654032 276664 654044
rect 276716 654032 276722 654084
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 10318 652780 10324 652792
rect 3108 652752 10324 652780
rect 3108 652740 3114 652752
rect 10318 652740 10324 652752
rect 10376 652740 10382 652792
rect 577498 650020 577504 650072
rect 577556 650060 577562 650072
rect 579614 650060 579620 650072
rect 577556 650032 579620 650060
rect 577556 650020 577562 650032
rect 579614 650020 579620 650032
rect 579672 650020 579678 650072
rect 113818 648864 113824 648916
rect 113876 648904 113882 648916
rect 116578 648904 116584 648916
rect 113876 648876 116584 648904
rect 113876 648864 113882 648876
rect 116578 648864 116584 648876
rect 116636 648864 116642 648916
rect 219066 647232 219072 647284
rect 219124 647272 219130 647284
rect 219250 647272 219256 647284
rect 219124 647244 219256 647272
rect 219124 647232 219130 647244
rect 219250 647232 219256 647244
rect 219308 647232 219314 647284
rect 283098 647232 283104 647284
rect 283156 647272 283162 647284
rect 283190 647272 283196 647284
rect 283156 647244 283196 647272
rect 283156 647232 283162 647244
rect 283190 647232 283196 647244
rect 283248 647232 283254 647284
rect 554406 647232 554412 647284
rect 554464 647272 554470 647284
rect 556246 647272 556252 647284
rect 554464 647244 556252 647272
rect 554464 647232 554470 647244
rect 556246 647232 556252 647244
rect 556304 647232 556310 647284
rect 219250 640404 219256 640416
rect 219084 640376 219256 640404
rect 219084 640280 219112 640376
rect 219250 640364 219256 640376
rect 219308 640364 219314 640416
rect 283098 640364 283104 640416
rect 283156 640404 283162 640416
rect 283190 640404 283196 640416
rect 283156 640376 283196 640404
rect 283156 640364 283162 640376
rect 283190 640364 283196 640376
rect 283248 640364 283254 640416
rect 219066 640228 219072 640280
rect 219124 640228 219130 640280
rect 219066 637508 219072 637560
rect 219124 637548 219130 637560
rect 219158 637548 219164 637560
rect 219124 637520 219164 637548
rect 219124 637508 219130 637520
rect 219158 637508 219164 637520
rect 219216 637508 219222 637560
rect 276658 635060 276664 635112
rect 276716 635100 276722 635112
rect 278038 635100 278044 635112
rect 276716 635072 278044 635100
rect 276716 635060 276722 635072
rect 278038 635060 278044 635072
rect 278096 635060 278102 635112
rect 110414 632408 110420 632460
rect 110472 632448 110478 632460
rect 113818 632448 113824 632460
rect 110472 632420 113824 632448
rect 110472 632408 110478 632420
rect 113818 632408 113824 632420
rect 113876 632408 113882 632460
rect 282914 630640 282920 630692
rect 282972 630680 282978 630692
rect 283190 630680 283196 630692
rect 282972 630652 283196 630680
rect 282972 630640 282978 630652
rect 283190 630640 283196 630652
rect 283248 630640 283254 630692
rect 105538 629280 105544 629332
rect 105596 629320 105602 629332
rect 110414 629320 110420 629332
rect 105596 629292 110420 629320
rect 105596 629280 105602 629292
rect 110414 629280 110420 629292
rect 110472 629280 110478 629332
rect 219158 627920 219164 627972
rect 219216 627960 219222 627972
rect 219342 627960 219348 627972
rect 219216 627932 219348 627960
rect 219216 627920 219222 627932
rect 219342 627920 219348 627932
rect 219400 627920 219406 627972
rect 41322 627172 41328 627224
rect 41380 627212 41386 627224
rect 312538 627212 312544 627224
rect 41380 627184 312544 627212
rect 41380 627172 41386 627184
rect 312538 627172 312544 627184
rect 312596 627172 312602 627224
rect 278038 626492 278044 626544
rect 278096 626532 278102 626544
rect 279142 626532 279148 626544
rect 278096 626504 279148 626532
rect 278096 626492 278102 626504
rect 279142 626492 279148 626504
rect 279200 626492 279206 626544
rect 95878 621732 95884 621784
rect 95936 621772 95942 621784
rect 105538 621772 105544 621784
rect 95936 621744 105544 621772
rect 95936 621732 95942 621744
rect 105538 621732 105544 621744
rect 105596 621732 105602 621784
rect 24762 621664 24768 621716
rect 24820 621704 24826 621716
rect 283006 621704 283012 621716
rect 24820 621676 283012 621704
rect 24820 621664 24826 621676
rect 283006 621664 283012 621676
rect 283064 621664 283070 621716
rect 219066 620984 219072 621036
rect 219124 621024 219130 621036
rect 219342 621024 219348 621036
rect 219124 620996 219348 621024
rect 219124 620984 219130 620996
rect 219342 620984 219348 620996
rect 219400 620984 219406 621036
rect 23382 619624 23388 619676
rect 23440 619664 23446 619676
rect 84102 619664 84108 619676
rect 23440 619636 84108 619664
rect 23440 619624 23446 619636
rect 84102 619624 84108 619636
rect 84160 619624 84166 619676
rect 219066 618876 219072 618928
rect 219124 618916 219130 618928
rect 284294 618916 284300 618928
rect 219124 618888 284300 618916
rect 219124 618876 219130 618888
rect 284294 618876 284300 618888
rect 284352 618876 284358 618928
rect 31478 617448 31484 617500
rect 31536 617448 31542 617500
rect 91094 617448 91100 617500
rect 91152 617448 91158 617500
rect 28626 616768 28632 616820
rect 28684 616808 28690 616820
rect 31496 616808 31524 617448
rect 28684 616780 31524 616808
rect 28684 616768 28690 616780
rect 28626 616564 28632 616616
rect 28684 616604 28690 616616
rect 30282 616604 30288 616616
rect 28684 616576 30288 616604
rect 28684 616564 28690 616576
rect 30282 616564 30288 616576
rect 30340 616564 30346 616616
rect 28626 616428 28632 616480
rect 28684 616468 28690 616480
rect 30190 616468 30196 616480
rect 28684 616440 30196 616468
rect 28684 616428 28690 616440
rect 30190 616428 30196 616440
rect 30248 616428 30254 616480
rect 28258 615680 28264 615732
rect 28316 615720 28322 615732
rect 91112 615720 91140 617448
rect 453298 616768 453304 616820
rect 453356 616808 453362 616820
rect 456794 616808 456800 616820
rect 453356 616780 456800 616808
rect 453356 616768 453362 616780
rect 456794 616768 456800 616780
rect 456852 616768 456858 616820
rect 551094 616156 551100 616208
rect 551152 616196 551158 616208
rect 551738 616196 551744 616208
rect 551152 616168 551744 616196
rect 551152 616156 551158 616168
rect 551738 616156 551744 616168
rect 551796 616156 551802 616208
rect 28316 615692 91140 615720
rect 28316 615680 28322 615692
rect 282914 611328 282920 611380
rect 282972 611368 282978 611380
rect 283282 611368 283288 611380
rect 282972 611340 283288 611368
rect 282972 611328 282978 611340
rect 283282 611328 283288 611340
rect 283340 611328 283346 611380
rect 3326 609968 3332 610020
rect 3384 610008 3390 610020
rect 11698 610008 11704 610020
rect 3384 609980 11704 610008
rect 3384 609968 3390 609980
rect 11698 609968 11704 609980
rect 11756 609968 11762 610020
rect 554130 609968 554136 610020
rect 554188 610008 554194 610020
rect 555510 610008 555516 610020
rect 554188 609980 555516 610008
rect 554188 609968 554194 609980
rect 555510 609968 555516 609980
rect 555568 609968 555574 610020
rect 551094 606500 551100 606552
rect 551152 606540 551158 606552
rect 551830 606540 551836 606552
rect 551152 606512 551836 606540
rect 551152 606500 551158 606512
rect 551830 606500 551836 606512
rect 551888 606500 551894 606552
rect 23290 605820 23296 605872
rect 23348 605860 23354 605872
rect 25222 605860 25228 605872
rect 23348 605832 25228 605860
rect 23348 605820 23354 605832
rect 25222 605820 25228 605832
rect 25280 605820 25286 605872
rect 24118 603440 24124 603492
rect 24176 603480 24182 603492
rect 28258 603480 28264 603492
rect 24176 603452 28264 603480
rect 24176 603440 24182 603452
rect 28258 603440 28264 603452
rect 28316 603440 28322 603492
rect 551922 603032 551928 603084
rect 551980 603072 551986 603084
rect 552658 603072 552664 603084
rect 551980 603044 552664 603072
rect 551980 603032 551986 603044
rect 552658 603032 552664 603044
rect 552716 603032 552722 603084
rect 551094 596844 551100 596896
rect 551152 596884 551158 596896
rect 551830 596884 551836 596896
rect 551152 596856 551836 596884
rect 551152 596844 551158 596856
rect 551830 596844 551836 596856
rect 551888 596844 551894 596896
rect 551830 596708 551836 596760
rect 551888 596748 551894 596760
rect 552658 596748 552664 596760
rect 551888 596720 552664 596748
rect 551888 596708 551894 596720
rect 552658 596708 552664 596720
rect 552716 596708 552722 596760
rect 3510 594804 3516 594856
rect 3568 594844 3574 594856
rect 9030 594844 9036 594856
rect 3568 594816 9036 594844
rect 3568 594804 3574 594816
rect 9030 594804 9036 594816
rect 9088 594804 9094 594856
rect 139210 594668 139216 594720
rect 139268 594708 139274 594720
rect 139578 594708 139584 594720
rect 139268 594680 139584 594708
rect 139268 594668 139274 594680
rect 139578 594668 139584 594680
rect 139636 594668 139642 594720
rect 28626 594192 28632 594244
rect 28684 594192 28690 594244
rect 28644 594040 28672 594192
rect 28626 593988 28632 594040
rect 28684 593988 28690 594040
rect 282914 591948 282920 592000
rect 282972 591988 282978 592000
rect 283190 591988 283196 592000
rect 282972 591960 283196 591988
rect 282972 591948 282978 591960
rect 283190 591948 283196 591960
rect 283248 591948 283254 592000
rect 554498 590656 554504 590708
rect 554556 590696 554562 590708
rect 555602 590696 555608 590708
rect 554556 590668 555608 590696
rect 554556 590656 554562 590668
rect 555602 590656 555608 590668
rect 555660 590656 555666 590708
rect 554498 589296 554504 589348
rect 554556 589336 554562 589348
rect 556154 589336 556160 589348
rect 554556 589308 556160 589336
rect 554556 589296 554562 589308
rect 556154 589296 556160 589308
rect 556212 589296 556218 589348
rect 554314 587868 554320 587920
rect 554372 587908 554378 587920
rect 557626 587908 557632 587920
rect 554372 587880 557632 587908
rect 554372 587868 554378 587880
rect 557626 587868 557632 587880
rect 557684 587868 557690 587920
rect 28626 587800 28632 587852
rect 28684 587800 28690 587852
rect 28718 587800 28724 587852
rect 28776 587800 28782 587852
rect 28644 587364 28672 587800
rect 28736 587432 28764 587800
rect 28736 587404 28948 587432
rect 28920 587376 28948 587404
rect 28810 587364 28816 587376
rect 28644 587336 28816 587364
rect 28810 587324 28816 587336
rect 28868 587324 28874 587376
rect 28902 587324 28908 587376
rect 28960 587324 28966 587376
rect 551094 587188 551100 587240
rect 551152 587228 551158 587240
rect 551830 587228 551836 587240
rect 551152 587200 551836 587228
rect 551152 587188 551158 587200
rect 551830 587188 551836 587200
rect 551888 587188 551894 587240
rect 554314 586984 554320 587036
rect 554372 587024 554378 587036
rect 556798 587024 556804 587036
rect 554372 586996 556804 587024
rect 554372 586984 554378 586996
rect 556798 586984 556804 586996
rect 556856 586984 556862 587036
rect 28074 586644 28080 586696
rect 28132 586684 28138 586696
rect 28902 586684 28908 586696
rect 28132 586656 28908 586684
rect 28132 586644 28138 586656
rect 28902 586644 28908 586656
rect 28960 586644 28966 586696
rect 28258 585556 28264 585608
rect 28316 585596 28322 585608
rect 28810 585596 28816 585608
rect 28316 585568 28816 585596
rect 28316 585556 28322 585568
rect 28810 585556 28816 585568
rect 28868 585556 28874 585608
rect 554498 585216 554504 585268
rect 554556 585256 554562 585268
rect 558914 585256 558920 585268
rect 554556 585228 558920 585256
rect 554556 585216 554562 585228
rect 558914 585216 558920 585228
rect 558972 585216 558978 585268
rect 554314 585148 554320 585200
rect 554372 585188 554378 585200
rect 560294 585188 560300 585200
rect 554372 585160 560300 585188
rect 554372 585148 554378 585160
rect 560294 585148 560300 585160
rect 560352 585148 560358 585200
rect 28534 583720 28540 583772
rect 28592 583760 28598 583772
rect 28994 583760 29000 583772
rect 28592 583732 29000 583760
rect 28592 583720 28598 583732
rect 28994 583720 29000 583732
rect 29052 583720 29058 583772
rect 554314 583720 554320 583772
rect 554372 583760 554378 583772
rect 561766 583760 561772 583772
rect 554372 583732 561772 583760
rect 554372 583720 554378 583732
rect 561766 583720 561772 583732
rect 561824 583720 561830 583772
rect 283190 582428 283196 582480
rect 283248 582428 283254 582480
rect 283208 582344 283236 582428
rect 283190 582292 283196 582344
rect 283248 582292 283254 582344
rect 554314 581000 554320 581052
rect 554372 581040 554378 581052
rect 563054 581040 563060 581052
rect 554372 581012 563060 581040
rect 554372 581000 554378 581012
rect 563054 581000 563060 581012
rect 563112 581000 563118 581052
rect 554314 579640 554320 579692
rect 554372 579680 554378 579692
rect 564434 579680 564440 579692
rect 554372 579652 564440 579680
rect 554372 579640 554378 579652
rect 564434 579640 564440 579652
rect 564492 579640 564498 579692
rect 26142 579164 26148 579216
rect 26200 579204 26206 579216
rect 28902 579204 28908 579216
rect 26200 579176 28908 579204
rect 26200 579164 26206 579176
rect 28902 579164 28908 579176
rect 28960 579164 28966 579216
rect 28534 578892 28540 578944
rect 28592 578932 28598 578944
rect 28718 578932 28724 578944
rect 28592 578904 28724 578932
rect 28592 578892 28598 578904
rect 28718 578892 28724 578904
rect 28776 578892 28782 578944
rect 28350 578756 28356 578808
rect 28408 578796 28414 578808
rect 28534 578796 28540 578808
rect 28408 578768 28540 578796
rect 28408 578756 28414 578768
rect 28534 578756 28540 578768
rect 28592 578756 28598 578808
rect 554314 578212 554320 578264
rect 554372 578252 554378 578264
rect 565814 578252 565820 578264
rect 554372 578224 565820 578252
rect 554372 578212 554378 578224
rect 565814 578212 565820 578224
rect 565872 578212 565878 578264
rect 551094 577532 551100 577584
rect 551152 577572 551158 577584
rect 551830 577572 551836 577584
rect 551152 577544 551836 577572
rect 551152 577532 551158 577544
rect 551830 577532 551836 577544
rect 551888 577532 551894 577584
rect 554314 576852 554320 576904
rect 554372 576892 554378 576904
rect 567286 576892 567292 576904
rect 554372 576864 567292 576892
rect 554372 576852 554378 576864
rect 567286 576852 567292 576864
rect 567344 576852 567350 576904
rect 28258 575560 28264 575612
rect 28316 575600 28322 575612
rect 28902 575600 28908 575612
rect 28316 575572 28908 575600
rect 28316 575560 28322 575572
rect 28902 575560 28908 575572
rect 28960 575560 28966 575612
rect 554406 575492 554412 575544
rect 554464 575532 554470 575544
rect 560938 575532 560944 575544
rect 554464 575504 560944 575532
rect 554464 575492 554470 575504
rect 560938 575492 560944 575504
rect 560996 575492 561002 575544
rect 554314 574132 554320 574184
rect 554372 574172 554378 574184
rect 568574 574172 568580 574184
rect 554372 574144 568580 574172
rect 554372 574132 554378 574144
rect 568574 574132 568580 574144
rect 568632 574132 568638 574184
rect 554406 574064 554412 574116
rect 554464 574104 554470 574116
rect 569954 574104 569960 574116
rect 554464 574076 569960 574104
rect 554464 574064 554470 574076
rect 569954 574064 569960 574076
rect 570012 574064 570018 574116
rect 29178 573452 29184 573504
rect 29236 573492 29242 573504
rect 29454 573492 29460 573504
rect 29236 573464 29460 573492
rect 29236 573452 29242 573464
rect 29454 573452 29460 573464
rect 29512 573452 29518 573504
rect 30282 573452 30288 573504
rect 30340 573492 30346 573504
rect 30340 573464 30420 573492
rect 30340 573452 30346 573464
rect 29546 573384 29552 573436
rect 29604 573424 29610 573436
rect 30392 573424 30420 573464
rect 29604 573396 30420 573424
rect 29604 573384 29610 573396
rect 28718 573248 28724 573300
rect 28776 573288 28782 573300
rect 30282 573288 30288 573300
rect 28776 573260 30288 573288
rect 28776 573248 28782 573260
rect 30282 573248 30288 573260
rect 30340 573248 30346 573300
rect 29546 572704 29552 572756
rect 29604 572744 29610 572756
rect 29730 572744 29736 572756
rect 29604 572716 29736 572744
rect 29604 572704 29610 572716
rect 29730 572704 29736 572716
rect 29788 572704 29794 572756
rect 283190 572704 283196 572756
rect 283248 572704 283254 572756
rect 554406 572704 554412 572756
rect 554464 572744 554470 572756
rect 571426 572744 571432 572756
rect 554464 572716 571432 572744
rect 554464 572704 554470 572716
rect 571426 572704 571432 572716
rect 571484 572704 571490 572756
rect 283208 572620 283236 572704
rect 551094 572636 551100 572688
rect 551152 572676 551158 572688
rect 551830 572676 551836 572688
rect 551152 572648 551836 572676
rect 551152 572636 551158 572648
rect 551830 572636 551836 572648
rect 551888 572636 551894 572688
rect 283190 572568 283196 572620
rect 283248 572568 283254 572620
rect 199286 572500 199292 572552
rect 199344 572540 199350 572552
rect 204254 572540 204260 572552
rect 199344 572512 204260 572540
rect 199344 572500 199350 572512
rect 204254 572500 204260 572512
rect 204312 572500 204318 572552
rect 198090 572364 198096 572416
rect 198148 572404 198154 572416
rect 202966 572404 202972 572416
rect 198148 572376 202972 572404
rect 198148 572364 198154 572376
rect 202966 572364 202972 572376
rect 203024 572364 203030 572416
rect 189534 572296 189540 572348
rect 189592 572336 189598 572348
rect 195974 572336 195980 572348
rect 189592 572308 195980 572336
rect 189592 572296 189598 572308
rect 195974 572296 195980 572308
rect 196032 572296 196038 572348
rect 196802 572296 196808 572348
rect 196860 572336 196866 572348
rect 202874 572336 202880 572348
rect 196860 572308 202880 572336
rect 196860 572296 196866 572308
rect 202874 572296 202880 572308
rect 202932 572296 202938 572348
rect 188338 572228 188344 572280
rect 188396 572268 188402 572280
rect 194594 572268 194600 572280
rect 188396 572240 194600 572268
rect 188396 572228 188402 572240
rect 194594 572228 194600 572240
rect 194652 572228 194658 572280
rect 206646 572160 206652 572212
rect 206704 572200 206710 572212
rect 211154 572200 211160 572212
rect 206704 572172 211160 572200
rect 206704 572160 206710 572172
rect 211154 572160 211160 572172
rect 211212 572160 211218 572212
rect 25130 572092 25136 572144
rect 25188 572132 25194 572144
rect 25188 572104 38700 572132
rect 25188 572092 25194 572104
rect 38672 571996 38700 572104
rect 195606 572092 195612 572144
rect 195664 572132 195670 572144
rect 201494 572132 201500 572144
rect 195664 572104 201500 572132
rect 195664 572092 195670 572104
rect 201494 572092 201500 572104
rect 201552 572092 201558 572144
rect 218882 572092 218888 572144
rect 218940 572132 218946 572144
rect 222194 572132 222200 572144
rect 218940 572104 222200 572132
rect 218940 572092 218946 572104
rect 222194 572092 222200 572104
rect 222252 572092 222258 572144
rect 277302 572092 277308 572144
rect 277360 572132 277366 572144
rect 279326 572132 279332 572144
rect 277360 572104 279332 572132
rect 277360 572092 277366 572104
rect 279326 572092 279332 572104
rect 279384 572092 279390 572144
rect 190270 572024 190276 572076
rect 190328 572064 190334 572076
rect 197354 572064 197360 572076
rect 190328 572036 197360 572064
rect 190328 572024 190334 572036
rect 197354 572024 197360 572036
rect 197412 572024 197418 572076
rect 207842 572024 207848 572076
rect 207900 572064 207906 572076
rect 212534 572064 212540 572076
rect 207900 572036 212540 572064
rect 207900 572024 207906 572036
rect 212534 572024 212540 572036
rect 212592 572024 212598 572076
rect 227438 572024 227444 572076
rect 227496 572064 227502 572076
rect 229094 572064 229100 572076
rect 227496 572036 229100 572064
rect 227496 572024 227502 572036
rect 229094 572024 229100 572036
rect 229152 572024 229158 572076
rect 267642 572024 267648 572076
rect 267700 572064 267706 572076
rect 268286 572064 268292 572076
rect 267700 572036 268292 572064
rect 267700 572024 267706 572036
rect 268286 572024 268292 572036
rect 268344 572024 268350 572076
rect 275922 572024 275928 572076
rect 275980 572064 275986 572076
rect 278038 572064 278044 572076
rect 275980 572036 278044 572064
rect 275980 572024 275986 572036
rect 278038 572024 278044 572036
rect 278096 572024 278102 572076
rect 38672 571968 41552 571996
rect 26786 571616 26792 571668
rect 26844 571656 26850 571668
rect 31846 571656 31852 571668
rect 26844 571628 31852 571656
rect 26844 571616 26850 571628
rect 31846 571616 31852 571628
rect 31904 571616 31910 571668
rect 26694 571548 26700 571600
rect 26752 571588 26758 571600
rect 33134 571588 33140 571600
rect 26752 571560 33140 571588
rect 26752 571548 26758 571560
rect 33134 571548 33140 571560
rect 33192 571548 33198 571600
rect 41414 571548 41420 571600
rect 41472 571588 41478 571600
rect 41524 571588 41552 571968
rect 209038 571956 209044 572008
rect 209096 571996 209102 572008
rect 214006 571996 214012 572008
rect 209096 571968 214012 571996
rect 209096 571956 209102 571968
rect 214006 571956 214012 571968
rect 214064 571956 214070 572008
rect 194410 571888 194416 571940
rect 194468 571928 194474 571940
rect 200114 571928 200120 571940
rect 194468 571900 200120 571928
rect 194468 571888 194474 571900
rect 200114 571888 200120 571900
rect 200172 571888 200178 571940
rect 216398 571888 216404 571940
rect 216456 571928 216462 571940
rect 219434 571928 219440 571940
rect 216456 571900 219440 571928
rect 216456 571888 216462 571900
rect 219434 571888 219440 571900
rect 219492 571888 219498 571940
rect 205358 571616 205364 571668
rect 205416 571656 205422 571668
rect 209774 571656 209780 571668
rect 205416 571628 209780 571656
rect 205416 571616 205422 571628
rect 209774 571616 209780 571628
rect 209832 571616 209838 571668
rect 217594 571616 217600 571668
rect 217652 571656 217658 571668
rect 220814 571656 220820 571668
rect 217652 571628 220820 571656
rect 217652 571616 217658 571628
rect 220814 571616 220820 571628
rect 220872 571616 220878 571668
rect 228634 571616 228640 571668
rect 228692 571656 228698 571668
rect 230474 571656 230480 571668
rect 228692 571628 230480 571656
rect 228692 571616 228698 571628
rect 230474 571616 230480 571628
rect 230532 571616 230538 571668
rect 41472 571560 41552 571588
rect 41472 571548 41478 571560
rect 202782 571548 202788 571600
rect 202840 571588 202846 571600
rect 208394 571588 208400 571600
rect 202840 571560 208400 571588
rect 202840 571548 202846 571560
rect 208394 571548 208400 571560
rect 208452 571548 208458 571600
rect 213822 571548 213828 571600
rect 213880 571588 213886 571600
rect 218054 571588 218060 571600
rect 213880 571560 218060 571588
rect 213880 571548 213886 571560
rect 218054 571548 218060 571560
rect 218112 571548 218118 571600
rect 220078 571548 220084 571600
rect 220136 571588 220142 571600
rect 223574 571588 223580 571600
rect 220136 571560 223580 571588
rect 220136 571548 220142 571560
rect 223574 571548 223580 571560
rect 223632 571548 223638 571600
rect 224862 571548 224868 571600
rect 224920 571588 224926 571600
rect 227806 571588 227812 571600
rect 224920 571560 227812 571588
rect 224920 571548 224926 571560
rect 227806 571548 227812 571560
rect 227864 571548 227870 571600
rect 26602 571480 26608 571532
rect 26660 571520 26666 571532
rect 26660 571492 30512 571520
rect 26660 571480 26666 571492
rect 28994 571412 29000 571464
rect 29052 571452 29058 571464
rect 30374 571452 30380 571464
rect 29052 571424 30380 571452
rect 29052 571412 29058 571424
rect 30374 571412 30380 571424
rect 30432 571412 30438 571464
rect 30484 571452 30512 571492
rect 201402 571480 201408 571532
rect 201460 571520 201466 571532
rect 207014 571520 207020 571532
rect 201460 571492 207020 571520
rect 201460 571480 201466 571492
rect 207014 571480 207020 571492
rect 207072 571480 207078 571532
rect 212442 571480 212448 571532
rect 212500 571520 212506 571532
rect 216674 571520 216680 571532
rect 212500 571492 216680 571520
rect 212500 571480 212506 571492
rect 216674 571480 216680 571492
rect 216732 571480 216738 571532
rect 223482 571480 223488 571532
rect 223540 571520 223546 571532
rect 226334 571520 226340 571532
rect 223540 571492 226340 571520
rect 223540 571480 223546 571492
rect 226334 571480 226340 571492
rect 226392 571480 226398 571532
rect 231026 571480 231032 571532
rect 231084 571520 231090 571532
rect 233326 571520 233332 571532
rect 231084 571492 233332 571520
rect 231084 571480 231090 571492
rect 233326 571480 233332 571492
rect 233384 571480 233390 571532
rect 273162 571480 273168 571532
rect 273220 571520 273226 571532
rect 275646 571520 275652 571532
rect 273220 571492 275652 571520
rect 273220 571480 273226 571492
rect 275646 571480 275652 571492
rect 275704 571480 275710 571532
rect 37274 571452 37280 571464
rect 30484 571424 37280 571452
rect 37274 571412 37280 571424
rect 37332 571412 37338 571464
rect 191742 571412 191748 571464
rect 191800 571452 191806 571464
rect 198826 571452 198832 571464
rect 191800 571424 198832 571452
rect 191800 571412 191806 571424
rect 198826 571412 198832 571424
rect 198884 571412 198890 571464
rect 200482 571412 200488 571464
rect 200540 571452 200546 571464
rect 205634 571452 205640 571464
rect 200540 571424 205640 571452
rect 200540 571412 200546 571424
rect 205634 571412 205640 571424
rect 205692 571412 205698 571464
rect 211522 571412 211528 571464
rect 211580 571452 211586 571464
rect 215294 571452 215300 571464
rect 211580 571424 215300 571452
rect 211580 571412 211586 571424
rect 215294 571412 215300 571424
rect 215352 571412 215358 571464
rect 222102 571412 222108 571464
rect 222160 571452 222166 571464
rect 224954 571452 224960 571464
rect 222160 571424 224960 571452
rect 222160 571412 222166 571424
rect 224954 571412 224960 571424
rect 225012 571412 225018 571464
rect 233142 571412 233148 571464
rect 233200 571452 233206 571464
rect 234614 571452 234620 571464
rect 233200 571424 234620 571452
rect 233200 571412 233206 571424
rect 234614 571412 234620 571424
rect 234672 571412 234678 571464
rect 235902 571412 235908 571464
rect 235960 571452 235966 571464
rect 235960 571424 237420 571452
rect 235960 571412 235966 571424
rect 23198 571344 23204 571396
rect 23256 571384 23262 571396
rect 25590 571384 25596 571396
rect 23256 571356 25596 571384
rect 23256 571344 23262 571356
rect 25590 571344 25596 571356
rect 25648 571344 25654 571396
rect 193122 571344 193128 571396
rect 193180 571384 193186 571396
rect 198734 571384 198740 571396
rect 193180 571356 198740 571384
rect 193180 571344 193186 571356
rect 198734 571344 198740 571356
rect 198792 571344 198798 571396
rect 204162 571344 204168 571396
rect 204220 571384 204226 571396
rect 208486 571384 208492 571396
rect 204220 571356 208492 571384
rect 204220 571344 204226 571356
rect 208486 571344 208492 571356
rect 208544 571344 208550 571396
rect 210326 571344 210332 571396
rect 210384 571384 210390 571396
rect 213914 571384 213920 571396
rect 210384 571356 213920 571384
rect 210384 571344 210390 571356
rect 213914 571344 213920 571356
rect 213972 571344 213978 571396
rect 215202 571344 215208 571396
rect 215260 571384 215266 571396
rect 218146 571384 218152 571396
rect 215260 571356 218152 571384
rect 215260 571344 215266 571356
rect 218146 571344 218152 571356
rect 218204 571344 218210 571396
rect 221274 571344 221280 571396
rect 221332 571384 221338 571396
rect 223666 571384 223672 571396
rect 221332 571356 223672 571384
rect 221332 571344 221338 571356
rect 223666 571344 223672 571356
rect 223724 571344 223730 571396
rect 226150 571344 226156 571396
rect 226208 571384 226214 571396
rect 227714 571384 227720 571396
rect 226208 571356 227720 571384
rect 226208 571344 226214 571356
rect 227714 571344 227720 571356
rect 227772 571344 227778 571396
rect 229830 571344 229836 571396
rect 229888 571384 229894 571396
rect 231854 571384 231860 571396
rect 229888 571356 231860 571384
rect 229888 571344 229894 571356
rect 231854 571344 231860 571356
rect 231912 571344 231918 571396
rect 232314 571344 232320 571396
rect 232372 571384 232378 571396
rect 233234 571384 233240 571396
rect 232372 571356 233240 571384
rect 232372 571344 232378 571356
rect 233234 571344 233240 571356
rect 233292 571344 233298 571396
rect 234522 571344 234528 571396
rect 234580 571384 234586 571396
rect 235994 571384 236000 571396
rect 234580 571356 236000 571384
rect 234580 571344 234586 571356
rect 235994 571344 236000 571356
rect 236052 571344 236058 571396
rect 237392 571328 237420 571424
rect 268930 571412 268936 571464
rect 268988 571452 268994 571464
rect 270770 571452 270776 571464
rect 268988 571424 270776 571452
rect 268988 571412 268994 571424
rect 270770 571412 270776 571424
rect 270828 571412 270834 571464
rect 271782 571412 271788 571464
rect 271840 571452 271846 571464
rect 273254 571452 273260 571464
rect 271840 571424 273260 571452
rect 271840 571412 271846 571424
rect 273254 571412 273260 571424
rect 273312 571412 273318 571464
rect 274542 571412 274548 571464
rect 274600 571452 274606 571464
rect 276842 571452 276848 571464
rect 274600 571424 276848 571452
rect 274600 571412 274606 571424
rect 276842 571412 276848 571424
rect 276900 571412 276906 571464
rect 278590 571412 278596 571464
rect 278648 571452 278654 571464
rect 281718 571452 281724 571464
rect 278648 571424 281724 571452
rect 278648 571412 278654 571424
rect 281718 571412 281724 571424
rect 281776 571412 281782 571464
rect 239582 571344 239588 571396
rect 239640 571384 239646 571396
rect 240134 571384 240140 571396
rect 239640 571356 240140 571384
rect 239640 571344 239646 571356
rect 240134 571344 240140 571356
rect 240192 571344 240198 571396
rect 240870 571344 240876 571396
rect 240928 571384 240934 571396
rect 241514 571384 241520 571396
rect 240928 571356 241520 571384
rect 240928 571344 240934 571356
rect 241514 571344 241520 571356
rect 241572 571344 241578 571396
rect 242066 571344 242072 571396
rect 242124 571384 242130 571396
rect 242986 571384 242992 571396
rect 242124 571356 242992 571384
rect 242124 571344 242130 571356
rect 242986 571344 242992 571356
rect 243044 571344 243050 571396
rect 254854 571384 254860 571396
rect 253952 571356 254860 571384
rect 253952 571328 253980 571356
rect 254854 571344 254860 571356
rect 254912 571344 254918 571396
rect 255314 571344 255320 571396
rect 255372 571384 255378 571396
rect 256050 571384 256056 571396
rect 255372 571356 256056 571384
rect 255372 571344 255378 571356
rect 256050 571344 256056 571356
rect 256108 571344 256114 571396
rect 256694 571344 256700 571396
rect 256752 571384 256758 571396
rect 257338 571384 257344 571396
rect 256752 571356 257344 571384
rect 256752 571344 256758 571356
rect 257338 571344 257344 571356
rect 257396 571344 257402 571396
rect 264606 571384 264612 571396
rect 263520 571356 264612 571384
rect 263520 571328 263548 571356
rect 264606 571344 264612 571356
rect 264664 571344 264670 571396
rect 264882 571344 264888 571396
rect 264940 571384 264946 571396
rect 265894 571384 265900 571396
rect 264940 571356 265900 571384
rect 264940 571344 264946 571356
rect 265894 571344 265900 571356
rect 265952 571344 265958 571396
rect 266262 571344 266268 571396
rect 266320 571384 266326 571396
rect 267090 571384 267096 571396
rect 266320 571356 267096 571384
rect 266320 571344 266326 571356
rect 267090 571344 267096 571356
rect 267148 571344 267154 571396
rect 269022 571344 269028 571396
rect 269080 571384 269086 571396
rect 269482 571384 269488 571396
rect 269080 571356 269488 571384
rect 269080 571344 269086 571356
rect 269482 571344 269488 571356
rect 269540 571344 269546 571396
rect 270402 571344 270408 571396
rect 270460 571384 270466 571396
rect 271966 571384 271972 571396
rect 270460 571356 271972 571384
rect 270460 571344 270466 571356
rect 271966 571344 271972 571356
rect 272024 571344 272030 571396
rect 273070 571344 273076 571396
rect 273128 571384 273134 571396
rect 274634 571384 274640 571396
rect 273128 571356 274640 571384
rect 273128 571344 273134 571356
rect 274634 571344 274640 571356
rect 274692 571344 274698 571396
rect 278682 571344 278688 571396
rect 278740 571384 278746 571396
rect 280522 571384 280528 571396
rect 278740 571356 280528 571384
rect 278740 571344 278746 571356
rect 280522 571344 280528 571356
rect 280580 571344 280586 571396
rect 554222 571344 554228 571396
rect 554280 571384 554286 571396
rect 558178 571384 558184 571396
rect 554280 571356 558184 571384
rect 554280 571344 554286 571356
rect 558178 571344 558184 571356
rect 558236 571344 558242 571396
rect 237374 571276 237380 571328
rect 237432 571276 237438 571328
rect 253934 571276 253940 571328
rect 253992 571276 253998 571328
rect 263502 571276 263508 571328
rect 263560 571276 263566 571328
rect 551922 571208 551928 571260
rect 551980 571248 551986 571260
rect 554590 571248 554596 571260
rect 551980 571220 554596 571248
rect 551980 571208 551986 571220
rect 554590 571208 554596 571220
rect 554648 571208 554654 571260
rect 28626 570800 28632 570852
rect 28684 570840 28690 570852
rect 45646 570840 45652 570852
rect 28684 570812 45652 570840
rect 28684 570800 28690 570812
rect 45646 570800 45652 570812
rect 45704 570800 45710 570852
rect 29178 570732 29184 570784
rect 29236 570772 29242 570784
rect 48314 570772 48320 570784
rect 29236 570744 48320 570772
rect 29236 570732 29242 570744
rect 48314 570732 48320 570744
rect 48372 570732 48378 570784
rect 29454 570664 29460 570716
rect 29512 570704 29518 570716
rect 52454 570704 52460 570716
rect 29512 570676 52460 570704
rect 29512 570664 29518 570676
rect 52454 570664 52460 570676
rect 52512 570664 52518 570716
rect 248414 570664 248420 570716
rect 248472 570704 248478 570716
rect 554314 570704 554320 570716
rect 248472 570676 248552 570704
rect 248472 570664 248478 570676
rect 28534 570596 28540 570648
rect 28592 570636 28598 570648
rect 53834 570636 53840 570648
rect 28592 570608 53840 570636
rect 28592 570596 28598 570608
rect 53834 570596 53840 570608
rect 53892 570596 53898 570648
rect 248524 570512 248552 570676
rect 550560 570676 554320 570704
rect 550560 570636 550588 570676
rect 554314 570664 554320 570676
rect 554372 570664 554378 570716
rect 525720 570608 550588 570636
rect 525720 570512 525748 570608
rect 248506 570460 248512 570512
rect 248564 570460 248570 570512
rect 525702 570460 525708 570512
rect 525760 570460 525766 570512
rect 543642 570392 543648 570444
rect 543700 570432 543706 570444
rect 554498 570432 554504 570444
rect 543700 570404 554504 570432
rect 543700 570392 543706 570404
rect 554498 570392 554504 570404
rect 554556 570392 554562 570444
rect 318518 569916 318524 569968
rect 318576 569956 318582 569968
rect 318702 569956 318708 569968
rect 318576 569928 318708 569956
rect 318576 569916 318582 569928
rect 318702 569916 318708 569928
rect 318760 569916 318766 569968
rect 354398 569916 354404 569968
rect 354456 569956 354462 569968
rect 354582 569956 354588 569968
rect 354456 569928 354588 569956
rect 354456 569916 354462 569928
rect 354582 569916 354588 569928
rect 354640 569916 354646 569968
rect 547782 569916 547788 569968
rect 547840 569956 547846 569968
rect 552934 569956 552940 569968
rect 547840 569928 552940 569956
rect 547840 569916 547846 569928
rect 552934 569916 552940 569928
rect 552992 569916 552998 569968
rect 554406 569916 554412 569968
rect 554464 569956 554470 569968
rect 572714 569956 572720 569968
rect 554464 569928 572720 569956
rect 554464 569916 554470 569928
rect 572714 569916 572720 569928
rect 572772 569916 572778 569968
rect 29178 569848 29184 569900
rect 29236 569888 29242 569900
rect 29730 569888 29736 569900
rect 29236 569860 29736 569888
rect 29236 569848 29242 569860
rect 29730 569848 29736 569860
rect 29788 569848 29794 569900
rect 112530 569848 112536 569900
rect 112588 569888 112594 569900
rect 138658 569888 138664 569900
rect 112588 569860 138664 569888
rect 112588 569848 112594 569860
rect 138658 569848 138664 569860
rect 138716 569848 138722 569900
rect 281534 569848 281540 569900
rect 281592 569888 281598 569900
rect 284386 569888 284392 569900
rect 281592 569860 284392 569888
rect 281592 569848 281598 569860
rect 284386 569848 284392 569860
rect 284444 569848 284450 569900
rect 28442 569304 28448 569356
rect 28500 569344 28506 569356
rect 71774 569344 71780 569356
rect 28500 569316 71780 569344
rect 28500 569304 28506 569316
rect 71774 569304 71780 569316
rect 71832 569304 71838 569356
rect 25774 569236 25780 569288
rect 25832 569276 25838 569288
rect 70394 569276 70400 569288
rect 25832 569248 70400 569276
rect 25832 569236 25838 569248
rect 70394 569236 70400 569248
rect 70452 569236 70458 569288
rect 56410 569168 56416 569220
rect 56468 569208 56474 569220
rect 281534 569208 281540 569220
rect 56468 569180 281540 569208
rect 56468 569168 56474 569180
rect 281534 569168 281540 569180
rect 281592 569168 281598 569220
rect 286318 569168 286324 569220
rect 286376 569208 286382 569220
rect 580534 569208 580540 569220
rect 286376 569180 580540 569208
rect 286376 569168 286382 569180
rect 580534 569168 580540 569180
rect 580592 569168 580598 569220
rect 549162 568556 549168 568608
rect 549220 568596 549226 568608
rect 553026 568596 553032 568608
rect 549220 568568 553032 568596
rect 549220 568556 549226 568568
rect 553026 568556 553032 568568
rect 553084 568556 553090 568608
rect 338298 568488 338304 568540
rect 338356 568528 338362 568540
rect 339310 568528 339316 568540
rect 338356 568500 339316 568528
rect 338356 568488 338362 568500
rect 339310 568488 339316 568500
rect 339368 568488 339374 568540
rect 340138 568488 340144 568540
rect 340196 568528 340202 568540
rect 385034 568528 385040 568540
rect 340196 568500 385040 568528
rect 340196 568488 340202 568500
rect 385034 568488 385040 568500
rect 385092 568488 385098 568540
rect 456058 568488 456064 568540
rect 456116 568528 456122 568540
rect 483658 568528 483664 568540
rect 456116 568500 483664 568528
rect 456116 568488 456122 568500
rect 483658 568488 483664 568500
rect 483716 568488 483722 568540
rect 336550 568420 336556 568472
rect 336608 568460 336614 568472
rect 387886 568460 387892 568472
rect 336608 568432 387892 568460
rect 336608 568420 336614 568432
rect 387886 568420 387892 568432
rect 387944 568420 387950 568472
rect 327534 568352 327540 568404
rect 327592 568392 327598 568404
rect 328270 568392 328276 568404
rect 327592 568364 328276 568392
rect 327592 568352 327598 568364
rect 328270 568352 328276 568364
rect 328328 568352 328334 568404
rect 332962 568352 332968 568404
rect 333020 568392 333026 568404
rect 389358 568392 389364 568404
rect 333020 568364 389364 568392
rect 333020 568352 333026 568364
rect 389358 568352 389364 568364
rect 389416 568352 389422 568404
rect 329374 568284 329380 568336
rect 329432 568324 329438 568336
rect 391934 568324 391940 568336
rect 329432 568296 391940 568324
rect 329432 568284 329438 568296
rect 391934 568284 391940 568296
rect 391992 568284 391998 568336
rect 325786 568216 325792 568268
rect 325844 568256 325850 568268
rect 394694 568256 394700 568268
rect 325844 568228 394700 568256
rect 325844 568216 325850 568228
rect 394694 568216 394700 568228
rect 394752 568216 394758 568268
rect 336642 568148 336648 568200
rect 336700 568188 336706 568200
rect 422570 568188 422576 568200
rect 336700 568160 422576 568188
rect 336700 568148 336706 568160
rect 422570 568148 422576 568160
rect 422628 568148 422634 568200
rect 335262 568080 335268 568132
rect 335320 568120 335326 568132
rect 426158 568120 426164 568132
rect 335320 568092 426164 568120
rect 335320 568080 335326 568092
rect 426158 568080 426164 568092
rect 426216 568080 426222 568132
rect 332502 568012 332508 568064
rect 332560 568052 332566 568064
rect 429746 568052 429752 568064
rect 332560 568024 429752 568052
rect 332560 568012 332566 568024
rect 429746 568012 429752 568024
rect 429804 568012 429810 568064
rect 331122 567944 331128 567996
rect 331180 567984 331186 567996
rect 433334 567984 433340 567996
rect 331180 567956 433340 567984
rect 331180 567944 331186 567956
rect 433334 567944 433340 567956
rect 433392 567944 433398 567996
rect 328362 567876 328368 567928
rect 328420 567916 328426 567928
rect 436922 567916 436928 567928
rect 328420 567888 436928 567916
rect 328420 567876 328426 567888
rect 436922 567876 436928 567888
rect 436980 567876 436986 567928
rect 326982 567808 326988 567860
rect 327040 567848 327046 567860
rect 440510 567848 440516 567860
rect 327040 567820 440516 567848
rect 327040 567808 327046 567820
rect 440510 567808 440516 567820
rect 440568 567808 440574 567860
rect 343726 567740 343732 567792
rect 343784 567780 343790 567792
rect 383746 567780 383752 567792
rect 343784 567752 383752 567780
rect 343784 567740 343790 567752
rect 383746 567740 383752 567752
rect 383804 567740 383810 567792
rect 345474 567672 345480 567724
rect 345532 567712 345538 567724
rect 346302 567712 346308 567724
rect 345532 567684 346308 567712
rect 345532 567672 345538 567684
rect 346302 567672 346308 567684
rect 346360 567672 346366 567724
rect 347314 567672 347320 567724
rect 347372 567712 347378 567724
rect 380894 567712 380900 567724
rect 347372 567684 380900 567712
rect 347372 567672 347378 567684
rect 380894 567672 380900 567684
rect 380952 567672 380958 567724
rect 29086 567604 29092 567656
rect 29144 567644 29150 567656
rect 29454 567644 29460 567656
rect 29144 567616 29460 567644
rect 29144 567604 29150 567616
rect 29454 567604 29460 567616
rect 29512 567604 29518 567656
rect 350902 567604 350908 567656
rect 350960 567644 350966 567656
rect 379514 567644 379520 567656
rect 350960 567616 379520 567644
rect 350960 567604 350966 567616
rect 379514 567604 379520 567616
rect 379572 567604 379578 567656
rect 361666 567536 361672 567588
rect 361724 567576 361730 567588
rect 362862 567576 362868 567588
rect 361724 567548 362868 567576
rect 361724 567536 361730 567548
rect 362862 567536 362868 567548
rect 362920 567536 362926 567588
rect 363414 567536 363420 567588
rect 363472 567576 363478 567588
rect 364242 567576 364248 567588
rect 363472 567548 364248 567576
rect 363472 567536 363478 567548
rect 364242 567536 364248 567548
rect 364300 567536 364306 567588
rect 3510 567196 3516 567248
rect 3568 567236 3574 567248
rect 9122 567236 9128 567248
rect 3568 567208 9128 567236
rect 3568 567196 3574 567208
rect 9122 567196 9128 567208
rect 9180 567196 9186 567248
rect 320358 567196 320364 567248
rect 320416 567236 320422 567248
rect 321462 567236 321468 567248
rect 320416 567208 321468 567236
rect 320416 567196 320422 567208
rect 321462 567196 321468 567208
rect 321520 567196 321526 567248
rect 356238 567196 356244 567248
rect 356296 567236 356302 567248
rect 357342 567236 357348 567248
rect 356296 567208 357348 567236
rect 356296 567196 356302 567208
rect 357342 567196 357348 567208
rect 357400 567196 357406 567248
rect 529014 567196 529020 567248
rect 529072 567236 529078 567248
rect 530578 567236 530584 567248
rect 529072 567208 530584 567236
rect 529072 567196 529078 567208
rect 530578 567196 530584 567208
rect 530636 567196 530642 567248
rect 355870 566448 355876 566500
rect 355928 566488 355934 566500
rect 389174 566488 389180 566500
rect 355928 566460 389180 566488
rect 355928 566448 355934 566460
rect 389174 566448 389180 566460
rect 389232 566448 389238 566500
rect 29270 565700 29276 565752
rect 29328 565740 29334 565752
rect 30006 565740 30012 565752
rect 29328 565712 30012 565740
rect 29328 565700 29334 565712
rect 30006 565700 30012 565712
rect 30064 565700 30070 565752
rect 339402 565088 339408 565140
rect 339460 565128 339466 565140
rect 418154 565128 418160 565140
rect 339460 565100 418160 565128
rect 339460 565088 339466 565100
rect 418154 565088 418160 565100
rect 418212 565088 418218 565140
rect 532602 565088 532608 565140
rect 532660 565128 532666 565140
rect 554774 565128 554780 565140
rect 532660 565100 554780 565128
rect 532660 565088 532666 565100
rect 554774 565088 554780 565100
rect 554832 565088 554838 565140
rect 342070 563660 342076 563712
rect 342128 563700 342134 563712
rect 415394 563700 415400 563712
rect 342128 563672 415400 563700
rect 342128 563660 342134 563672
rect 415394 563660 415400 563672
rect 415452 563660 415458 563712
rect 528462 563660 528468 563712
rect 528520 563700 528526 563712
rect 555142 563700 555148 563712
rect 528520 563672 555148 563700
rect 528520 563660 528526 563672
rect 555142 563660 555148 563672
rect 555200 563660 555206 563712
rect 29546 563184 29552 563236
rect 29604 563224 29610 563236
rect 30282 563224 30288 563236
rect 29604 563196 30288 563224
rect 29604 563184 29610 563196
rect 30282 563184 30288 563196
rect 30340 563184 30346 563236
rect 551094 563048 551100 563100
rect 551152 563088 551158 563100
rect 551830 563088 551836 563100
rect 551152 563060 551836 563088
rect 551152 563048 551158 563060
rect 551830 563048 551836 563060
rect 551888 563048 551894 563100
rect 346210 562300 346216 562352
rect 346268 562340 346274 562352
rect 407114 562340 407120 562352
rect 346268 562312 407120 562340
rect 346268 562300 346274 562312
rect 407114 562300 407120 562312
rect 407172 562300 407178 562352
rect 538122 562300 538128 562352
rect 538180 562340 538186 562352
rect 555510 562340 555516 562352
rect 538180 562312 555516 562340
rect 538180 562300 538186 562312
rect 555510 562300 555516 562312
rect 555568 562300 555574 562352
rect 347682 560940 347688 560992
rect 347740 560980 347746 560992
rect 404354 560980 404360 560992
rect 347740 560952 404360 560980
rect 347740 560940 347746 560952
rect 404354 560940 404360 560952
rect 404412 560940 404418 560992
rect 533982 560940 533988 560992
rect 534040 560980 534046 560992
rect 555326 560980 555332 560992
rect 534040 560952 555332 560980
rect 534040 560940 534046 560952
rect 555326 560940 555332 560952
rect 555384 560940 555390 560992
rect 29178 560260 29184 560312
rect 29236 560300 29242 560312
rect 29730 560300 29736 560312
rect 29236 560272 29736 560300
rect 29236 560260 29242 560272
rect 29730 560260 29736 560272
rect 29788 560260 29794 560312
rect 350442 559512 350448 559564
rect 350500 559552 350506 559564
rect 400214 559552 400220 559564
rect 350500 559524 400220 559552
rect 350500 559512 350506 559524
rect 400214 559512 400220 559524
rect 400272 559512 400278 559564
rect 529842 559512 529848 559564
rect 529900 559552 529906 559564
rect 555050 559552 555056 559564
rect 529900 559524 555056 559552
rect 529900 559512 529906 559524
rect 555050 559512 555056 559524
rect 555108 559512 555114 559564
rect 283190 558900 283196 558952
rect 283248 558940 283254 558952
rect 283374 558940 283380 558952
rect 283248 558912 283380 558940
rect 283248 558900 283254 558912
rect 283374 558900 283380 558912
rect 283432 558900 283438 558952
rect 29362 558492 29368 558544
rect 29420 558532 29426 558544
rect 29638 558532 29644 558544
rect 29420 558504 29644 558532
rect 29420 558492 29426 558504
rect 29638 558492 29644 558504
rect 29696 558492 29702 558544
rect 29546 558152 29552 558204
rect 29604 558192 29610 558204
rect 30282 558192 30288 558204
rect 29604 558164 30288 558192
rect 29604 558152 29610 558164
rect 30282 558152 30288 558164
rect 30340 558152 30346 558204
rect 351730 558152 351736 558204
rect 351788 558192 351794 558204
rect 397454 558192 397460 558204
rect 351788 558164 397460 558192
rect 351788 558152 351794 558164
rect 397454 558152 397460 558164
rect 397512 558152 397518 558204
rect 483658 556452 483664 556504
rect 483716 556492 483722 556504
rect 485774 556492 485780 556504
rect 483716 556464 485780 556492
rect 483716 556452 483722 556464
rect 485774 556452 485780 556464
rect 485832 556452 485838 556504
rect 304258 556180 304264 556232
rect 304316 556220 304322 556232
rect 579798 556220 579804 556232
rect 304316 556192 579804 556220
rect 304316 556180 304322 556192
rect 579798 556180 579804 556192
rect 579856 556180 579862 556232
rect 354490 555432 354496 555484
rect 354548 555472 354554 555484
rect 393314 555472 393320 555484
rect 354548 555444 393320 555472
rect 354548 555432 354554 555444
rect 393314 555432 393320 555444
rect 393372 555432 393378 555484
rect 358630 554004 358636 554056
rect 358688 554044 358694 554056
rect 386414 554044 386420 554056
rect 358688 554016 386420 554044
rect 358688 554004 358694 554016
rect 386414 554004 386420 554016
rect 386472 554004 386478 554056
rect 485774 554004 485780 554056
rect 485832 554044 485838 554056
rect 498194 554044 498200 554056
rect 485832 554016 498200 554044
rect 485832 554004 485838 554016
rect 498194 554004 498200 554016
rect 498252 554004 498258 554056
rect 29270 553392 29276 553444
rect 29328 553432 29334 553444
rect 30006 553432 30012 553444
rect 29328 553404 30012 553432
rect 29328 553392 29334 553404
rect 30006 553392 30012 553404
rect 30064 553392 30070 553444
rect 283190 553392 283196 553444
rect 283248 553392 283254 553444
rect 551002 553392 551008 553444
rect 551060 553432 551066 553444
rect 551060 553404 551140 553432
rect 551060 553392 551066 553404
rect 283208 553296 283236 553392
rect 551112 553376 551140 553404
rect 551094 553324 551100 553376
rect 551152 553324 551158 553376
rect 283282 553296 283288 553308
rect 283208 553268 283288 553296
rect 283282 553256 283288 553268
rect 283340 553256 283346 553308
rect 324130 552644 324136 552696
rect 324188 552684 324194 552696
rect 442994 552684 443000 552696
rect 324188 552656 443000 552684
rect 324188 552644 324194 552656
rect 442994 552644 443000 552656
rect 443052 552644 443058 552696
rect 540882 552644 540888 552696
rect 540940 552684 540946 552696
rect 555234 552684 555240 552696
rect 540940 552656 555240 552684
rect 540940 552644 540946 552656
rect 555234 552644 555240 552656
rect 555292 552644 555298 552696
rect 3142 552032 3148 552084
rect 3200 552072 3206 552084
rect 312538 552072 312544 552084
rect 3200 552044 312544 552072
rect 3200 552032 3206 552044
rect 312538 552032 312544 552044
rect 312596 552032 312602 552084
rect 329742 551284 329748 551336
rect 329800 551324 329806 551336
rect 434714 551324 434720 551336
rect 329800 551296 434720 551324
rect 329800 551284 329806 551296
rect 434714 551284 434720 551296
rect 434772 551284 434778 551336
rect 498194 551284 498200 551336
rect 498252 551324 498258 551336
rect 504358 551324 504364 551336
rect 498252 551296 504364 551324
rect 498252 551284 498258 551296
rect 504358 551284 504364 551296
rect 504416 551284 504422 551336
rect 536742 551284 536748 551336
rect 536800 551324 536806 551336
rect 554958 551324 554964 551336
rect 536800 551296 554964 551324
rect 536800 551284 536806 551296
rect 554958 551284 554964 551296
rect 555016 551284 555022 551336
rect 29454 550536 29460 550588
rect 29512 550576 29518 550588
rect 29730 550576 29736 550588
rect 29512 550548 29736 550576
rect 29512 550536 29518 550548
rect 29730 550536 29736 550548
rect 29788 550536 29794 550588
rect 332410 549856 332416 549908
rect 332468 549896 332474 549908
rect 430574 549896 430580 549908
rect 332468 549868 430580 549896
rect 332468 549856 332474 549868
rect 430574 549856 430580 549868
rect 430632 549856 430638 549908
rect 551002 549244 551008 549296
rect 551060 549284 551066 549296
rect 551094 549284 551100 549296
rect 551060 549256 551100 549284
rect 551060 549244 551066 549256
rect 551094 549244 551100 549256
rect 551152 549244 551158 549296
rect 333882 548496 333888 548548
rect 333940 548536 333946 548548
rect 427814 548536 427820 548548
rect 333940 548508 427820 548536
rect 333940 548496 333946 548508
rect 427814 548496 427820 548508
rect 427872 548496 427878 548548
rect 549070 547680 549076 547732
rect 549128 547720 549134 547732
rect 552750 547720 552756 547732
rect 549128 547692 552756 547720
rect 549128 547680 549134 547692
rect 552750 547680 552756 547692
rect 552808 547680 552814 547732
rect 26142 547476 26148 547528
rect 26200 547516 26206 547528
rect 35894 547516 35900 547528
rect 26200 547488 35900 547516
rect 26200 547476 26206 547488
rect 35894 547476 35900 547488
rect 35952 547476 35958 547528
rect 26878 547408 26884 547460
rect 26936 547448 26942 547460
rect 46934 547448 46940 547460
rect 26936 547420 46940 547448
rect 26936 547408 26942 547420
rect 46934 547408 46940 547420
rect 46992 547408 46998 547460
rect 26970 547340 26976 547392
rect 27028 547380 27034 547392
rect 55306 547380 55312 547392
rect 27028 547352 55312 547380
rect 27028 547340 27034 547352
rect 55306 547340 55312 547352
rect 55364 547340 55370 547392
rect 28166 547272 28172 547324
rect 28224 547312 28230 547324
rect 62114 547312 62120 547324
rect 28224 547284 62120 547312
rect 28224 547272 28230 547284
rect 62114 547272 62120 547284
rect 62172 547272 62178 547324
rect 27062 547204 27068 547256
rect 27120 547244 27126 547256
rect 64874 547244 64880 547256
rect 27120 547216 64880 547244
rect 27120 547204 27126 547216
rect 64874 547204 64880 547216
rect 64932 547204 64938 547256
rect 531222 547204 531228 547256
rect 531280 547244 531286 547256
rect 551646 547244 551652 547256
rect 531280 547216 551652 547244
rect 531280 547204 531286 547216
rect 551646 547204 551652 547216
rect 551704 547204 551710 547256
rect 27982 547136 27988 547188
rect 28040 547176 28046 547188
rect 80054 547176 80060 547188
rect 28040 547148 80060 547176
rect 28040 547136 28046 547148
rect 80054 547136 80060 547148
rect 80112 547136 80118 547188
rect 336550 547136 336556 547188
rect 336608 547176 336614 547188
rect 423674 547176 423680 547188
rect 336608 547148 423680 547176
rect 336608 547136 336614 547148
rect 423674 547136 423680 547148
rect 423732 547136 423738 547188
rect 527082 547136 527088 547188
rect 527140 547176 527146 547188
rect 551554 547176 551560 547188
rect 527140 547148 551560 547176
rect 527140 547136 527146 547148
rect 551554 547136 551560 547148
rect 551612 547136 551618 547188
rect 550542 547068 550548 547120
rect 550600 547108 550606 547120
rect 552842 547108 552848 547120
rect 550600 547080 552848 547108
rect 550600 547068 550606 547080
rect 552842 547068 552848 547080
rect 552900 547068 552906 547120
rect 366910 545776 366916 545828
rect 366968 545816 366974 545828
rect 373994 545816 374000 545828
rect 366968 545788 374000 545816
rect 366968 545776 366974 545788
rect 373994 545776 374000 545788
rect 374052 545776 374058 545828
rect 322842 545708 322848 545760
rect 322900 545748 322906 545760
rect 396074 545748 396080 545760
rect 322900 545720 396080 545748
rect 322900 545708 322906 545720
rect 396074 545708 396080 545720
rect 396132 545708 396138 545760
rect 326890 544348 326896 544400
rect 326948 544388 326954 544400
rect 437474 544388 437480 544400
rect 326948 544360 437480 544388
rect 326948 544348 326954 544360
rect 437474 544348 437480 544360
rect 437532 544348 437538 544400
rect 283282 543844 283288 543856
rect 283116 543816 283288 543844
rect 283116 543720 283144 543816
rect 283282 543804 283288 543816
rect 283340 543804 283346 543856
rect 368382 543736 368388 543788
rect 368440 543776 368446 543788
rect 369854 543776 369860 543788
rect 368440 543748 369860 543776
rect 368440 543736 368446 543748
rect 369854 543736 369860 543748
rect 369912 543736 369918 543788
rect 29362 543668 29368 543720
rect 29420 543708 29426 543720
rect 30006 543708 30012 543720
rect 29420 543680 30012 543708
rect 29420 543668 29426 543680
rect 30006 543668 30012 543680
rect 30064 543668 30070 543720
rect 283098 543668 283104 543720
rect 283156 543668 283162 543720
rect 367002 543260 367008 543312
rect 367060 543300 367066 543312
rect 369854 543300 369860 543312
rect 367060 543272 369860 543300
rect 367060 543260 367066 543272
rect 369854 543260 369860 543272
rect 369912 543260 369918 543312
rect 324222 542988 324228 543040
rect 324280 543028 324286 543040
rect 394878 543028 394884 543040
rect 324280 543000 394884 543028
rect 324280 542988 324286 543000
rect 394878 542988 394884 543000
rect 394936 542988 394942 543040
rect 364242 541696 364248 541748
rect 364300 541736 364306 541748
rect 371326 541736 371332 541748
rect 364300 541708 371332 541736
rect 364300 541696 364306 541708
rect 371326 541696 371332 541708
rect 371384 541696 371390 541748
rect 325602 541628 325608 541680
rect 325660 541668 325666 541680
rect 441614 541668 441620 541680
rect 325660 541640 441620 541668
rect 325660 541628 325666 541640
rect 441614 541628 441620 541640
rect 441672 541628 441678 541680
rect 29454 540948 29460 541000
rect 29512 540988 29518 541000
rect 29730 540988 29736 541000
rect 29512 540960 29736 540988
rect 29512 540948 29518 540960
rect 29730 540948 29736 540960
rect 29788 540948 29794 541000
rect 360102 540268 360108 540320
rect 360160 540308 360166 540320
rect 373994 540308 374000 540320
rect 360160 540280 374000 540308
rect 360160 540268 360166 540280
rect 373994 540268 374000 540280
rect 374052 540268 374058 540320
rect 343542 540200 343548 540252
rect 343600 540240 343606 540252
rect 411254 540240 411260 540252
rect 343600 540212 411260 540240
rect 343600 540200 343606 540212
rect 411254 540200 411260 540212
rect 411312 540200 411318 540252
rect 29270 538840 29276 538892
rect 29328 538880 29334 538892
rect 29546 538880 29552 538892
rect 29328 538852 29552 538880
rect 29328 538840 29334 538852
rect 29546 538840 29552 538852
rect 29604 538840 29610 538892
rect 357342 538840 357348 538892
rect 357400 538880 357406 538892
rect 375466 538880 375472 538892
rect 357400 538852 375472 538880
rect 357400 538840 357406 538852
rect 375466 538840 375472 538852
rect 375524 538840 375530 538892
rect 524322 538840 524328 538892
rect 524380 538880 524386 538892
rect 554866 538880 554872 538892
rect 524380 538852 554872 538880
rect 524380 538840 524386 538852
rect 554866 538840 554872 538852
rect 554924 538840 554930 538892
rect 3510 538228 3516 538280
rect 3568 538268 3574 538280
rect 10410 538268 10416 538280
rect 3568 538240 10416 538268
rect 3568 538228 3574 538240
rect 10410 538228 10416 538240
rect 10468 538228 10474 538280
rect 353202 537480 353208 537532
rect 353260 537520 353266 537532
rect 378226 537520 378232 537532
rect 353260 537492 378232 537520
rect 353260 537480 353266 537492
rect 378226 537480 378232 537492
rect 378284 537480 378290 537532
rect 165430 537344 165436 537396
rect 165488 537384 165494 537396
rect 431034 537384 431040 537396
rect 165488 537356 431040 537384
rect 165488 537344 165494 537356
rect 431034 537344 431040 537356
rect 431092 537344 431098 537396
rect 163222 537276 163228 537328
rect 163280 537316 163286 537328
rect 433334 537316 433340 537328
rect 163280 537288 433340 537316
rect 163280 537276 163286 537288
rect 433334 537276 433340 537288
rect 433392 537276 433398 537328
rect 158898 537208 158904 537260
rect 158956 537248 158962 537260
rect 437566 537248 437572 537260
rect 158956 537220 437572 537248
rect 158956 537208 158962 537220
rect 437566 537208 437572 537220
rect 437624 537208 437630 537260
rect 156782 537140 156788 537192
rect 156840 537180 156846 537192
rect 439682 537180 439688 537192
rect 156840 537152 439688 537180
rect 156840 537140 156846 537152
rect 439682 537140 439688 537152
rect 439740 537140 439746 537192
rect 152458 537072 152464 537124
rect 152516 537112 152522 537124
rect 444374 537112 444380 537124
rect 152516 537084 444380 537112
rect 152516 537072 152522 537084
rect 444374 537072 444380 537084
rect 444432 537072 444438 537124
rect 150342 537004 150348 537056
rect 150400 537044 150406 537056
rect 446122 537044 446128 537056
rect 150400 537016 446128 537044
rect 150400 537004 150406 537016
rect 446122 537004 446128 537016
rect 446180 537004 446186 537056
rect 148134 536936 148140 536988
rect 148192 536976 148198 536988
rect 448698 536976 448704 536988
rect 148192 536948 448704 536976
rect 148192 536936 148198 536948
rect 448698 536936 448704 536948
rect 448756 536936 448762 536988
rect 146018 536868 146024 536920
rect 146076 536908 146082 536920
rect 450446 536908 450452 536920
rect 146076 536880 450452 536908
rect 146076 536868 146082 536880
rect 450446 536868 450452 536880
rect 450504 536868 450510 536920
rect 112622 536800 112628 536852
rect 112680 536840 112686 536852
rect 483842 536840 483848 536852
rect 112680 536812 483848 536840
rect 112680 536800 112686 536812
rect 483842 536800 483848 536812
rect 483900 536800 483906 536852
rect 363782 536256 363788 536308
rect 363840 536296 363846 536308
rect 376754 536296 376760 536308
rect 363840 536268 376760 536296
rect 363840 536256 363846 536268
rect 376754 536256 376760 536268
rect 376812 536256 376818 536308
rect 317322 536188 317328 536240
rect 317380 536228 317386 536240
rect 400214 536228 400220 536240
rect 317380 536200 400220 536228
rect 317380 536188 317386 536200
rect 400214 536188 400220 536200
rect 400272 536188 400278 536240
rect 194502 536120 194508 536172
rect 194560 536160 194566 536172
rect 401962 536160 401968 536172
rect 194560 536132 401968 536160
rect 194560 536120 194566 536132
rect 401962 536120 401968 536132
rect 402020 536120 402026 536172
rect 193398 536052 193404 536104
rect 193456 536092 193462 536104
rect 403158 536092 403164 536104
rect 193456 536064 403164 536092
rect 193456 536052 193462 536064
rect 403158 536052 403164 536064
rect 403216 536052 403222 536104
rect 154666 535984 154672 536036
rect 154724 536024 154730 536036
rect 441798 536024 441804 536036
rect 154724 535996 441804 536024
rect 154724 535984 154730 535996
rect 441798 535984 441804 535996
rect 441856 535984 441862 536036
rect 139486 535916 139492 535968
rect 139544 535956 139550 535968
rect 456978 535956 456984 535968
rect 139544 535928 456984 535956
rect 139544 535916 139550 535928
rect 456978 535916 456984 535928
rect 457036 535916 457042 535968
rect 137370 535848 137376 535900
rect 137428 535888 137434 535900
rect 459094 535888 459100 535900
rect 137428 535860 459100 535888
rect 137428 535848 137434 535860
rect 459094 535848 459100 535860
rect 459152 535848 459158 535900
rect 127710 535780 127716 535832
rect 127768 535820 127774 535832
rect 468754 535820 468760 535832
rect 127768 535792 468760 535820
rect 127768 535780 127774 535792
rect 468754 535780 468760 535792
rect 468812 535780 468818 535832
rect 125502 535712 125508 535764
rect 125560 535752 125566 535764
rect 470962 535752 470968 535764
rect 125560 535724 470968 535752
rect 125560 535712 125566 535724
rect 470962 535712 470968 535724
rect 471020 535712 471026 535764
rect 123386 535644 123392 535696
rect 123444 535684 123450 535696
rect 473446 535684 473452 535696
rect 123444 535656 473452 535684
rect 123444 535644 123450 535656
rect 473446 535644 473452 535656
rect 473504 535644 473510 535696
rect 121178 535576 121184 535628
rect 121236 535616 121242 535628
rect 475286 535616 475292 535628
rect 121236 535588 475292 535616
rect 121236 535576 121242 535588
rect 475286 535576 475292 535588
rect 475344 535576 475350 535628
rect 117958 535508 117964 535560
rect 118016 535548 118022 535560
rect 478874 535548 478880 535560
rect 118016 535520 478880 535548
rect 118016 535508 118022 535520
rect 478874 535508 478880 535520
rect 478932 535508 478938 535560
rect 109310 535440 109316 535492
rect 109368 535480 109374 535492
rect 483658 535480 483664 535492
rect 109368 535452 483664 535480
rect 109368 535440 109374 535452
rect 483658 535440 483664 535452
rect 483716 535440 483722 535492
rect 364886 535100 364892 535152
rect 364944 535140 364950 535152
rect 364944 535112 373028 535140
rect 364944 535100 364950 535112
rect 372890 535072 372896 535084
rect 365548 535044 372896 535072
rect 28350 534964 28356 535016
rect 28408 535004 28414 535016
rect 37182 535004 37188 535016
rect 28408 534976 37188 535004
rect 28408 534964 28414 534976
rect 37182 534964 37188 534976
rect 37240 534964 37246 535016
rect 25406 534896 25412 534948
rect 25464 534936 25470 534948
rect 34974 534936 34980 534948
rect 25464 534908 34980 534936
rect 25464 534896 25470 534908
rect 34974 534896 34980 534908
rect 35032 534896 35038 534948
rect 362862 534896 362868 534948
rect 362920 534936 362926 534948
rect 365548 534936 365576 535044
rect 372890 535032 372896 535044
rect 372948 535032 372954 535084
rect 365622 534964 365628 535016
rect 365680 535004 365686 535016
rect 370682 535004 370688 535016
rect 365680 534976 370688 535004
rect 365680 534964 365686 534976
rect 370682 534964 370688 534976
rect 370740 534964 370746 535016
rect 373000 535004 373028 535112
rect 375374 535004 375380 535016
rect 373000 534976 375380 535004
rect 375374 534964 375380 534976
rect 375432 534964 375438 535016
rect 362920 534908 365576 534936
rect 362920 534896 362926 534908
rect 367002 534896 367008 534948
rect 367060 534936 367066 534948
rect 371234 534936 371240 534948
rect 367060 534908 371240 534936
rect 367060 534896 367066 534908
rect 371234 534896 371240 534908
rect 371292 534896 371298 534948
rect 25682 534828 25688 534880
rect 25740 534868 25746 534880
rect 39298 534868 39304 534880
rect 25740 534840 39304 534868
rect 25740 534828 25746 534840
rect 39298 534828 39304 534840
rect 39356 534828 39362 534880
rect 358722 534828 358728 534880
rect 358780 534868 358786 534880
rect 375374 534868 375380 534880
rect 358780 534840 375380 534868
rect 358780 534828 358786 534840
rect 375374 534828 375380 534840
rect 375432 534828 375438 534880
rect 28074 534760 28080 534812
rect 28132 534800 28138 534812
rect 41414 534800 41420 534812
rect 28132 534772 41420 534800
rect 28132 534760 28138 534772
rect 41414 534760 41420 534772
rect 41472 534760 41478 534812
rect 362770 534760 362776 534812
rect 362828 534800 362834 534812
rect 379606 534800 379612 534812
rect 362828 534772 379612 534800
rect 362828 534760 362834 534772
rect 379606 534760 379612 534772
rect 379664 534760 379670 534812
rect 25866 534692 25872 534744
rect 25924 534732 25930 534744
rect 43622 534732 43628 534744
rect 25924 534704 43628 534732
rect 25924 534692 25930 534704
rect 43622 534692 43628 534704
rect 43680 534692 43686 534744
rect 360562 534692 360568 534744
rect 360620 534732 360626 534744
rect 382274 534732 382280 534744
rect 360620 534704 382280 534732
rect 360620 534692 360626 534704
rect 382274 534692 382280 534704
rect 382332 534692 382338 534744
rect 192386 534624 192392 534676
rect 192444 534664 192450 534676
rect 404446 534664 404452 534676
rect 192444 534636 404452 534664
rect 192444 534624 192450 534636
rect 404446 534624 404452 534636
rect 404504 534624 404510 534676
rect 189074 534556 189080 534608
rect 189132 534596 189138 534608
rect 407390 534596 407396 534608
rect 189132 534568 407396 534596
rect 189132 534556 189138 534568
rect 407390 534556 407396 534568
rect 407448 534556 407454 534608
rect 185854 534488 185860 534540
rect 185912 534528 185918 534540
rect 410610 534528 410616 534540
rect 185912 534500 410616 534528
rect 185912 534488 185918 534500
rect 410610 534488 410616 534500
rect 410668 534488 410674 534540
rect 179414 534420 179420 534472
rect 179472 534460 179478 534472
rect 417050 534460 417056 534472
rect 179472 534432 417056 534460
rect 179472 534420 179478 534432
rect 417050 534420 417056 534432
rect 417108 534420 417114 534472
rect 177298 534352 177304 534404
rect 177356 534392 177362 534404
rect 419626 534392 419632 534404
rect 177356 534364 419632 534392
rect 177356 534352 177362 534364
rect 419626 534352 419632 534364
rect 419684 534352 419690 534404
rect 172974 534284 172980 534336
rect 173032 534324 173038 534336
rect 423674 534324 423680 534336
rect 173032 534296 423680 534324
rect 173032 534284 173038 534296
rect 423674 534284 423680 534296
rect 423732 534284 423738 534336
rect 170766 534216 170772 534268
rect 170824 534256 170830 534268
rect 425698 534256 425704 534268
rect 170824 534228 425704 534256
rect 170824 534216 170830 534228
rect 425698 534216 425704 534228
rect 425756 534216 425762 534268
rect 166442 534148 166448 534200
rect 166500 534188 166506 534200
rect 430022 534188 430028 534200
rect 166500 534160 430028 534188
rect 166500 534148 166506 534160
rect 430022 534148 430028 534160
rect 430080 534148 430086 534200
rect 29362 534080 29368 534132
rect 29420 534120 29426 534132
rect 30006 534120 30012 534132
rect 29420 534092 30012 534120
rect 29420 534080 29426 534092
rect 30006 534080 30012 534092
rect 30064 534080 30070 534132
rect 164326 534080 164332 534132
rect 164384 534120 164390 534132
rect 432138 534120 432144 534132
rect 164384 534092 432144 534120
rect 164384 534080 164390 534092
rect 432138 534080 432144 534092
rect 432196 534080 432202 534132
rect 342162 534012 342168 534064
rect 342220 534052 342226 534064
rect 385126 534052 385132 534064
rect 342220 534024 385132 534052
rect 342220 534012 342226 534024
rect 385126 534012 385132 534024
rect 385184 534012 385190 534064
rect 339310 533944 339316 533996
rect 339368 533984 339374 533996
rect 386874 533984 386880 533996
rect 339368 533956 386880 533984
rect 339368 533944 339374 533956
rect 386874 533944 386880 533956
rect 386932 533944 386938 533996
rect 335170 533876 335176 533928
rect 335228 533916 335234 533928
rect 389174 533916 389180 533928
rect 335228 533888 389180 533916
rect 335228 533876 335234 533888
rect 389174 533876 389180 533888
rect 389232 533876 389238 533928
rect 30190 533808 30196 533860
rect 30248 533848 30254 533860
rect 52270 533848 52276 533860
rect 30248 533820 52276 533848
rect 30248 533808 30254 533820
rect 52270 533808 52276 533820
rect 52328 533808 52334 533860
rect 331030 533808 331036 533860
rect 331088 533848 331094 533860
rect 391198 533848 391204 533860
rect 331088 533820 391204 533848
rect 331088 533808 331094 533820
rect 391198 533808 391204 533820
rect 391256 533808 391262 533860
rect 518710 533808 518716 533860
rect 518768 533848 518774 533860
rect 553854 533848 553860 533860
rect 518768 533820 553860 533848
rect 518768 533808 518774 533820
rect 553854 533808 553860 533820
rect 553912 533808 553918 533860
rect 25958 533740 25964 533792
rect 26016 533780 26022 533792
rect 50062 533780 50068 533792
rect 26016 533752 50068 533780
rect 26016 533740 26022 533752
rect 50062 533740 50068 533752
rect 50120 533740 50126 533792
rect 328270 533740 328276 533792
rect 328328 533780 328334 533792
rect 393314 533780 393320 533792
rect 328328 533752 393320 533780
rect 328328 533740 328334 533752
rect 393314 533740 393320 533752
rect 393372 533740 393378 533792
rect 516870 533740 516876 533792
rect 516928 533780 516934 533792
rect 553762 533780 553768 533792
rect 516928 533752 553768 533780
rect 516928 533740 516934 533752
rect 553762 533740 553768 533752
rect 553820 533740 553826 533792
rect 30006 533672 30012 533724
rect 30064 533712 30070 533724
rect 60826 533712 60832 533724
rect 30064 533684 60832 533712
rect 30064 533672 30070 533684
rect 60826 533672 60832 533684
rect 60884 533672 60890 533724
rect 318702 533672 318708 533724
rect 318760 533712 318766 533724
rect 398926 533712 398932 533724
rect 318760 533684 398932 533712
rect 318760 533672 318766 533684
rect 398926 533672 398932 533684
rect 398984 533672 398990 533724
rect 514662 533672 514668 533724
rect 514720 533712 514726 533724
rect 551186 533712 551192 533724
rect 514720 533684 551192 533712
rect 514720 533672 514726 533684
rect 551186 533672 551192 533684
rect 551244 533672 551250 533724
rect 26050 533604 26056 533656
rect 26108 533644 26114 533656
rect 58710 533644 58716 533656
rect 26108 533616 58716 533644
rect 26108 533604 26114 533616
rect 58710 533604 58716 533616
rect 58768 533604 58774 533656
rect 322842 533604 322848 533656
rect 322900 533644 322906 533656
rect 445754 533644 445760 533656
rect 322900 533616 445760 533644
rect 322900 533604 322906 533616
rect 445754 533604 445760 533616
rect 445812 533604 445818 533656
rect 512546 533604 512552 533656
rect 512604 533644 512610 533656
rect 553670 533644 553676 533656
rect 512604 533616 553676 533644
rect 512604 533604 512610 533616
rect 553670 533604 553676 533616
rect 553728 533604 553734 533656
rect 27154 533536 27160 533588
rect 27212 533576 27218 533588
rect 69474 533576 69480 533588
rect 27212 533548 69480 533576
rect 27212 533536 27218 533548
rect 69474 533536 69480 533548
rect 69532 533536 69538 533588
rect 321278 533536 321284 533588
rect 321336 533576 321342 533588
rect 447134 533576 447140 533588
rect 321336 533548 447140 533576
rect 321336 533536 321342 533548
rect 447134 533536 447140 533548
rect 447192 533536 447198 533588
rect 510430 533536 510436 533588
rect 510488 533576 510494 533588
rect 553578 533576 553584 533588
rect 510488 533548 553584 533576
rect 510488 533536 510494 533548
rect 553578 533536 553584 533548
rect 553636 533536 553642 533588
rect 27246 533468 27252 533520
rect 27304 533508 27310 533520
rect 73798 533508 73804 533520
rect 27304 533480 73804 533508
rect 27304 533468 27310 533480
rect 73798 533468 73804 533480
rect 73856 533468 73862 533520
rect 320726 533468 320732 533520
rect 320784 533508 320790 533520
rect 448514 533508 448520 533520
rect 320784 533480 448520 533508
rect 320784 533468 320790 533480
rect 448514 533468 448520 533480
rect 448572 533468 448578 533520
rect 530578 533468 530584 533520
rect 530636 533508 530642 533520
rect 574370 533508 574376 533520
rect 530636 533480 574376 533508
rect 530636 533468 530642 533480
rect 574370 533468 574376 533480
rect 574428 533468 574434 533520
rect 27338 533400 27344 533452
rect 27396 533440 27402 533452
rect 78122 533440 78128 533452
rect 27396 533412 78128 533440
rect 27396 533400 27402 533412
rect 78122 533400 78128 533412
rect 78180 533400 78186 533452
rect 319622 533400 319628 533452
rect 319680 533440 319686 533452
rect 451274 533440 451280 533452
rect 319680 533412 451280 533440
rect 319680 533400 319686 533412
rect 451274 533400 451280 533412
rect 451332 533400 451338 533452
rect 508222 533400 508228 533452
rect 508280 533440 508286 533452
rect 553486 533440 553492 533452
rect 508280 533412 553492 533440
rect 508280 533400 508286 533412
rect 553486 533400 553492 533412
rect 553544 533400 553550 533452
rect 27614 533332 27620 533384
rect 27672 533372 27678 533384
rect 80238 533372 80244 533384
rect 27672 533344 80244 533372
rect 27672 533332 27678 533344
rect 80238 533332 80244 533344
rect 80296 533332 80302 533384
rect 318518 533332 318524 533384
rect 318576 533372 318582 533384
rect 452654 533372 452660 533384
rect 318576 533344 452660 533372
rect 318576 533332 318582 533344
rect 452654 533332 452660 533344
rect 452712 533332 452718 533384
rect 503622 533332 503628 533384
rect 503680 533372 503686 533384
rect 553394 533372 553400 533384
rect 503680 533344 553400 533372
rect 503680 533332 503686 533344
rect 553394 533332 553400 533344
rect 553452 533332 553458 533384
rect 346302 533264 346308 533316
rect 346360 533304 346366 533316
rect 382550 533304 382556 533316
rect 346360 533276 382556 533304
rect 346360 533264 346366 533276
rect 382550 533264 382556 533276
rect 382608 533264 382614 533316
rect 349062 533196 349068 533248
rect 349120 533236 349126 533248
rect 380434 533236 380440 533248
rect 349120 533208 380440 533236
rect 349120 533196 349126 533208
rect 380434 533196 380440 533208
rect 380492 533196 380498 533248
rect 354582 533128 354588 533180
rect 354640 533168 354646 533180
rect 377214 533168 377220 533180
rect 354640 533140 377220 533168
rect 354640 533128 354646 533140
rect 377214 533128 377220 533140
rect 377272 533128 377278 533180
rect 188062 532788 188068 532840
rect 188120 532828 188126 532840
rect 408586 532828 408592 532840
rect 188120 532800 408592 532828
rect 188120 532788 188126 532800
rect 408586 532788 408592 532800
rect 408644 532788 408650 532840
rect 168650 532720 168656 532772
rect 168708 532760 168714 532772
rect 427906 532760 427912 532772
rect 168708 532732 427912 532760
rect 168708 532720 168714 532732
rect 427906 532720 427912 532732
rect 427964 532720 427970 532772
rect 357250 532652 357256 532704
rect 357308 532692 357314 532704
rect 387794 532692 387800 532704
rect 357308 532664 387800 532692
rect 357308 532652 357314 532664
rect 387794 532652 387800 532664
rect 387852 532652 387858 532704
rect 504358 532652 504364 532704
rect 504416 532692 504422 532704
rect 508498 532692 508504 532704
rect 504416 532664 508504 532692
rect 504416 532652 504422 532664
rect 508498 532652 508504 532664
rect 508556 532652 508562 532704
rect 355226 532584 355232 532636
rect 355284 532624 355290 532636
rect 392026 532624 392032 532636
rect 355284 532596 392032 532624
rect 355284 532584 355290 532596
rect 392026 532584 392032 532596
rect 392084 532584 392090 532636
rect 353018 532516 353024 532568
rect 353076 532556 353082 532568
rect 394786 532556 394792 532568
rect 353076 532528 394792 532556
rect 353076 532516 353082 532528
rect 394786 532516 394792 532528
rect 394844 532516 394850 532568
rect 261294 532448 261300 532500
rect 261352 532488 261358 532500
rect 262122 532488 262128 532500
rect 261352 532460 262128 532488
rect 261352 532448 261358 532460
rect 262122 532448 262128 532460
rect 262180 532448 262186 532500
rect 262398 532448 262404 532500
rect 262456 532488 262462 532500
rect 263410 532488 263416 532500
rect 262456 532460 263416 532488
rect 262456 532448 262462 532460
rect 263410 532448 263416 532460
rect 263468 532448 263474 532500
rect 350902 532448 350908 532500
rect 350960 532488 350966 532500
rect 398834 532488 398840 532500
rect 350960 532460 398840 532488
rect 350960 532448 350966 532460
rect 398834 532448 398840 532460
rect 398892 532448 398898 532500
rect 348694 532380 348700 532432
rect 348752 532420 348758 532432
rect 401594 532420 401600 532432
rect 348752 532392 401600 532420
rect 348752 532380 348758 532392
rect 401594 532380 401600 532392
rect 401652 532380 401658 532432
rect 346302 532312 346308 532364
rect 346360 532352 346366 532364
rect 405734 532352 405740 532364
rect 346360 532324 405740 532352
rect 346360 532312 346366 532324
rect 405734 532312 405740 532324
rect 405792 532312 405798 532364
rect 344370 532244 344376 532296
rect 344428 532284 344434 532296
rect 409874 532284 409880 532296
rect 344428 532256 409880 532284
rect 344428 532244 344434 532256
rect 409874 532244 409880 532256
rect 409932 532244 409938 532296
rect 342162 532176 342168 532228
rect 342220 532216 342226 532228
rect 412634 532216 412640 532228
rect 342220 532188 412640 532216
rect 342220 532176 342226 532188
rect 412634 532176 412640 532188
rect 412692 532176 412698 532228
rect 30282 532108 30288 532160
rect 30340 532148 30346 532160
rect 40402 532148 40408 532160
rect 30340 532120 40408 532148
rect 30340 532108 30346 532120
rect 40402 532108 40408 532120
rect 40460 532108 40466 532160
rect 340046 532108 340052 532160
rect 340104 532148 340110 532160
rect 416774 532148 416780 532160
rect 340104 532120 416780 532148
rect 340104 532108 340110 532120
rect 416774 532108 416780 532120
rect 416832 532108 416838 532160
rect 521194 532108 521200 532160
rect 521252 532148 521258 532160
rect 553946 532148 553952 532160
rect 521252 532120 553952 532148
rect 521252 532108 521258 532120
rect 553946 532108 553952 532120
rect 554004 532108 554010 532160
rect 27430 532040 27436 532092
rect 27488 532080 27494 532092
rect 87782 532080 87788 532092
rect 27488 532052 87788 532080
rect 27488 532040 27494 532052
rect 87782 532040 87788 532052
rect 87840 532040 87846 532092
rect 321462 532040 321468 532092
rect 321520 532080 321526 532092
rect 397638 532080 397644 532092
rect 321520 532052 397644 532080
rect 321520 532040 321526 532052
rect 397638 532040 397644 532052
rect 397696 532040 397702 532092
rect 401502 532040 401508 532092
rect 401560 532080 401566 532092
rect 455414 532080 455420 532092
rect 401560 532052 455420 532080
rect 401560 532040 401566 532052
rect 455414 532040 455420 532052
rect 455472 532040 455478 532092
rect 517974 532040 517980 532092
rect 518032 532080 518038 532092
rect 551278 532080 551284 532092
rect 518032 532052 551284 532080
rect 518032 532040 518038 532052
rect 551278 532040 551284 532052
rect 551336 532040 551342 532092
rect 27522 531972 27528 532024
rect 27580 532012 27586 532024
rect 89990 532012 89996 532024
rect 27580 531984 89996 532012
rect 27580 531972 27586 531984
rect 89990 531972 89996 531984
rect 90048 531972 90054 532024
rect 337930 531972 337936 532024
rect 337988 532012 337994 532024
rect 419534 532012 419540 532024
rect 337988 531984 419540 532012
rect 337988 531972 337994 531984
rect 419534 531972 419540 531984
rect 419592 531972 419598 532024
rect 513650 531972 513656 532024
rect 513708 532012 513714 532024
rect 550726 532012 550732 532024
rect 513708 531984 550732 532012
rect 513708 531972 513714 531984
rect 550726 531972 550732 531984
rect 550784 531972 550790 532024
rect 359458 531904 359464 531956
rect 359516 531944 359522 531956
rect 383654 531944 383660 531956
rect 359516 531916 383660 531944
rect 359516 531904 359522 531916
rect 383654 531904 383660 531916
rect 383712 531904 383718 531956
rect 361482 531836 361488 531888
rect 361540 531876 361546 531888
rect 380986 531876 380992 531888
rect 361540 531848 380992 531876
rect 361540 531836 361546 531848
rect 380986 531836 380992 531848
rect 381044 531836 381050 531888
rect 178310 531768 178316 531820
rect 178368 531808 178374 531820
rect 340138 531808 340144 531820
rect 178368 531780 340144 531808
rect 178368 531768 178374 531780
rect 340138 531768 340144 531780
rect 340196 531768 340202 531820
rect 176194 531700 176200 531752
rect 176252 531740 176258 531752
rect 343634 531740 343640 531752
rect 176252 531712 343640 531740
rect 176252 531700 176258 531712
rect 343634 531700 343640 531712
rect 343692 531700 343698 531752
rect 173986 531632 173992 531684
rect 174044 531672 174050 531684
rect 349062 531672 349068 531684
rect 174044 531644 349068 531672
rect 174044 531632 174050 531644
rect 349062 531632 349068 531644
rect 349120 531632 349126 531684
rect 171870 531564 171876 531616
rect 171928 531604 171934 531616
rect 351914 531604 351920 531616
rect 171928 531576 351920 531604
rect 171928 531564 171934 531576
rect 351914 531564 351920 531576
rect 351972 531564 351978 531616
rect 169754 531496 169760 531548
rect 169812 531536 169818 531548
rect 357342 531536 357348 531548
rect 169812 531508 357348 531536
rect 169812 531496 169818 531508
rect 357342 531496 357348 531508
rect 357400 531496 357406 531548
rect 183738 531428 183744 531480
rect 183796 531468 183802 531480
rect 412726 531468 412732 531480
rect 183796 531440 412732 531468
rect 183796 531428 183802 531440
rect 412726 531428 412732 531440
rect 412784 531428 412790 531480
rect 147030 531360 147036 531412
rect 147088 531400 147094 531412
rect 449434 531400 449440 531412
rect 147088 531372 449440 531400
rect 147088 531360 147094 531372
rect 449434 531360 449440 531372
rect 449492 531360 449498 531412
rect 142798 531292 142804 531344
rect 142856 531332 142862 531344
rect 454034 531332 454040 531344
rect 142856 531304 454040 531332
rect 142856 531292 142862 531304
rect 454034 531292 454040 531304
rect 454092 531292 454098 531344
rect 544838 531292 544844 531344
rect 544896 531332 544902 531344
rect 551738 531332 551744 531344
rect 544896 531304 551744 531332
rect 544896 531292 544902 531304
rect 551738 531292 551744 531304
rect 551796 531292 551802 531344
rect 30098 531224 30104 531276
rect 30156 531264 30162 531276
rect 51166 531264 51172 531276
rect 30156 531236 51172 531264
rect 30156 531224 30162 531236
rect 51166 531224 51172 531236
rect 51224 531224 51230 531276
rect 331490 531224 331496 531276
rect 331548 531264 331554 531276
rect 332410 531264 332416 531276
rect 331548 531236 332416 531264
rect 331548 531224 331554 531236
rect 332410 531224 332416 531236
rect 332468 531224 332474 531276
rect 334710 531224 334716 531276
rect 334768 531264 334774 531276
rect 335262 531264 335268 531276
rect 334768 531236 335268 531264
rect 334768 531224 334774 531236
rect 335262 531224 335268 531236
rect 335320 531224 335326 531276
rect 335814 531224 335820 531276
rect 335872 531264 335878 531276
rect 336550 531264 336556 531276
rect 335872 531236 336556 531264
rect 335872 531224 335878 531236
rect 336550 531224 336556 531236
rect 336608 531224 336614 531276
rect 341150 531224 341156 531276
rect 341208 531264 341214 531276
rect 342070 531264 342076 531276
rect 341208 531236 342076 531264
rect 341208 531224 341214 531236
rect 342070 531224 342076 531236
rect 342128 531224 342134 531276
rect 345474 531224 345480 531276
rect 345532 531264 345538 531276
rect 346210 531264 346216 531276
rect 345532 531236 346216 531264
rect 345532 531224 345538 531236
rect 346210 531224 346216 531236
rect 346268 531224 346274 531276
rect 349798 531224 349804 531276
rect 349856 531264 349862 531276
rect 350442 531264 350448 531276
rect 349856 531236 350448 531264
rect 349856 531224 349862 531236
rect 350442 531224 350448 531236
rect 350500 531224 350506 531276
rect 354030 531224 354036 531276
rect 354088 531264 354094 531276
rect 354490 531264 354496 531276
rect 354088 531236 354496 531264
rect 354088 531224 354094 531236
rect 354490 531224 354496 531236
rect 354548 531224 354554 531276
rect 365990 531224 365996 531276
rect 366048 531264 366054 531276
rect 366910 531264 366916 531276
rect 366048 531236 366916 531264
rect 366048 531224 366054 531236
rect 366910 531224 366916 531236
rect 366968 531224 366974 531276
rect 483658 531224 483664 531276
rect 483716 531264 483722 531276
rect 487154 531264 487160 531276
rect 483716 531236 487160 531264
rect 483716 531224 483722 531236
rect 487154 531224 487160 531236
rect 487212 531224 487218 531276
rect 526530 531224 526536 531276
rect 526588 531264 526594 531276
rect 527082 531264 527088 531276
rect 526588 531236 527088 531264
rect 526588 531224 526594 531236
rect 527082 531224 527088 531236
rect 527140 531224 527146 531276
rect 527634 531224 527640 531276
rect 527692 531264 527698 531276
rect 528462 531264 528468 531276
rect 527692 531236 528468 531264
rect 527692 531224 527698 531236
rect 528462 531224 528468 531236
rect 528520 531224 528526 531276
rect 530854 531224 530860 531276
rect 530912 531264 530918 531276
rect 531222 531264 531228 531276
rect 530912 531236 531228 531264
rect 530912 531224 530918 531236
rect 531222 531224 531228 531236
rect 531280 531224 531286 531276
rect 531958 531224 531964 531276
rect 532016 531264 532022 531276
rect 532602 531264 532608 531276
rect 532016 531236 532608 531264
rect 532016 531224 532022 531236
rect 532602 531224 532608 531236
rect 532660 531224 532666 531276
rect 536282 531224 536288 531276
rect 536340 531264 536346 531276
rect 536742 531264 536748 531276
rect 536340 531236 536748 531264
rect 536340 531224 536346 531236
rect 536742 531224 536748 531236
rect 536800 531224 536806 531276
rect 545574 531224 545580 531276
rect 545632 531264 545638 531276
rect 552014 531264 552020 531276
rect 545632 531236 552020 531264
rect 545632 531224 545638 531236
rect 552014 531224 552020 531236
rect 552072 531224 552078 531276
rect 553210 531224 553216 531276
rect 553268 531264 553274 531276
rect 554038 531264 554044 531276
rect 553268 531236 554044 531264
rect 553268 531224 553274 531236
rect 554038 531224 554044 531236
rect 554096 531224 554102 531276
rect 29914 531156 29920 531208
rect 29972 531196 29978 531208
rect 55490 531196 55496 531208
rect 29972 531168 55496 531196
rect 29972 531156 29978 531168
rect 55490 531156 55496 531168
rect 55548 531156 55554 531208
rect 552474 531196 552480 531208
rect 548076 531168 552480 531196
rect 24578 531088 24584 531140
rect 24636 531128 24642 531140
rect 25314 531128 25320 531140
rect 24636 531100 25320 531128
rect 24636 531088 24642 531100
rect 25314 531088 25320 531100
rect 25372 531088 25378 531140
rect 25498 531088 25504 531140
rect 25556 531128 25562 531140
rect 27430 531128 27436 531140
rect 25556 531100 27436 531128
rect 25556 531088 25562 531100
rect 27430 531088 27436 531100
rect 27488 531088 27494 531140
rect 27890 531088 27896 531140
rect 27948 531128 27954 531140
rect 57606 531128 57612 531140
rect 27948 531100 57612 531128
rect 27948 531088 27954 531100
rect 57606 531088 57612 531100
rect 57664 531088 57670 531140
rect 119062 531088 119068 531140
rect 119120 531128 119126 531140
rect 477494 531128 477500 531140
rect 119120 531100 477500 531128
rect 119120 531088 119126 531100
rect 477494 531088 477500 531100
rect 477552 531088 477558 531140
rect 543550 531088 543556 531140
rect 543608 531128 543614 531140
rect 548076 531128 548104 531168
rect 552474 531156 552480 531168
rect 552532 531156 552538 531208
rect 543608 531100 548104 531128
rect 543608 531088 543614 531100
rect 551370 531088 551376 531140
rect 551428 531128 551434 531140
rect 551922 531128 551928 531140
rect 551428 531100 551928 531128
rect 551428 531088 551434 531100
rect 551922 531088 551928 531100
rect 551980 531088 551986 531140
rect 29822 531020 29828 531072
rect 29880 531060 29886 531072
rect 59814 531060 59820 531072
rect 29880 531032 59820 531060
rect 29880 531020 29886 531032
rect 59814 531020 59820 531032
rect 59872 531020 59878 531072
rect 198734 531020 198740 531072
rect 198792 531060 198798 531072
rect 199654 531060 199660 531072
rect 198792 531032 199660 531060
rect 198792 531020 198798 531032
rect 199654 531020 199660 531032
rect 199712 531020 199718 531072
rect 213914 531020 213920 531072
rect 213972 531060 213978 531072
rect 214742 531060 214748 531072
rect 213972 531032 214748 531060
rect 213972 531020 213978 531032
rect 214742 531020 214748 531032
rect 214800 531020 214806 531072
rect 227714 531020 227720 531072
rect 227772 531060 227778 531072
rect 228726 531060 228732 531072
rect 227772 531032 228732 531060
rect 227772 531020 227778 531032
rect 228726 531020 228732 531032
rect 228784 531020 228790 531072
rect 233234 531020 233240 531072
rect 233292 531060 233298 531072
rect 234062 531060 234068 531072
rect 233292 531032 234068 531060
rect 233292 531020 233298 531032
rect 234062 531020 234068 531032
rect 234120 531020 234126 531072
rect 242894 531020 242900 531072
rect 242952 531060 242958 531072
rect 243814 531060 243820 531072
rect 242952 531032 243820 531060
rect 242952 531020 242958 531032
rect 243814 531020 243820 531032
rect 243872 531020 243878 531072
rect 248414 531020 248420 531072
rect 248472 531060 248478 531072
rect 249150 531060 249156 531072
rect 248472 531032 249156 531060
rect 248472 531020 248478 531032
rect 249150 531020 249156 531032
rect 249208 531020 249214 531072
rect 266722 531020 266728 531072
rect 266780 531060 266786 531072
rect 267642 531060 267648 531072
rect 266780 531032 267648 531060
rect 266780 531020 266786 531032
rect 267642 531020 267648 531032
rect 267700 531020 267706 531072
rect 267826 531020 267832 531072
rect 267884 531060 267890 531072
rect 269022 531060 269028 531072
rect 267884 531032 269028 531060
rect 267884 531020 267890 531032
rect 269022 531020 269028 531032
rect 269080 531020 269086 531072
rect 272058 531020 272064 531072
rect 272116 531060 272122 531072
rect 273070 531060 273076 531072
rect 272116 531032 273076 531060
rect 272116 531020 272122 531032
rect 273070 531020 273076 531032
rect 273128 531020 273134 531072
rect 276382 531020 276388 531072
rect 276440 531060 276446 531072
rect 277302 531060 277308 531072
rect 276440 531032 277308 531060
rect 276440 531020 276446 531032
rect 277302 531020 277308 531032
rect 277360 531020 277366 531072
rect 277486 531020 277492 531072
rect 277544 531060 277550 531072
rect 278682 531060 278688 531072
rect 277544 531032 278688 531060
rect 277544 531020 277550 531032
rect 278682 531020 278688 531032
rect 278740 531020 278746 531072
rect 325050 531020 325056 531072
rect 325108 531060 325114 531072
rect 325602 531060 325608 531072
rect 325108 531032 325608 531060
rect 325108 531020 325114 531032
rect 325602 531020 325608 531032
rect 325660 531020 325666 531072
rect 329282 531020 329288 531072
rect 329340 531060 329346 531072
rect 329742 531060 329748 531072
rect 329340 531032 329748 531060
rect 329340 531020 329346 531032
rect 329742 531020 329748 531032
rect 329800 531020 329806 531072
rect 330386 531020 330392 531072
rect 330444 531060 330450 531072
rect 331122 531060 331128 531072
rect 330444 531032 331128 531060
rect 330444 531020 330450 531032
rect 331122 531020 331128 531032
rect 331180 531020 331186 531072
rect 357342 531020 357348 531072
rect 357400 531060 357406 531072
rect 426710 531060 426716 531072
rect 357400 531032 426716 531060
rect 357400 531020 357406 531032
rect 426710 531020 426716 531032
rect 426768 531020 426774 531072
rect 541618 531020 541624 531072
rect 541676 531060 541682 531072
rect 541676 531032 545896 531060
rect 541676 531020 541682 531032
rect 27798 530952 27804 531004
rect 27856 530992 27862 531004
rect 61930 530992 61936 531004
rect 27856 530964 61936 530992
rect 27856 530952 27862 530964
rect 61930 530952 61936 530964
rect 61988 530952 61994 531004
rect 271046 530952 271052 531004
rect 271104 530992 271110 531004
rect 271782 530992 271788 531004
rect 271104 530964 271788 530992
rect 271104 530952 271110 530964
rect 271782 530952 271788 530964
rect 271840 530952 271846 531004
rect 351914 530952 351920 531004
rect 351972 530992 351978 531004
rect 424594 530992 424600 531004
rect 351972 530964 424600 530992
rect 351972 530952 351978 530964
rect 424594 530952 424600 530964
rect 424652 530952 424658 531004
rect 539502 530952 539508 531004
rect 539560 530992 539566 531004
rect 545758 530992 545764 531004
rect 539560 530964 545764 530992
rect 539560 530952 539566 530964
rect 545758 530952 545764 530964
rect 545816 530952 545822 531004
rect 545868 530992 545896 531032
rect 545942 531020 545948 531072
rect 546000 531060 546006 531072
rect 552566 531060 552572 531072
rect 546000 531032 552572 531060
rect 546000 531020 546006 531032
rect 552566 531020 552572 531032
rect 552624 531020 552630 531072
rect 552382 530992 552388 531004
rect 545868 530964 552388 530992
rect 552382 530952 552388 530964
rect 552440 530952 552446 531004
rect 29730 530884 29736 530936
rect 29788 530924 29794 530936
rect 64046 530924 64052 530936
rect 29788 530896 64052 530924
rect 29788 530884 29794 530896
rect 64046 530884 64052 530896
rect 64104 530884 64110 530936
rect 326062 530884 326068 530936
rect 326120 530924 326126 530936
rect 326982 530924 326988 530936
rect 326120 530896 326988 530924
rect 326120 530884 326126 530896
rect 326982 530884 326988 530896
rect 327040 530884 327046 530936
rect 349062 530884 349068 530936
rect 349120 530924 349126 530936
rect 422478 530924 422484 530936
rect 349120 530896 422484 530924
rect 349120 530884 349126 530896
rect 422478 530884 422484 530896
rect 422536 530884 422542 530936
rect 537294 530884 537300 530936
rect 537352 530924 537358 530936
rect 552198 530924 552204 530936
rect 537352 530896 552204 530924
rect 537352 530884 537358 530896
rect 552198 530884 552204 530896
rect 552256 530884 552262 530936
rect 29546 530816 29552 530868
rect 29604 530856 29610 530868
rect 66254 530856 66260 530868
rect 29604 530828 66260 530856
rect 29604 530816 29610 530828
rect 66254 530816 66260 530828
rect 66312 530816 66318 530868
rect 343634 530816 343640 530868
rect 343692 530856 343698 530868
rect 420270 530856 420276 530868
rect 343692 530828 420276 530856
rect 343692 530816 343698 530828
rect 420270 530816 420276 530828
rect 420328 530816 420334 530868
rect 523310 530816 523316 530868
rect 523368 530856 523374 530868
rect 524322 530856 524328 530868
rect 523368 530828 524328 530856
rect 523368 530816 523374 530828
rect 524322 530816 524328 530828
rect 524380 530816 524386 530868
rect 535178 530816 535184 530868
rect 535236 530856 535242 530868
rect 545666 530856 545672 530868
rect 535236 530828 545672 530856
rect 535236 530816 535242 530828
rect 545666 530816 545672 530828
rect 545724 530816 545730 530868
rect 545758 530816 545764 530868
rect 545816 530856 545822 530868
rect 552290 530856 552296 530868
rect 545816 530828 552296 530856
rect 545816 530816 545822 530828
rect 552290 530816 552296 530828
rect 552348 530816 552354 530868
rect 27706 530748 27712 530800
rect 27764 530788 27770 530800
rect 68370 530788 68376 530800
rect 27764 530760 68376 530788
rect 27764 530748 27770 530760
rect 68370 530748 68376 530760
rect 68428 530748 68434 530800
rect 340138 530748 340144 530800
rect 340196 530788 340202 530800
rect 418246 530788 418252 530800
rect 340196 530760 418252 530788
rect 340196 530748 340202 530760
rect 418246 530748 418252 530760
rect 418304 530748 418310 530800
rect 533062 530748 533068 530800
rect 533120 530788 533126 530800
rect 551462 530788 551468 530800
rect 533120 530760 551468 530788
rect 533120 530748 533126 530760
rect 551462 530748 551468 530760
rect 551520 530748 551526 530800
rect 25222 530680 25228 530732
rect 25280 530720 25286 530732
rect 67358 530720 67364 530732
rect 25280 530692 67364 530720
rect 25280 530680 25286 530692
rect 67358 530680 67364 530692
rect 67416 530680 67422 530732
rect 186958 530680 186964 530732
rect 187016 530720 187022 530732
rect 409874 530720 409880 530732
rect 187016 530692 409880 530720
rect 187016 530680 187022 530692
rect 409874 530680 409880 530692
rect 409932 530680 409938 530732
rect 528462 530680 528468 530732
rect 528520 530720 528526 530732
rect 545574 530720 545580 530732
rect 528520 530692 545580 530720
rect 528520 530680 528526 530692
rect 545574 530680 545580 530692
rect 545632 530680 545638 530732
rect 545666 530680 545672 530732
rect 545724 530720 545730 530732
rect 552106 530720 552112 530732
rect 545724 530692 552112 530720
rect 545724 530680 545730 530692
rect 552106 530680 552112 530692
rect 552164 530680 552170 530732
rect 555418 530680 555424 530732
rect 555476 530720 555482 530732
rect 562594 530720 562600 530732
rect 555476 530692 562600 530720
rect 555476 530680 555482 530692
rect 562594 530680 562600 530692
rect 562652 530680 562658 530732
rect 23290 530612 23296 530664
rect 23348 530652 23354 530664
rect 23348 530624 23520 530652
rect 23348 530612 23354 530624
rect 22094 530544 22100 530596
rect 22152 530584 22158 530596
rect 23382 530584 23388 530596
rect 22152 530556 23388 530584
rect 22152 530544 22158 530556
rect 23382 530544 23388 530556
rect 23440 530544 23446 530596
rect 23492 530584 23520 530624
rect 24762 530612 24768 530664
rect 24820 530652 24826 530664
rect 77018 530652 77024 530664
rect 24820 530624 77024 530652
rect 24820 530612 24826 530624
rect 77018 530612 77024 530624
rect 77076 530612 77082 530664
rect 184842 530612 184848 530664
rect 184900 530652 184906 530664
rect 411622 530652 411628 530664
rect 184900 530624 411628 530652
rect 184900 530612 184906 530624
rect 411622 530612 411628 530624
rect 411680 530612 411686 530664
rect 522206 530612 522212 530664
rect 522264 530652 522270 530664
rect 551278 530652 551284 530664
rect 522264 530624 551284 530652
rect 522264 530612 522270 530624
rect 551278 530612 551284 530624
rect 551336 530612 551342 530664
rect 85666 530584 85672 530596
rect 23492 530556 85672 530584
rect 85666 530544 85672 530556
rect 85724 530544 85730 530596
rect 182634 530544 182640 530596
rect 182692 530584 182698 530596
rect 414014 530584 414020 530596
rect 182692 530556 414020 530584
rect 182692 530544 182698 530556
rect 414014 530544 414020 530556
rect 414072 530544 414078 530596
rect 505002 530544 505008 530596
rect 505060 530584 505066 530596
rect 556246 530584 556252 530596
rect 505060 530556 556252 530584
rect 505060 530544 505066 530556
rect 556246 530544 556252 530556
rect 556304 530544 556310 530596
rect 558178 530544 558184 530596
rect 558236 530584 558242 530596
rect 572254 530584 572260 530596
rect 558236 530556 572260 530584
rect 558236 530544 558242 530556
rect 572254 530544 572260 530556
rect 572312 530544 572318 530596
rect 24670 530476 24676 530528
rect 24728 530516 24734 530528
rect 44726 530516 44732 530528
rect 24728 530488 44732 530516
rect 24728 530476 24734 530488
rect 44726 530476 44732 530488
rect 44784 530476 44790 530528
rect 115842 530476 115848 530528
rect 115900 530516 115906 530528
rect 348878 530516 348884 530528
rect 115900 530488 348884 530516
rect 115900 530476 115906 530488
rect 348878 530476 348884 530488
rect 348936 530476 348942 530528
rect 29270 530408 29276 530460
rect 29328 530448 29334 530460
rect 46842 530448 46848 530460
rect 29328 530420 46848 530448
rect 29328 530408 29334 530420
rect 46842 530408 46848 530420
rect 46900 530408 46906 530460
rect 180518 530408 180524 530460
rect 180576 530448 180582 530460
rect 415946 530448 415952 530460
rect 180576 530420 415952 530448
rect 180576 530408 180582 530420
rect 415946 530408 415952 530420
rect 416004 530408 416010 530460
rect 25038 530340 25044 530392
rect 25096 530380 25102 530392
rect 32858 530380 32864 530392
rect 25096 530352 32864 530380
rect 25096 530340 25102 530352
rect 32858 530340 32864 530352
rect 32916 530340 32922 530392
rect 133046 530340 133052 530392
rect 133104 530380 133110 530392
rect 463786 530380 463792 530392
rect 133104 530352 463792 530380
rect 133104 530340 133110 530352
rect 463786 530340 463792 530352
rect 463844 530340 463850 530392
rect 130930 530272 130936 530324
rect 130988 530312 130994 530324
rect 465534 530312 465540 530324
rect 130988 530284 465540 530312
rect 130988 530272 130994 530284
rect 465534 530272 465540 530284
rect 465592 530272 465598 530324
rect 128722 530204 128728 530256
rect 128780 530244 128786 530256
rect 467834 530244 467840 530256
rect 128780 530216 467840 530244
rect 128780 530204 128786 530216
rect 467834 530204 467840 530216
rect 467892 530204 467898 530256
rect 24946 530136 24952 530188
rect 25004 530176 25010 530188
rect 29638 530176 29644 530188
rect 25004 530148 29644 530176
rect 25004 530136 25010 530148
rect 29638 530136 29644 530148
rect 29696 530136 29702 530188
rect 126606 530136 126612 530188
rect 126664 530176 126670 530188
rect 469858 530176 469864 530188
rect 126664 530148 469864 530176
rect 126664 530136 126670 530148
rect 469858 530136 469864 530148
rect 469916 530136 469922 530188
rect 542722 530136 542728 530188
rect 542780 530176 542786 530188
rect 543642 530176 543648 530188
rect 542780 530148 543648 530176
rect 542780 530136 542786 530148
rect 543642 530136 543648 530148
rect 543700 530136 543706 530188
rect 547046 530136 547052 530188
rect 547104 530176 547110 530188
rect 547782 530176 547788 530188
rect 547104 530148 547788 530176
rect 547104 530136 547110 530148
rect 547782 530136 547788 530148
rect 547840 530136 547846 530188
rect 548150 530136 548156 530188
rect 548208 530176 548214 530188
rect 549070 530176 549076 530188
rect 548208 530148 549076 530176
rect 548208 530136 548214 530148
rect 549070 530136 549076 530148
rect 549128 530136 549134 530188
rect 124398 530068 124404 530120
rect 124456 530108 124462 530120
rect 472066 530108 472072 530120
rect 124456 530080 472072 530108
rect 124456 530068 124462 530080
rect 472066 530068 472072 530080
rect 472124 530068 472130 530120
rect 122282 530000 122288 530052
rect 122340 530040 122346 530052
rect 474182 530040 474188 530052
rect 122340 530012 474188 530040
rect 122340 530000 122346 530012
rect 474182 530000 474188 530012
rect 474240 530000 474246 530052
rect 419442 529932 419448 529984
rect 419500 529972 419506 529984
rect 429286 529972 429292 529984
rect 419500 529944 429292 529972
rect 419500 529932 419506 529944
rect 429286 529932 429292 529944
rect 429344 529932 429350 529984
rect 556798 529932 556804 529984
rect 556856 529972 556862 529984
rect 558270 529972 558276 529984
rect 556856 529944 558276 529972
rect 556856 529932 556862 529944
rect 558270 529932 558276 529944
rect 558328 529932 558334 529984
rect 560938 529932 560944 529984
rect 560996 529972 561002 529984
rect 567930 529972 567936 529984
rect 560996 529944 567936 529972
rect 560996 529932 561002 529944
rect 567930 529932 567936 529944
rect 567988 529932 567994 529984
rect 348878 529592 348884 529644
rect 348936 529632 348942 529644
rect 480622 529632 480628 529644
rect 348936 529604 480628 529632
rect 348936 529592 348942 529604
rect 480622 529592 480628 529604
rect 480680 529592 480686 529644
rect 191282 529524 191288 529576
rect 191340 529564 191346 529576
rect 405182 529564 405188 529576
rect 191340 529536 405188 529564
rect 191340 529524 191346 529536
rect 405182 529524 405188 529536
rect 405240 529524 405246 529576
rect 175090 529456 175096 529508
rect 175148 529496 175154 529508
rect 421374 529496 421380 529508
rect 175148 529468 421380 529496
rect 175148 529456 175154 529468
rect 421374 529456 421380 529468
rect 421432 529456 421438 529508
rect 167546 529388 167552 529440
rect 167604 529428 167610 529440
rect 419442 529428 419448 529440
rect 167604 529400 419448 529428
rect 167604 529388 167610 529400
rect 419442 529388 419448 529400
rect 419500 529388 419506 529440
rect 155678 529320 155684 529372
rect 155736 529360 155742 529372
rect 440786 529360 440792 529372
rect 155736 529332 440792 529360
rect 155736 529320 155742 529332
rect 440786 529320 440792 529332
rect 440844 529320 440850 529372
rect 149238 529252 149244 529304
rect 149296 529292 149302 529304
rect 447226 529292 447232 529304
rect 149296 529264 447232 529292
rect 149296 529252 149302 529264
rect 447226 529252 447232 529264
rect 447284 529252 447290 529304
rect 144914 529184 144920 529236
rect 144972 529224 144978 529236
rect 451550 529224 451556 529236
rect 144972 529196 451556 529224
rect 144972 529184 144978 529196
rect 451550 529184 451556 529196
rect 451608 529184 451614 529236
rect 140590 529116 140596 529168
rect 140648 529156 140654 529168
rect 455874 529156 455880 529168
rect 140648 529128 455880 529156
rect 140648 529116 140654 529128
rect 455874 529116 455880 529128
rect 455932 529116 455938 529168
rect 136266 529048 136272 529100
rect 136324 529088 136330 529100
rect 460520 529088 460526 529100
rect 136324 529060 460526 529088
rect 136324 529048 136330 529060
rect 460520 529048 460526 529060
rect 460578 529048 460584 529100
rect 134150 528980 134156 529032
rect 134208 529020 134214 529032
rect 462636 529020 462642 529032
rect 134208 528992 462642 529020
rect 134208 528980 134214 528992
rect 462636 528980 462642 528992
rect 462694 528980 462700 529032
rect 120442 528912 120448 528964
rect 120500 528952 120506 528964
rect 476298 528952 476304 528964
rect 120500 528924 476304 528952
rect 120500 528912 120506 528924
rect 476298 528912 476304 528924
rect 476356 528912 476362 528964
rect 117130 528844 117136 528896
rect 117188 528884 117194 528896
rect 479610 528884 479616 528896
rect 117188 528856 479616 528884
rect 117188 528844 117194 528856
rect 479610 528844 479616 528856
rect 479668 528844 479674 528896
rect 114002 528776 114008 528828
rect 114060 528816 114066 528828
rect 483014 528816 483020 528828
rect 114060 528788 483020 528816
rect 114060 528776 114066 528788
rect 483014 528776 483020 528788
rect 483072 528776 483078 528828
rect 110690 528708 110696 528760
rect 110748 528748 110754 528760
rect 398834 528748 398840 528760
rect 110748 528720 398840 528748
rect 110748 528708 110754 528720
rect 398834 528708 398840 528720
rect 398892 528708 398898 528760
rect 399202 528708 399208 528760
rect 399260 528748 399266 528760
rect 486050 528748 486056 528760
rect 399260 528720 486056 528748
rect 399260 528708 399266 528720
rect 486050 528708 486056 528720
rect 486108 528708 486114 528760
rect 108666 528640 108672 528692
rect 108724 528680 108730 528692
rect 398926 528680 398932 528692
rect 108724 528652 398932 528680
rect 108724 528640 108730 528652
rect 398926 528640 398932 528652
rect 398984 528640 398990 528692
rect 403618 528640 403624 528692
rect 403676 528680 403682 528692
rect 488350 528680 488356 528692
rect 403676 528652 488356 528680
rect 403676 528640 403682 528652
rect 488350 528640 488356 528652
rect 488408 528640 488414 528692
rect 107562 528572 107568 528624
rect 107620 528612 107626 528624
rect 411254 528612 411260 528624
rect 107620 528584 398972 528612
rect 107620 528572 107626 528584
rect 251910 528504 251916 528556
rect 251968 528544 251974 528556
rect 254210 528544 254216 528556
rect 251968 528516 254216 528544
rect 251968 528504 251974 528516
rect 254210 528504 254216 528516
rect 254268 528504 254274 528556
rect 315390 528504 315396 528556
rect 315448 528544 315454 528556
rect 319622 528544 319628 528556
rect 315448 528516 319628 528544
rect 315448 528504 315454 528516
rect 319622 528504 319628 528516
rect 319680 528504 319686 528556
rect 398834 528544 398840 528556
rect 386156 528516 398840 528544
rect 184198 528476 184204 528488
rect 182284 528448 184204 528476
rect 153930 528368 153936 528420
rect 153988 528408 153994 528420
rect 159358 528408 159364 528420
rect 153988 528380 159364 528408
rect 153988 528368 153994 528380
rect 159358 528368 159364 528380
rect 159416 528368 159422 528420
rect 175182 528368 175188 528420
rect 175240 528408 175246 528420
rect 175240 528380 177988 528408
rect 175240 528368 175246 528380
rect 151464 528244 159312 528272
rect 144178 528164 144184 528216
rect 144236 528164 144242 528216
rect 144196 528000 144224 528164
rect 151464 528000 151492 528244
rect 151722 528164 151728 528216
rect 151780 528204 151786 528216
rect 151780 528176 158944 528204
rect 151780 528164 151786 528176
rect 144196 527972 151492 528000
rect 158916 528000 158944 528176
rect 159284 528000 159312 528244
rect 162762 528232 162768 528284
rect 162820 528272 162826 528284
rect 175182 528272 175188 528284
rect 162820 528244 175188 528272
rect 162820 528232 162826 528244
rect 175182 528232 175188 528244
rect 175240 528232 175246 528284
rect 177960 528272 177988 528380
rect 182174 528272 182180 528284
rect 176028 528244 177804 528272
rect 177960 528244 182180 528272
rect 159358 528164 159364 528216
rect 159416 528164 159422 528216
rect 160370 528164 160376 528216
rect 160428 528204 160434 528216
rect 175918 528204 175924 528216
rect 160428 528176 175924 528204
rect 160428 528164 160434 528176
rect 175918 528164 175924 528176
rect 175976 528164 175982 528216
rect 159376 528136 159404 528164
rect 176028 528136 176056 528244
rect 159376 528108 176056 528136
rect 177776 528136 177804 528244
rect 182174 528232 182180 528244
rect 182232 528232 182238 528284
rect 177942 528164 177948 528216
rect 178000 528204 178006 528216
rect 182284 528204 182312 528448
rect 184198 528436 184204 528448
rect 184256 528436 184262 528488
rect 195422 528436 195428 528488
rect 195480 528476 195486 528488
rect 197998 528476 198004 528488
rect 195480 528448 198004 528476
rect 195480 528436 195486 528448
rect 197998 528436 198004 528448
rect 198056 528436 198062 528488
rect 234154 528436 234160 528488
rect 234212 528476 234218 528488
rect 235074 528476 235080 528488
rect 234212 528448 235080 528476
rect 234212 528436 234218 528448
rect 235074 528436 235080 528448
rect 235132 528436 235138 528488
rect 262214 528436 262220 528488
rect 262272 528476 262278 528488
rect 263042 528476 263048 528488
rect 262272 528448 263048 528476
rect 262272 528436 262278 528448
rect 263042 528436 263048 528448
rect 263100 528436 263106 528488
rect 318058 528436 318064 528488
rect 318116 528476 318122 528488
rect 322014 528476 322020 528488
rect 318116 528448 322020 528476
rect 318116 528436 318122 528448
rect 322014 528436 322020 528448
rect 322072 528436 322078 528488
rect 190362 528368 190368 528420
rect 190420 528408 190426 528420
rect 251818 528408 251824 528420
rect 190420 528380 251824 528408
rect 190420 528368 190426 528380
rect 251818 528368 251824 528380
rect 251876 528368 251882 528420
rect 253842 528368 253848 528420
rect 253900 528408 253906 528420
rect 324130 528408 324136 528420
rect 253900 528380 324136 528408
rect 253900 528368 253906 528380
rect 324130 528368 324136 528380
rect 324188 528368 324194 528420
rect 324222 528368 324228 528420
rect 324280 528408 324286 528420
rect 385678 528408 385684 528420
rect 324280 528380 385684 528408
rect 324280 528368 324286 528380
rect 385678 528368 385684 528380
rect 385736 528368 385742 528420
rect 184106 528340 184112 528352
rect 178000 528176 182312 528204
rect 182652 528312 184112 528340
rect 178000 528164 178006 528176
rect 182652 528136 182680 528312
rect 184106 528300 184112 528312
rect 184164 528300 184170 528352
rect 185946 528300 185952 528352
rect 186004 528340 186010 528352
rect 385770 528340 385776 528352
rect 186004 528312 385776 528340
rect 186004 528300 186010 528312
rect 385770 528300 385776 528312
rect 385828 528300 385834 528352
rect 177776 528108 182680 528136
rect 182744 528244 183692 528272
rect 182744 528000 182772 528244
rect 158916 527972 159036 528000
rect 159284 527972 182772 528000
rect 182836 528176 183600 528204
rect 159008 527932 159036 527972
rect 182836 527932 182864 528176
rect 159008 527904 168420 527932
rect 168392 527864 168420 527904
rect 177960 527904 182864 527932
rect 177960 527864 177988 527904
rect 168392 527836 177988 527864
rect 183572 527864 183600 528176
rect 183664 528000 183692 528244
rect 183922 528232 183928 528284
rect 183980 528272 183986 528284
rect 315206 528272 315212 528284
rect 183980 528244 315212 528272
rect 183980 528232 183986 528244
rect 315206 528232 315212 528244
rect 315264 528232 315270 528284
rect 319622 528232 319628 528284
rect 319680 528272 319686 528284
rect 323946 528272 323952 528284
rect 319680 528244 323952 528272
rect 319680 528232 319686 528244
rect 323946 528232 323952 528244
rect 324004 528232 324010 528284
rect 324222 528232 324228 528284
rect 324280 528272 324286 528284
rect 385954 528272 385960 528284
rect 324280 528244 385960 528272
rect 324280 528232 324286 528244
rect 385954 528232 385960 528244
rect 386012 528232 386018 528284
rect 184106 528164 184112 528216
rect 184164 528164 184170 528216
rect 184198 528164 184204 528216
rect 184256 528204 184262 528216
rect 195422 528204 195428 528216
rect 184256 528176 195428 528204
rect 184256 528164 184262 528176
rect 195422 528164 195428 528176
rect 195480 528164 195486 528216
rect 195716 528176 196112 528204
rect 184124 528136 184152 528164
rect 195716 528136 195744 528176
rect 184124 528108 195744 528136
rect 196084 528136 196112 528176
rect 197998 528164 198004 528216
rect 198056 528204 198062 528216
rect 207014 528204 207020 528216
rect 198056 528176 207020 528204
rect 198056 528164 198062 528176
rect 207014 528164 207020 528176
rect 207072 528164 207078 528216
rect 207566 528164 207572 528216
rect 207624 528204 207630 528216
rect 234154 528204 234160 528216
rect 207624 528176 234160 528204
rect 207624 528164 207630 528176
rect 234154 528164 234160 528176
rect 234212 528164 234218 528216
rect 234356 528176 234844 528204
rect 234356 528136 234384 528176
rect 196084 528108 234384 528136
rect 234816 528136 234844 528176
rect 235074 528164 235080 528216
rect 235132 528204 235138 528216
rect 251818 528204 251824 528216
rect 235132 528176 251824 528204
rect 235132 528164 235138 528176
rect 251818 528164 251824 528176
rect 251876 528164 251882 528216
rect 251910 528164 251916 528216
rect 251968 528164 251974 528216
rect 254210 528164 254216 528216
rect 254268 528164 254274 528216
rect 254302 528164 254308 528216
rect 254360 528204 254366 528216
rect 262214 528204 262220 528216
rect 254360 528176 262220 528204
rect 254360 528164 254366 528176
rect 262214 528164 262220 528176
rect 262272 528164 262278 528216
rect 262508 528176 262996 528204
rect 251928 528136 251956 528164
rect 234816 528108 251956 528136
rect 254228 528136 254256 528164
rect 262508 528136 262536 528176
rect 254228 528108 262536 528136
rect 262968 528136 262996 528176
rect 263042 528164 263048 528216
rect 263100 528204 263106 528216
rect 315390 528204 315396 528216
rect 263100 528176 315396 528204
rect 263100 528164 263106 528176
rect 315390 528164 315396 528176
rect 315448 528164 315454 528216
rect 320082 528164 320088 528216
rect 320140 528164 320146 528216
rect 322014 528164 322020 528216
rect 322072 528164 322078 528216
rect 324130 528164 324136 528216
rect 324188 528204 324194 528216
rect 385402 528204 385408 528216
rect 324188 528176 385408 528204
rect 324188 528164 324194 528176
rect 385402 528164 385408 528176
rect 385460 528164 385466 528216
rect 385862 528164 385868 528216
rect 385920 528164 385926 528216
rect 318058 528136 318064 528148
rect 262968 528108 318064 528136
rect 318058 528096 318064 528108
rect 318116 528096 318122 528148
rect 263612 528040 265480 528068
rect 263612 528000 263640 528040
rect 183664 527972 234568 528000
rect 202800 527904 210004 527932
rect 183572 527836 193168 527864
rect 193140 527660 193168 527836
rect 202800 527660 202828 527904
rect 209976 527864 210004 527904
rect 210160 527904 229692 527932
rect 210160 527864 210188 527904
rect 209976 527836 210188 527864
rect 193140 527632 202828 527660
rect 229664 527592 229692 527904
rect 234540 527660 234568 527972
rect 234908 527972 260972 528000
rect 234908 527660 234936 527972
rect 260944 527932 260972 527972
rect 261128 527972 263640 528000
rect 261128 527932 261156 527972
rect 234540 527632 234936 527660
rect 235000 527904 244320 527932
rect 235000 527592 235028 527904
rect 244292 527728 244320 527904
rect 252204 527904 260880 527932
rect 260944 527904 261156 527932
rect 265452 527932 265480 528040
rect 302142 528028 302148 528080
rect 302200 528068 302206 528080
rect 320100 528068 320128 528164
rect 322032 528136 322060 528164
rect 385880 528136 385908 528164
rect 322032 528108 385908 528136
rect 386156 528068 386184 528516
rect 398834 528504 398840 528516
rect 398892 528504 398898 528556
rect 398944 528544 398972 528584
rect 399128 528584 411260 528612
rect 399128 528544 399156 528584
rect 411254 528572 411260 528584
rect 411312 528572 411318 528624
rect 411438 528572 411444 528624
rect 411496 528612 411502 528624
rect 489270 528612 489276 528624
rect 411496 528584 489276 528612
rect 411496 528572 411502 528584
rect 489270 528572 489276 528584
rect 489328 528572 489334 528624
rect 398944 528516 399156 528544
rect 398926 528436 398932 528488
rect 398984 528476 398990 528488
rect 403618 528476 403624 528488
rect 398984 528448 403624 528476
rect 398984 528436 398990 528448
rect 403618 528436 403624 528448
rect 403676 528436 403682 528488
rect 403710 528436 403716 528488
rect 403768 528476 403774 528488
rect 408218 528476 408224 528488
rect 403768 528448 408224 528476
rect 403768 528436 403774 528448
rect 408218 528436 408224 528448
rect 408276 528436 408282 528488
rect 443362 528476 443368 528488
rect 442920 528448 443368 528476
rect 386230 528368 386236 528420
rect 386288 528408 386294 528420
rect 406286 528408 406292 528420
rect 386288 528380 406292 528408
rect 386288 528368 386294 528380
rect 406286 528368 406292 528380
rect 406344 528368 406350 528420
rect 422294 528408 422300 528420
rect 422220 528380 422300 528408
rect 422220 528352 422248 528380
rect 422294 528368 422300 528380
rect 422352 528368 422358 528420
rect 431862 528368 431868 528420
rect 431920 528408 431926 528420
rect 434714 528408 434720 528420
rect 431920 528380 434720 528408
rect 431920 528368 431926 528380
rect 434714 528368 434720 528380
rect 434772 528368 434778 528420
rect 434806 528368 434812 528420
rect 434864 528408 434870 528420
rect 442920 528408 442948 528448
rect 443362 528436 443368 528448
rect 443420 528436 443426 528488
rect 434864 528380 442948 528408
rect 434864 528368 434870 528380
rect 386322 528300 386328 528352
rect 386380 528340 386386 528352
rect 414934 528340 414940 528352
rect 386380 528312 414940 528340
rect 386380 528300 386386 528312
rect 414934 528300 414940 528312
rect 414992 528300 414998 528352
rect 422202 528300 422208 528352
rect 422260 528300 422266 528352
rect 386506 528232 386512 528284
rect 386564 528272 386570 528284
rect 434254 528272 434260 528284
rect 386564 528244 434260 528272
rect 386564 528232 386570 528244
rect 434254 528232 434260 528244
rect 434312 528232 434318 528284
rect 386414 528164 386420 528216
rect 386472 528164 386478 528216
rect 387334 528164 387340 528216
rect 387392 528204 387398 528216
rect 436462 528204 436468 528216
rect 387392 528176 436468 528204
rect 387392 528164 387398 528176
rect 436462 528164 436468 528176
rect 436520 528164 436526 528216
rect 442810 528164 442816 528216
rect 442868 528164 442874 528216
rect 443362 528164 443368 528216
rect 443420 528164 443426 528216
rect 444926 528164 444932 528216
rect 444984 528164 444990 528216
rect 452746 528164 452752 528216
rect 452804 528164 452810 528216
rect 386432 528136 386460 528164
rect 442828 528136 442856 528164
rect 386432 528108 386828 528136
rect 302200 528040 302372 528068
rect 320100 528040 386184 528068
rect 386800 528068 386828 528108
rect 405752 528108 442856 528136
rect 405752 528068 405780 528108
rect 386800 528040 405780 528068
rect 443380 528068 443408 528164
rect 444944 528068 444972 528164
rect 443380 528040 444972 528068
rect 302200 528028 302206 528040
rect 282822 527960 282828 528012
rect 282880 528000 282886 528012
rect 302234 528000 302240 528012
rect 282880 527972 302240 528000
rect 282880 527960 282886 527972
rect 302234 527960 302240 527972
rect 302292 527960 302298 528012
rect 265452 527904 274036 527932
rect 252204 527728 252232 527904
rect 260852 527864 260880 527904
rect 260852 527836 263640 527864
rect 244292 527700 252232 527728
rect 229664 527564 235028 527592
rect 263612 527592 263640 527836
rect 263612 527564 273944 527592
rect 273916 527388 273944 527564
rect 274008 527524 274036 527904
rect 278682 527892 278688 527944
rect 278740 527932 278746 527944
rect 288526 527932 288532 527944
rect 278740 527904 288532 527932
rect 278740 527892 278746 527904
rect 288526 527892 288532 527904
rect 288584 527892 288590 527944
rect 302142 527864 302148 527876
rect 292684 527836 302148 527864
rect 288526 527756 288532 527808
rect 288584 527796 288590 527808
rect 292684 527796 292712 527836
rect 302142 527824 302148 527836
rect 302200 527824 302206 527876
rect 302344 527864 302372 528040
rect 302418 527960 302424 528012
rect 302476 528000 302482 528012
rect 452764 528000 452792 528164
rect 302476 527972 452792 528000
rect 302476 527960 302482 527972
rect 315298 527864 315304 527876
rect 302344 527836 315304 527864
rect 315298 527824 315304 527836
rect 315356 527824 315362 527876
rect 288584 527768 292712 527796
rect 288584 527756 288590 527768
rect 282822 527524 282828 527536
rect 274008 527496 282828 527524
rect 282822 527484 282828 527496
rect 282880 527484 282886 527536
rect 278682 527388 278688 527400
rect 273916 527360 278688 527388
rect 278682 527348 278688 527360
rect 278740 527348 278746 527400
rect 282822 527076 282828 527128
rect 282880 527116 282886 527128
rect 283098 527116 283104 527128
rect 282880 527088 283104 527116
rect 282880 527076 282886 527088
rect 283098 527076 283104 527088
rect 283156 527076 283162 527128
rect 283006 511980 283012 512032
rect 283064 512020 283070 512032
rect 283098 512020 283104 512032
rect 283064 511992 283104 512020
rect 283064 511980 283070 511992
rect 283098 511980 283104 511992
rect 283156 511980 283162 512032
rect 2866 509260 2872 509312
rect 2924 509300 2930 509312
rect 15838 509300 15844 509312
rect 2924 509272 15844 509300
rect 2924 509260 2930 509272
rect 15838 509260 15844 509272
rect 15896 509260 15902 509312
rect 416590 503004 416596 503056
rect 416648 503044 416654 503056
rect 418154 503044 418160 503056
rect 416648 503016 418160 503044
rect 416648 503004 416654 503016
rect 418154 503004 418160 503016
rect 418212 503004 418218 503056
rect 418798 503004 418804 503056
rect 418856 503044 418862 503056
rect 420270 503044 420276 503056
rect 418856 503016 420276 503044
rect 418856 503004 418862 503016
rect 420270 503004 420276 503016
rect 420328 503004 420334 503056
rect 574002 503004 574008 503056
rect 574060 503044 574066 503056
rect 580442 503044 580448 503056
rect 574060 503016 580448 503044
rect 574060 503004 574066 503016
rect 580442 503004 580448 503016
rect 580500 503004 580506 503056
rect 412082 502936 412088 502988
rect 412140 502976 412146 502988
rect 580350 502976 580356 502988
rect 412140 502948 580356 502976
rect 412140 502936 412146 502948
rect 580350 502936 580356 502948
rect 580408 502936 580414 502988
rect 481266 502868 481272 502920
rect 481324 502908 481330 502920
rect 484302 502908 484308 502920
rect 481324 502880 484308 502908
rect 481324 502868 481330 502880
rect 484302 502868 484308 502880
rect 484360 502908 484366 502920
rect 487154 502908 487160 502920
rect 484360 502880 487160 502908
rect 484360 502868 484366 502880
rect 487154 502868 487160 502880
rect 487212 502868 487218 502920
rect 459462 502664 459468 502716
rect 459520 502704 459526 502716
rect 461210 502704 461216 502716
rect 459520 502676 461216 502704
rect 459520 502664 459526 502676
rect 461210 502664 461216 502676
rect 461268 502664 461274 502716
rect 282914 502324 282920 502376
rect 282972 502364 282978 502376
rect 283190 502364 283196 502376
rect 282972 502336 283196 502364
rect 282972 502324 282978 502336
rect 283190 502324 283196 502336
rect 283248 502324 283254 502376
rect 573358 502324 573364 502376
rect 573416 502364 573422 502376
rect 574002 502364 574008 502376
rect 573416 502336 574008 502364
rect 573416 502324 573422 502336
rect 574002 502324 574008 502336
rect 574060 502324 574066 502376
rect 417418 501576 417424 501628
rect 417476 501616 417482 501628
rect 580534 501616 580540 501628
rect 417476 501588 580540 501616
rect 417476 501576 417482 501588
rect 580534 501576 580540 501588
rect 580592 501576 580598 501628
rect 173894 501168 173900 501220
rect 173952 501208 173958 501220
rect 174814 501208 174820 501220
rect 173952 501180 174820 501208
rect 173952 501168 173958 501180
rect 174814 501168 174820 501180
rect 174872 501168 174878 501220
rect 183646 501168 183652 501220
rect 183704 501208 183710 501220
rect 184566 501208 184572 501220
rect 183704 501180 184572 501208
rect 183704 501168 183710 501180
rect 184566 501168 184572 501180
rect 184624 501168 184630 501220
rect 561674 501168 561680 501220
rect 561732 501208 561738 501220
rect 562594 501208 562600 501220
rect 561732 501180 562600 501208
rect 561732 501168 561738 501180
rect 562594 501168 562600 501180
rect 562652 501168 562658 501220
rect 27522 500896 27528 500948
rect 27580 500936 27586 500948
rect 29638 500936 29644 500948
rect 27580 500908 29644 500936
rect 27580 500896 27586 500908
rect 29638 500896 29644 500908
rect 29696 500896 29702 500948
rect 31662 500896 31668 500948
rect 31720 500936 31726 500948
rect 31754 500936 31760 500948
rect 31720 500908 31760 500936
rect 31720 500896 31726 500908
rect 31754 500896 31760 500908
rect 31812 500896 31818 500948
rect 51166 500896 51172 500948
rect 51224 500936 51230 500948
rect 52362 500936 52368 500948
rect 51224 500908 52368 500936
rect 51224 500896 51230 500908
rect 52362 500896 52368 500908
rect 52420 500896 52426 500948
rect 55490 500896 55496 500948
rect 55548 500936 55554 500948
rect 56502 500936 56508 500948
rect 55548 500908 56508 500936
rect 55548 500896 55554 500908
rect 56502 500896 56508 500908
rect 56560 500896 56566 500948
rect 95418 500896 95424 500948
rect 95476 500936 95482 500948
rect 96430 500936 96436 500948
rect 95476 500908 96436 500936
rect 95476 500896 95482 500908
rect 96430 500896 96436 500908
rect 96488 500896 96494 500948
rect 99650 500896 99656 500948
rect 99708 500936 99714 500948
rect 100662 500936 100668 500948
rect 99708 500908 100668 500936
rect 99708 500896 99714 500908
rect 100662 500896 100668 500908
rect 100720 500896 100726 500948
rect 100754 500896 100760 500948
rect 100812 500936 100818 500948
rect 102042 500936 102048 500948
rect 100812 500908 102048 500936
rect 100812 500896 100818 500908
rect 102042 500896 102048 500908
rect 102100 500896 102106 500948
rect 103974 500896 103980 500948
rect 104032 500936 104038 500948
rect 104802 500936 104808 500948
rect 104032 500908 104808 500936
rect 104032 500896 104038 500908
rect 104802 500896 104808 500908
rect 104860 500896 104866 500948
rect 105078 500896 105084 500948
rect 105136 500936 105142 500948
rect 106918 500936 106924 500948
rect 105136 500908 106924 500936
rect 105136 500896 105142 500908
rect 106918 500896 106924 500908
rect 106976 500896 106982 500948
rect 136266 500896 136272 500948
rect 136324 500936 136330 500948
rect 153654 500936 153660 500948
rect 136324 500908 153660 500936
rect 136324 500896 136330 500908
rect 153654 500896 153660 500908
rect 153712 500896 153718 500948
rect 194594 500896 194600 500948
rect 194652 500936 194658 500948
rect 195606 500936 195612 500948
rect 194652 500908 195612 500936
rect 194652 500896 194658 500908
rect 195606 500896 195612 500908
rect 195664 500896 195670 500948
rect 201494 500896 201500 500948
rect 201552 500936 201558 500948
rect 203150 500936 203156 500948
rect 201552 500908 203156 500936
rect 201552 500896 201558 500908
rect 203150 500896 203156 500908
rect 203208 500896 203214 500948
rect 204898 500896 204904 500948
rect 204956 500936 204962 500948
rect 208486 500936 208492 500948
rect 204956 500908 208492 500936
rect 204956 500896 204962 500908
rect 208486 500896 208492 500908
rect 208544 500896 208550 500948
rect 213822 500896 213828 500948
rect 213880 500936 213886 500948
rect 216030 500936 216036 500948
rect 213880 500908 216036 500936
rect 213880 500896 213886 500908
rect 216030 500896 216036 500908
rect 216088 500896 216094 500948
rect 223482 500896 223488 500948
rect 223540 500936 223546 500948
rect 224678 500936 224684 500948
rect 223540 500908 224684 500936
rect 223540 500896 223546 500908
rect 224678 500896 224684 500908
rect 224736 500896 224742 500948
rect 229094 500896 229100 500948
rect 229152 500936 229158 500948
rect 230106 500936 230112 500948
rect 229152 500908 230112 500936
rect 229152 500896 229158 500908
rect 230106 500896 230112 500908
rect 230164 500896 230170 500948
rect 233050 500896 233056 500948
rect 233108 500936 233114 500948
rect 234338 500936 234344 500948
rect 233108 500908 234344 500936
rect 233108 500896 233114 500908
rect 234338 500896 234344 500908
rect 234396 500896 234402 500948
rect 235902 500896 235908 500948
rect 235960 500936 235966 500948
rect 236546 500936 236552 500948
rect 235960 500908 236552 500936
rect 235960 500896 235966 500908
rect 236546 500896 236552 500908
rect 236604 500896 236610 500948
rect 251174 500896 251180 500948
rect 251232 500936 251238 500948
rect 253750 500936 253756 500948
rect 251232 500908 253756 500936
rect 251232 500896 251238 500908
rect 253750 500896 253756 500908
rect 253808 500896 253814 500948
rect 253934 500896 253940 500948
rect 253992 500936 253998 500948
rect 255958 500936 255964 500948
rect 253992 500908 255964 500936
rect 253992 500896 253998 500908
rect 255958 500896 255964 500908
rect 256016 500896 256022 500948
rect 262214 500896 262220 500948
rect 262272 500936 262278 500948
rect 263502 500936 263508 500948
rect 262272 500908 263508 500936
rect 262272 500896 262278 500908
rect 263502 500896 263508 500908
rect 263560 500896 263566 500948
rect 263594 500896 263600 500948
rect 263652 500936 263658 500948
rect 264514 500936 264520 500948
rect 263652 500908 264520 500936
rect 263652 500896 263658 500908
rect 264514 500896 264520 500908
rect 264572 500896 264578 500948
rect 269114 500896 269120 500948
rect 269172 500936 269178 500948
rect 269942 500936 269948 500948
rect 269172 500908 269948 500936
rect 269172 500896 269178 500908
rect 269942 500896 269948 500908
rect 270000 500896 270006 500948
rect 271966 500896 271972 500948
rect 272024 500936 272030 500948
rect 273162 500936 273168 500948
rect 272024 500908 273168 500936
rect 272024 500896 272030 500908
rect 273162 500896 273168 500908
rect 273220 500896 273226 500948
rect 277578 500896 277584 500948
rect 277636 500936 277642 500948
rect 278590 500936 278596 500948
rect 277636 500908 278596 500936
rect 277636 500896 277642 500908
rect 278590 500896 278596 500908
rect 278648 500896 278654 500948
rect 317322 500896 317328 500948
rect 317380 500936 317386 500948
rect 317874 500936 317880 500948
rect 317380 500908 317880 500936
rect 317380 500896 317386 500908
rect 317874 500896 317880 500908
rect 317932 500896 317938 500948
rect 340138 500896 340144 500948
rect 340196 500936 340202 500948
rect 340782 500936 340788 500948
rect 340196 500908 340788 500936
rect 340196 500896 340202 500908
rect 340782 500896 340788 500908
rect 340840 500896 340846 500948
rect 341150 500896 341156 500948
rect 341208 500936 341214 500948
rect 342070 500936 342076 500948
rect 341208 500908 342076 500936
rect 341208 500896 341214 500908
rect 342070 500896 342076 500908
rect 342128 500896 342134 500948
rect 343174 500896 343180 500948
rect 343232 500936 343238 500948
rect 343726 500936 343732 500948
rect 343232 500908 343732 500936
rect 343232 500896 343238 500908
rect 343726 500896 343732 500908
rect 343784 500896 343790 500948
rect 345474 500896 345480 500948
rect 345532 500936 345538 500948
rect 346210 500936 346216 500948
rect 345532 500908 346216 500936
rect 345532 500896 345538 500908
rect 346210 500896 346216 500908
rect 346268 500896 346274 500948
rect 349798 500896 349804 500948
rect 349856 500936 349862 500948
rect 350442 500936 350448 500948
rect 349856 500908 350448 500936
rect 349856 500896 349862 500908
rect 350442 500896 350448 500908
rect 350500 500896 350506 500948
rect 350902 500896 350908 500948
rect 350960 500936 350966 500948
rect 351822 500936 351828 500948
rect 350960 500908 351828 500936
rect 350960 500896 350966 500908
rect 351822 500896 351828 500908
rect 351880 500896 351886 500948
rect 354122 500896 354128 500948
rect 354180 500936 354186 500948
rect 354582 500936 354588 500948
rect 354180 500908 354588 500936
rect 354180 500896 354186 500908
rect 354582 500896 354588 500908
rect 354640 500896 354646 500948
rect 359458 500896 359464 500948
rect 359516 500936 359522 500948
rect 360102 500936 360108 500948
rect 359516 500908 360108 500936
rect 359516 500896 359522 500908
rect 360102 500896 360108 500908
rect 360160 500896 360166 500948
rect 364886 500896 364892 500948
rect 364944 500936 364950 500948
rect 365622 500936 365628 500948
rect 364944 500908 365628 500936
rect 364944 500896 364950 500908
rect 365622 500896 365628 500908
rect 365680 500896 365686 500948
rect 365990 500896 365996 500948
rect 366048 500936 366054 500948
rect 367002 500936 367008 500948
rect 366048 500908 367008 500936
rect 366048 500896 366054 500908
rect 367002 500896 367008 500908
rect 367060 500896 367066 500948
rect 375650 500896 375656 500948
rect 375708 500936 375714 500948
rect 376570 500936 376576 500948
rect 375708 500908 376576 500936
rect 375708 500896 375714 500908
rect 376570 500896 376576 500908
rect 376628 500896 376634 500948
rect 379974 500896 379980 500948
rect 380032 500936 380038 500948
rect 380710 500936 380716 500948
rect 380032 500908 380716 500936
rect 380032 500896 380038 500908
rect 380710 500896 380716 500908
rect 380768 500896 380774 500948
rect 384298 500896 384304 500948
rect 384356 500936 384362 500948
rect 384942 500936 384948 500948
rect 384356 500908 384948 500936
rect 384356 500896 384362 500908
rect 384942 500896 384948 500908
rect 385000 500896 385006 500948
rect 385402 500896 385408 500948
rect 385460 500936 385466 500948
rect 386322 500936 386328 500948
rect 385460 500908 386328 500936
rect 385460 500896 385466 500908
rect 386322 500896 386328 500908
rect 386380 500896 386386 500948
rect 400490 500896 400496 500948
rect 400548 500936 400554 500948
rect 401502 500936 401508 500948
rect 400548 500908 401508 500936
rect 400548 500896 400554 500908
rect 401502 500896 401508 500908
rect 401560 500896 401566 500948
rect 404722 500896 404728 500948
rect 404780 500936 404786 500948
rect 411622 500936 411628 500948
rect 404780 500908 411628 500936
rect 404780 500896 404786 500908
rect 411622 500896 411628 500908
rect 411680 500896 411686 500948
rect 420822 500896 420828 500948
rect 420880 500936 420886 500948
rect 423122 500936 423128 500948
rect 420880 500908 423128 500936
rect 420880 500896 420886 500908
rect 423122 500896 423128 500908
rect 423180 500936 423186 500948
rect 424962 500936 424968 500948
rect 423180 500908 424968 500936
rect 423180 500896 423186 500908
rect 424962 500896 424968 500908
rect 425020 500936 425026 500948
rect 427078 500936 427084 500948
rect 425020 500908 427084 500936
rect 425020 500896 425026 500908
rect 427078 500896 427084 500908
rect 427136 500936 427142 500948
rect 429286 500936 429292 500948
rect 427136 500908 429292 500936
rect 427136 500896 427142 500908
rect 429286 500896 429292 500908
rect 429344 500936 429350 500948
rect 431402 500936 431408 500948
rect 429344 500908 431408 500936
rect 429344 500896 429350 500908
rect 431402 500896 431408 500908
rect 431460 500936 431466 500948
rect 433426 500936 433432 500948
rect 431460 500908 433432 500936
rect 431460 500896 431466 500908
rect 433426 500896 433432 500908
rect 433484 500936 433490 500948
rect 435542 500936 435548 500948
rect 433484 500908 435548 500936
rect 433484 500896 433490 500908
rect 435542 500896 435548 500908
rect 435600 500936 435606 500948
rect 437566 500936 437572 500948
rect 435600 500908 437572 500936
rect 435600 500896 435606 500908
rect 437566 500896 437572 500908
rect 437624 500936 437630 500948
rect 439682 500936 439688 500948
rect 437624 500908 439688 500936
rect 437624 500896 437630 500908
rect 439682 500896 439688 500908
rect 439740 500936 439746 500948
rect 441982 500936 441988 500948
rect 439740 500908 441988 500936
rect 439740 500896 439746 500908
rect 441982 500896 441988 500908
rect 442040 500936 442046 500948
rect 444374 500936 444380 500948
rect 442040 500908 444380 500936
rect 442040 500896 442046 500908
rect 444374 500896 444380 500908
rect 444432 500936 444438 500948
rect 446306 500936 446312 500948
rect 444432 500908 446312 500936
rect 444432 500896 444438 500908
rect 446306 500896 446312 500908
rect 446364 500936 446370 500948
rect 448514 500936 448520 500948
rect 446364 500908 448520 500936
rect 446364 500896 446370 500908
rect 448514 500896 448520 500908
rect 448572 500936 448578 500948
rect 450446 500936 450452 500948
rect 448572 500908 450452 500936
rect 448572 500896 448578 500908
rect 450446 500896 450452 500908
rect 450504 500936 450510 500948
rect 453298 500936 453304 500948
rect 450504 500908 453304 500936
rect 450504 500896 450510 500908
rect 453298 500896 453304 500908
rect 453356 500936 453362 500948
rect 455322 500936 455328 500948
rect 453356 500908 455328 500936
rect 453356 500896 453362 500908
rect 455322 500896 455328 500908
rect 455380 500936 455386 500948
rect 457346 500936 457352 500948
rect 455380 500908 457352 500936
rect 455380 500896 455386 500908
rect 457346 500896 457352 500908
rect 457404 500936 457410 500948
rect 461854 500936 461860 500948
rect 457404 500908 461860 500936
rect 457404 500896 457410 500908
rect 461854 500896 461860 500908
rect 461912 500936 461918 500948
rect 464062 500936 464068 500948
rect 461912 500908 464068 500936
rect 461912 500896 461918 500908
rect 464062 500896 464068 500908
rect 464120 500936 464126 500948
rect 465902 500936 465908 500948
rect 464120 500908 465908 500936
rect 464120 500896 464126 500908
rect 465902 500896 465908 500908
rect 465960 500936 465966 500948
rect 468110 500936 468116 500948
rect 465960 500908 468116 500936
rect 465960 500896 465966 500908
rect 468110 500896 468116 500908
rect 468168 500936 468174 500948
rect 470226 500936 470232 500948
rect 468168 500908 470232 500936
rect 468168 500896 468174 500908
rect 470226 500896 470232 500908
rect 470284 500936 470290 500948
rect 472710 500936 472716 500948
rect 470284 500908 472716 500936
rect 470284 500896 470290 500908
rect 472710 500896 472716 500908
rect 472768 500936 472774 500948
rect 474642 500936 474648 500948
rect 472768 500908 474648 500936
rect 472768 500896 472774 500908
rect 474642 500896 474648 500908
rect 474700 500936 474706 500948
rect 477770 500936 477776 500948
rect 474700 500908 477776 500936
rect 474700 500896 474706 500908
rect 477770 500896 477776 500908
rect 477828 500936 477834 500948
rect 480806 500936 480812 500948
rect 477828 500908 480812 500936
rect 477828 500896 477834 500908
rect 480806 500896 480812 500908
rect 480864 500896 480870 500948
rect 502886 500896 502892 500948
rect 502944 500936 502950 500948
rect 503622 500936 503628 500948
rect 502944 500908 503628 500936
rect 502944 500896 502950 500908
rect 503622 500896 503628 500908
rect 503680 500896 503686 500948
rect 511442 500896 511448 500948
rect 511500 500936 511506 500948
rect 511902 500936 511908 500948
rect 511500 500908 511908 500936
rect 511500 500896 511506 500908
rect 511902 500896 511908 500908
rect 511960 500896 511966 500948
rect 516870 500896 516876 500948
rect 516928 500936 516934 500948
rect 517422 500936 517428 500948
rect 516928 500908 517428 500936
rect 516928 500896 516934 500908
rect 517422 500896 517428 500908
rect 517480 500896 517486 500948
rect 523310 500896 523316 500948
rect 523368 500936 523374 500948
rect 524322 500936 524328 500948
rect 523368 500908 524328 500936
rect 523368 500896 523374 500908
rect 524322 500896 524328 500908
rect 524380 500896 524386 500948
rect 545942 500896 545948 500948
rect 546000 500936 546006 500948
rect 552106 500936 552112 500948
rect 546000 500908 552112 500936
rect 546000 500896 546006 500908
rect 552106 500896 552112 500908
rect 552164 500896 552170 500948
rect 552382 500896 552388 500948
rect 552440 500936 552446 500948
rect 553486 500936 553492 500948
rect 552440 500908 553492 500936
rect 552440 500896 552446 500908
rect 553486 500896 553492 500908
rect 553544 500896 553550 500948
rect 45738 500828 45744 500880
rect 45796 500868 45802 500880
rect 53926 500868 53932 500880
rect 45796 500840 53932 500868
rect 45796 500828 45802 500840
rect 53926 500828 53932 500840
rect 53984 500828 53990 500880
rect 95326 500828 95332 500880
rect 95384 500868 95390 500880
rect 96522 500868 96528 500880
rect 95384 500840 96528 500868
rect 95384 500828 95390 500840
rect 96522 500828 96528 500840
rect 96580 500828 96586 500880
rect 137370 500828 137376 500880
rect 137428 500868 137434 500880
rect 155126 500868 155132 500880
rect 137428 500840 155132 500868
rect 137428 500828 137434 500840
rect 155126 500828 155132 500840
rect 155184 500828 155190 500880
rect 195054 500828 195060 500880
rect 195112 500868 195118 500880
rect 197722 500868 197728 500880
rect 195112 500840 197728 500868
rect 195112 500828 195118 500840
rect 197722 500828 197728 500840
rect 197780 500828 197786 500880
rect 205634 500828 205640 500880
rect 205692 500868 205698 500880
rect 209590 500868 209596 500880
rect 205692 500840 209596 500868
rect 205692 500828 205698 500840
rect 209590 500828 209596 500840
rect 209648 500828 209654 500880
rect 214650 500828 214656 500880
rect 214708 500868 214714 500880
rect 217134 500868 217140 500880
rect 214708 500840 217140 500868
rect 214708 500828 214714 500840
rect 217134 500828 217140 500840
rect 217192 500828 217198 500880
rect 403710 500828 403716 500880
rect 403768 500868 403774 500880
rect 409874 500868 409880 500880
rect 403768 500840 409880 500868
rect 403768 500828 403774 500840
rect 409874 500828 409880 500840
rect 409932 500828 409938 500880
rect 543642 500828 543648 500880
rect 543700 500868 543706 500880
rect 553762 500868 553768 500880
rect 543700 500840 553768 500868
rect 543700 500828 543706 500840
rect 553762 500828 553768 500840
rect 553820 500828 553826 500880
rect 80054 500760 80060 500812
rect 80112 500800 80118 500812
rect 81342 500800 81348 500812
rect 80112 500772 81348 500800
rect 80112 500760 80118 500772
rect 81342 500760 81348 500772
rect 81400 500760 81406 500812
rect 134150 500760 134156 500812
rect 134208 500800 134214 500812
rect 153838 500800 153844 500812
rect 134208 500772 153844 500800
rect 134208 500760 134214 500772
rect 153838 500760 153844 500772
rect 153896 500760 153902 500812
rect 191834 500760 191840 500812
rect 191892 500800 191898 500812
rect 199930 500800 199936 500812
rect 191892 500772 199936 500800
rect 191892 500760 191898 500772
rect 199930 500760 199936 500772
rect 199988 500760 199994 500812
rect 267734 500760 267740 500812
rect 267792 500800 267798 500812
rect 268838 500800 268844 500812
rect 267792 500772 268844 500800
rect 267792 500760 267798 500772
rect 268838 500760 268844 500772
rect 268896 500760 268902 500812
rect 355226 500760 355232 500812
rect 355284 500800 355290 500812
rect 355962 500800 355968 500812
rect 355284 500772 355968 500800
rect 355284 500760 355290 500772
rect 355962 500760 355968 500772
rect 356020 500760 356026 500812
rect 541618 500760 541624 500812
rect 541676 500800 541682 500812
rect 553854 500800 553860 500812
rect 541676 500772 553860 500800
rect 541676 500760 541682 500772
rect 553854 500760 553860 500772
rect 553912 500760 553918 500812
rect 41414 500692 41420 500744
rect 41472 500732 41478 500744
rect 47026 500732 47032 500744
rect 41472 500704 47032 500732
rect 41472 500692 41478 500704
rect 47026 500692 47032 500704
rect 47084 500692 47090 500744
rect 135254 500692 135260 500744
rect 135312 500732 135318 500744
rect 155310 500732 155316 500744
rect 135312 500704 155316 500732
rect 135312 500692 135318 500704
rect 155310 500692 155316 500704
rect 155368 500692 155374 500744
rect 224862 500692 224868 500744
rect 224920 500732 224926 500744
rect 225782 500732 225788 500744
rect 224920 500704 225788 500732
rect 224920 500692 224926 500704
rect 225782 500692 225788 500704
rect 225840 500692 225846 500744
rect 230474 500692 230480 500744
rect 230532 500732 230538 500744
rect 232222 500732 232228 500744
rect 230532 500704 232228 500732
rect 230532 500692 230538 500704
rect 232222 500692 232228 500704
rect 232280 500692 232286 500744
rect 320266 500692 320272 500744
rect 320324 500732 320330 500744
rect 321094 500732 321100 500744
rect 320324 500704 321100 500732
rect 320324 500692 320330 500704
rect 321094 500692 321100 500704
rect 321152 500692 321158 500744
rect 539502 500692 539508 500744
rect 539560 500732 539566 500744
rect 552014 500732 552020 500744
rect 539560 500704 552020 500732
rect 539560 500692 539566 500704
rect 552014 500692 552020 500704
rect 552072 500692 552078 500744
rect 552106 500692 552112 500744
rect 552164 500732 552170 500744
rect 553670 500732 553676 500744
rect 552164 500704 553676 500732
rect 552164 500692 552170 500704
rect 553670 500692 553676 500704
rect 553728 500692 553734 500744
rect 131942 500624 131948 500676
rect 132000 500664 132006 500676
rect 155494 500664 155500 500676
rect 132000 500636 155500 500664
rect 132000 500624 132006 500636
rect 155494 500624 155500 500636
rect 155552 500624 155558 500676
rect 191926 500624 191932 500676
rect 191984 500664 191990 500676
rect 196618 500664 196624 500676
rect 191984 500636 196624 500664
rect 191984 500624 191990 500636
rect 196618 500624 196624 500636
rect 196676 500624 196682 500676
rect 197170 500624 197176 500676
rect 197228 500664 197234 500676
rect 202046 500664 202052 500676
rect 197228 500636 202052 500664
rect 197228 500624 197234 500636
rect 202046 500624 202052 500636
rect 202104 500624 202110 500676
rect 258258 500624 258264 500676
rect 258316 500664 258322 500676
rect 260282 500664 260288 500676
rect 258316 500636 260288 500664
rect 258316 500624 258322 500636
rect 260282 500624 260288 500636
rect 260340 500624 260346 500676
rect 260834 500624 260840 500676
rect 260892 500664 260898 500676
rect 262398 500664 262404 500676
rect 260892 500636 262404 500664
rect 260892 500624 260898 500636
rect 262398 500624 262404 500636
rect 262456 500624 262462 500676
rect 360562 500624 360568 500676
rect 360620 500664 360626 500676
rect 361390 500664 361396 500676
rect 360620 500636 361396 500664
rect 360620 500624 360626 500636
rect 361390 500624 361396 500636
rect 361448 500624 361454 500676
rect 370314 500624 370320 500676
rect 370372 500664 370378 500676
rect 371050 500664 371056 500676
rect 370372 500636 371056 500664
rect 370372 500624 370378 500636
rect 371050 500624 371056 500636
rect 371108 500624 371114 500676
rect 512546 500624 512552 500676
rect 512604 500664 512610 500676
rect 513282 500664 513288 500676
rect 512604 500636 513288 500664
rect 512604 500624 512610 500636
rect 513282 500624 513288 500636
rect 513340 500624 513346 500676
rect 513650 500624 513656 500676
rect 513708 500664 513714 500676
rect 514662 500664 514668 500676
rect 513708 500636 514668 500664
rect 513708 500624 513714 500636
rect 514662 500624 514668 500636
rect 514720 500624 514726 500676
rect 537294 500624 537300 500676
rect 537352 500664 537358 500676
rect 553946 500664 553952 500676
rect 537352 500636 553952 500664
rect 537352 500624 537358 500636
rect 553946 500624 553952 500636
rect 554004 500624 554010 500676
rect 129826 500556 129832 500608
rect 129884 500596 129890 500608
rect 154758 500596 154764 500608
rect 129884 500568 154764 500596
rect 129884 500556 129890 500568
rect 154758 500556 154764 500568
rect 154816 500556 154822 500608
rect 201586 500556 201592 500608
rect 201644 500596 201650 500608
rect 206370 500596 206376 500608
rect 201644 500568 206376 500596
rect 201644 500556 201650 500568
rect 206370 500556 206376 500568
rect 206428 500556 206434 500608
rect 207106 500556 207112 500608
rect 207164 500596 207170 500608
rect 211706 500596 211712 500608
rect 207164 500568 211712 500596
rect 207164 500556 207170 500568
rect 211706 500556 211712 500568
rect 211764 500556 211770 500608
rect 215386 500556 215392 500608
rect 215444 500596 215450 500608
rect 219250 500596 219256 500608
rect 215444 500568 219256 500596
rect 215444 500556 215450 500568
rect 219250 500556 219256 500568
rect 219308 500556 219314 500608
rect 219526 500556 219532 500608
rect 219584 500596 219590 500608
rect 222562 500596 222568 500608
rect 219584 500568 222568 500596
rect 219584 500556 219590 500568
rect 222562 500556 222568 500568
rect 222620 500556 222626 500608
rect 535178 500556 535184 500608
rect 535236 500596 535242 500608
rect 554038 500596 554044 500608
rect 535236 500568 554044 500596
rect 535236 500556 535242 500568
rect 554038 500556 554044 500568
rect 554096 500556 554102 500608
rect 20622 500488 20628 500540
rect 20680 500528 20686 500540
rect 25314 500528 25320 500540
rect 20680 500500 25320 500528
rect 20680 500488 20686 500500
rect 25314 500488 25320 500500
rect 25372 500488 25378 500540
rect 97534 500488 97540 500540
rect 97592 500528 97598 500540
rect 115198 500528 115204 500540
rect 97592 500500 115204 500528
rect 97592 500488 97598 500500
rect 115198 500488 115204 500500
rect 115256 500488 115262 500540
rect 127710 500488 127716 500540
rect 127768 500528 127774 500540
rect 154850 500528 154856 500540
rect 127768 500500 154856 500528
rect 127768 500488 127774 500500
rect 154850 500488 154856 500500
rect 154908 500488 154914 500540
rect 196434 500488 196440 500540
rect 196492 500528 196498 500540
rect 200942 500528 200948 500540
rect 196492 500500 200948 500528
rect 196492 500488 196498 500500
rect 200942 500488 200948 500500
rect 201000 500488 201006 500540
rect 257522 500488 257528 500540
rect 257580 500528 257586 500540
rect 259178 500528 259184 500540
rect 257580 500500 259184 500528
rect 257580 500488 257586 500500
rect 259178 500488 259184 500500
rect 259236 500488 259242 500540
rect 363782 500488 363788 500540
rect 363840 500528 363846 500540
rect 364242 500528 364248 500540
rect 363840 500500 364248 500528
rect 363840 500488 363846 500500
rect 364242 500488 364248 500500
rect 364300 500488 364306 500540
rect 369210 500488 369216 500540
rect 369268 500528 369274 500540
rect 369762 500528 369768 500540
rect 369268 500500 369768 500528
rect 369268 500488 369274 500500
rect 369762 500488 369768 500500
rect 369820 500488 369826 500540
rect 531958 500488 531964 500540
rect 532016 500528 532022 500540
rect 532602 500528 532608 500540
rect 532016 500500 532608 500528
rect 532016 500488 532022 500500
rect 532602 500488 532608 500500
rect 532660 500488 532666 500540
rect 533062 500488 533068 500540
rect 533120 500528 533126 500540
rect 551186 500528 551192 500540
rect 533120 500500 551192 500528
rect 533120 500488 533126 500500
rect 551186 500488 551192 500500
rect 551244 500488 551250 500540
rect 551370 500488 551376 500540
rect 551428 500528 551434 500540
rect 551922 500528 551928 500540
rect 551428 500500 551928 500528
rect 551428 500488 551434 500500
rect 551922 500488 551928 500500
rect 551980 500488 551986 500540
rect 22094 500420 22100 500472
rect 22152 500460 22158 500472
rect 23382 500460 23388 500472
rect 22152 500432 23388 500460
rect 22152 500420 22158 500432
rect 23382 500420 23388 500432
rect 23440 500420 23446 500472
rect 42518 500420 42524 500472
rect 42576 500460 42582 500472
rect 47578 500460 47584 500472
rect 42576 500432 47584 500460
rect 42576 500420 42582 500432
rect 47578 500420 47584 500432
rect 47636 500420 47642 500472
rect 93210 500420 93216 500472
rect 93268 500460 93274 500472
rect 113818 500460 113824 500472
rect 93268 500432 113824 500460
rect 93268 500420 93274 500432
rect 113818 500420 113824 500432
rect 113876 500420 113882 500472
rect 125502 500420 125508 500472
rect 125560 500460 125566 500472
rect 155218 500460 155224 500472
rect 125560 500432 155224 500460
rect 125560 500420 125566 500432
rect 155218 500420 155224 500432
rect 155276 500420 155282 500472
rect 187418 500420 187424 500472
rect 187476 500460 187482 500472
rect 192386 500460 192392 500472
rect 187476 500432 192392 500460
rect 187476 500420 187482 500432
rect 192386 500420 192392 500432
rect 192444 500420 192450 500472
rect 203886 500420 203892 500472
rect 203944 500460 203950 500472
rect 207474 500460 207480 500472
rect 203944 500432 207480 500460
rect 203944 500420 203950 500432
rect 207474 500420 207480 500432
rect 207532 500420 207538 500472
rect 211154 500420 211160 500472
rect 211212 500460 211218 500472
rect 215018 500460 215024 500472
rect 211212 500432 215024 500460
rect 211212 500420 211218 500432
rect 215018 500420 215024 500432
rect 215076 500420 215082 500472
rect 218146 500420 218152 500472
rect 218204 500460 218210 500472
rect 221458 500460 221464 500472
rect 218204 500432 221464 500460
rect 218204 500420 218210 500432
rect 221458 500420 221464 500432
rect 221516 500420 221522 500472
rect 224218 500420 224224 500472
rect 224276 500460 224282 500472
rect 226794 500460 226800 500472
rect 224276 500432 226800 500460
rect 224276 500420 224282 500432
rect 226794 500420 226800 500432
rect 226852 500420 226858 500472
rect 528462 500420 528468 500472
rect 528520 500460 528526 500472
rect 528520 500432 551416 500460
rect 528520 500420 528526 500432
rect 551388 500404 551416 500432
rect 43622 500352 43628 500404
rect 43680 500392 43686 500404
rect 48958 500392 48964 500404
rect 43680 500364 48964 500392
rect 43680 500352 43686 500364
rect 48958 500352 48964 500364
rect 49016 500352 49022 500404
rect 88886 500352 88892 500404
rect 88944 500392 88950 500404
rect 112438 500392 112444 500404
rect 88944 500364 112444 500392
rect 88944 500352 88950 500364
rect 112438 500352 112444 500364
rect 112496 500352 112502 500404
rect 123386 500352 123392 500404
rect 123444 500392 123450 500404
rect 154942 500392 154948 500404
rect 123444 500364 154948 500392
rect 123444 500352 123450 500364
rect 154942 500352 154948 500364
rect 155000 500352 155006 500404
rect 187602 500352 187608 500404
rect 187660 500392 187666 500404
rect 193398 500392 193404 500404
rect 187660 500364 193404 500392
rect 187660 500352 187666 500364
rect 193398 500352 193404 500364
rect 193456 500352 193462 500404
rect 209130 500352 209136 500404
rect 209188 500392 209194 500404
rect 212810 500392 212816 500404
rect 209188 500364 212816 500392
rect 209188 500352 209194 500364
rect 212810 500352 212816 500364
rect 212868 500352 212874 500404
rect 215202 500352 215208 500404
rect 215260 500392 215266 500404
rect 218238 500392 218244 500404
rect 215260 500364 218244 500392
rect 215260 500352 215266 500364
rect 218238 500352 218244 500364
rect 218296 500352 218302 500404
rect 322842 500352 322848 500404
rect 322900 500392 322906 500404
rect 323302 500392 323308 500404
rect 322900 500364 323308 500392
rect 322900 500352 322906 500364
rect 323302 500352 323308 500364
rect 323360 500352 323366 500404
rect 398282 500352 398288 500404
rect 398340 500392 398346 500404
rect 398742 500392 398748 500404
rect 398340 500364 398748 500392
rect 398340 500352 398346 500364
rect 398742 500352 398748 500364
rect 398800 500352 398806 500404
rect 497458 500352 497464 500404
rect 497516 500392 497522 500404
rect 498102 500392 498108 500404
rect 497516 500364 498108 500392
rect 497516 500352 497522 500364
rect 498102 500352 498108 500364
rect 498160 500352 498166 500404
rect 507118 500352 507124 500404
rect 507176 500392 507182 500404
rect 507762 500392 507768 500404
rect 507176 500364 507768 500392
rect 507176 500352 507182 500364
rect 507762 500352 507768 500364
rect 507820 500352 507826 500404
rect 526530 500352 526536 500404
rect 526588 500392 526594 500404
rect 551278 500392 551284 500404
rect 526588 500364 551284 500392
rect 526588 500352 526594 500364
rect 551278 500352 551284 500364
rect 551336 500352 551342 500404
rect 551370 500352 551376 500404
rect 551428 500352 551434 500404
rect 555050 500392 555056 500404
rect 551480 500364 555056 500392
rect 44726 500284 44732 500336
rect 44784 500324 44790 500336
rect 52546 500324 52552 500336
rect 44784 500296 52552 500324
rect 44784 500284 44790 500296
rect 52546 500284 52552 500296
rect 52604 500284 52610 500336
rect 84562 500284 84568 500336
rect 84620 500324 84626 500336
rect 109678 500324 109684 500336
rect 84620 500296 109684 500324
rect 84620 500284 84626 500296
rect 109678 500284 109684 500296
rect 109736 500284 109742 500336
rect 121178 500284 121184 500336
rect 121236 500324 121242 500336
rect 153286 500324 153292 500336
rect 121236 500296 153292 500324
rect 121236 500284 121242 500296
rect 153286 500284 153292 500296
rect 153344 500284 153350 500336
rect 195882 500284 195888 500336
rect 195940 500324 195946 500336
rect 198826 500324 198832 500336
rect 195940 500296 198832 500324
rect 195940 500284 195946 500296
rect 198826 500284 198832 500296
rect 198884 500284 198890 500336
rect 199470 500284 199476 500336
rect 199528 500324 199534 500336
rect 204162 500324 204168 500336
rect 199528 500296 204168 500324
rect 199528 500284 199534 500296
rect 204162 500284 204168 500296
rect 204220 500284 204226 500336
rect 209866 500284 209872 500336
rect 209924 500324 209930 500336
rect 213914 500324 213920 500336
rect 209924 500296 213920 500324
rect 209924 500284 209930 500296
rect 213914 500284 213920 500296
rect 213972 500284 213978 500336
rect 255314 500284 255320 500336
rect 255372 500324 255378 500336
rect 256970 500324 256976 500336
rect 255372 500296 256976 500324
rect 255372 500284 255378 500296
rect 256970 500284 256976 500296
rect 257028 500284 257034 500336
rect 524230 500284 524236 500336
rect 524288 500324 524294 500336
rect 547966 500324 547972 500336
rect 524288 500296 547972 500324
rect 524288 500284 524294 500296
rect 547966 500284 547972 500296
rect 548024 500284 548030 500336
rect 551480 500324 551508 500364
rect 555050 500352 555056 500364
rect 555108 500352 555114 500404
rect 548076 500296 551508 500324
rect 80238 500216 80244 500268
rect 80296 500256 80302 500268
rect 108298 500256 108304 500268
rect 80296 500228 108304 500256
rect 80296 500216 80302 500228
rect 108298 500216 108304 500228
rect 108356 500216 108362 500268
rect 120166 500216 120172 500268
rect 120224 500256 120230 500268
rect 153378 500256 153384 500268
rect 120224 500228 153384 500256
rect 120224 500216 120230 500228
rect 153378 500216 153384 500228
rect 153436 500216 153442 500268
rect 187510 500216 187516 500268
rect 187568 500256 187574 500268
rect 194502 500256 194508 500268
rect 187568 500228 194508 500256
rect 187568 500216 187574 500228
rect 194502 500216 194508 500228
rect 194560 500216 194566 500268
rect 259454 500216 259460 500268
rect 259512 500256 259518 500268
rect 261294 500256 261300 500268
rect 259512 500228 261300 500256
rect 259512 500216 259518 500228
rect 261294 500216 261300 500228
rect 261352 500216 261358 500268
rect 289722 500216 289728 500268
rect 289780 500256 289786 500268
rect 416130 500256 416136 500268
rect 289780 500228 416136 500256
rect 289780 500216 289786 500228
rect 416130 500216 416136 500228
rect 416188 500216 416194 500268
rect 498562 500216 498568 500268
rect 498620 500256 498626 500268
rect 499482 500256 499488 500268
rect 498620 500228 499488 500256
rect 498620 500216 498626 500228
rect 499482 500216 499488 500228
rect 499540 500216 499546 500268
rect 522206 500216 522212 500268
rect 522264 500256 522270 500268
rect 548076 500256 548104 500296
rect 553302 500284 553308 500336
rect 553360 500324 553366 500336
rect 554222 500324 554228 500336
rect 553360 500296 554228 500324
rect 553360 500284 553366 500296
rect 554222 500284 554228 500296
rect 554280 500284 554286 500336
rect 522264 500228 548104 500256
rect 522264 500216 522270 500228
rect 548150 500216 548156 500268
rect 548208 500256 548214 500268
rect 553578 500256 553584 500268
rect 548208 500228 553584 500256
rect 548208 500216 548214 500228
rect 553578 500216 553584 500228
rect 553636 500216 553642 500268
rect 556798 500216 556804 500268
rect 556856 500256 556862 500268
rect 571334 500256 571340 500268
rect 556856 500228 571340 500256
rect 556856 500216 556862 500228
rect 571334 500216 571340 500228
rect 571392 500216 571398 500268
rect 61930 500148 61936 500200
rect 61988 500188 61994 500200
rect 61988 500160 70440 500188
rect 61988 500148 61994 500160
rect 70412 500120 70440 500160
rect 138474 500148 138480 500200
rect 138532 500188 138538 500200
rect 146846 500188 146852 500200
rect 138532 500160 146852 500188
rect 138532 500148 138538 500160
rect 146846 500148 146852 500160
rect 146904 500148 146910 500200
rect 527634 500148 527640 500200
rect 527692 500188 527698 500200
rect 528462 500188 528468 500200
rect 527692 500160 528468 500188
rect 527692 500148 527698 500160
rect 528462 500148 528468 500160
rect 528520 500148 528526 500200
rect 536282 500148 536288 500200
rect 536340 500188 536346 500200
rect 536742 500188 536748 500200
rect 536340 500160 536748 500188
rect 536340 500148 536346 500160
rect 536742 500148 536748 500160
rect 536800 500148 536806 500200
rect 547046 500148 547052 500200
rect 547104 500188 547110 500200
rect 552658 500188 552664 500200
rect 547104 500160 552664 500188
rect 547104 500148 547110 500160
rect 552658 500148 552664 500160
rect 552716 500148 552722 500200
rect 80238 500120 80244 500132
rect 70412 500092 80244 500120
rect 80238 500080 80244 500092
rect 80296 500080 80302 500132
rect 139486 500080 139492 500132
rect 139544 500120 139550 500132
rect 155034 500120 155040 500132
rect 139544 500092 155040 500120
rect 139544 500080 139550 500092
rect 155034 500080 155040 500092
rect 155092 500080 155098 500132
rect 220814 500080 220820 500132
rect 220872 500120 220878 500132
rect 223574 500120 223580 500132
rect 220872 500092 223580 500120
rect 220872 500080 220878 500092
rect 223574 500080 223580 500092
rect 223632 500080 223638 500132
rect 547966 500080 547972 500132
rect 548024 500120 548030 500132
rect 554958 500120 554964 500132
rect 548024 500092 554964 500120
rect 548024 500080 548030 500092
rect 554958 500080 554964 500092
rect 555016 500080 555022 500132
rect 140590 500012 140596 500064
rect 140648 500052 140654 500064
rect 153746 500052 153752 500064
rect 140648 500024 153752 500052
rect 140648 500012 140654 500024
rect 153746 500012 153752 500024
rect 153804 500012 153810 500064
rect 551186 500012 551192 500064
rect 551244 500052 551250 500064
rect 555418 500052 555424 500064
rect 551244 500024 555424 500052
rect 551244 500012 551250 500024
rect 555418 500012 555424 500024
rect 555476 500012 555482 500064
rect 142798 499944 142804 499996
rect 142856 499984 142862 499996
rect 154022 499984 154028 499996
rect 142856 499956 154028 499984
rect 142856 499944 142862 499956
rect 154022 499944 154028 499956
rect 154080 499944 154086 499996
rect 223574 499944 223580 499996
rect 223632 499984 223638 499996
rect 229002 499984 229008 499996
rect 223632 499956 229008 499984
rect 223632 499944 223638 499956
rect 229002 499944 229008 499956
rect 229060 499944 229066 499996
rect 374546 499944 374552 499996
rect 374604 499984 374610 499996
rect 375282 499984 375288 499996
rect 374604 499956 375288 499984
rect 374604 499944 374610 499956
rect 375282 499944 375288 499956
rect 375340 499944 375346 499996
rect 378870 499944 378876 499996
rect 378928 499984 378934 499996
rect 379422 499984 379428 499996
rect 378928 499956 379428 499984
rect 378928 499944 378934 499956
rect 379422 499944 379428 499956
rect 379480 499944 379486 499996
rect 389634 499944 389640 499996
rect 389692 499984 389698 499996
rect 390462 499984 390468 499996
rect 389692 499956 390468 499984
rect 389692 499944 389698 499956
rect 390462 499944 390468 499956
rect 390520 499944 390526 499996
rect 393958 499944 393964 499996
rect 394016 499984 394022 499996
rect 394602 499984 394608 499996
rect 394016 499956 394608 499984
rect 394016 499944 394022 499956
rect 394602 499944 394608 499956
rect 394660 499944 394666 499996
rect 395062 499944 395068 499996
rect 395120 499984 395126 499996
rect 395890 499984 395896 499996
rect 395120 499956 395896 499984
rect 395120 499944 395126 499956
rect 395890 499944 395896 499956
rect 395948 499944 395954 499996
rect 399386 499944 399392 499996
rect 399444 499984 399450 499996
rect 400122 499984 400128 499996
rect 399444 499956 400128 499984
rect 399444 499944 399450 499956
rect 400122 499944 400128 499956
rect 400180 499944 400186 499996
rect 501782 499944 501788 499996
rect 501840 499984 501846 499996
rect 502242 499984 502248 499996
rect 501840 499956 502248 499984
rect 501840 499944 501846 499956
rect 502242 499944 502248 499956
rect 502300 499944 502306 499996
rect 388622 499876 388628 499928
rect 388680 499916 388686 499928
rect 389082 499916 389088 499928
rect 388680 499888 389088 499916
rect 388680 499876 388686 499888
rect 389082 499876 389088 499888
rect 389140 499876 389146 499928
rect 92106 499808 92112 499860
rect 92164 499848 92170 499860
rect 93762 499848 93768 499860
rect 92164 499820 93768 499848
rect 92164 499808 92170 499820
rect 93762 499808 93768 499820
rect 93820 499808 93826 499860
rect 344370 499808 344376 499860
rect 344428 499848 344434 499860
rect 344922 499848 344928 499860
rect 344428 499820 344928 499848
rect 344428 499808 344434 499820
rect 344922 499808 344928 499820
rect 344980 499808 344986 499860
rect 50062 499740 50068 499792
rect 50120 499780 50126 499792
rect 50982 499780 50988 499792
rect 50120 499752 50988 499780
rect 50120 499740 50126 499752
rect 50982 499740 50988 499752
rect 51040 499740 51046 499792
rect 144914 499740 144920 499792
rect 144972 499780 144978 499792
rect 153930 499780 153936 499792
rect 144972 499752 153936 499780
rect 144972 499740 144978 499752
rect 153930 499740 153936 499752
rect 153988 499740 153994 499792
rect 200114 499740 200120 499792
rect 200172 499780 200178 499792
rect 205266 499780 205272 499792
rect 200172 499752 205272 499780
rect 200172 499740 200178 499752
rect 205266 499740 205272 499752
rect 205324 499740 205330 499792
rect 234522 499740 234528 499792
rect 234580 499780 234586 499792
rect 235442 499780 235448 499792
rect 234580 499752 235448 499780
rect 234580 499740 234586 499752
rect 235442 499740 235448 499752
rect 235500 499740 235506 499792
rect 206370 499672 206376 499724
rect 206428 499712 206434 499724
rect 210694 499712 210700 499724
rect 206428 499684 210700 499712
rect 206428 499672 206434 499684
rect 210694 499672 210700 499684
rect 210752 499672 210758 499724
rect 216674 499604 216680 499656
rect 216732 499644 216738 499656
rect 220354 499644 220360 499656
rect 216732 499616 220360 499644
rect 216732 499604 216738 499616
rect 220354 499604 220360 499616
rect 220412 499604 220418 499656
rect 252646 499604 252652 499656
rect 252704 499644 252710 499656
rect 254854 499644 254860 499656
rect 252704 499616 254860 499644
rect 252704 499604 252710 499616
rect 254854 499604 254860 499616
rect 254912 499604 254918 499656
rect 24762 499536 24768 499588
rect 24820 499576 24826 499588
rect 27430 499576 27436 499588
rect 24820 499548 27436 499576
rect 24820 499536 24826 499548
rect 27430 499536 27436 499548
rect 27488 499536 27494 499588
rect 32030 499536 32036 499588
rect 32088 499576 32094 499588
rect 32858 499576 32864 499588
rect 32088 499548 32864 499576
rect 32088 499536 32094 499548
rect 32858 499536 32864 499548
rect 32916 499536 32922 499588
rect 34974 499536 34980 499588
rect 35032 499576 35038 499588
rect 35802 499576 35808 499588
rect 35032 499548 35808 499576
rect 35032 499536 35038 499548
rect 35802 499536 35808 499548
rect 35860 499536 35866 499588
rect 36078 499536 36084 499588
rect 36136 499576 36142 499588
rect 37182 499576 37188 499588
rect 36136 499548 37188 499576
rect 36136 499536 36142 499548
rect 37182 499536 37188 499548
rect 37240 499536 37246 499588
rect 40402 499536 40408 499588
rect 40460 499576 40466 499588
rect 41322 499576 41328 499588
rect 40460 499548 41328 499576
rect 40460 499536 40466 499548
rect 41322 499536 41328 499548
rect 41380 499536 41386 499588
rect 60826 499536 60832 499588
rect 60884 499576 60890 499588
rect 62022 499576 62028 499588
rect 60884 499548 62028 499576
rect 60884 499536 60890 499548
rect 62022 499536 62028 499548
rect 62080 499536 62086 499588
rect 65150 499536 65156 499588
rect 65208 499576 65214 499588
rect 66162 499576 66168 499588
rect 65208 499548 66168 499576
rect 65208 499536 65214 499548
rect 66162 499536 66168 499548
rect 66220 499536 66226 499588
rect 69474 499536 69480 499588
rect 69532 499576 69538 499588
rect 70302 499576 70308 499588
rect 69532 499548 70308 499576
rect 69532 499536 69538 499548
rect 70302 499536 70308 499548
rect 70360 499536 70366 499588
rect 71774 499536 71780 499588
rect 71832 499576 71838 499588
rect 72694 499576 72700 499588
rect 71832 499548 72700 499576
rect 71832 499536 71838 499548
rect 72694 499536 72700 499548
rect 72752 499536 72758 499588
rect 75914 499536 75920 499588
rect 75972 499576 75978 499588
rect 77202 499576 77208 499588
rect 75972 499548 77208 499576
rect 75972 499536 75978 499548
rect 77202 499536 77208 499548
rect 77260 499536 77266 499588
rect 247034 499536 247040 499588
rect 247092 499576 247098 499588
rect 249426 499576 249432 499588
rect 247092 499548 249432 499576
rect 247092 499536 247098 499548
rect 249426 499536 249432 499548
rect 249484 499536 249490 499588
rect 256786 499536 256792 499588
rect 256844 499576 256850 499588
rect 258074 499576 258080 499588
rect 256844 499548 258080 499576
rect 256844 499536 256850 499548
rect 258074 499536 258080 499548
rect 258132 499536 258138 499588
rect 266538 499536 266544 499588
rect 266596 499576 266602 499588
rect 267826 499576 267832 499588
rect 266596 499548 267832 499576
rect 266596 499536 266602 499548
rect 267826 499536 267832 499548
rect 267884 499536 267890 499588
rect 560938 499536 560944 499588
rect 560996 499576 561002 499588
rect 567194 499576 567200 499588
rect 560996 499548 567200 499576
rect 560996 499536 561002 499548
rect 567194 499536 567200 499548
rect 567252 499536 567258 499588
rect 164234 499128 164240 499180
rect 164292 499168 164298 499180
rect 165062 499168 165068 499180
rect 164292 499140 165068 499168
rect 164292 499128 164298 499140
rect 165062 499128 165068 499140
rect 165120 499128 165126 499180
rect 80054 498856 80060 498908
rect 80112 498896 80118 498908
rect 113174 498896 113180 498908
rect 80112 498868 113180 498896
rect 80112 498856 80118 498868
rect 113174 498856 113180 498868
rect 113232 498856 113238 498908
rect 66254 498788 66260 498840
rect 66312 498828 66318 498840
rect 88334 498828 88340 498840
rect 66312 498800 88340 498828
rect 66312 498788 66318 498800
rect 88334 498788 88340 498800
rect 88392 498788 88398 498840
rect 89806 498788 89812 498840
rect 89864 498828 89870 498840
rect 126974 498828 126980 498840
rect 89864 498800 126980 498828
rect 89864 498788 89870 498800
rect 126974 498788 126980 498800
rect 127032 498788 127038 498840
rect 194594 498788 194600 498840
rect 194652 498828 194658 498840
rect 280154 498828 280160 498840
rect 194652 498800 280160 498828
rect 194652 498788 194658 498800
rect 280154 498788 280160 498800
rect 280212 498788 280218 498840
rect 501598 498788 501604 498840
rect 501656 498828 501662 498840
rect 574094 498828 574100 498840
rect 501656 498800 574100 498828
rect 501656 498788 501662 498800
rect 574094 498788 574100 498800
rect 574152 498788 574158 498840
rect 104894 498108 104900 498160
rect 104952 498148 104958 498160
rect 153194 498148 153200 498160
rect 104952 498120 153200 498148
rect 104952 498108 104958 498120
rect 153194 498108 153200 498120
rect 153252 498108 153258 498160
rect 132494 497632 132500 497684
rect 132552 497672 132558 497684
rect 157426 497672 157432 497684
rect 132552 497644 157432 497672
rect 132552 497632 132558 497644
rect 157426 497632 157432 497644
rect 157484 497632 157490 497684
rect 70578 497564 70584 497616
rect 70636 497604 70642 497616
rect 95234 497604 95240 497616
rect 70636 497576 95240 497604
rect 70636 497564 70642 497576
rect 95234 497564 95240 497576
rect 95292 497564 95298 497616
rect 121454 497564 121460 497616
rect 121512 497604 121518 497616
rect 155586 497604 155592 497616
rect 121512 497576 155592 497604
rect 121512 497564 121518 497576
rect 155586 497564 155592 497576
rect 155644 497564 155650 497616
rect 82814 497496 82820 497548
rect 82872 497536 82878 497548
rect 115934 497536 115940 497548
rect 82872 497508 115940 497536
rect 82872 497496 82878 497508
rect 115934 497496 115940 497508
rect 115992 497496 115998 497548
rect 118694 497496 118700 497548
rect 118752 497536 118758 497548
rect 153470 497536 153476 497548
rect 118752 497508 153476 497536
rect 118752 497496 118758 497508
rect 153470 497496 153476 497508
rect 153528 497496 153534 497548
rect 93854 497428 93860 497480
rect 93912 497468 93918 497480
rect 133874 497468 133880 497480
rect 93912 497440 133880 497468
rect 93912 497428 93918 497440
rect 133874 497428 133880 497440
rect 133932 497428 133938 497480
rect 299382 496068 299388 496120
rect 299440 496108 299446 496120
rect 414014 496108 414020 496120
rect 299440 496080 414020 496108
rect 299440 496068 299446 496080
rect 414014 496068 414020 496080
rect 414072 496068 414078 496120
rect 3510 495456 3516 495508
rect 3568 495496 3574 495508
rect 298094 495496 298100 495508
rect 3568 495468 298100 495496
rect 3568 495456 3574 495468
rect 298094 495456 298100 495468
rect 298152 495496 298158 495508
rect 299382 495496 299388 495508
rect 298152 495468 299388 495496
rect 298152 495456 298158 495468
rect 299382 495456 299388 495468
rect 299440 495456 299446 495508
rect 571334 495456 571340 495508
rect 571392 495496 571398 495508
rect 573450 495496 573456 495508
rect 571392 495468 573456 495496
rect 571392 495456 571398 495468
rect 573450 495456 573456 495468
rect 573508 495456 573514 495508
rect 74534 494844 74540 494896
rect 74592 494884 74598 494896
rect 102134 494884 102140 494896
rect 74592 494856 102140 494884
rect 74592 494844 74598 494856
rect 102134 494844 102140 494856
rect 102192 494844 102198 494896
rect 85666 494776 85672 494828
rect 85724 494816 85730 494828
rect 120074 494816 120080 494828
rect 85724 494788 120080 494816
rect 85724 494776 85730 494788
rect 120074 494776 120080 494788
rect 120132 494776 120138 494828
rect 63494 494708 63500 494760
rect 63552 494748 63558 494760
rect 84194 494748 84200 494760
rect 63552 494720 84200 494748
rect 63552 494708 63558 494720
rect 84194 494708 84200 494720
rect 84252 494708 84258 494760
rect 95418 494708 95424 494760
rect 95476 494748 95482 494760
rect 138658 494748 138664 494760
rect 95476 494720 138664 494748
rect 95476 494708 95482 494720
rect 138658 494708 138664 494720
rect 138716 494708 138722 494760
rect 194502 493960 194508 494012
rect 194560 494000 194566 494012
rect 197170 494000 197176 494012
rect 194560 493972 197176 494000
rect 194560 493960 194566 493972
rect 197170 493960 197176 493972
rect 197228 493960 197234 494012
rect 202874 493960 202880 494012
rect 202932 494000 202938 494012
rect 205634 494000 205640 494012
rect 202932 493972 205640 494000
rect 202932 493960 202938 493972
rect 205634 493960 205640 493972
rect 205692 493960 205698 494012
rect 208854 493960 208860 494012
rect 208912 494000 208918 494012
rect 211154 494000 211160 494012
rect 208912 493972 211160 494000
rect 208912 493960 208918 493972
rect 211154 493960 211160 493972
rect 211212 493960 211218 494012
rect 213638 493960 213644 494012
rect 213696 494000 213702 494012
rect 215386 494000 215392 494012
rect 213696 493972 215392 494000
rect 213696 493960 213702 493972
rect 215386 493960 215392 493972
rect 215444 493960 215450 494012
rect 218422 493960 218428 494012
rect 218480 494000 218486 494012
rect 220814 494000 220820 494012
rect 218480 493972 220820 494000
rect 218480 493960 218486 493972
rect 220814 493960 220820 493972
rect 220872 493960 220878 494012
rect 235166 493960 235172 494012
rect 235224 494000 235230 494012
rect 237558 494000 237564 494012
rect 235224 493972 237564 494000
rect 235224 493960 235230 493972
rect 237558 493960 237564 493972
rect 237616 493960 237622 494012
rect 241146 493960 241152 494012
rect 241204 494000 241210 494012
rect 243078 494000 243084 494012
rect 241204 493972 243084 494000
rect 241204 493960 241210 493972
rect 243078 493960 243084 493972
rect 243136 493960 243142 494012
rect 245930 493960 245936 494012
rect 245988 494000 245994 494012
rect 248414 494000 248420 494012
rect 245988 493972 248420 494000
rect 245988 493960 245994 493972
rect 248414 493960 248420 493972
rect 248472 493960 248478 494012
rect 258258 493960 258264 494012
rect 258316 494000 258322 494012
rect 259086 494000 259092 494012
rect 258316 493972 259092 494000
rect 258316 493960 258322 493972
rect 259086 493960 259092 493972
rect 259144 493960 259150 494012
rect 259454 493960 259460 494012
rect 259512 494000 259518 494012
rect 260282 494000 260288 494012
rect 259512 493972 260288 494000
rect 259512 493960 259518 493972
rect 260282 493960 260288 493972
rect 260340 493960 260346 494012
rect 232774 493892 232780 493944
rect 232832 493932 232838 493944
rect 235902 493932 235908 493944
rect 232832 493904 235908 493932
rect 232832 493892 232838 493904
rect 235902 493892 235908 493904
rect 235960 493892 235966 493944
rect 249794 493932 249800 493944
rect 248432 493904 249800 493932
rect 198090 493824 198096 493876
rect 198148 493864 198154 493876
rect 200114 493864 200120 493876
rect 198148 493836 200120 493864
rect 198148 493824 198154 493836
rect 200114 493824 200120 493836
rect 200172 493824 200178 493876
rect 220814 493824 220820 493876
rect 220872 493864 220878 493876
rect 224862 493864 224868 493876
rect 220872 493836 224868 493864
rect 220872 493824 220878 493836
rect 224862 493824 224868 493836
rect 224920 493824 224926 493876
rect 227990 493824 227996 493876
rect 228048 493864 228054 493876
rect 230474 493864 230480 493876
rect 228048 493836 230480 493864
rect 228048 493824 228054 493836
rect 230474 493824 230480 493836
rect 230532 493824 230538 493876
rect 237558 493824 237564 493876
rect 237616 493864 237622 493876
rect 240134 493864 240140 493876
rect 237616 493836 240140 493864
rect 237616 493824 237622 493836
rect 240134 493824 240140 493836
rect 240192 493824 240198 493876
rect 193306 493756 193312 493808
rect 193364 493796 193370 493808
rect 196434 493796 196440 493808
rect 193364 493768 196440 493796
rect 193364 493756 193370 493768
rect 196434 493756 196440 493768
rect 196492 493756 196498 493808
rect 199286 493756 199292 493808
rect 199344 493796 199350 493808
rect 201586 493796 201592 493808
rect 199344 493768 201592 493796
rect 199344 493756 199350 493768
rect 201586 493756 201592 493768
rect 201644 493756 201650 493808
rect 201678 493756 201684 493808
rect 201736 493796 201742 493808
rect 204898 493796 204904 493808
rect 201736 493768 204904 493796
rect 201736 493756 201742 493768
rect 204898 493756 204904 493768
rect 204956 493756 204962 493808
rect 211246 493756 211252 493808
rect 211304 493796 211310 493808
rect 214650 493796 214656 493808
rect 211304 493768 214656 493796
rect 211304 493756 211310 493768
rect 214650 493756 214656 493768
rect 214708 493756 214714 493808
rect 236362 493756 236368 493808
rect 236420 493796 236426 493808
rect 238754 493796 238760 493808
rect 236420 493768 238760 493796
rect 236420 493756 236426 493768
rect 238754 493756 238760 493768
rect 238812 493756 238818 493808
rect 248322 493756 248328 493808
rect 248380 493796 248386 493808
rect 248432 493796 248460 493904
rect 249794 493892 249800 493904
rect 249852 493892 249858 493944
rect 248380 493768 248460 493796
rect 248380 493756 248386 493768
rect 249518 493756 249524 493808
rect 249576 493796 249582 493808
rect 251266 493796 251272 493808
rect 249576 493768 251272 493796
rect 249576 493756 249582 493768
rect 251266 493756 251272 493768
rect 251324 493756 251330 493808
rect 188614 493688 188620 493740
rect 188672 493728 188678 493740
rect 191926 493728 191932 493740
rect 188672 493700 191932 493728
rect 188672 493688 188678 493700
rect 191926 493688 191932 493700
rect 191984 493688 191990 493740
rect 200482 493688 200488 493740
rect 200540 493728 200546 493740
rect 203886 493728 203892 493740
rect 200540 493700 203892 493728
rect 200540 493688 200546 493700
rect 203886 493688 203892 493700
rect 203944 493688 203950 493740
rect 210050 493688 210056 493740
rect 210108 493728 210114 493740
rect 213822 493728 213828 493740
rect 210108 493700 213828 493728
rect 210108 493688 210114 493700
rect 213822 493688 213828 493700
rect 213880 493688 213886 493740
rect 195698 493620 195704 493672
rect 195756 493660 195762 493672
rect 201494 493660 201500 493672
rect 195756 493632 201500 493660
rect 195756 493620 195762 493632
rect 201494 493620 201500 493632
rect 201552 493620 201558 493672
rect 204070 493620 204076 493672
rect 204128 493660 204134 493672
rect 206370 493660 206376 493672
rect 204128 493632 206376 493660
rect 204128 493620 204134 493632
rect 206370 493620 206376 493632
rect 206428 493620 206434 493672
rect 206462 493620 206468 493672
rect 206520 493660 206526 493672
rect 209130 493660 209136 493672
rect 206520 493632 209136 493660
rect 206520 493620 206526 493632
rect 209130 493620 209136 493632
rect 209188 493620 209194 493672
rect 222010 493620 222016 493672
rect 222068 493660 222074 493672
rect 224218 493660 224224 493672
rect 222068 493632 224224 493660
rect 222068 493620 222074 493632
rect 224218 493620 224224 493632
rect 224276 493620 224282 493672
rect 231578 493620 231584 493672
rect 231636 493660 231642 493672
rect 234522 493660 234528 493672
rect 231636 493632 234528 493660
rect 231636 493620 231642 493632
rect 234522 493620 234528 493632
rect 234580 493620 234586 493672
rect 196894 493552 196900 493604
rect 196952 493592 196958 493604
rect 199470 493592 199476 493604
rect 196952 493564 199476 493592
rect 196952 493552 196958 493564
rect 199470 493552 199476 493564
rect 199528 493552 199534 493604
rect 217226 493552 217232 493604
rect 217284 493592 217290 493604
rect 219526 493592 219532 493604
rect 217284 493564 219532 493592
rect 217284 493552 217290 493564
rect 219526 493552 219532 493564
rect 219584 493552 219590 493604
rect 219618 493552 219624 493604
rect 219676 493592 219682 493604
rect 223482 493592 223488 493604
rect 219676 493564 223488 493592
rect 219676 493552 219682 493564
rect 223482 493552 223488 493564
rect 223540 493552 223546 493604
rect 225598 493552 225604 493604
rect 225656 493592 225662 493604
rect 229002 493592 229008 493604
rect 225656 493564 229008 493592
rect 225656 493552 225662 493564
rect 229002 493552 229008 493564
rect 229060 493552 229066 493604
rect 233970 493552 233976 493604
rect 234028 493592 234034 493604
rect 237282 493592 237288 493604
rect 234028 493564 237288 493592
rect 234028 493552 234034 493564
rect 237282 493552 237288 493564
rect 237340 493552 237346 493604
rect 205266 493484 205272 493536
rect 205324 493524 205330 493536
rect 207106 493524 207112 493536
rect 205324 493496 207112 493524
rect 205324 493484 205330 493496
rect 207106 493484 207112 493496
rect 207164 493484 207170 493536
rect 212442 493484 212448 493536
rect 212500 493524 212506 493536
rect 215202 493524 215208 493536
rect 212500 493496 215208 493524
rect 212500 493484 212506 493496
rect 215202 493484 215208 493496
rect 215260 493484 215266 493536
rect 216030 493484 216036 493536
rect 216088 493524 216094 493536
rect 218146 493524 218152 493536
rect 216088 493496 218152 493524
rect 216088 493484 216094 493496
rect 218146 493484 218152 493496
rect 218204 493484 218210 493536
rect 239950 493484 239956 493536
rect 240008 493524 240014 493536
rect 242802 493524 242808 493536
rect 240008 493496 242808 493524
rect 240008 493484 240014 493496
rect 242802 493484 242808 493496
rect 242860 493484 242866 493536
rect 71774 493416 71780 493468
rect 71832 493456 71838 493468
rect 97994 493456 98000 493468
rect 71832 493428 98000 493456
rect 71832 493416 71838 493428
rect 97994 493416 98000 493428
rect 98052 493416 98058 493468
rect 229186 493416 229192 493468
rect 229244 493456 229250 493468
rect 233142 493456 233148 493468
rect 229244 493428 233148 493456
rect 229244 493416 229250 493428
rect 233142 493416 233148 493428
rect 233200 493416 233206 493468
rect 238754 493416 238760 493468
rect 238812 493456 238818 493468
rect 241514 493456 241520 493468
rect 238812 493428 241520 493456
rect 238812 493416 238818 493428
rect 241514 493416 241520 493428
rect 241572 493416 241578 493468
rect 243538 493416 243544 493468
rect 243596 493456 243602 493468
rect 245654 493456 245660 493468
rect 243596 493428 245660 493456
rect 243596 493416 243602 493428
rect 245654 493416 245660 493428
rect 245712 493416 245718 493468
rect 78674 493348 78680 493400
rect 78732 493388 78738 493400
rect 109034 493388 109040 493400
rect 78732 493360 109040 493388
rect 78732 493348 78738 493360
rect 109034 493348 109040 493360
rect 109092 493348 109098 493400
rect 189718 493348 189724 493400
rect 189776 493388 189782 493400
rect 195054 493388 195060 493400
rect 189776 493360 195060 493388
rect 189776 493348 189782 493360
rect 195054 493348 195060 493360
rect 195112 493348 195118 493400
rect 59354 493280 59360 493332
rect 59412 493320 59418 493332
rect 77294 493320 77300 493332
rect 59412 493292 77300 493320
rect 59412 493280 59418 493292
rect 77294 493280 77300 493292
rect 77352 493280 77358 493332
rect 93762 493280 93768 493332
rect 93820 493320 93826 493332
rect 131114 493320 131120 493332
rect 93820 493292 131120 493320
rect 93820 493280 93826 493292
rect 131114 493280 131120 493292
rect 131172 493280 131178 493332
rect 207658 493280 207664 493332
rect 207716 493320 207722 493332
rect 209866 493320 209872 493332
rect 207716 493292 209872 493320
rect 207716 493280 207722 493292
rect 209866 493280 209872 493292
rect 209924 493280 209930 493332
rect 244734 493280 244740 493332
rect 244792 493320 244798 493332
rect 247218 493320 247224 493332
rect 244792 493292 247224 493320
rect 244792 493280 244798 493292
rect 247218 493280 247224 493292
rect 247276 493280 247282 493332
rect 563698 493280 563704 493332
rect 563756 493320 563762 493332
rect 571334 493320 571340 493332
rect 563756 493292 571340 493320
rect 563756 493280 563762 493292
rect 571334 493280 571340 493292
rect 571392 493280 571398 493332
rect 214834 493212 214840 493264
rect 214892 493252 214898 493264
rect 216674 493252 216680 493264
rect 214892 493224 216680 493252
rect 214892 493212 214898 493224
rect 216674 493212 216680 493224
rect 216732 493212 216738 493264
rect 226794 493212 226800 493264
rect 226852 493252 226858 493264
rect 230382 493252 230388 493264
rect 226852 493224 230388 493252
rect 226852 493212 226858 493224
rect 230382 493212 230388 493224
rect 230440 493212 230446 493264
rect 242342 493212 242348 493264
rect 242400 493252 242406 493264
rect 244274 493252 244280 493264
rect 242400 493224 244280 493252
rect 242400 493212 242406 493224
rect 244274 493212 244280 493224
rect 244332 493212 244338 493264
rect 277578 493144 277584 493196
rect 277636 493184 277642 493196
rect 279418 493184 279424 493196
rect 277636 493156 279424 493184
rect 277636 493144 277642 493156
rect 279418 493144 279424 493156
rect 279476 493144 279482 493196
rect 230382 493076 230388 493128
rect 230440 493116 230446 493128
rect 233050 493116 233056 493128
rect 230440 493088 233056 493116
rect 230440 493076 230446 493088
rect 233050 493076 233056 493088
rect 233108 493076 233114 493128
rect 266446 493076 266452 493128
rect 266504 493116 266510 493128
rect 267458 493116 267464 493128
rect 266504 493088 267464 493116
rect 266504 493076 266510 493088
rect 267458 493076 267464 493088
rect 267516 493076 267522 493128
rect 250714 492940 250720 492992
rect 250772 492980 250778 492992
rect 252738 492980 252744 492992
rect 250772 492952 252744 492980
rect 250772 492940 250778 492952
rect 252738 492940 252744 492952
rect 252796 492940 252802 492992
rect 223206 492872 223212 492924
rect 223264 492912 223270 492924
rect 227898 492912 227904 492924
rect 223264 492884 227904 492912
rect 223264 492872 223270 492884
rect 227898 492872 227904 492884
rect 227956 492872 227962 492924
rect 190914 492804 190920 492856
rect 190972 492844 190978 492856
rect 195882 492844 195888 492856
rect 190972 492816 195888 492844
rect 190972 492804 190978 492816
rect 195882 492804 195888 492816
rect 195940 492804 195946 492856
rect 271966 492804 271972 492856
rect 272024 492844 272030 492856
rect 273438 492844 273444 492856
rect 272024 492816 273444 492844
rect 272024 492804 272030 492816
rect 273438 492804 273444 492816
rect 273496 492804 273502 492856
rect 223574 492736 223580 492788
rect 223632 492776 223638 492788
rect 224402 492776 224408 492788
rect 223632 492748 224408 492776
rect 223632 492736 223638 492748
rect 224402 492736 224408 492748
rect 224460 492736 224466 492788
rect 146018 492668 146024 492720
rect 146076 492708 146082 492720
rect 154114 492708 154120 492720
rect 146076 492680 154120 492708
rect 146076 492668 146082 492680
rect 154114 492668 154120 492680
rect 154172 492668 154178 492720
rect 154298 492668 154304 492720
rect 154356 492708 154362 492720
rect 154390 492708 154396 492720
rect 154356 492680 154396 492708
rect 154356 492668 154362 492680
rect 154390 492668 154396 492680
rect 154448 492668 154454 492720
rect 155678 492600 155684 492652
rect 155736 492640 155742 492652
rect 156138 492640 156144 492652
rect 155736 492612 156144 492640
rect 155736 492600 155742 492612
rect 156138 492600 156144 492612
rect 156196 492600 156202 492652
rect 158898 492600 158904 492652
rect 158956 492640 158962 492652
rect 158990 492640 158996 492652
rect 158956 492612 158996 492640
rect 158956 492600 158962 492612
rect 158990 492600 158996 492612
rect 159048 492600 159054 492652
rect 68922 492056 68928 492108
rect 68980 492096 68986 492108
rect 92106 492096 92112 492108
rect 68980 492068 92112 492096
rect 68980 492056 68986 492068
rect 92106 492056 92112 492068
rect 92164 492056 92170 492108
rect 77110 491988 77116 492040
rect 77168 492028 77174 492040
rect 106458 492028 106464 492040
rect 77168 492000 106464 492028
rect 77168 491988 77174 492000
rect 106458 491988 106464 492000
rect 106516 491988 106522 492040
rect 57882 491920 57888 491972
rect 57940 491960 57946 491972
rect 74166 491960 74172 491972
rect 57940 491932 74172 491960
rect 57940 491920 57946 491932
rect 74166 491920 74172 491932
rect 74224 491920 74230 491972
rect 88242 491920 88248 491972
rect 88300 491960 88306 491972
rect 124306 491960 124312 491972
rect 88300 491932 124312 491960
rect 88300 491920 88306 491932
rect 124306 491920 124312 491932
rect 124364 491920 124370 491972
rect 154298 491240 154304 491292
rect 154356 491280 154362 491292
rect 154482 491280 154488 491292
rect 154356 491252 154488 491280
rect 154356 491240 154362 491252
rect 154482 491240 154488 491252
rect 154540 491240 154546 491292
rect 11698 490560 11704 490612
rect 11756 490600 11762 490612
rect 443638 490600 443644 490612
rect 11756 490572 443644 490600
rect 11756 490560 11762 490572
rect 443638 490560 443644 490572
rect 443696 490560 443702 490612
rect 35802 489812 35808 489864
rect 35860 489852 35866 489864
rect 36538 489852 36544 489864
rect 35860 489824 36544 489852
rect 35860 489812 35866 489824
rect 36538 489812 36544 489824
rect 36596 489812 36602 489864
rect 82722 489812 82728 489864
rect 82780 489852 82786 489864
rect 115014 489852 115020 489864
rect 82780 489824 115020 489852
rect 82780 489812 82786 489824
rect 115014 489812 115020 489824
rect 115072 489812 115078 489864
rect 115198 489812 115204 489864
rect 115256 489852 115262 489864
rect 140498 489852 140504 489864
rect 115256 489824 140504 489852
rect 115256 489812 115262 489824
rect 140498 489812 140504 489824
rect 140556 489812 140562 489864
rect 52362 489744 52368 489796
rect 52420 489784 52426 489796
rect 63126 489784 63132 489796
rect 52420 489756 63132 489784
rect 52420 489744 52426 489756
rect 63126 489744 63132 489756
rect 63184 489744 63190 489796
rect 86862 489744 86868 489796
rect 86920 489784 86926 489796
rect 122558 489784 122564 489796
rect 86920 489756 122564 489784
rect 86920 489744 86926 489756
rect 122558 489744 122564 489756
rect 122616 489744 122622 489796
rect 55122 489676 55128 489728
rect 55180 489716 55186 489728
rect 68738 489716 68744 489728
rect 55180 489688 68744 489716
rect 55180 489676 55186 489688
rect 68738 489676 68744 489688
rect 68796 489676 68802 489728
rect 90910 489676 90916 489728
rect 90968 489716 90974 489728
rect 129734 489716 129740 489728
rect 90968 489688 129740 489716
rect 90968 489676 90974 489688
rect 129734 489676 129740 489688
rect 129792 489676 129798 489728
rect 62022 489608 62028 489660
rect 62080 489648 62086 489660
rect 79502 489648 79508 489660
rect 62080 489620 79508 489648
rect 62080 489608 62086 489620
rect 79502 489608 79508 489620
rect 79560 489608 79566 489660
rect 96522 489608 96528 489660
rect 96580 489648 96586 489660
rect 136910 489648 136916 489660
rect 96580 489620 136916 489648
rect 96580 489608 96586 489620
rect 136910 489608 136916 489620
rect 136968 489608 136974 489660
rect 49602 489540 49608 489592
rect 49660 489580 49666 489592
rect 59814 489580 59820 489592
rect 49660 489552 59820 489580
rect 49660 489540 49666 489552
rect 59814 489540 59820 489552
rect 59872 489540 59878 489592
rect 63402 489540 63408 489592
rect 63460 489580 63466 489592
rect 83090 489580 83096 489592
rect 63460 489552 83096 489580
rect 63460 489540 63466 489552
rect 83090 489540 83096 489552
rect 83148 489540 83154 489592
rect 100662 489540 100668 489592
rect 100720 489580 100726 489592
rect 144086 489580 144092 489592
rect 100720 489552 144092 489580
rect 100720 489540 100726 489552
rect 144086 489540 144092 489552
rect 144144 489540 144150 489592
rect 22186 489472 22192 489524
rect 22244 489512 22250 489524
rect 26326 489512 26332 489524
rect 22244 489484 26332 489512
rect 22244 489472 22250 489484
rect 26326 489472 26332 489484
rect 26384 489472 26390 489524
rect 50982 489472 50988 489524
rect 51040 489512 51046 489524
rect 61654 489512 61660 489524
rect 51040 489484 61660 489512
rect 51040 489472 51046 489484
rect 61654 489472 61660 489484
rect 61712 489472 61718 489524
rect 66162 489472 66168 489524
rect 66220 489512 66226 489524
rect 86678 489512 86684 489524
rect 66220 489484 86684 489512
rect 66220 489472 66226 489484
rect 86678 489472 86684 489484
rect 86736 489472 86742 489524
rect 99282 489472 99288 489524
rect 99340 489512 99346 489524
rect 142246 489512 142252 489524
rect 99340 489484 142252 489512
rect 99340 489472 99346 489484
rect 142246 489472 142252 489484
rect 142304 489472 142310 489524
rect 53742 489404 53748 489456
rect 53800 489444 53806 489456
rect 66990 489444 66996 489456
rect 53800 489416 66996 489444
rect 53800 489404 53806 489416
rect 66990 489404 66996 489416
rect 67048 489404 67054 489456
rect 67450 489404 67456 489456
rect 67508 489444 67514 489456
rect 90266 489444 90272 489456
rect 67508 489416 90272 489444
rect 67508 489404 67514 489416
rect 90266 489404 90272 489416
rect 90324 489404 90330 489456
rect 102042 489404 102048 489456
rect 102100 489444 102106 489456
rect 145834 489444 145840 489456
rect 102100 489416 145840 489444
rect 102100 489404 102106 489416
rect 145834 489404 145840 489416
rect 145892 489404 145898 489456
rect 25774 489336 25780 489388
rect 25832 489376 25838 489388
rect 27614 489376 27620 489388
rect 25832 489348 27620 489376
rect 25832 489336 25838 489348
rect 27614 489336 27620 489348
rect 27672 489336 27678 489388
rect 52270 489336 52276 489388
rect 52328 489376 52334 489388
rect 65150 489376 65156 489388
rect 52328 489348 65156 489376
rect 52328 489336 52334 489348
rect 65150 489336 65156 489348
rect 65208 489336 65214 489388
rect 70302 489336 70308 489388
rect 70360 489376 70366 489388
rect 93854 489376 93860 489388
rect 70360 489348 93860 489376
rect 70360 489336 70366 489348
rect 93854 489336 93860 489348
rect 93912 489336 93918 489388
rect 106918 489336 106924 489388
rect 106976 489376 106982 489388
rect 153010 489376 153016 489388
rect 106976 489348 153016 489376
rect 106976 489336 106982 489348
rect 153010 489336 153016 489348
rect 153068 489336 153074 489388
rect 48222 489268 48228 489320
rect 48280 489308 48286 489320
rect 58066 489308 58072 489320
rect 48280 489280 58072 489308
rect 48280 489268 48286 489280
rect 58066 489268 58072 489280
rect 58124 489268 58130 489320
rect 59262 489268 59268 489320
rect 59320 489308 59326 489320
rect 75914 489308 75920 489320
rect 59320 489280 75920 489308
rect 59320 489268 59326 489280
rect 75914 489268 75920 489280
rect 75972 489268 75978 489320
rect 77202 489268 77208 489320
rect 77260 489308 77266 489320
rect 104618 489308 104624 489320
rect 77260 489280 104624 489308
rect 77260 489268 77266 489280
rect 104618 489268 104624 489280
rect 104676 489268 104682 489320
rect 104802 489268 104808 489320
rect 104860 489308 104866 489320
rect 151262 489308 151268 489320
rect 104860 489280 151268 489308
rect 104860 489268 104866 489280
rect 151262 489268 151268 489280
rect 151320 489268 151326 489320
rect 37090 489200 37096 489252
rect 37148 489240 37154 489252
rect 40126 489240 40132 489252
rect 37148 489212 40132 489240
rect 37148 489200 37154 489212
rect 40126 489200 40132 489212
rect 40184 489200 40190 489252
rect 56502 489200 56508 489252
rect 56560 489240 56566 489252
rect 70578 489240 70584 489252
rect 56560 489212 70584 489240
rect 56560 489200 56566 489212
rect 70578 489200 70584 489212
rect 70636 489200 70642 489252
rect 71682 489200 71688 489252
rect 71740 489240 71746 489252
rect 97442 489240 97448 489252
rect 71740 489212 97448 489240
rect 71740 489200 71746 489212
rect 97442 489200 97448 489212
rect 97500 489200 97506 489252
rect 103422 489200 103428 489252
rect 103480 489240 103486 489252
rect 149422 489240 149428 489252
rect 103480 489212 149428 489240
rect 103480 489200 103486 489212
rect 149422 489200 149428 489212
rect 149480 489200 149486 489252
rect 37182 489132 37188 489184
rect 37240 489172 37246 489184
rect 38286 489172 38292 489184
rect 37240 489144 38292 489172
rect 37240 489132 37246 489144
rect 38286 489132 38292 489144
rect 38344 489132 38350 489184
rect 46842 489132 46848 489184
rect 46900 489172 46906 489184
rect 56226 489172 56232 489184
rect 46900 489144 56232 489172
rect 46900 489132 46906 489144
rect 56226 489132 56232 489144
rect 56284 489132 56290 489184
rect 56410 489132 56416 489184
rect 56468 489172 56474 489184
rect 72326 489172 72332 489184
rect 56468 489144 72332 489172
rect 56468 489132 56474 489144
rect 72326 489132 72332 489144
rect 72384 489132 72390 489184
rect 74442 489132 74448 489184
rect 74500 489172 74506 489184
rect 101030 489172 101036 489184
rect 74500 489144 101036 489172
rect 74500 489132 74506 489144
rect 101030 489132 101036 489144
rect 101088 489132 101094 489184
rect 101950 489132 101956 489184
rect 102008 489172 102014 489184
rect 147674 489172 147680 489184
rect 102008 489144 147680 489172
rect 102008 489132 102014 489144
rect 147674 489132 147680 489144
rect 147732 489132 147738 489184
rect 78582 489064 78588 489116
rect 78640 489104 78646 489116
rect 108206 489104 108212 489116
rect 78640 489076 108212 489104
rect 78640 489064 78646 489076
rect 108206 489064 108212 489076
rect 108264 489064 108270 489116
rect 113818 489064 113824 489116
rect 113876 489104 113882 489116
rect 133322 489104 133328 489116
rect 113876 489076 133328 489104
rect 113876 489064 113882 489076
rect 133322 489064 133328 489076
rect 133380 489064 133386 489116
rect 112438 488996 112444 489048
rect 112496 489036 112502 489048
rect 126146 489036 126152 489048
rect 112496 489008 126152 489036
rect 112496 488996 112502 489008
rect 126146 488996 126152 489008
rect 126204 488996 126210 489048
rect 109678 488928 109684 488980
rect 109736 488968 109742 488980
rect 118970 488968 118976 488980
rect 109736 488940 118976 488968
rect 109736 488928 109742 488940
rect 118970 488928 118976 488940
rect 119028 488928 119034 488980
rect 39942 488656 39948 488708
rect 40000 488696 40006 488708
rect 43714 488696 43720 488708
rect 40000 488668 43720 488696
rect 40000 488656 40006 488668
rect 43714 488656 43720 488668
rect 43772 488656 43778 488708
rect 18598 488588 18604 488640
rect 18656 488628 18662 488640
rect 23566 488628 23572 488640
rect 18656 488600 23572 488628
rect 18656 488588 18662 488600
rect 23566 488588 23572 488600
rect 23624 488588 23630 488640
rect 38562 488588 38568 488640
rect 38620 488628 38626 488640
rect 41874 488628 41880 488640
rect 38620 488600 41880 488628
rect 38620 488588 38626 488600
rect 41874 488588 41880 488600
rect 41932 488588 41938 488640
rect 48958 488588 48964 488640
rect 49016 488628 49022 488640
rect 50890 488628 50896 488640
rect 49016 488600 50896 488628
rect 49016 488588 49022 488600
rect 50890 488588 50896 488600
rect 50948 488588 50954 488640
rect 16850 488520 16856 488572
rect 16908 488560 16914 488572
rect 22278 488560 22284 488572
rect 16908 488532 22284 488560
rect 16908 488520 16914 488532
rect 22278 488520 22284 488532
rect 22336 488520 22342 488572
rect 23934 488520 23940 488572
rect 23992 488560 23998 488572
rect 24762 488560 24768 488572
rect 23992 488532 24768 488560
rect 23992 488520 23998 488532
rect 24762 488520 24768 488532
rect 24820 488520 24826 488572
rect 29362 488520 29368 488572
rect 29420 488560 29426 488572
rect 30282 488560 30288 488572
rect 29420 488532 30288 488560
rect 29420 488520 29426 488532
rect 30282 488520 30288 488532
rect 30340 488520 30346 488572
rect 41322 488520 41328 488572
rect 41380 488560 41386 488572
rect 45462 488560 45468 488572
rect 41380 488532 45468 488560
rect 41380 488520 41386 488532
rect 45462 488520 45468 488532
rect 45520 488520 45526 488572
rect 47578 488520 47584 488572
rect 47636 488560 47642 488572
rect 49050 488560 49056 488572
rect 47636 488532 49056 488560
rect 47636 488520 47642 488532
rect 49050 488520 49056 488532
rect 49108 488520 49114 488572
rect 108298 488520 108304 488572
rect 108356 488560 108362 488572
rect 111794 488560 111800 488572
rect 108356 488532 111800 488560
rect 108356 488520 108362 488532
rect 111794 488520 111800 488532
rect 111852 488520 111858 488572
rect 23382 486412 23388 486464
rect 23440 486452 23446 486464
rect 156046 486452 156052 486464
rect 23440 486424 156052 486452
rect 23440 486412 23446 486424
rect 156046 486412 156052 486424
rect 156104 486412 156110 486464
rect 283006 485800 283012 485852
rect 283064 485800 283070 485852
rect 158898 485732 158904 485784
rect 158956 485772 158962 485784
rect 158990 485772 158996 485784
rect 158956 485744 158996 485772
rect 158956 485732 158962 485744
rect 158990 485732 158996 485744
rect 159048 485732 159054 485784
rect 283024 485772 283052 485800
rect 283098 485772 283104 485784
rect 283024 485744 283104 485772
rect 283098 485732 283104 485744
rect 283156 485732 283162 485784
rect 3418 485052 3424 485104
rect 3476 485092 3482 485104
rect 185578 485092 185584 485104
rect 3476 485064 185584 485092
rect 3476 485052 3482 485064
rect 185578 485052 185584 485064
rect 185636 485052 185642 485104
rect 283098 482944 283104 482996
rect 283156 482984 283162 482996
rect 283282 482984 283288 482996
rect 283156 482956 283288 482984
rect 283156 482944 283162 482956
rect 283282 482944 283288 482956
rect 283340 482944 283346 482996
rect 560386 482808 560392 482860
rect 560444 482848 560450 482860
rect 563698 482848 563704 482860
rect 560444 482820 563704 482848
rect 560444 482808 560450 482820
rect 563698 482808 563704 482820
rect 563756 482808 563762 482860
rect 154298 481652 154304 481704
rect 154356 481692 154362 481704
rect 154482 481692 154488 481704
rect 154356 481664 154488 481692
rect 154356 481652 154362 481664
rect 154482 481652 154488 481664
rect 154540 481652 154546 481704
rect 3142 480224 3148 480276
rect 3200 480264 3206 480276
rect 11698 480264 11704 480276
rect 3200 480236 11704 480264
rect 3200 480224 3206 480236
rect 11698 480224 11704 480236
rect 11756 480224 11762 480276
rect 183646 480224 183652 480276
rect 183704 480264 183710 480276
rect 183830 480264 183836 480276
rect 183704 480236 183836 480264
rect 183704 480224 183710 480236
rect 183830 480224 183836 480236
rect 183888 480224 183894 480276
rect 559558 479476 559564 479528
rect 559616 479516 559622 479528
rect 560386 479516 560392 479528
rect 559616 479488 560392 479516
rect 559616 479476 559622 479488
rect 560386 479476 560392 479488
rect 560444 479476 560450 479528
rect 344922 477436 344928 477488
rect 344980 477476 344986 477488
rect 346026 477476 346032 477488
rect 344980 477448 346032 477476
rect 344980 477436 344986 477448
rect 346026 477436 346032 477448
rect 346084 477436 346090 477488
rect 353202 477436 353208 477488
rect 353260 477476 353266 477488
rect 355778 477476 355784 477488
rect 353260 477448 355784 477476
rect 353260 477436 353266 477448
rect 355778 477436 355784 477448
rect 355836 477436 355842 477488
rect 362862 477436 362868 477488
rect 362920 477476 362926 477488
rect 366726 477476 366732 477488
rect 362920 477448 366732 477476
rect 362920 477436 362926 477448
rect 366726 477436 366732 477448
rect 366784 477436 366790 477488
rect 369762 477436 369768 477488
rect 369820 477476 369826 477488
rect 374086 477476 374092 477488
rect 369820 477448 374092 477476
rect 369820 477436 369826 477448
rect 374086 477436 374092 477448
rect 374144 477436 374150 477488
rect 354582 477368 354588 477420
rect 354640 477408 354646 477420
rect 356974 477408 356980 477420
rect 354640 477380 356980 477408
rect 354640 477368 354646 477380
rect 356974 477368 356980 477380
rect 357032 477368 357038 477420
rect 390462 477300 390468 477352
rect 390520 477340 390526 477352
rect 397270 477340 397276 477352
rect 390520 477312 397276 477340
rect 390520 477300 390526 477312
rect 397270 477300 397276 477312
rect 397328 477300 397334 477352
rect 382182 477164 382188 477216
rect 382240 477204 382246 477216
rect 388714 477204 388720 477216
rect 382240 477176 388720 477204
rect 382240 477164 382246 477176
rect 388714 477164 388720 477176
rect 388772 477164 388778 477216
rect 391842 477164 391848 477216
rect 391900 477204 391906 477216
rect 399754 477204 399760 477216
rect 391900 477176 399760 477204
rect 391900 477164 391906 477176
rect 399754 477164 399760 477176
rect 399812 477164 399818 477216
rect 400122 477164 400128 477216
rect 400180 477204 400186 477216
rect 408310 477204 408316 477216
rect 400180 477176 408316 477204
rect 400180 477164 400186 477176
rect 408310 477164 408316 477176
rect 408368 477164 408374 477216
rect 393222 477096 393228 477148
rect 393280 477136 393286 477148
rect 400950 477136 400956 477148
rect 393280 477108 400956 477136
rect 393280 477096 393286 477108
rect 400950 477096 400956 477108
rect 401008 477096 401014 477148
rect 401502 477096 401508 477148
rect 401560 477136 401566 477148
rect 409506 477136 409512 477148
rect 401560 477108 409512 477136
rect 401560 477096 401566 477108
rect 409506 477096 409512 477108
rect 409564 477096 409570 477148
rect 531222 477096 531228 477148
rect 531280 477136 531286 477148
rect 552750 477136 552756 477148
rect 531280 477108 552756 477136
rect 531280 477096 531286 477108
rect 552750 477096 552756 477108
rect 552808 477096 552814 477148
rect 364242 477028 364248 477080
rect 364300 477068 364306 477080
rect 368014 477068 368020 477080
rect 364300 477040 368020 477068
rect 364300 477028 364306 477040
rect 368014 477028 368020 477040
rect 368072 477028 368078 477080
rect 375282 477028 375288 477080
rect 375340 477068 375346 477080
rect 380158 477068 380164 477080
rect 375340 477040 380164 477068
rect 375340 477028 375346 477040
rect 380158 477028 380164 477040
rect 380216 477028 380222 477080
rect 386230 477028 386236 477080
rect 386288 477068 386294 477080
rect 392486 477068 392492 477080
rect 386288 477040 392492 477068
rect 386288 477028 386294 477040
rect 392486 477028 392492 477040
rect 392544 477028 392550 477080
rect 395890 477028 395896 477080
rect 395948 477068 395954 477080
rect 403434 477068 403440 477080
rect 395948 477040 403440 477068
rect 395948 477028 395954 477040
rect 403434 477028 403440 477040
rect 403492 477028 403498 477080
rect 521562 477028 521568 477080
rect 521620 477068 521626 477080
rect 553210 477068 553216 477080
rect 521620 477040 553216 477068
rect 521620 477028 521626 477040
rect 553210 477028 553216 477040
rect 553268 477028 553274 477080
rect 361482 476960 361488 477012
rect 361540 477000 361546 477012
rect 365530 477000 365536 477012
rect 361540 476972 365536 477000
rect 361540 476960 361546 476972
rect 365530 476960 365536 476972
rect 365588 476960 365594 477012
rect 372522 476960 372528 477012
rect 372580 477000 372586 477012
rect 377766 477000 377772 477012
rect 372580 476972 377772 477000
rect 372580 476960 372586 476972
rect 377766 476960 377772 476972
rect 377824 476960 377830 477012
rect 395982 476960 395988 477012
rect 396040 477000 396046 477012
rect 404630 477000 404636 477012
rect 396040 476972 404636 477000
rect 396040 476960 396046 476972
rect 404630 476960 404636 476972
rect 404688 476960 404694 477012
rect 518802 476960 518808 477012
rect 518860 477000 518866 477012
rect 518860 476972 549668 477000
rect 518860 476960 518866 476972
rect 351822 476892 351828 476944
rect 351880 476932 351886 476944
rect 353294 476932 353300 476944
rect 351880 476904 353300 476932
rect 351880 476892 351886 476904
rect 353294 476892 353300 476904
rect 353352 476892 353358 476944
rect 355870 476892 355876 476944
rect 355928 476932 355934 476944
rect 359458 476932 359464 476944
rect 355928 476904 359464 476932
rect 355928 476892 355934 476904
rect 359458 476892 359464 476904
rect 359516 476892 359522 476944
rect 368382 476892 368388 476944
rect 368440 476932 368446 476944
rect 372890 476932 372896 476944
rect 368440 476904 372896 476932
rect 368440 476892 368446 476904
rect 372890 476892 372896 476904
rect 372948 476892 372954 476944
rect 373902 476892 373908 476944
rect 373960 476932 373966 476944
rect 378962 476932 378968 476944
rect 373960 476904 378968 476932
rect 373960 476892 373966 476904
rect 378962 476892 378968 476904
rect 379020 476892 379026 476944
rect 380802 476892 380808 476944
rect 380860 476932 380866 476944
rect 387518 476932 387524 476944
rect 380860 476904 387524 476932
rect 380860 476892 380866 476904
rect 387518 476892 387524 476904
rect 387576 476892 387582 476944
rect 389082 476892 389088 476944
rect 389140 476932 389146 476944
rect 396074 476932 396080 476944
rect 389140 476904 396080 476932
rect 389140 476892 389146 476904
rect 396074 476892 396080 476904
rect 396132 476892 396138 476944
rect 397362 476892 397368 476944
rect 397420 476932 397426 476944
rect 405826 476932 405832 476944
rect 397420 476904 405832 476932
rect 397420 476892 397426 476904
rect 405826 476892 405832 476904
rect 405884 476892 405890 476944
rect 517422 476892 517428 476944
rect 517480 476932 517486 476944
rect 547322 476932 547328 476944
rect 517480 476904 547328 476932
rect 517480 476892 517486 476904
rect 547322 476892 547328 476904
rect 547380 476892 547386 476944
rect 549640 476932 549668 476972
rect 551922 476960 551928 477012
rect 551980 477000 551986 477012
rect 554130 477000 554136 477012
rect 551980 476972 554136 477000
rect 551980 476960 551986 476972
rect 554130 476960 554136 476972
rect 554188 476960 554194 477012
rect 552106 476932 552112 476944
rect 549640 476904 552112 476932
rect 552106 476892 552112 476904
rect 552164 476892 552170 476944
rect 316678 476824 316684 476876
rect 316736 476864 316742 476876
rect 317322 476864 317328 476876
rect 316736 476836 317328 476864
rect 316736 476824 316742 476836
rect 317322 476824 317328 476836
rect 317380 476824 317386 476876
rect 317874 476824 317880 476876
rect 317932 476864 317938 476876
rect 318702 476864 318708 476876
rect 317932 476836 318708 476864
rect 317932 476824 317938 476836
rect 318702 476824 318708 476836
rect 318760 476824 318766 476876
rect 319070 476824 319076 476876
rect 319128 476864 319134 476876
rect 320082 476864 320088 476876
rect 319128 476836 320088 476864
rect 319128 476824 319134 476836
rect 320082 476824 320088 476836
rect 320140 476824 320146 476876
rect 332594 476824 332600 476876
rect 332652 476864 332658 476876
rect 333790 476864 333796 476876
rect 332652 476836 333796 476864
rect 332652 476824 332658 476836
rect 333790 476824 333796 476836
rect 333848 476824 333854 476876
rect 335354 476824 335360 476876
rect 335412 476864 335418 476876
rect 336182 476864 336188 476876
rect 335412 476836 336188 476864
rect 335412 476824 335418 476836
rect 336182 476824 336188 476836
rect 336240 476824 336246 476876
rect 336642 476824 336648 476876
rect 336700 476864 336706 476876
rect 337470 476864 337476 476876
rect 336700 476836 337476 476864
rect 336700 476824 336706 476836
rect 337470 476824 337476 476836
rect 337528 476824 337534 476876
rect 342162 476824 342168 476876
rect 342220 476864 342226 476876
rect 343542 476864 343548 476876
rect 342220 476836 343548 476864
rect 342220 476824 342226 476836
rect 343542 476824 343548 476836
rect 343600 476824 343606 476876
rect 346210 476824 346216 476876
rect 346268 476864 346274 476876
rect 347222 476864 347228 476876
rect 346268 476836 347228 476864
rect 346268 476824 346274 476836
rect 347222 476824 347228 476836
rect 347280 476824 347286 476876
rect 350442 476824 350448 476876
rect 350500 476864 350506 476876
rect 352098 476864 352104 476876
rect 350500 476836 352104 476864
rect 350500 476824 350506 476836
rect 352098 476824 352104 476836
rect 352156 476824 352162 476876
rect 355962 476824 355968 476876
rect 356020 476864 356026 476876
rect 358170 476864 358176 476876
rect 356020 476836 358176 476864
rect 356020 476824 356026 476836
rect 358170 476824 358176 476836
rect 358228 476824 358234 476876
rect 358722 476824 358728 476876
rect 358780 476864 358786 476876
rect 361850 476864 361856 476876
rect 358780 476836 361856 476864
rect 358780 476824 358786 476836
rect 361850 476824 361856 476836
rect 361908 476824 361914 476876
rect 371050 476824 371056 476876
rect 371108 476864 371114 476876
rect 375282 476864 375288 476876
rect 371108 476836 375288 476864
rect 371108 476824 371114 476836
rect 375282 476824 375288 476836
rect 375340 476824 375346 476876
rect 376570 476824 376576 476876
rect 376628 476864 376634 476876
rect 381446 476864 381452 476876
rect 376628 476836 381452 476864
rect 376628 476824 376634 476836
rect 381446 476824 381452 476836
rect 381504 476824 381510 476876
rect 386322 476824 386328 476876
rect 386380 476864 386386 476876
rect 392394 476864 392400 476876
rect 386380 476836 392400 476864
rect 386380 476824 386386 476836
rect 392394 476824 392400 476836
rect 392452 476824 392458 476876
rect 392486 476824 392492 476876
rect 392544 476864 392550 476876
rect 393682 476864 393688 476876
rect 392544 476836 393688 476864
rect 392544 476824 392550 476836
rect 393682 476824 393688 476836
rect 393740 476824 393746 476876
rect 398742 476824 398748 476876
rect 398800 476864 398806 476876
rect 407114 476864 407120 476876
rect 398800 476836 407120 476864
rect 398800 476824 398806 476836
rect 407114 476824 407120 476836
rect 407172 476824 407178 476876
rect 514570 476824 514576 476876
rect 514628 476864 514634 476876
rect 551922 476864 551928 476876
rect 514628 476836 551928 476864
rect 514628 476824 514634 476836
rect 551922 476824 551928 476836
rect 551980 476824 551986 476876
rect 351730 476756 351736 476808
rect 351788 476796 351794 476808
rect 354582 476796 354588 476808
rect 351788 476768 354588 476796
rect 351788 476756 351794 476768
rect 354582 476756 354588 476768
rect 354640 476756 354646 476808
rect 383562 476756 383568 476808
rect 383620 476796 383626 476808
rect 390002 476796 390008 476808
rect 383620 476768 390008 476796
rect 383620 476756 383626 476768
rect 390002 476756 390008 476768
rect 390060 476756 390066 476808
rect 390370 476756 390376 476808
rect 390428 476796 390434 476808
rect 398558 476796 398564 476808
rect 390428 476768 398564 476796
rect 390428 476756 390434 476768
rect 398558 476756 398564 476768
rect 398616 476756 398622 476808
rect 401410 476756 401416 476808
rect 401468 476796 401474 476808
rect 410702 476796 410708 476808
rect 401468 476768 410708 476796
rect 401468 476756 401474 476768
rect 410702 476756 410708 476768
rect 410760 476756 410766 476808
rect 510522 476756 510528 476808
rect 510580 476796 510586 476808
rect 553118 476796 553124 476808
rect 510580 476768 553124 476796
rect 510580 476756 510586 476768
rect 553118 476756 553124 476768
rect 553176 476756 553182 476808
rect 361390 476688 361396 476740
rect 361448 476728 361454 476740
rect 364334 476728 364340 476740
rect 361448 476700 364340 476728
rect 361448 476688 361454 476700
rect 364334 476688 364340 476700
rect 364392 476688 364398 476740
rect 371142 476688 371148 476740
rect 371200 476728 371206 476740
rect 376570 476728 376576 476740
rect 371200 476700 376576 476728
rect 371200 476688 371206 476700
rect 376570 476688 376576 476700
rect 376628 476688 376634 476740
rect 394602 476688 394608 476740
rect 394660 476728 394666 476740
rect 402238 476728 402244 476740
rect 394660 476700 402244 476728
rect 394660 476688 394666 476700
rect 402238 476688 402244 476700
rect 402296 476688 402302 476740
rect 365622 476620 365628 476672
rect 365680 476660 365686 476672
rect 369210 476660 369216 476672
rect 365680 476632 369216 476660
rect 365680 476620 365686 476632
rect 369210 476620 369216 476632
rect 369268 476620 369274 476672
rect 333974 476552 333980 476604
rect 334032 476592 334038 476604
rect 334986 476592 334992 476604
rect 334032 476564 334992 476592
rect 334032 476552 334038 476564
rect 334986 476552 334992 476564
rect 335044 476552 335050 476604
rect 349062 476552 349068 476604
rect 349120 476592 349126 476604
rect 350902 476592 350908 476604
rect 349120 476564 350908 476592
rect 349120 476552 349126 476564
rect 350902 476552 350908 476564
rect 350960 476552 350966 476604
rect 357342 476552 357348 476604
rect 357400 476592 357406 476604
rect 360654 476592 360660 476604
rect 357400 476564 360660 476592
rect 357400 476552 357406 476564
rect 360654 476552 360660 476564
rect 360712 476552 360718 476604
rect 366910 476552 366916 476604
rect 366968 476592 366974 476604
rect 371602 476592 371608 476604
rect 366968 476564 371608 476592
rect 366968 476552 366974 476564
rect 371602 476552 371608 476564
rect 371660 476552 371666 476604
rect 547322 476552 547328 476604
rect 547380 476592 547386 476604
rect 553302 476592 553308 476604
rect 547380 476564 553308 476592
rect 547380 476552 547386 476564
rect 553302 476552 553308 476564
rect 553360 476552 553366 476604
rect 360102 476484 360108 476536
rect 360160 476524 360166 476536
rect 363046 476524 363052 476536
rect 360160 476496 363052 476524
rect 360160 476484 360166 476496
rect 363046 476484 363052 476496
rect 363104 476484 363110 476536
rect 331398 476416 331404 476468
rect 331456 476456 331462 476468
rect 332502 476456 332508 476468
rect 331456 476428 332508 476456
rect 331456 476416 331462 476428
rect 332502 476416 332508 476428
rect 332560 476416 332566 476468
rect 378042 476416 378048 476468
rect 378100 476456 378106 476468
rect 383838 476456 383844 476468
rect 378100 476428 383844 476456
rect 378100 476416 378106 476428
rect 383838 476416 383844 476428
rect 383896 476416 383902 476468
rect 387702 476416 387708 476468
rect 387760 476456 387766 476468
rect 394878 476456 394884 476468
rect 387760 476428 394884 476456
rect 387760 476416 387766 476428
rect 394878 476416 394884 476428
rect 394936 476416 394942 476468
rect 347682 476348 347688 476400
rect 347740 476388 347746 476400
rect 349614 476388 349620 476400
rect 347740 476360 349620 476388
rect 347740 476348 347746 476360
rect 349614 476348 349620 476360
rect 349672 476348 349678 476400
rect 367002 476348 367008 476400
rect 367060 476388 367066 476400
rect 370406 476388 370412 476400
rect 367060 476360 370412 476388
rect 367060 476348 367066 476360
rect 370406 476348 370412 476360
rect 370464 476348 370470 476400
rect 379422 476348 379428 476400
rect 379480 476388 379486 476400
rect 385126 476388 385132 476400
rect 379480 476360 385132 476388
rect 379480 476348 379486 476360
rect 385126 476348 385132 476360
rect 385184 476348 385190 476400
rect 346302 476280 346308 476332
rect 346360 476320 346366 476332
rect 348418 476320 348424 476332
rect 346360 476292 348424 476320
rect 346360 476280 346366 476292
rect 348418 476280 348424 476292
rect 348476 476280 348482 476332
rect 552658 476280 552664 476332
rect 552716 476320 552722 476332
rect 555234 476320 555240 476332
rect 552716 476292 555240 476320
rect 552716 476280 552722 476292
rect 555234 476280 555240 476292
rect 555292 476280 555298 476332
rect 380710 476212 380716 476264
rect 380768 476252 380774 476264
rect 386322 476252 386328 476264
rect 380768 476224 386328 476252
rect 380768 476212 380774 476224
rect 386322 476212 386328 476224
rect 386380 476212 386386 476264
rect 376662 476144 376668 476196
rect 376720 476184 376726 476196
rect 382642 476184 382648 476196
rect 376720 476156 382648 476184
rect 376720 476144 376726 476156
rect 382642 476144 382648 476156
rect 382700 476144 382706 476196
rect 384942 476144 384948 476196
rect 385000 476184 385006 476196
rect 391198 476184 391204 476196
rect 385000 476156 391204 476184
rect 385000 476144 385006 476156
rect 391198 476144 391204 476156
rect 391256 476144 391262 476196
rect 158806 476076 158812 476128
rect 158864 476116 158870 476128
rect 158990 476116 158996 476128
rect 158864 476088 158996 476116
rect 158864 476076 158870 476088
rect 158990 476076 158996 476088
rect 159048 476076 159054 476128
rect 538122 475736 538128 475788
rect 538180 475776 538186 475788
rect 551738 475776 551744 475788
rect 538180 475748 551744 475776
rect 538180 475736 538186 475748
rect 551738 475736 551744 475748
rect 551796 475736 551802 475788
rect 536742 475668 536748 475720
rect 536800 475708 536806 475720
rect 554314 475708 554320 475720
rect 536800 475680 554320 475708
rect 536800 475668 536806 475680
rect 554314 475668 554320 475680
rect 554372 475668 554378 475720
rect 532602 475600 532608 475652
rect 532660 475640 532666 475652
rect 551646 475640 551652 475652
rect 532660 475612 551652 475640
rect 532660 475600 532666 475612
rect 551646 475600 551652 475612
rect 551704 475600 551710 475652
rect 528462 475532 528468 475584
rect 528520 475572 528526 475584
rect 528520 475544 549116 475572
rect 528520 475532 528526 475544
rect 525702 475464 525708 475516
rect 525760 475504 525766 475516
rect 549088 475504 549116 475544
rect 549162 475532 549168 475584
rect 549220 475572 549226 475584
rect 551554 475572 551560 475584
rect 549220 475544 551560 475572
rect 549220 475532 549226 475544
rect 551554 475532 551560 475544
rect 551612 475532 551618 475584
rect 552842 475504 552848 475516
rect 525760 475476 549024 475504
rect 549088 475476 552848 475504
rect 525760 475464 525766 475476
rect 524322 475396 524328 475448
rect 524380 475436 524386 475448
rect 547414 475436 547420 475448
rect 524380 475408 547420 475436
rect 524380 475396 524386 475408
rect 547414 475396 547420 475408
rect 547472 475396 547478 475448
rect 548996 475436 549024 475476
rect 552842 475464 552848 475476
rect 552900 475464 552906 475516
rect 552934 475436 552940 475448
rect 548996 475408 552940 475436
rect 552934 475396 552940 475408
rect 552992 475396 552998 475448
rect 499482 475328 499488 475380
rect 499540 475368 499546 475380
rect 552566 475368 552572 475380
rect 499540 475340 552572 475368
rect 499540 475328 499546 475340
rect 552566 475328 552572 475340
rect 552624 475328 552630 475380
rect 499298 474716 499304 474768
rect 499356 474756 499362 474768
rect 501598 474756 501604 474768
rect 499356 474728 501604 474756
rect 499356 474716 499362 474728
rect 501598 474716 501604 474728
rect 501656 474716 501662 474768
rect 547414 474512 547420 474564
rect 547472 474552 547478 474564
rect 555326 474552 555332 474564
rect 547472 474524 555332 474552
rect 547472 474512 547478 474524
rect 555326 474512 555332 474524
rect 555384 474512 555390 474564
rect 545022 474444 545028 474496
rect 545080 474484 545086 474496
rect 553394 474484 553400 474496
rect 545080 474456 553400 474484
rect 545080 474444 545086 474456
rect 553394 474444 553400 474456
rect 553452 474444 553458 474496
rect 540882 474376 540888 474428
rect 540940 474416 540946 474428
rect 555602 474416 555608 474428
rect 540940 474388 555608 474416
rect 540940 474376 540946 474388
rect 555602 474376 555608 474388
rect 555660 474376 555666 474428
rect 533982 474308 533988 474360
rect 534040 474348 534046 474360
rect 551830 474348 551836 474360
rect 534040 474320 551836 474348
rect 534040 474308 534046 474320
rect 551830 474308 551836 474320
rect 551888 474308 551894 474360
rect 529842 474240 529848 474292
rect 529900 474280 529906 474292
rect 555786 474280 555792 474292
rect 529900 474252 555792 474280
rect 529900 474240 529906 474252
rect 555786 474240 555792 474252
rect 555844 474240 555850 474292
rect 516042 474172 516048 474224
rect 516100 474212 516106 474224
rect 552658 474212 552664 474224
rect 516100 474184 552664 474212
rect 516100 474172 516106 474184
rect 552658 474172 552664 474184
rect 552716 474172 552722 474224
rect 514662 474104 514668 474156
rect 514720 474144 514726 474156
rect 555878 474144 555884 474156
rect 514720 474116 555884 474144
rect 514720 474104 514726 474116
rect 555878 474104 555884 474116
rect 555936 474104 555942 474156
rect 511902 474036 511908 474088
rect 511960 474076 511966 474088
rect 511960 474048 552520 474076
rect 511960 474036 511966 474048
rect 498102 473968 498108 474020
rect 498160 474008 498166 474020
rect 552382 474008 552388 474020
rect 498160 473980 552388 474008
rect 498160 473968 498166 473980
rect 552382 473968 552388 473980
rect 552440 473968 552446 474020
rect 552492 474008 552520 474048
rect 554682 474036 554688 474088
rect 554740 474076 554746 474088
rect 555142 474076 555148 474088
rect 554740 474048 555148 474076
rect 554740 474036 554746 474048
rect 555142 474036 555148 474048
rect 555200 474036 555206 474088
rect 556062 474008 556068 474020
rect 552492 473980 556068 474008
rect 556062 473968 556068 473980
rect 556120 473968 556126 474020
rect 481634 473696 481640 473748
rect 481692 473736 481698 473748
rect 490650 473736 490656 473748
rect 481692 473708 490656 473736
rect 481692 473696 481698 473708
rect 490650 473696 490656 473708
rect 490708 473696 490714 473748
rect 520550 473628 520556 473680
rect 520608 473668 520614 473680
rect 522666 473668 522672 473680
rect 520608 473640 522672 473668
rect 520608 473628 520614 473640
rect 522666 473628 522672 473640
rect 522724 473628 522730 473680
rect 505002 473560 505008 473612
rect 505060 473600 505066 473612
rect 512638 473600 512644 473612
rect 505060 473572 512644 473600
rect 505060 473560 505066 473572
rect 512638 473560 512644 473572
rect 512696 473560 512702 473612
rect 520458 473560 520464 473612
rect 520516 473600 520522 473612
rect 522850 473600 522856 473612
rect 520516 473572 522856 473600
rect 520516 473560 520522 473572
rect 522850 473560 522856 473572
rect 522908 473560 522914 473612
rect 154298 473492 154304 473544
rect 154356 473492 154362 473544
rect 520384 473504 524460 473532
rect 154316 473408 154344 473492
rect 491846 473424 491852 473476
rect 491904 473424 491910 473476
rect 493134 473424 493140 473476
rect 493192 473424 493198 473476
rect 508498 473424 508504 473476
rect 508556 473424 508562 473476
rect 154298 473356 154304 473408
rect 154356 473356 154362 473408
rect 283006 473356 283012 473408
rect 283064 473396 283070 473408
rect 283282 473396 283288 473408
rect 283064 473368 283288 473396
rect 283064 473356 283070 473368
rect 283282 473356 283288 473368
rect 283340 473356 283346 473408
rect 314654 473356 314660 473408
rect 314712 473396 314718 473408
rect 315942 473396 315948 473408
rect 314712 473368 315948 473396
rect 314712 473356 314718 473368
rect 315942 473356 315948 473368
rect 316000 473396 316006 473408
rect 447778 473396 447784 473408
rect 316000 473368 447784 473396
rect 316000 473356 316006 473368
rect 447778 473356 447784 473368
rect 447836 473356 447842 473408
rect 155770 473288 155776 473340
rect 155828 473328 155834 473340
rect 156138 473328 156144 473340
rect 155828 473300 156144 473328
rect 155828 473288 155834 473300
rect 156138 473288 156144 473300
rect 156196 473288 156202 473340
rect 158898 473288 158904 473340
rect 158956 473328 158962 473340
rect 158990 473328 158996 473340
rect 158956 473300 158996 473328
rect 158956 473288 158962 473300
rect 158990 473288 158996 473300
rect 159048 473288 159054 473340
rect 283006 473220 283012 473272
rect 283064 473260 283070 473272
rect 283190 473260 283196 473272
rect 283064 473232 283196 473260
rect 283064 473220 283070 473232
rect 283190 473220 283196 473232
rect 283248 473220 283254 473272
rect 491864 472852 491892 473424
rect 493152 472988 493180 473424
rect 508516 473328 508544 473424
rect 520384 473328 520412 473504
rect 520458 473424 520464 473476
rect 520516 473424 520522 473476
rect 520550 473424 520556 473476
rect 520608 473424 520614 473476
rect 520734 473424 520740 473476
rect 520792 473424 520798 473476
rect 522666 473424 522672 473476
rect 522724 473424 522730 473476
rect 522850 473424 522856 473476
rect 522908 473424 522914 473476
rect 524432 473464 524460 473504
rect 524432 473436 528508 473464
rect 508516 473300 520412 473328
rect 520476 473056 520504 473424
rect 508056 473028 520504 473056
rect 508056 472988 508084 473028
rect 493152 472960 499344 472988
rect 499316 472852 499344 472960
rect 507872 472960 508084 472988
rect 507872 472852 507900 472960
rect 491864 472824 495388 472852
rect 499316 472824 507900 472852
rect 495360 472716 495388 472824
rect 520568 472716 520596 473424
rect 495360 472688 502380 472716
rect 502352 472580 502380 472688
rect 519556 472688 520596 472716
rect 519556 472580 519584 472688
rect 520752 472580 520780 473424
rect 522684 472784 522712 473424
rect 522868 472852 522896 473424
rect 528480 472920 528508 473436
rect 542906 473424 542912 473476
rect 542964 473424 542970 473476
rect 542924 473328 542952 473424
rect 551462 473328 551468 473340
rect 542924 473300 551468 473328
rect 551462 473288 551468 473300
rect 551520 473288 551526 473340
rect 553026 472920 553032 472932
rect 528480 472892 553032 472920
rect 553026 472880 553032 472892
rect 553084 472880 553090 472932
rect 552198 472852 552204 472864
rect 522868 472824 552204 472852
rect 552198 472812 552204 472824
rect 552256 472812 552262 472864
rect 522684 472756 525104 472784
rect 502352 472552 519584 472580
rect 520660 472552 520780 472580
rect 520660 472172 520688 472552
rect 525076 472376 525104 472756
rect 552106 472608 552112 472660
rect 552164 472648 552170 472660
rect 552164 472620 553072 472648
rect 552164 472608 552170 472620
rect 553044 472592 553072 472620
rect 553026 472540 553032 472592
rect 553084 472540 553090 472592
rect 552106 472444 552112 472456
rect 536760 472416 552112 472444
rect 536760 472376 536788 472416
rect 552106 472404 552112 472416
rect 552164 472404 552170 472456
rect 525076 472348 536788 472376
rect 551554 472268 551560 472320
rect 551612 472308 551618 472320
rect 552106 472308 552112 472320
rect 551612 472280 552112 472308
rect 551612 472268 551618 472280
rect 552106 472268 552112 472280
rect 552164 472268 552170 472320
rect 551462 472200 551468 472252
rect 551520 472240 551526 472252
rect 552198 472240 552204 472252
rect 551520 472212 552204 472240
rect 551520 472200 551526 472212
rect 552198 472200 552204 472212
rect 552256 472200 552262 472252
rect 520660 472144 520780 472172
rect 520752 472036 520780 472144
rect 551554 472132 551560 472184
rect 551612 472172 551618 472184
rect 551738 472172 551744 472184
rect 551612 472144 551744 472172
rect 551612 472132 551618 472144
rect 551738 472132 551744 472144
rect 551796 472132 551802 472184
rect 520752 472008 547460 472036
rect 154298 471928 154304 471980
rect 154356 471968 154362 471980
rect 154482 471968 154488 471980
rect 154356 471940 154488 471968
rect 154356 471928 154362 471940
rect 154482 471928 154488 471940
rect 154540 471928 154546 471980
rect 547432 471968 547460 472008
rect 551738 471996 551744 472048
rect 551796 472036 551802 472048
rect 552750 472036 552756 472048
rect 551796 472008 552756 472036
rect 551796 471996 551802 472008
rect 552750 471996 552756 472008
rect 552808 471996 552814 472048
rect 555694 471968 555700 471980
rect 547432 471940 555700 471968
rect 555694 471928 555700 471940
rect 555752 471928 555758 471980
rect 552750 471860 552756 471912
rect 552808 471900 552814 471912
rect 553210 471900 553216 471912
rect 552808 471872 553216 471900
rect 552808 471860 552814 471872
rect 553210 471860 553216 471872
rect 553268 471860 553274 471912
rect 551646 471792 551652 471844
rect 551704 471832 551710 471844
rect 551704 471804 551784 471832
rect 551704 471792 551710 471804
rect 551756 471232 551784 471804
rect 552474 471724 552480 471776
rect 552532 471764 552538 471776
rect 552934 471764 552940 471776
rect 552532 471736 552940 471764
rect 552532 471724 552538 471736
rect 552934 471724 552940 471736
rect 552992 471724 552998 471776
rect 552934 471520 552940 471572
rect 552992 471560 552998 471572
rect 553026 471560 553032 471572
rect 552992 471532 553032 471560
rect 552992 471520 552998 471532
rect 553026 471520 553032 471532
rect 553084 471520 553090 471572
rect 551738 471180 551744 471232
rect 551796 471180 551802 471232
rect 551830 470636 551836 470688
rect 551888 470676 551894 470688
rect 552290 470676 552296 470688
rect 551888 470648 552296 470676
rect 551888 470636 551894 470648
rect 552290 470636 552296 470648
rect 552348 470636 552354 470688
rect 552382 469956 552388 470008
rect 552440 469996 552446 470008
rect 552842 469996 552848 470008
rect 552440 469968 552848 469996
rect 552440 469956 552446 469968
rect 552842 469956 552848 469968
rect 552900 469956 552906 470008
rect 554866 469140 554872 469192
rect 554924 469180 554930 469192
rect 555326 469180 555332 469192
rect 554924 469152 555332 469180
rect 554924 469140 554930 469152
rect 555326 469140 555332 469152
rect 555384 469140 555390 469192
rect 555326 469004 555332 469056
rect 555384 469044 555390 469056
rect 555602 469044 555608 469056
rect 555384 469016 555608 469044
rect 555384 469004 555390 469016
rect 555602 469004 555608 469016
rect 555660 469004 555666 469056
rect 555602 468868 555608 468920
rect 555660 468908 555666 468920
rect 555786 468908 555792 468920
rect 555660 468880 555792 468908
rect 555660 468868 555666 468880
rect 555786 468868 555792 468880
rect 555844 468868 555850 468920
rect 552934 468392 552940 468444
rect 552992 468432 552998 468444
rect 553210 468432 553216 468444
rect 552992 468404 553216 468432
rect 552992 468392 552998 468404
rect 553210 468392 553216 468404
rect 553268 468392 553274 468444
rect 558546 467780 558552 467832
rect 558604 467820 558610 467832
rect 559558 467820 559564 467832
rect 558604 467792 559564 467820
rect 558604 467780 558610 467792
rect 559558 467780 559564 467792
rect 559616 467780 559622 467832
rect 158990 466460 158996 466472
rect 158916 466432 158996 466460
rect 158916 466404 158944 466432
rect 158990 466420 158996 466432
rect 159048 466420 159054 466472
rect 552658 466420 552664 466472
rect 552716 466460 552722 466472
rect 552750 466460 552756 466472
rect 552716 466432 552756 466460
rect 552716 466420 552722 466432
rect 552750 466420 552756 466432
rect 552808 466420 552814 466472
rect 158898 466352 158904 466404
rect 158956 466352 158962 466404
rect 551738 466352 551744 466404
rect 551796 466352 551802 466404
rect 552474 466352 552480 466404
rect 552532 466392 552538 466404
rect 553118 466392 553124 466404
rect 552532 466364 553124 466392
rect 552532 466352 552538 466364
rect 553118 466352 553124 466364
rect 553176 466352 553182 466404
rect 551756 466200 551784 466352
rect 551738 466148 551744 466200
rect 551796 466148 551802 466200
rect 552658 463700 552664 463752
rect 552716 463740 552722 463752
rect 552750 463740 552756 463752
rect 552716 463712 552756 463740
rect 552716 463700 552722 463712
rect 552750 463700 552756 463712
rect 552808 463700 552814 463752
rect 154298 462340 154304 462392
rect 154356 462380 154362 462392
rect 154482 462380 154488 462392
rect 154356 462352 154488 462380
rect 154356 462340 154362 462352
rect 154482 462340 154488 462352
rect 154540 462340 154546 462392
rect 556890 462340 556896 462392
rect 556948 462380 556954 462392
rect 558546 462380 558552 462392
rect 556948 462352 558552 462380
rect 556948 462340 556954 462352
rect 558546 462340 558552 462352
rect 558604 462340 558610 462392
rect 563698 462340 563704 462392
rect 563756 462380 563762 462392
rect 580166 462380 580172 462392
rect 563756 462352 580172 462380
rect 563756 462340 563762 462352
rect 580166 462340 580172 462352
rect 580224 462340 580230 462392
rect 552382 461592 552388 461644
rect 552440 461632 552446 461644
rect 552566 461632 552572 461644
rect 552440 461604 552572 461632
rect 552440 461592 552446 461604
rect 552566 461592 552572 461604
rect 552624 461592 552630 461644
rect 183646 460912 183652 460964
rect 183704 460952 183710 460964
rect 183830 460952 183836 460964
rect 183704 460924 183836 460952
rect 183704 460912 183710 460924
rect 183830 460912 183836 460924
rect 183888 460912 183894 460964
rect 551830 460844 551836 460896
rect 551888 460884 551894 460896
rect 553026 460884 553032 460896
rect 551888 460856 553032 460884
rect 551888 460844 551894 460856
rect 553026 460844 553032 460856
rect 553084 460844 553090 460896
rect 551738 460708 551744 460760
rect 551796 460748 551802 460760
rect 552382 460748 552388 460760
rect 551796 460720 552388 460748
rect 551796 460708 551802 460720
rect 552382 460708 552388 460720
rect 552440 460708 552446 460760
rect 552382 460572 552388 460624
rect 552440 460612 552446 460624
rect 553118 460612 553124 460624
rect 552440 460584 553124 460612
rect 552440 460572 552446 460584
rect 553118 460572 553124 460584
rect 553176 460572 553182 460624
rect 551738 459824 551744 459876
rect 551796 459864 551802 459876
rect 551922 459864 551928 459876
rect 551796 459836 551928 459864
rect 551796 459824 551802 459836
rect 551922 459824 551928 459836
rect 551980 459824 551986 459876
rect 551738 459280 551744 459332
rect 551796 459320 551802 459332
rect 552474 459320 552480 459332
rect 551796 459292 552480 459320
rect 551796 459280 551802 459292
rect 552474 459280 552480 459292
rect 552532 459280 552538 459332
rect 158806 456764 158812 456816
rect 158864 456804 158870 456816
rect 158990 456804 158996 456816
rect 158864 456776 158996 456804
rect 158864 456764 158870 456776
rect 158990 456764 158996 456776
rect 159048 456764 159054 456816
rect 551738 456764 551744 456816
rect 551796 456804 551802 456816
rect 552658 456804 552664 456816
rect 551796 456776 552664 456804
rect 551796 456764 551802 456776
rect 552658 456764 552664 456776
rect 552716 456764 552722 456816
rect 551738 456288 551744 456340
rect 551796 456328 551802 456340
rect 552750 456328 552756 456340
rect 551796 456300 552756 456328
rect 551796 456288 551802 456300
rect 552750 456288 552756 456300
rect 552808 456288 552814 456340
rect 551738 454860 551744 454912
rect 551796 454900 551802 454912
rect 552474 454900 552480 454912
rect 551796 454872 552480 454900
rect 551796 454860 551802 454872
rect 552474 454860 552480 454872
rect 552532 454860 552538 454912
rect 551738 454724 551744 454776
rect 551796 454764 551802 454776
rect 553026 454764 553032 454776
rect 551796 454736 553032 454764
rect 551796 454724 551802 454736
rect 553026 454724 553032 454736
rect 553084 454724 553090 454776
rect 552014 454112 552020 454164
rect 552072 454152 552078 454164
rect 552474 454152 552480 454164
rect 552072 454124 552480 454152
rect 552072 454112 552078 454124
rect 552474 454112 552480 454124
rect 552532 454112 552538 454164
rect 155770 453976 155776 454028
rect 155828 454016 155834 454028
rect 155862 454016 155868 454028
rect 155828 453988 155868 454016
rect 155828 453976 155834 453988
rect 155862 453976 155868 453988
rect 155920 453976 155926 454028
rect 158898 453976 158904 454028
rect 158956 454016 158962 454028
rect 158990 454016 158996 454028
rect 158956 453988 158996 454016
rect 158956 453976 158962 453988
rect 158990 453976 158996 453988
rect 159048 453976 159054 454028
rect 154298 452548 154304 452600
rect 154356 452588 154362 452600
rect 154482 452588 154488 452600
rect 154356 452560 154488 452588
rect 154356 452548 154362 452560
rect 154482 452548 154488 452560
rect 154540 452548 154546 452600
rect 552198 452004 552204 452056
rect 552256 452044 552262 452056
rect 552566 452044 552572 452056
rect 552256 452016 552572 452044
rect 552256 452004 552262 452016
rect 552566 452004 552572 452016
rect 552624 452004 552630 452056
rect 552198 451868 552204 451920
rect 552256 451908 552262 451920
rect 552474 451908 552480 451920
rect 552256 451880 552480 451908
rect 552256 451868 552262 451880
rect 552474 451868 552480 451880
rect 552532 451868 552538 451920
rect 3418 451256 3424 451308
rect 3476 451296 3482 451308
rect 11790 451296 11796 451308
rect 3476 451268 11796 451296
rect 3476 451256 3482 451268
rect 11790 451256 11796 451268
rect 11848 451256 11854 451308
rect 155862 447108 155868 447160
rect 155920 447108 155926 447160
rect 158990 447148 158996 447160
rect 158916 447120 158996 447148
rect 155770 447040 155776 447092
rect 155828 447080 155834 447092
rect 155880 447080 155908 447108
rect 158916 447092 158944 447120
rect 158990 447108 158996 447120
rect 159048 447108 159054 447160
rect 282914 447108 282920 447160
rect 282972 447108 282978 447160
rect 155828 447052 155908 447080
rect 155828 447040 155834 447052
rect 158898 447040 158904 447092
rect 158956 447040 158962 447092
rect 282932 447080 282960 447108
rect 283006 447080 283012 447092
rect 282932 447052 283012 447080
rect 283006 447040 283012 447052
rect 283064 447040 283070 447092
rect 9122 444320 9128 444372
rect 9180 444360 9186 444372
rect 12618 444360 12624 444372
rect 9180 444332 12624 444360
rect 9180 444320 9186 444332
rect 12618 444320 12624 444332
rect 12676 444320 12682 444372
rect 282730 444320 282736 444372
rect 282788 444360 282794 444372
rect 283006 444360 283012 444372
rect 282788 444332 283012 444360
rect 282788 444320 282794 444332
rect 283006 444320 283012 444332
rect 283064 444320 283070 444372
rect 154298 442960 154304 443012
rect 154356 443000 154362 443012
rect 154482 443000 154488 443012
rect 154356 442972 154488 443000
rect 154356 442960 154362 442972
rect 154482 442960 154488 442972
rect 154540 442960 154546 443012
rect 183646 441600 183652 441652
rect 183704 441640 183710 441652
rect 183830 441640 183836 441652
rect 183704 441612 183836 441640
rect 183704 441600 183710 441612
rect 183830 441600 183836 441612
rect 183888 441600 183894 441652
rect 289630 438880 289636 438932
rect 289688 438920 289694 438932
rect 313274 438920 313280 438932
rect 289688 438892 313280 438920
rect 289688 438880 289694 438892
rect 313274 438880 313280 438892
rect 313332 438880 313338 438932
rect 554866 438880 554872 438932
rect 554924 438920 554930 438932
rect 556890 438920 556896 438932
rect 554924 438892 556896 438920
rect 554924 438880 554930 438892
rect 556890 438880 556896 438892
rect 556948 438880 556954 438932
rect 3510 437452 3516 437504
rect 3568 437492 3574 437504
rect 13078 437492 13084 437504
rect 3568 437464 13084 437492
rect 3568 437452 3574 437464
rect 13078 437452 13084 437464
rect 13136 437452 13142 437504
rect 158806 437452 158812 437504
rect 158864 437492 158870 437504
rect 158990 437492 158996 437504
rect 158864 437464 158996 437492
rect 158864 437452 158870 437464
rect 158990 437452 158996 437464
rect 159048 437452 159054 437504
rect 554774 437248 554780 437300
rect 554832 437288 554838 437300
rect 557626 437288 557632 437300
rect 554832 437260 557632 437288
rect 554832 437248 554838 437260
rect 557626 437248 557632 437260
rect 557684 437248 557690 437300
rect 551738 436908 551744 436960
rect 551796 436948 551802 436960
rect 554866 436948 554872 436960
rect 551796 436920 554872 436948
rect 551796 436908 551802 436920
rect 554866 436908 554872 436920
rect 554924 436908 554930 436960
rect 554774 436500 554780 436552
rect 554832 436540 554838 436552
rect 557718 436540 557724 436552
rect 554832 436512 557724 436540
rect 554832 436500 554838 436512
rect 557718 436500 557724 436512
rect 557776 436500 557782 436552
rect 554866 436024 554872 436076
rect 554924 436064 554930 436076
rect 560294 436064 560300 436076
rect 554924 436036 560300 436064
rect 554924 436024 554930 436036
rect 560294 436024 560300 436036
rect 560352 436024 560358 436076
rect 554774 435956 554780 436008
rect 554832 435996 554838 436008
rect 558914 435996 558920 436008
rect 554832 435968 558920 435996
rect 554832 435956 554838 435968
rect 558914 435956 558920 435968
rect 558972 435956 558978 436008
rect 158898 434664 158904 434716
rect 158956 434704 158962 434716
rect 158990 434704 158996 434716
rect 158956 434676 158996 434704
rect 158956 434664 158962 434676
rect 158990 434664 158996 434676
rect 159048 434664 159054 434716
rect 554866 434664 554872 434716
rect 554924 434704 554930 434716
rect 561674 434704 561680 434716
rect 554924 434676 561680 434704
rect 554924 434664 554930 434676
rect 561674 434664 561680 434676
rect 561732 434664 561738 434716
rect 554774 434596 554780 434648
rect 554832 434636 554838 434648
rect 561766 434636 561772 434648
rect 554832 434608 561772 434636
rect 554832 434596 554838 434608
rect 561766 434596 561772 434608
rect 561824 434596 561830 434648
rect 154298 433236 154304 433288
rect 154356 433276 154362 433288
rect 154482 433276 154488 433288
rect 154356 433248 154488 433276
rect 154356 433236 154362 433248
rect 154482 433236 154488 433248
rect 154540 433236 154546 433288
rect 554866 433236 554872 433288
rect 554924 433276 554930 433288
rect 564434 433276 564440 433288
rect 554924 433248 564440 433276
rect 554924 433236 554930 433248
rect 564434 433236 564440 433248
rect 564492 433236 564498 433288
rect 554774 433168 554780 433220
rect 554832 433208 554838 433220
rect 563054 433208 563060 433220
rect 554832 433180 563060 433208
rect 554832 433168 554838 433180
rect 563054 433168 563060 433180
rect 563112 433168 563118 433220
rect 554958 431876 554964 431928
rect 555016 431916 555022 431928
rect 567286 431916 567292 431928
rect 555016 431888 567292 431916
rect 555016 431876 555022 431888
rect 567286 431876 567292 431888
rect 567344 431876 567350 431928
rect 554774 431808 554780 431860
rect 554832 431848 554838 431860
rect 565814 431848 565820 431860
rect 554832 431820 565820 431848
rect 554832 431808 554838 431820
rect 565814 431808 565820 431820
rect 565872 431808 565878 431860
rect 554866 431740 554872 431792
rect 554924 431780 554930 431792
rect 560938 431780 560944 431792
rect 554924 431752 560944 431780
rect 554924 431740 554930 431752
rect 560938 431740 560944 431752
rect 560996 431740 561002 431792
rect 554866 430516 554872 430568
rect 554924 430556 554930 430568
rect 569954 430556 569960 430568
rect 554924 430528 569960 430556
rect 554924 430516 554930 430528
rect 569954 430516 569960 430528
rect 570012 430516 570018 430568
rect 554774 430448 554780 430500
rect 554832 430488 554838 430500
rect 568574 430488 568580 430500
rect 554832 430460 568580 430488
rect 554832 430448 554838 430460
rect 568574 430448 568580 430460
rect 568632 430448 568638 430500
rect 155770 429836 155776 429888
rect 155828 429876 155834 429888
rect 156046 429876 156052 429888
rect 155828 429848 156052 429876
rect 155828 429836 155834 429848
rect 156046 429836 156052 429848
rect 156104 429836 156110 429888
rect 554774 429088 554780 429140
rect 554832 429128 554838 429140
rect 571610 429128 571616 429140
rect 554832 429100 571616 429128
rect 554832 429088 554838 429100
rect 571610 429088 571616 429100
rect 571668 429088 571674 429140
rect 554866 428884 554872 428936
rect 554924 428924 554930 428936
rect 556798 428924 556804 428936
rect 554924 428896 556804 428924
rect 554924 428884 554930 428896
rect 556798 428884 556804 428896
rect 556856 428884 556862 428936
rect 158990 427836 158996 427848
rect 158916 427808 158996 427836
rect 158916 427780 158944 427808
rect 158990 427796 158996 427808
rect 159048 427796 159054 427848
rect 282914 427796 282920 427848
rect 282972 427796 282978 427848
rect 158898 427728 158904 427780
rect 158956 427728 158962 427780
rect 282932 427768 282960 427796
rect 283006 427768 283012 427780
rect 282932 427740 283012 427768
rect 283006 427728 283012 427740
rect 283064 427728 283070 427780
rect 554774 427728 554780 427780
rect 554832 427768 554838 427780
rect 572714 427768 572720 427780
rect 554832 427740 572720 427768
rect 554832 427728 554838 427740
rect 572714 427728 572720 427740
rect 572772 427728 572778 427780
rect 447778 426368 447784 426420
rect 447836 426408 447842 426420
rect 499298 426408 499304 426420
rect 447836 426380 499304 426408
rect 447836 426368 447842 426380
rect 499298 426368 499304 426380
rect 499356 426408 499362 426420
rect 551462 426408 551468 426420
rect 499356 426380 551468 426408
rect 499356 426368 499362 426380
rect 551462 426368 551468 426380
rect 551520 426368 551526 426420
rect 155770 425144 155776 425196
rect 155828 425184 155834 425196
rect 156046 425184 156052 425196
rect 155828 425156 156052 425184
rect 155828 425144 155834 425156
rect 156046 425144 156052 425156
rect 156104 425144 156110 425196
rect 155770 425008 155776 425060
rect 155828 425048 155834 425060
rect 155862 425048 155868 425060
rect 155828 425020 155868 425048
rect 155828 425008 155834 425020
rect 155862 425008 155868 425020
rect 155920 425008 155926 425060
rect 3418 423648 3424 423700
rect 3476 423688 3482 423700
rect 14458 423688 14464 423700
rect 3476 423660 14464 423688
rect 3476 423648 3482 423660
rect 14458 423648 14464 423660
rect 14516 423648 14522 423700
rect 154298 423648 154304 423700
rect 154356 423688 154362 423700
rect 154482 423688 154488 423700
rect 154356 423660 154488 423688
rect 154356 423648 154362 423660
rect 154482 423648 154488 423660
rect 154540 423648 154546 423700
rect 183646 422288 183652 422340
rect 183704 422328 183710 422340
rect 183830 422328 183836 422340
rect 183704 422300 183836 422328
rect 183704 422288 183710 422300
rect 183830 422288 183836 422300
rect 183888 422288 183894 422340
rect 281626 421540 281632 421592
rect 281684 421580 281690 421592
rect 282178 421580 282184 421592
rect 281684 421552 282184 421580
rect 281684 421540 281690 421552
rect 282178 421540 282184 421552
rect 282236 421580 282242 421592
rect 292574 421580 292580 421592
rect 282236 421552 292580 421580
rect 282236 421540 282242 421552
rect 292574 421540 292580 421552
rect 292632 421540 292638 421592
rect 155862 418180 155868 418192
rect 155788 418152 155868 418180
rect 155788 418124 155816 418152
rect 155862 418140 155868 418152
rect 155920 418140 155926 418192
rect 158806 418140 158812 418192
rect 158864 418180 158870 418192
rect 158990 418180 158996 418192
rect 158864 418152 158996 418180
rect 158864 418140 158870 418152
rect 158990 418140 158996 418152
rect 159048 418140 159054 418192
rect 155770 418072 155776 418124
rect 155828 418072 155834 418124
rect 304350 415420 304356 415472
rect 304408 415460 304414 415472
rect 580166 415460 580172 415472
rect 304408 415432 580172 415460
rect 304408 415420 304414 415432
rect 580166 415420 580172 415432
rect 580224 415420 580230 415472
rect 155862 415352 155868 415404
rect 155920 415392 155926 415404
rect 156138 415392 156144 415404
rect 155920 415364 156144 415392
rect 155920 415352 155926 415364
rect 156138 415352 156144 415364
rect 156196 415352 156202 415404
rect 158898 415352 158904 415404
rect 158956 415392 158962 415404
rect 159174 415392 159180 415404
rect 158956 415364 159180 415392
rect 158956 415352 158962 415364
rect 159174 415352 159180 415364
rect 159232 415352 159238 415404
rect 282914 415352 282920 415404
rect 282972 415392 282978 415404
rect 283098 415392 283104 415404
rect 282972 415364 283104 415392
rect 282972 415352 282978 415364
rect 283098 415352 283104 415364
rect 283156 415352 283162 415404
rect 154298 413924 154304 413976
rect 154356 413964 154362 413976
rect 154482 413964 154488 413976
rect 154356 413936 154488 413964
rect 154356 413924 154362 413936
rect 154482 413924 154488 413936
rect 154540 413924 154546 413976
rect 158990 405696 158996 405748
rect 159048 405736 159054 405748
rect 159174 405736 159180 405748
rect 159048 405708 159180 405736
rect 159048 405696 159054 405708
rect 159174 405696 159180 405708
rect 159232 405696 159238 405748
rect 282914 405696 282920 405748
rect 282972 405736 282978 405748
rect 283190 405736 283196 405748
rect 282972 405708 283196 405736
rect 282972 405696 282978 405708
rect 283190 405696 283196 405708
rect 283248 405696 283254 405748
rect 154298 404336 154304 404388
rect 154356 404376 154362 404388
rect 154482 404376 154488 404388
rect 154356 404348 154488 404376
rect 154356 404336 154362 404348
rect 154482 404336 154488 404348
rect 154540 404336 154546 404388
rect 183646 402976 183652 403028
rect 183704 403016 183710 403028
rect 183830 403016 183836 403028
rect 183704 402988 183836 403016
rect 183704 402976 183710 402988
rect 183830 402976 183836 402988
rect 183888 402976 183894 403028
rect 140682 401548 140688 401600
rect 140740 401588 140746 401600
rect 153746 401588 153752 401600
rect 140740 401560 153752 401588
rect 140740 401548 140746 401560
rect 153746 401548 153752 401560
rect 153804 401548 153810 401600
rect 140590 401480 140596 401532
rect 140648 401520 140654 401532
rect 155034 401520 155040 401532
rect 140648 401492 155040 401520
rect 140648 401480 140654 401492
rect 155034 401480 155040 401492
rect 155092 401480 155098 401532
rect 139302 401412 139308 401464
rect 139360 401452 139366 401464
rect 154206 401452 154212 401464
rect 139360 401424 154212 401452
rect 139360 401412 139366 401424
rect 154206 401412 154212 401424
rect 154264 401412 154270 401464
rect 136542 401344 136548 401396
rect 136600 401384 136606 401396
rect 153654 401384 153660 401396
rect 136600 401356 153660 401384
rect 136600 401344 136606 401356
rect 153654 401344 153660 401356
rect 153712 401344 153718 401396
rect 137922 401276 137928 401328
rect 137980 401316 137986 401328
rect 155126 401316 155132 401328
rect 137980 401288 155132 401316
rect 137980 401276 137986 401288
rect 155126 401276 155132 401288
rect 155184 401276 155190 401328
rect 135162 401208 135168 401260
rect 135220 401248 135226 401260
rect 153838 401248 153844 401260
rect 135220 401220 153844 401248
rect 135220 401208 135226 401220
rect 153838 401208 153844 401220
rect 153896 401208 153902 401260
rect 136450 401140 136456 401192
rect 136508 401180 136514 401192
rect 155310 401180 155316 401192
rect 136508 401152 155316 401180
rect 136508 401140 136514 401152
rect 155310 401140 155316 401152
rect 155368 401140 155374 401192
rect 132402 401072 132408 401124
rect 132460 401112 132466 401124
rect 155494 401112 155500 401124
rect 132460 401084 155500 401112
rect 132460 401072 132466 401084
rect 155494 401072 155500 401084
rect 155552 401072 155558 401124
rect 133782 401004 133788 401056
rect 133840 401044 133846 401056
rect 157426 401044 157432 401056
rect 133840 401016 157432 401044
rect 133840 401004 133846 401016
rect 157426 401004 157432 401016
rect 157484 401004 157490 401056
rect 125410 400936 125416 400988
rect 125468 400976 125474 400988
rect 155218 400976 155224 400988
rect 125468 400948 155224 400976
rect 125468 400936 125474 400948
rect 155218 400936 155224 400948
rect 155276 400936 155282 400988
rect 122742 400868 122748 400920
rect 122800 400908 122806 400920
rect 155586 400908 155592 400920
rect 122800 400880 155592 400908
rect 122800 400868 122806 400880
rect 155586 400868 155592 400880
rect 155644 400868 155650 400920
rect 142062 400800 142068 400852
rect 142120 400840 142126 400852
rect 153562 400840 153568 400852
rect 142120 400812 153568 400840
rect 142120 400800 142126 400812
rect 153562 400800 153568 400812
rect 153620 400800 153626 400852
rect 143442 400732 143448 400784
rect 143500 400772 143506 400784
rect 154022 400772 154028 400784
rect 143500 400744 154028 400772
rect 143500 400732 143506 400744
rect 154022 400732 154028 400744
rect 154080 400732 154086 400784
rect 144822 400664 144828 400716
rect 144880 400704 144886 400716
rect 155402 400704 155408 400716
rect 144880 400676 155408 400704
rect 144880 400664 144886 400676
rect 155402 400664 155408 400676
rect 155460 400664 155466 400716
rect 146202 400596 146208 400648
rect 146260 400636 146266 400648
rect 154114 400636 154120 400648
rect 146260 400608 154120 400636
rect 146260 400596 146266 400608
rect 154114 400596 154120 400608
rect 154172 400596 154178 400648
rect 146110 400256 146116 400308
rect 146168 400296 146174 400308
rect 153930 400296 153936 400308
rect 146168 400268 153936 400296
rect 146168 400256 146174 400268
rect 153930 400256 153936 400268
rect 153988 400256 153994 400308
rect 154114 394612 154120 394664
rect 154172 394652 154178 394664
rect 154298 394652 154304 394664
rect 154172 394624 154304 394652
rect 154172 394612 154178 394624
rect 154298 394612 154304 394624
rect 154356 394612 154362 394664
rect 155770 394612 155776 394664
rect 155828 394652 155834 394664
rect 155862 394652 155868 394664
rect 155828 394624 155868 394652
rect 155828 394612 155834 394624
rect 155862 394612 155868 394624
rect 155920 394612 155926 394664
rect 158806 386316 158812 386368
rect 158864 386356 158870 386368
rect 158990 386356 158996 386368
rect 158864 386328 158996 386356
rect 158864 386316 158870 386328
rect 158990 386316 158996 386328
rect 159048 386316 159054 386368
rect 154114 385024 154120 385076
rect 154172 385064 154178 385076
rect 154298 385064 154304 385076
rect 154172 385036 154304 385064
rect 154172 385024 154178 385036
rect 154298 385024 154304 385036
rect 154356 385024 154362 385076
rect 183646 383664 183652 383716
rect 183704 383704 183710 383716
rect 183830 383704 183836 383716
rect 183704 383676 183836 383704
rect 183704 383664 183710 383676
rect 183830 383664 183836 383676
rect 183888 383664 183894 383716
rect 155862 379556 155868 379568
rect 155696 379528 155868 379556
rect 155696 379500 155724 379528
rect 155862 379516 155868 379528
rect 155920 379516 155926 379568
rect 155678 379448 155684 379500
rect 155736 379448 155742 379500
rect 282178 377204 282184 377256
rect 282236 377244 282242 377256
rect 284386 377244 284392 377256
rect 282236 377216 284392 377244
rect 282236 377204 282242 377216
rect 284386 377204 284392 377216
rect 284444 377204 284450 377256
rect 78582 376728 78588 376780
rect 78640 376768 78646 376780
rect 186958 376768 186964 376780
rect 78640 376740 186964 376768
rect 78640 376728 78646 376740
rect 186958 376728 186964 376740
rect 187016 376728 187022 376780
rect 154114 375300 154120 375352
rect 154172 375340 154178 375352
rect 154298 375340 154304 375352
rect 154172 375312 154304 375340
rect 154172 375300 154178 375312
rect 154298 375300 154304 375312
rect 154356 375300 154362 375352
rect 304442 368500 304448 368552
rect 304500 368540 304506 368552
rect 580166 368540 580172 368552
rect 304500 368512 580172 368540
rect 304500 368500 304506 368512
rect 580166 368500 580172 368512
rect 580224 368500 580230 368552
rect 153838 365712 153844 365764
rect 153896 365752 153902 365764
rect 154114 365752 154120 365764
rect 153896 365724 154120 365752
rect 153896 365712 153902 365724
rect 154114 365712 154120 365724
rect 154172 365712 154178 365764
rect 183646 364352 183652 364404
rect 183704 364392 183710 364404
rect 183830 364392 183836 364404
rect 183704 364364 183836 364392
rect 183704 364352 183710 364364
rect 183830 364352 183836 364364
rect 183888 364352 183894 364404
rect 155494 362244 155500 362296
rect 155552 362284 155558 362296
rect 155770 362284 155776 362296
rect 155552 362256 155776 362284
rect 155552 362244 155558 362256
rect 155770 362244 155776 362256
rect 155828 362244 155834 362296
rect 186958 360136 186964 360188
rect 187016 360176 187022 360188
rect 282178 360176 282184 360188
rect 187016 360148 282184 360176
rect 187016 360136 187022 360148
rect 282178 360136 282184 360148
rect 282236 360136 282242 360188
rect 187418 357484 187424 357536
rect 187476 357524 187482 357536
rect 191926 357524 191932 357536
rect 187476 357496 191932 357524
rect 187476 357484 187482 357496
rect 191926 357484 191932 357496
rect 191984 357484 191990 357536
rect 153838 357416 153844 357468
rect 153896 357456 153902 357468
rect 153930 357456 153936 357468
rect 153896 357428 153936 357456
rect 153896 357416 153902 357428
rect 153930 357416 153936 357428
rect 153988 357416 153994 357468
rect 155494 357416 155500 357468
rect 155552 357456 155558 357468
rect 155586 357456 155592 357468
rect 155552 357428 155592 357456
rect 155552 357416 155558 357428
rect 155586 357416 155592 357428
rect 155644 357416 155650 357468
rect 274634 356396 274640 356448
rect 274692 356436 274698 356448
rect 275646 356436 275652 356448
rect 274692 356408 275652 356436
rect 274692 356396 274698 356408
rect 275646 356396 275652 356408
rect 275704 356396 275710 356448
rect 194410 355988 194416 356040
rect 194468 356028 194474 356040
rect 198918 356028 198924 356040
rect 194468 356000 198924 356028
rect 194468 355988 194474 356000
rect 198918 355988 198924 356000
rect 198976 355988 198982 356040
rect 201402 355988 201408 356040
rect 201460 356028 201466 356040
rect 206922 356028 206928 356040
rect 201460 356000 206928 356028
rect 201460 355988 201466 356000
rect 206922 355988 206928 356000
rect 206980 355988 206986 356040
rect 210326 355988 210332 356040
rect 210384 356028 210390 356040
rect 214742 356028 214748 356040
rect 210384 356000 214748 356028
rect 210384 355988 210390 356000
rect 214742 355988 214748 356000
rect 214800 355988 214806 356040
rect 215202 355988 215208 356040
rect 215260 356028 215266 356040
rect 218974 356028 218980 356040
rect 215260 356000 218980 356028
rect 215260 355988 215266 356000
rect 218974 355988 218980 356000
rect 219032 355988 219038 356040
rect 221274 355988 221280 356040
rect 221332 356028 221338 356040
rect 222838 356028 222844 356040
rect 221332 356000 222844 356028
rect 221332 355988 221338 356000
rect 222838 355988 222844 356000
rect 222896 355988 222902 356040
rect 226150 355988 226156 356040
rect 226208 356028 226214 356040
rect 226978 356028 226984 356040
rect 226208 356000 226984 356028
rect 226208 355988 226214 356000
rect 226978 355988 226984 356000
rect 227036 355988 227042 356040
rect 227438 355988 227444 356040
rect 227496 356028 227502 356040
rect 228174 356028 228180 356040
rect 227496 356000 228180 356028
rect 227496 355988 227502 356000
rect 228174 355988 228180 356000
rect 228232 355988 228238 356040
rect 229830 355988 229836 356040
rect 229888 356028 229894 356040
rect 230474 356028 230480 356040
rect 229888 356000 230480 356028
rect 229888 355988 229894 356000
rect 230474 355988 230480 356000
rect 230532 355988 230538 356040
rect 233142 355988 233148 356040
rect 233200 356028 233206 356040
rect 233694 356028 233700 356040
rect 233200 356000 233700 356028
rect 233200 355988 233206 356000
rect 233694 355988 233700 356000
rect 233752 355988 233758 356040
rect 234522 355988 234528 356040
rect 234580 356028 234586 356040
rect 235902 356028 235908 356040
rect 234580 356000 235908 356028
rect 234580 355988 234586 356000
rect 235902 355988 235908 356000
rect 235960 355988 235966 356040
rect 237190 355988 237196 356040
rect 237248 356028 237254 356040
rect 238294 356028 238300 356040
rect 237248 356000 238300 356028
rect 237248 355988 237254 356000
rect 238294 355988 238300 356000
rect 238352 355988 238358 356040
rect 239582 355988 239588 356040
rect 239640 356028 239646 356040
rect 240502 356028 240508 356040
rect 239640 356000 240508 356028
rect 239640 355988 239646 356000
rect 240502 355988 240508 356000
rect 240560 355988 240566 356040
rect 258074 355988 258080 356040
rect 258132 356028 258138 356040
rect 258534 356028 258540 356040
rect 258132 356000 258540 356028
rect 258132 355988 258138 356000
rect 258534 355988 258540 356000
rect 258592 355988 258598 356040
rect 261570 355988 261576 356040
rect 261628 356028 261634 356040
rect 262214 356028 262220 356040
rect 261628 356000 262220 356028
rect 261628 355988 261634 356000
rect 262214 355988 262220 356000
rect 262272 355988 262278 356040
rect 262674 355988 262680 356040
rect 262732 356028 262738 356040
rect 263594 356028 263600 356040
rect 262732 356000 263600 356028
rect 262732 355988 262738 356000
rect 263594 355988 263600 356000
rect 263652 355988 263658 356040
rect 193122 355920 193128 355972
rect 193180 355960 193186 355972
rect 199654 355960 199660 355972
rect 193180 355932 199660 355960
rect 193180 355920 193186 355932
rect 199654 355920 199660 355932
rect 199712 355920 199718 355972
rect 213822 355920 213828 355972
rect 213880 355960 213886 355972
rect 218054 355960 218060 355972
rect 213880 355932 218060 355960
rect 213880 355920 213886 355932
rect 218054 355920 218060 355932
rect 218112 355920 218118 355972
rect 232314 355920 232320 355972
rect 232372 355960 232378 355972
rect 234062 355960 234068 355972
rect 232372 355932 234068 355960
rect 232372 355920 232378 355932
rect 234062 355920 234068 355932
rect 234120 355920 234126 355972
rect 235810 355920 235816 355972
rect 235868 355960 235874 355972
rect 237282 355960 237288 355972
rect 235868 355932 237288 355960
rect 235868 355920 235874 355932
rect 237282 355920 237288 355932
rect 237340 355920 237346 355972
rect 211522 355852 211528 355904
rect 211580 355892 211586 355904
rect 215662 355892 215668 355904
rect 211580 355864 215668 355892
rect 211580 355852 211586 355864
rect 215662 355852 215668 355864
rect 215720 355852 215726 355904
rect 224862 355852 224868 355904
rect 224920 355892 224926 355904
rect 227714 355892 227720 355904
rect 224920 355864 227720 355892
rect 224920 355852 224926 355864
rect 227714 355852 227720 355864
rect 227772 355852 227778 355904
rect 204162 355784 204168 355836
rect 204220 355824 204226 355836
rect 209222 355824 209228 355836
rect 204220 355796 209228 355824
rect 204220 355784 204226 355796
rect 209222 355784 209228 355796
rect 209280 355784 209286 355836
rect 222102 355784 222108 355836
rect 222160 355824 222166 355836
rect 225414 355824 225420 355836
rect 222160 355796 225420 355824
rect 222160 355784 222166 355796
rect 225414 355784 225420 355796
rect 225472 355784 225478 355836
rect 242066 355784 242072 355836
rect 242124 355824 242130 355836
rect 242802 355824 242808 355836
rect 242124 355796 242808 355824
rect 242124 355784 242130 355796
rect 242802 355784 242808 355796
rect 242860 355784 242866 355836
rect 281442 355784 281448 355836
rect 281500 355824 281506 355836
rect 281718 355824 281724 355836
rect 281500 355796 281724 355824
rect 281500 355784 281506 355796
rect 281718 355784 281724 355796
rect 281776 355784 281782 355836
rect 199286 355716 199292 355768
rect 199344 355756 199350 355768
rect 204990 355756 204996 355768
rect 199344 355728 204996 355756
rect 199344 355716 199350 355728
rect 204990 355716 204996 355728
rect 205048 355716 205054 355768
rect 198090 355648 198096 355700
rect 198148 355688 198154 355700
rect 203886 355688 203892 355700
rect 198148 355660 203892 355688
rect 198148 355648 198154 355660
rect 203886 355648 203892 355660
rect 203944 355648 203950 355700
rect 240870 355648 240876 355700
rect 240928 355688 240934 355700
rect 241698 355688 241704 355700
rect 240928 355660 241704 355688
rect 240928 355648 240934 355660
rect 241698 355648 241704 355660
rect 241756 355648 241762 355700
rect 255314 355648 255320 355700
rect 255372 355688 255378 355700
rect 256050 355688 256056 355700
rect 255372 355660 256056 355688
rect 255372 355648 255378 355660
rect 256050 355648 256056 355660
rect 256108 355648 256114 355700
rect 217594 355580 217600 355632
rect 217652 355620 217658 355632
rect 221182 355620 221188 355632
rect 217652 355592 221188 355620
rect 217652 355580 217658 355592
rect 221182 355580 221188 355592
rect 221240 355580 221246 355632
rect 200482 355512 200488 355564
rect 200540 355552 200546 355564
rect 206094 355552 206100 355564
rect 200540 355524 206100 355552
rect 200540 355512 200546 355524
rect 206094 355512 206100 355524
rect 206152 355512 206158 355564
rect 263410 355512 263416 355564
rect 263468 355552 263474 355564
rect 264606 355552 264612 355564
rect 263468 355524 264612 355552
rect 263468 355512 263474 355524
rect 264606 355512 264612 355524
rect 264664 355512 264670 355564
rect 189534 355444 189540 355496
rect 189592 355484 189598 355496
rect 196342 355484 196348 355496
rect 189592 355456 196348 355484
rect 189592 355444 189598 355456
rect 196342 355444 196348 355456
rect 196400 355444 196406 355496
rect 207842 355376 207848 355428
rect 207900 355416 207906 355428
rect 212626 355416 212632 355428
rect 207900 355388 212632 355416
rect 207900 355376 207906 355388
rect 212626 355376 212632 355388
rect 212684 355376 212690 355428
rect 218882 355376 218888 355428
rect 218940 355416 218946 355428
rect 222378 355416 222384 355428
rect 218940 355388 222384 355416
rect 218940 355376 218946 355388
rect 222378 355376 222384 355388
rect 222436 355376 222442 355428
rect 231026 355376 231032 355428
rect 231084 355416 231090 355428
rect 233142 355416 233148 355428
rect 231084 355388 233148 355416
rect 231084 355376 231090 355388
rect 233142 355376 233148 355388
rect 233200 355376 233206 355428
rect 256694 355376 256700 355428
rect 256752 355416 256758 355428
rect 257338 355416 257344 355428
rect 256752 355388 257344 355416
rect 256752 355376 256758 355388
rect 257338 355376 257344 355388
rect 257396 355376 257402 355428
rect 266078 355376 266084 355428
rect 266136 355416 266142 355428
rect 267090 355416 267096 355428
rect 266136 355388 267096 355416
rect 266136 355376 266142 355388
rect 267090 355376 267096 355388
rect 267148 355376 267154 355428
rect 190362 355308 190368 355360
rect 190420 355348 190426 355360
rect 197262 355348 197268 355360
rect 190420 355320 197268 355348
rect 190420 355308 190426 355320
rect 197262 355308 197268 355320
rect 197320 355308 197326 355360
rect 209038 355308 209044 355360
rect 209096 355348 209102 355360
rect 214006 355348 214012 355360
rect 209096 355320 214012 355348
rect 209096 355308 209102 355320
rect 214006 355308 214012 355320
rect 214064 355308 214070 355360
rect 243262 355308 243268 355360
rect 243320 355348 243326 355360
rect 243814 355348 243820 355360
rect 243320 355320 243820 355348
rect 243320 355308 243326 355320
rect 243814 355308 243820 355320
rect 243872 355308 243878 355360
rect 244090 355308 244096 355360
rect 244148 355348 244154 355360
rect 244918 355348 244924 355360
rect 244148 355320 244924 355348
rect 244148 355308 244154 355320
rect 244918 355308 244924 355320
rect 244976 355308 244982 355360
rect 220078 355240 220084 355292
rect 220136 355280 220142 355292
rect 223666 355280 223672 355292
rect 220136 355252 223672 355280
rect 220136 355240 220142 355252
rect 223666 355240 223672 355252
rect 223724 355240 223730 355292
rect 264882 355240 264888 355292
rect 264940 355280 264946 355292
rect 265894 355280 265900 355292
rect 264940 355252 265900 355280
rect 264940 355240 264946 355252
rect 265894 355240 265900 355252
rect 265952 355240 265958 355292
rect 202782 355172 202788 355224
rect 202840 355212 202846 355224
rect 208302 355212 208308 355224
rect 202840 355184 208308 355212
rect 202840 355172 202846 355184
rect 208302 355172 208308 355184
rect 208360 355172 208366 355224
rect 254118 355104 254124 355156
rect 254176 355144 254182 355156
rect 254854 355144 254860 355156
rect 254176 355116 254860 355144
rect 254176 355104 254182 355116
rect 254854 355104 254860 355116
rect 254912 355104 254918 355156
rect 268194 355104 268200 355156
rect 268252 355144 268258 355156
rect 269482 355144 269488 355156
rect 268252 355116 269488 355144
rect 268252 355104 268258 355116
rect 269482 355104 269488 355116
rect 269540 355104 269546 355156
rect 212350 354968 212356 355020
rect 212408 355008 212414 355020
rect 216766 355008 216772 355020
rect 212408 354980 216772 355008
rect 212408 354968 212414 354980
rect 216766 354968 216772 354980
rect 216824 354968 216830 355020
rect 191742 354832 191748 354884
rect 191800 354872 191806 354884
rect 194962 354872 194968 354884
rect 191800 354844 194968 354872
rect 191800 354832 191806 354844
rect 194962 354832 194968 354844
rect 195020 354832 195026 354884
rect 196802 354832 196808 354884
rect 196860 354872 196866 354884
rect 201494 354872 201500 354884
rect 196860 354844 201500 354872
rect 196860 354832 196866 354844
rect 201494 354832 201500 354844
rect 201552 354832 201558 354884
rect 223390 354832 223396 354884
rect 223448 354872 223454 354884
rect 226518 354872 226524 354884
rect 223448 354844 226524 354872
rect 223448 354832 223454 354844
rect 226518 354832 226524 354844
rect 226576 354832 226582 354884
rect 206646 354764 206652 354816
rect 206704 354804 206710 354816
rect 211430 354804 211436 354816
rect 206704 354776 211436 354804
rect 206704 354764 206710 354776
rect 211430 354764 211436 354776
rect 211488 354764 211494 354816
rect 238386 354764 238392 354816
rect 238444 354804 238450 354816
rect 239398 354804 239404 354816
rect 238444 354776 239404 354804
rect 238444 354764 238450 354776
rect 239398 354764 239404 354776
rect 239456 354764 239462 354816
rect 248046 354764 248052 354816
rect 248104 354804 248110 354816
rect 248506 354804 248512 354816
rect 248104 354776 248512 354804
rect 248104 354764 248110 354776
rect 248506 354764 248512 354776
rect 248564 354764 248570 354816
rect 188338 354696 188344 354748
rect 188396 354736 188402 354748
rect 193214 354736 193220 354748
rect 188396 354708 193220 354736
rect 188396 354696 188402 354708
rect 193214 354696 193220 354708
rect 193272 354696 193278 354748
rect 195606 354696 195612 354748
rect 195664 354736 195670 354748
rect 201402 354736 201408 354748
rect 195664 354708 201408 354736
rect 195664 354696 195670 354708
rect 201402 354696 201408 354708
rect 201460 354696 201466 354748
rect 205358 354696 205364 354748
rect 205416 354736 205422 354748
rect 210326 354736 210332 354748
rect 205416 354708 210332 354736
rect 205416 354696 205422 354708
rect 210326 354696 210332 354708
rect 210384 354696 210390 354748
rect 216398 354696 216404 354748
rect 216456 354736 216462 354748
rect 220078 354736 220084 354748
rect 216456 354708 220084 354736
rect 216456 354696 216462 354708
rect 220078 354696 220084 354708
rect 220136 354696 220142 354748
rect 228634 354696 228640 354748
rect 228692 354736 228698 354748
rect 230382 354736 230388 354748
rect 228692 354708 230388 354736
rect 228692 354696 228698 354708
rect 230382 354696 230388 354708
rect 230440 354696 230446 354748
rect 260558 354696 260564 354748
rect 260616 354736 260622 354748
rect 261018 354736 261024 354748
rect 260616 354708 261024 354736
rect 260616 354696 260622 354708
rect 261018 354696 261024 354708
rect 261076 354696 261082 354748
rect 267090 354696 267096 354748
rect 267148 354736 267154 354748
rect 268286 354736 268292 354748
rect 267148 354708 268292 354736
rect 267148 354696 267154 354708
rect 268286 354696 268292 354708
rect 268344 354696 268350 354748
rect 39942 354628 39948 354680
rect 40000 354668 40006 354680
rect 50982 354668 50988 354680
rect 40000 354640 50988 354668
rect 40000 354628 40006 354640
rect 50982 354628 50988 354640
rect 51040 354628 51046 354680
rect 51442 354628 51448 354680
rect 51500 354668 51506 354680
rect 63586 354668 63592 354680
rect 51500 354640 63592 354668
rect 51500 354628 51506 354640
rect 63586 354628 63592 354640
rect 63644 354628 63650 354680
rect 48314 354560 48320 354612
rect 48372 354600 48378 354612
rect 59630 354600 59636 354612
rect 48372 354572 59636 354600
rect 48372 354560 48378 354572
rect 59630 354560 59636 354572
rect 59688 354560 59694 354612
rect 61562 354560 61568 354612
rect 61620 354600 61626 354612
rect 70394 354600 70400 354612
rect 61620 354572 70400 354600
rect 61620 354560 61626 354572
rect 70394 354560 70400 354572
rect 70452 354560 70458 354612
rect 33502 354492 33508 354544
rect 33560 354532 33566 354544
rect 38654 354532 38660 354544
rect 33560 354504 38660 354532
rect 33560 354492 33566 354504
rect 38654 354492 38660 354504
rect 38712 354492 38718 354544
rect 45002 354492 45008 354544
rect 45060 354532 45066 354544
rect 56962 354532 56968 354544
rect 45060 354504 56968 354532
rect 45060 354492 45066 354504
rect 56962 354492 56968 354504
rect 57020 354492 57026 354544
rect 58618 354492 58624 354544
rect 58676 354532 58682 354544
rect 68922 354532 68928 354544
rect 58676 354504 68928 354532
rect 58676 354492 58682 354504
rect 68922 354492 68928 354504
rect 68980 354492 68986 354544
rect 70854 354492 70860 354544
rect 70912 354532 70918 354544
rect 80054 354532 80060 354544
rect 70912 354504 80060 354532
rect 70912 354492 70918 354504
rect 80054 354492 80060 354504
rect 80112 354492 80118 354544
rect 35618 354424 35624 354476
rect 35676 354464 35682 354476
rect 40310 354464 40316 354476
rect 35676 354436 40316 354464
rect 35676 354424 35682 354436
rect 40310 354424 40316 354436
rect 40368 354424 40374 354476
rect 46474 354424 46480 354476
rect 46532 354464 46538 354476
rect 58066 354464 58072 354476
rect 46532 354436 58072 354464
rect 46532 354424 46538 354436
rect 58066 354424 58072 354436
rect 58124 354424 58130 354476
rect 68002 354424 68008 354476
rect 68060 354464 68066 354476
rect 80146 354464 80152 354476
rect 68060 354436 80152 354464
rect 68060 354424 68066 354436
rect 80146 354424 80152 354436
rect 80204 354424 80210 354476
rect 39298 354356 39304 354408
rect 39356 354396 39362 354408
rect 49694 354396 49700 354408
rect 39356 354368 49700 354396
rect 39356 354356 39362 354368
rect 49694 354356 49700 354368
rect 49752 354356 49758 354408
rect 50706 354356 50712 354408
rect 50764 354396 50770 354408
rect 62206 354396 62212 354408
rect 50764 354368 62212 354396
rect 50764 354356 50770 354368
rect 62206 354356 62212 354368
rect 62264 354356 62270 354408
rect 64782 354356 64788 354408
rect 64840 354396 64846 354408
rect 79318 354396 79324 354408
rect 64840 354368 79324 354396
rect 64840 354356 64846 354368
rect 79318 354356 79324 354368
rect 79376 354356 79382 354408
rect 46842 354288 46848 354340
rect 46900 354328 46906 354340
rect 58618 354328 58624 354340
rect 46900 354300 58624 354328
rect 46900 354288 46906 354300
rect 58618 354288 58624 354300
rect 58676 354288 58682 354340
rect 62022 354288 62028 354340
rect 62080 354328 62086 354340
rect 78582 354328 78588 354340
rect 62080 354300 78588 354328
rect 62080 354288 62086 354300
rect 78582 354288 78588 354300
rect 78640 354288 78646 354340
rect 25590 354220 25596 354272
rect 25648 354260 25654 354272
rect 29270 354260 29276 354272
rect 25648 354232 29276 354260
rect 25648 354220 25654 354232
rect 29270 354220 29276 354232
rect 29328 354220 29334 354272
rect 45462 354220 45468 354272
rect 45520 354260 45526 354272
rect 57146 354260 57152 354272
rect 45520 354232 57152 354260
rect 45520 354220 45526 354232
rect 57146 354220 57152 354232
rect 57204 354220 57210 354272
rect 59262 354220 59268 354272
rect 59320 354260 59326 354272
rect 77202 354260 77208 354272
rect 59320 354232 77208 354260
rect 59320 354220 59326 354232
rect 77202 354220 77208 354232
rect 77260 354220 77266 354272
rect 34238 354152 34244 354204
rect 34296 354192 34302 354204
rect 39206 354192 39212 354204
rect 34296 354164 39212 354192
rect 34296 354152 34302 354164
rect 39206 354152 39212 354164
rect 39264 354152 39270 354204
rect 42702 354152 42708 354204
rect 42760 354192 42766 354204
rect 55122 354192 55128 354204
rect 42760 354164 55128 354192
rect 42760 354152 42766 354164
rect 55122 354152 55128 354164
rect 55180 354152 55186 354204
rect 56502 354152 56508 354204
rect 56560 354192 56566 354204
rect 76006 354192 76012 354204
rect 56560 354164 76012 354192
rect 56560 354152 56566 354164
rect 76006 354152 76012 354164
rect 76064 354152 76070 354204
rect 37826 354084 37832 354136
rect 37884 354124 37890 354136
rect 42794 354124 42800 354136
rect 37884 354096 42800 354124
rect 37884 354084 37890 354096
rect 42794 354084 42800 354096
rect 42852 354084 42858 354136
rect 47854 354084 47860 354136
rect 47912 354124 47918 354136
rect 59354 354124 59360 354136
rect 47912 354096 59360 354124
rect 47912 354084 47918 354096
rect 59354 354084 59360 354096
rect 59412 354084 59418 354136
rect 64414 354084 64420 354136
rect 64472 354124 64478 354136
rect 87414 354124 87420 354136
rect 64472 354096 87420 354124
rect 64472 354084 64478 354096
rect 87414 354084 87420 354096
rect 87472 354084 87478 354136
rect 34974 354016 34980 354068
rect 35032 354056 35038 354068
rect 40034 354056 40040 354068
rect 35032 354028 40040 354056
rect 35032 354016 35038 354028
rect 40034 354016 40040 354028
rect 40092 354016 40098 354068
rect 44082 354016 44088 354068
rect 44140 354056 44146 354068
rect 57238 354056 57244 354068
rect 44140 354028 57244 354056
rect 44140 354016 44146 354028
rect 57238 354016 57244 354028
rect 57296 354016 57302 354068
rect 67266 354016 67272 354068
rect 67324 354056 67330 354068
rect 91830 354056 91836 354068
rect 67324 354028 91836 354056
rect 67324 354016 67330 354028
rect 91830 354016 91836 354028
rect 91888 354016 91894 354068
rect 26142 353948 26148 354000
rect 26200 353988 26206 354000
rect 30374 353988 30380 354000
rect 26200 353960 30380 353988
rect 26200 353948 26206 353960
rect 30374 353948 30380 353960
rect 30432 353948 30438 354000
rect 31662 353948 31668 354000
rect 31720 353988 31726 354000
rect 36722 353988 36728 354000
rect 31720 353960 36728 353988
rect 31720 353948 31726 353960
rect 36722 353948 36728 353960
rect 36780 353948 36786 354000
rect 38378 353948 38384 354000
rect 38436 353988 38442 354000
rect 48590 353988 48596 354000
rect 38436 353960 48596 353988
rect 38436 353948 38442 353960
rect 48590 353948 48596 353960
rect 48648 353948 48654 354000
rect 49326 353948 49332 354000
rect 49384 353988 49390 354000
rect 64966 353988 64972 354000
rect 49384 353960 64972 353988
rect 49384 353948 49390 353960
rect 64966 353948 64972 353960
rect 65024 353948 65030 354000
rect 70118 353948 70124 354000
rect 70176 353988 70182 354000
rect 96062 353988 96068 354000
rect 70176 353960 96068 353988
rect 70176 353948 70182 353960
rect 96062 353948 96068 353960
rect 96120 353948 96126 354000
rect 50062 353880 50068 353932
rect 50120 353920 50126 353932
rect 62114 353920 62120 353932
rect 50120 353892 62120 353920
rect 50120 353880 50126 353892
rect 62114 353880 62120 353892
rect 62172 353880 62178 353932
rect 32766 353812 32772 353864
rect 32824 353852 32830 353864
rect 37826 353852 37832 353864
rect 32824 353824 37832 353852
rect 32824 353812 32830 353824
rect 37826 353812 37832 353824
rect 37884 353812 37890 353864
rect 55766 353812 55772 353864
rect 55824 353852 55830 353864
rect 67542 353852 67548 353864
rect 55824 353824 67548 353852
rect 55824 353812 55830 353824
rect 67542 353812 67548 353824
rect 67600 353812 67606 353864
rect 29914 353744 29920 353796
rect 29972 353784 29978 353796
rect 35802 353784 35808 353796
rect 29972 353756 35808 353784
rect 29972 353744 29978 353756
rect 35802 353744 35808 353756
rect 35860 353744 35866 353796
rect 41322 353744 41328 353796
rect 41380 353784 41386 353796
rect 53006 353784 53012 353796
rect 41380 353756 53012 353784
rect 41380 353744 41386 353756
rect 53006 353744 53012 353756
rect 53064 353744 53070 353796
rect 54294 353744 54300 353796
rect 54352 353784 54358 353796
rect 63494 353784 63500 353796
rect 54352 353756 63500 353784
rect 54352 353744 54358 353756
rect 63494 353744 63500 353756
rect 63552 353744 63558 353796
rect 30282 353676 30288 353728
rect 30340 353716 30346 353728
rect 34514 353716 34520 353728
rect 30340 353688 34520 353716
rect 30340 353676 30346 353688
rect 34514 353676 34520 353688
rect 34572 353676 34578 353728
rect 42150 353676 42156 353728
rect 42208 353716 42214 353728
rect 54110 353716 54116 353728
rect 42208 353688 54116 353716
rect 42208 353676 42214 353688
rect 54110 353676 54116 353688
rect 54168 353676 54174 353728
rect 40678 353608 40684 353660
rect 40736 353648 40742 353660
rect 51902 353648 51908 353660
rect 40736 353620 51908 353648
rect 40736 353608 40742 353620
rect 51902 353608 51908 353620
rect 51960 353608 51966 353660
rect 27062 353540 27068 353592
rect 27120 353580 27126 353592
rect 31846 353580 31852 353592
rect 27120 353552 31852 353580
rect 27120 353540 27126 353552
rect 31846 353540 31852 353552
rect 31904 353540 31910 353592
rect 37090 353540 37096 353592
rect 37148 353580 37154 353592
rect 42242 353580 42248 353592
rect 37148 353552 42248 353580
rect 37148 353540 37154 353552
rect 42242 353540 42248 353552
rect 42300 353540 42306 353592
rect 43530 353540 43536 353592
rect 43588 353580 43594 353592
rect 56134 353580 56140 353592
rect 43588 353552 56140 353580
rect 43588 353540 43594 353552
rect 56134 353540 56140 353552
rect 56192 353540 56198 353592
rect 24762 353472 24768 353524
rect 24820 353512 24826 353524
rect 28166 353512 28172 353524
rect 24820 353484 28172 353512
rect 24820 353472 24826 353484
rect 28166 353472 28172 353484
rect 28224 353472 28230 353524
rect 28902 353472 28908 353524
rect 28960 353512 28966 353524
rect 34422 353512 34428 353524
rect 28960 353484 34428 353512
rect 28960 353472 28966 353484
rect 34422 353472 34428 353484
rect 34480 353472 34486 353524
rect 22002 353404 22008 353456
rect 22060 353444 22066 353456
rect 23934 353444 23940 353456
rect 22060 353416 23940 353444
rect 22060 353404 22066 353416
rect 23934 353404 23940 353416
rect 23992 353404 23998 353456
rect 24210 353404 24216 353456
rect 24268 353444 24274 353456
rect 27062 353444 27068 353456
rect 24268 353416 27068 353444
rect 24268 353404 24274 353416
rect 27062 353404 27068 353416
rect 27120 353404 27126 353456
rect 31386 353404 31392 353456
rect 31444 353444 31450 353456
rect 37090 353444 37096 353456
rect 31444 353416 37096 353444
rect 31444 353404 31450 353416
rect 37090 353404 37096 353416
rect 37148 353404 37154 353456
rect 21266 353336 21272 353388
rect 21324 353376 21330 353388
rect 22830 353376 22836 353388
rect 21324 353348 22836 353376
rect 21324 353336 21330 353348
rect 22830 353336 22836 353348
rect 22888 353336 22894 353388
rect 23382 353336 23388 353388
rect 23440 353376 23446 353388
rect 26234 353376 26240 353388
rect 23440 353348 26240 353376
rect 23440 353336 23446 353348
rect 26234 353336 26240 353348
rect 26292 353336 26298 353388
rect 28442 353336 28448 353388
rect 28500 353376 28506 353388
rect 33502 353376 33508 353388
rect 28500 353348 33508 353376
rect 28500 353336 28506 353348
rect 33502 353336 33508 353348
rect 33560 353336 33566 353388
rect 20622 353268 20628 353320
rect 20680 353308 20686 353320
rect 22186 353308 22192 353320
rect 20680 353280 22192 353308
rect 20680 353268 20686 353280
rect 22186 353268 22192 353280
rect 22244 353268 22250 353320
rect 22738 353268 22744 353320
rect 22796 353308 22802 353320
rect 25038 353308 25044 353320
rect 22796 353280 25044 353308
rect 22796 353268 22802 353280
rect 25038 353268 25044 353280
rect 25096 353268 25102 353320
rect 27522 353268 27528 353320
rect 27580 353308 27586 353320
rect 32582 353308 32588 353320
rect 27580 353280 32588 353308
rect 27580 353268 27586 353280
rect 32582 353268 32588 353280
rect 32640 353268 32646 353320
rect 36354 353268 36360 353320
rect 36412 353308 36418 353320
rect 41414 353308 41420 353320
rect 36412 353280 41420 353308
rect 36412 353268 36418 353280
rect 41414 353268 41420 353280
rect 41472 353268 41478 353320
rect 63494 353132 63500 353184
rect 63552 353172 63558 353184
rect 72326 353172 72332 353184
rect 63552 353144 72332 353172
rect 63552 353132 63558 353144
rect 72326 353132 72332 353144
rect 72384 353132 72390 353184
rect 67542 353064 67548 353116
rect 67600 353104 67606 353116
rect 74718 353104 74724 353116
rect 67600 353076 74724 353104
rect 67600 353064 67606 353076
rect 74718 353064 74724 353076
rect 74776 353064 74782 353116
rect 68922 352996 68928 353048
rect 68980 353036 68986 353048
rect 78766 353036 78772 353048
rect 68980 353008 78772 353036
rect 68980 352996 68986 353008
rect 78766 352996 78772 353008
rect 78824 352996 78830 353048
rect 70394 352928 70400 352980
rect 70452 352968 70458 352980
rect 83182 352968 83188 352980
rect 70452 352940 83188 352968
rect 70452 352928 70458 352940
rect 83182 352928 83188 352940
rect 83240 352928 83246 352980
rect 57054 352860 57060 352912
rect 57112 352900 57118 352912
rect 76742 352900 76748 352912
rect 57112 352872 76748 352900
rect 57112 352860 57118 352872
rect 76742 352860 76748 352872
rect 76800 352860 76806 352912
rect 60090 352792 60096 352844
rect 60148 352832 60154 352844
rect 80974 352832 80980 352844
rect 60148 352804 80980 352832
rect 60148 352792 60154 352804
rect 80974 352792 80980 352804
rect 81032 352792 81038 352844
rect 62942 352724 62948 352776
rect 63000 352764 63006 352776
rect 85574 352764 85580 352776
rect 63000 352736 85580 352764
rect 63000 352724 63006 352736
rect 85574 352724 85580 352736
rect 85632 352724 85638 352776
rect 65794 352656 65800 352708
rect 65852 352696 65858 352708
rect 89714 352696 89720 352708
rect 65852 352668 89720 352696
rect 65852 352656 65858 352668
rect 89714 352656 89720 352668
rect 89772 352656 89778 352708
rect 68738 352588 68744 352640
rect 68796 352628 68802 352640
rect 94038 352628 94044 352640
rect 68796 352600 94044 352628
rect 68796 352588 68802 352600
rect 94038 352588 94044 352600
rect 94096 352588 94102 352640
rect 52914 352520 52920 352572
rect 52972 352560 52978 352572
rect 70394 352560 70400 352572
rect 52972 352532 70400 352560
rect 52972 352520 52978 352532
rect 70394 352520 70400 352532
rect 70452 352520 70458 352572
rect 71590 352520 71596 352572
rect 71648 352560 71654 352572
rect 98270 352560 98276 352572
rect 71648 352532 98276 352560
rect 71648 352520 71654 352532
rect 98270 352520 98276 352532
rect 98328 352520 98334 352572
rect 58066 351840 58072 351892
rect 58124 351880 58130 351892
rect 60734 351880 60740 351892
rect 58124 351852 60740 351880
rect 58124 351840 58130 351852
rect 60734 351840 60740 351852
rect 60792 351840 60798 351892
rect 77846 351880 77852 351892
rect 60844 351852 77852 351880
rect 36722 351772 36728 351824
rect 36780 351812 36786 351824
rect 39022 351812 39028 351824
rect 36780 351784 39028 351812
rect 36780 351772 36786 351784
rect 39022 351772 39028 351784
rect 39080 351772 39086 351824
rect 57790 351704 57796 351756
rect 57848 351744 57854 351756
rect 60844 351744 60872 351852
rect 77846 351840 77852 351852
rect 77904 351840 77910 351892
rect 80054 351840 80060 351892
rect 80112 351880 80118 351892
rect 97166 351880 97172 351892
rect 80112 351852 97172 351880
rect 80112 351840 80118 351852
rect 97166 351840 97172 351852
rect 97224 351840 97230 351892
rect 138842 351840 138848 351892
rect 138900 351880 138906 351892
rect 139302 351880 139308 351892
rect 138900 351852 139308 351880
rect 138900 351840 138906 351852
rect 139302 351840 139308 351852
rect 139360 351840 139366 351892
rect 139762 351840 139768 351892
rect 139820 351880 139826 351892
rect 140590 351880 140596 351892
rect 139820 351852 140596 351880
rect 139820 351840 139826 351852
rect 140590 351840 140596 351852
rect 140648 351840 140654 351892
rect 142982 351840 142988 351892
rect 143040 351880 143046 351892
rect 143442 351880 143448 351892
rect 143040 351852 143448 351880
rect 143040 351840 143046 351852
rect 143442 351840 143448 351852
rect 143500 351840 143506 351892
rect 144178 351840 144184 351892
rect 144236 351880 144242 351892
rect 144822 351880 144828 351892
rect 144236 351852 144828 351880
rect 144236 351840 144242 351852
rect 144822 351840 144828 351852
rect 144880 351840 144886 351892
rect 145282 351840 145288 351892
rect 145340 351880 145346 351892
rect 146110 351880 146116 351892
rect 145340 351852 146116 351880
rect 145340 351840 145346 351852
rect 146110 351840 146116 351852
rect 146168 351840 146174 351892
rect 155954 351840 155960 351892
rect 156012 351880 156018 351892
rect 156414 351880 156420 351892
rect 156012 351852 156420 351880
rect 156012 351840 156018 351852
rect 156414 351840 156420 351852
rect 156472 351840 156478 351892
rect 158806 351840 158812 351892
rect 158864 351880 158870 351892
rect 159726 351880 159732 351892
rect 158864 351852 159732 351880
rect 158864 351840 158870 351852
rect 159726 351840 159732 351852
rect 159784 351840 159790 351892
rect 160094 351840 160100 351892
rect 160152 351880 160158 351892
rect 160830 351880 160836 351892
rect 160152 351852 160836 351880
rect 160152 351840 160158 351852
rect 160830 351840 160836 351852
rect 160888 351840 160894 351892
rect 161474 351840 161480 351892
rect 161532 351880 161538 351892
rect 161934 351880 161940 351892
rect 161532 351852 161940 351880
rect 161532 351840 161538 351852
rect 161934 351840 161940 351852
rect 161992 351840 161998 351892
rect 164234 351840 164240 351892
rect 164292 351880 164298 351892
rect 165062 351880 165068 351892
rect 164292 351852 165068 351880
rect 164292 351840 164298 351852
rect 165062 351840 165068 351852
rect 165120 351840 165126 351892
rect 165614 351840 165620 351892
rect 165672 351880 165678 351892
rect 166166 351880 166172 351892
rect 165672 351852 166172 351880
rect 165672 351840 165678 351852
rect 166166 351840 166172 351852
rect 166224 351840 166230 351892
rect 187510 351840 187516 351892
rect 187568 351880 187574 351892
rect 194134 351880 194140 351892
rect 187568 351852 194140 351880
rect 187568 351840 187574 351852
rect 194134 351840 194140 351852
rect 194192 351840 194198 351892
rect 198918 351840 198924 351892
rect 198976 351880 198982 351892
rect 200574 351880 200580 351892
rect 198976 351852 200580 351880
rect 198976 351840 198982 351852
rect 200574 351840 200580 351852
rect 200632 351840 200638 351892
rect 275738 351840 275744 351892
rect 275796 351880 275802 351892
rect 277394 351880 277400 351892
rect 275796 351852 277400 351880
rect 275796 351840 275802 351852
rect 277394 351840 277400 351852
rect 277452 351840 277458 351892
rect 82078 351812 82084 351824
rect 57848 351716 60872 351744
rect 60936 351784 82084 351812
rect 57848 351704 57854 351716
rect 60642 351636 60648 351688
rect 60700 351676 60706 351688
rect 60936 351676 60964 351784
rect 82078 351772 82084 351784
rect 82136 351772 82142 351824
rect 63402 351704 63408 351756
rect 63460 351744 63466 351756
rect 86310 351744 86316 351756
rect 63460 351716 86316 351744
rect 63460 351704 63466 351716
rect 86310 351704 86316 351716
rect 86368 351704 86374 351756
rect 60700 351648 60964 351676
rect 60700 351636 60706 351648
rect 66162 351636 66168 351688
rect 66220 351676 66226 351688
rect 90726 351676 90732 351688
rect 66220 351648 90732 351676
rect 66220 351636 66226 351648
rect 90726 351636 90732 351648
rect 90784 351636 90790 351688
rect 38654 351568 38660 351620
rect 38712 351608 38718 351620
rect 41506 351608 41512 351620
rect 38712 351580 41512 351608
rect 38712 351568 38718 351580
rect 41506 351568 41512 351580
rect 41564 351568 41570 351620
rect 59630 351568 59636 351620
rect 59688 351608 59694 351620
rect 63678 351608 63684 351620
rect 59688 351580 63684 351608
rect 59688 351568 59694 351580
rect 63678 351568 63684 351580
rect 63736 351568 63742 351620
rect 63770 351568 63776 351620
rect 63828 351608 63834 351620
rect 66990 351608 66996 351620
rect 63828 351580 66996 351608
rect 63828 351568 63834 351580
rect 66990 351568 66996 351580
rect 67048 351568 67054 351620
rect 69382 351568 69388 351620
rect 69440 351608 69446 351620
rect 95234 351608 95240 351620
rect 69440 351580 95240 351608
rect 69440 351568 69446 351580
rect 95234 351568 95240 351580
rect 95292 351568 95298 351620
rect 127986 351568 127992 351620
rect 128044 351608 128050 351620
rect 128044 351580 129964 351608
rect 128044 351568 128050 351580
rect 34514 351500 34520 351552
rect 34572 351540 34578 351552
rect 36814 351540 36820 351552
rect 34572 351512 36820 351540
rect 34572 351500 34578 351512
rect 36814 351500 36820 351512
rect 36872 351500 36878 351552
rect 37826 351500 37832 351552
rect 37884 351540 37890 351552
rect 40126 351540 40132 351552
rect 37884 351512 40132 351540
rect 37884 351500 37890 351512
rect 40126 351500 40132 351512
rect 40184 351500 40190 351552
rect 73706 351500 73712 351552
rect 73764 351540 73770 351552
rect 101398 351540 101404 351552
rect 73764 351512 101404 351540
rect 73764 351500 73770 351512
rect 101398 351500 101404 351512
rect 101456 351500 101462 351552
rect 123754 351500 123760 351552
rect 123812 351540 123818 351552
rect 123812 351512 129872 351540
rect 123812 351500 123818 351512
rect 40310 351432 40316 351484
rect 40368 351472 40374 351484
rect 44358 351472 44364 351484
rect 40368 351444 44364 351472
rect 40368 351432 40374 351444
rect 44358 351432 44364 351444
rect 44416 351432 44422 351484
rect 56962 351432 56968 351484
rect 57020 351472 57026 351484
rect 58342 351472 58348 351484
rect 57020 351444 58348 351472
rect 57020 351432 57026 351444
rect 58342 351432 58348 351444
rect 58400 351432 58406 351484
rect 59354 351432 59360 351484
rect 59412 351472 59418 351484
rect 62758 351472 62764 351484
rect 59412 351444 62764 351472
rect 59412 351432 59418 351444
rect 62758 351432 62764 351444
rect 62816 351432 62822 351484
rect 63586 351432 63592 351484
rect 63644 351472 63650 351484
rect 68094 351472 68100 351484
rect 63644 351444 68100 351472
rect 63644 351432 63650 351444
rect 68094 351432 68100 351444
rect 68152 351432 68158 351484
rect 72234 351432 72240 351484
rect 72292 351472 72298 351484
rect 99374 351472 99380 351484
rect 72292 351444 99380 351472
rect 72292 351432 72298 351444
rect 99374 351432 99380 351444
rect 99432 351432 99438 351484
rect 129090 351432 129096 351484
rect 129148 351472 129154 351484
rect 129642 351472 129648 351484
rect 129148 351444 129648 351472
rect 129148 351432 129154 351444
rect 129642 351432 129648 351444
rect 129700 351432 129706 351484
rect 41414 351364 41420 351416
rect 41472 351404 41478 351416
rect 43438 351404 43444 351416
rect 41472 351376 43444 351404
rect 41472 351364 41478 351376
rect 43438 351364 43444 351376
rect 43496 351364 43502 351416
rect 58618 351364 58624 351416
rect 58676 351404 58682 351416
rect 61654 351404 61660 351416
rect 58676 351376 61660 351404
rect 58676 351364 58682 351376
rect 61654 351364 61660 351376
rect 61712 351364 61718 351416
rect 62206 351364 62212 351416
rect 62264 351404 62270 351416
rect 63770 351404 63776 351416
rect 62264 351376 63776 351404
rect 62264 351364 62270 351376
rect 63770 351364 63776 351376
rect 63828 351364 63834 351416
rect 75178 351364 75184 351416
rect 75236 351404 75242 351416
rect 103698 351404 103704 351416
rect 75236 351376 103704 351404
rect 75236 351364 75242 351376
rect 103698 351364 103704 351376
rect 103756 351364 103762 351416
rect 129844 351404 129872 351512
rect 129936 351472 129964 351580
rect 133322 351568 133328 351620
rect 133380 351608 133386 351620
rect 133782 351608 133788 351620
rect 133380 351580 133788 351608
rect 133380 351568 133386 351580
rect 133782 351568 133788 351580
rect 133840 351568 133846 351620
rect 135530 351568 135536 351620
rect 135588 351608 135594 351620
rect 136450 351608 136456 351620
rect 135588 351580 136456 351608
rect 135588 351568 135594 351580
rect 136450 351568 136456 351580
rect 136508 351568 136514 351620
rect 130194 351500 130200 351552
rect 130252 351540 130258 351552
rect 154758 351540 154764 351552
rect 130252 351512 154764 351540
rect 130252 351500 130258 351512
rect 154758 351500 154764 351512
rect 154816 351500 154822 351552
rect 271322 351500 271328 351552
rect 271380 351540 271386 351552
rect 273254 351540 273260 351552
rect 271380 351512 273260 351540
rect 271380 351500 271386 351512
rect 273254 351500 273260 351512
rect 273312 351500 273318 351552
rect 154850 351472 154856 351484
rect 129936 351444 154856 351472
rect 154850 351432 154856 351444
rect 154908 351432 154914 351484
rect 169938 351432 169944 351484
rect 169996 351472 170002 351484
rect 170398 351472 170404 351484
rect 169996 351444 170404 351472
rect 169996 351432 170002 351444
rect 170398 351432 170404 351444
rect 170456 351432 170462 351484
rect 171134 351432 171140 351484
rect 171192 351472 171198 351484
rect 171594 351472 171600 351484
rect 171192 351444 171600 351472
rect 171192 351432 171198 351444
rect 171594 351432 171600 351444
rect 171652 351432 171658 351484
rect 175274 351432 175280 351484
rect 175332 351472 175338 351484
rect 175918 351472 175924 351484
rect 175332 351444 175924 351472
rect 175332 351432 175338 351444
rect 175918 351432 175924 351444
rect 175976 351432 175982 351484
rect 176654 351432 176660 351484
rect 176712 351472 176718 351484
rect 177114 351472 177120 351484
rect 176712 351444 177120 351472
rect 176712 351432 176718 351444
rect 177114 351432 177120 351444
rect 177172 351432 177178 351484
rect 179506 351432 179512 351484
rect 179564 351472 179570 351484
rect 180150 351472 180156 351484
rect 179564 351444 180156 351472
rect 179564 351432 179570 351444
rect 180150 351432 180156 351444
rect 180208 351432 180214 351484
rect 180794 351432 180800 351484
rect 180852 351472 180858 351484
rect 181254 351472 181260 351484
rect 180852 351444 181260 351472
rect 180852 351432 180858 351444
rect 181254 351432 181260 351444
rect 181312 351432 181318 351484
rect 184934 351432 184940 351484
rect 184992 351472 184998 351484
rect 185486 351472 185492 351484
rect 184992 351444 185492 351472
rect 184992 351432 184998 351444
rect 185486 351432 185492 351444
rect 185544 351432 185550 351484
rect 194962 351432 194968 351484
rect 195020 351472 195026 351484
rect 198734 351472 198740 351484
rect 195020 351444 198740 351472
rect 195020 351432 195026 351444
rect 198734 351432 198740 351444
rect 198792 351432 198798 351484
rect 269022 351432 269028 351484
rect 269080 351472 269086 351484
rect 270494 351472 270500 351484
rect 269080 351444 270500 351472
rect 269080 351432 269086 351444
rect 270494 351432 270500 351444
rect 270552 351432 270558 351484
rect 273070 351432 273076 351484
rect 273128 351472 273134 351484
rect 274634 351472 274640 351484
rect 273128 351444 274640 351472
rect 273128 351432 273134 351444
rect 274634 351432 274640 351444
rect 274692 351432 274698 351484
rect 278682 351432 278688 351484
rect 278740 351472 278746 351484
rect 281442 351472 281448 351484
rect 278740 351444 281448 351472
rect 278740 351432 278746 351444
rect 281442 351432 281448 351444
rect 281500 351432 281506 351484
rect 154942 351404 154948 351416
rect 129844 351376 154948 351404
rect 154942 351364 154948 351376
rect 155000 351364 155006 351416
rect 270218 351364 270224 351416
rect 270276 351404 270282 351416
rect 271874 351404 271880 351416
rect 270276 351376 271880 351404
rect 270276 351364 270282 351376
rect 271874 351364 271880 351376
rect 271932 351364 271938 351416
rect 274542 351364 274548 351416
rect 274600 351404 274606 351416
rect 276198 351404 276204 351416
rect 274600 351376 276204 351404
rect 274600 351364 274606 351376
rect 276198 351364 276204 351376
rect 276256 351364 276262 351416
rect 277762 351364 277768 351416
rect 277820 351404 277826 351416
rect 280154 351404 280160 351416
rect 277820 351376 280160 351404
rect 277820 351364 277826 351376
rect 280154 351364 280160 351376
rect 280212 351364 280218 351416
rect 42794 351296 42800 351348
rect 42852 351336 42858 351348
rect 47670 351336 47676 351348
rect 42852 351308 47676 351336
rect 42852 351296 42858 351308
rect 47670 351296 47676 351308
rect 47728 351296 47734 351348
rect 52178 351296 52184 351348
rect 52236 351336 52242 351348
rect 69198 351336 69204 351348
rect 52236 351308 69204 351336
rect 52236 351296 52242 351308
rect 69198 351296 69204 351308
rect 69256 351296 69262 351348
rect 72970 351296 72976 351348
rect 73028 351336 73034 351348
rect 100846 351336 100852 351348
rect 73028 351308 100852 351336
rect 73028 351296 73034 351308
rect 100846 351296 100852 351308
rect 100904 351296 100910 351348
rect 121362 351296 121368 351348
rect 121420 351336 121426 351348
rect 153286 351336 153292 351348
rect 121420 351308 153292 351336
rect 121420 351296 121426 351308
rect 153286 351296 153292 351308
rect 153344 351296 153350 351348
rect 276658 351296 276664 351348
rect 276716 351336 276722 351348
rect 278774 351336 278780 351348
rect 276716 351308 278780 351336
rect 276716 351296 276722 351308
rect 278774 351296 278780 351308
rect 278832 351296 278838 351348
rect 40034 351228 40040 351280
rect 40092 351268 40098 351280
rect 43254 351268 43260 351280
rect 40092 351240 43260 351268
rect 40092 351228 40098 351240
rect 43254 351228 43260 351240
rect 43312 351228 43318 351280
rect 46566 351268 46572 351280
rect 43364 351240 46572 351268
rect 39206 351160 39212 351212
rect 39264 351200 39270 351212
rect 42150 351200 42156 351212
rect 39264 351172 42156 351200
rect 39264 351160 39270 351172
rect 42150 351160 42156 351172
rect 42208 351160 42214 351212
rect 42242 351160 42248 351212
rect 42300 351200 42306 351212
rect 43364 351200 43392 351240
rect 46566 351228 46572 351240
rect 46624 351228 46630 351280
rect 53650 351228 53656 351280
rect 53708 351268 53714 351280
rect 71222 351268 71228 351280
rect 53708 351240 71228 351268
rect 53708 351228 53714 351240
rect 71222 351228 71228 351240
rect 71280 351228 71286 351280
rect 74442 351228 74448 351280
rect 74500 351268 74506 351280
rect 102502 351268 102508 351280
rect 74500 351240 102508 351268
rect 74500 351228 74506 351240
rect 102502 351228 102508 351240
rect 102560 351228 102566 351280
rect 120442 351228 120448 351280
rect 120500 351268 120506 351280
rect 153378 351268 153384 351280
rect 120500 351240 153384 351268
rect 120500 351228 120506 351240
rect 153378 351228 153384 351240
rect 153436 351228 153442 351280
rect 42300 351172 43392 351200
rect 42300 351160 42306 351172
rect 43438 351160 43444 351212
rect 43496 351200 43502 351212
rect 45646 351200 45652 351212
rect 43496 351172 45652 351200
rect 43496 351160 43502 351172
rect 45646 351160 45652 351172
rect 45704 351160 45710 351212
rect 55030 351160 55036 351212
rect 55088 351200 55094 351212
rect 73430 351200 73436 351212
rect 55088 351172 73436 351200
rect 55088 351160 55094 351172
rect 73430 351160 73436 351172
rect 73488 351160 73494 351212
rect 75822 351160 75828 351212
rect 75880 351200 75886 351212
rect 104894 351200 104900 351212
rect 75880 351172 104900 351200
rect 75880 351160 75886 351172
rect 104894 351160 104900 351172
rect 104952 351160 104958 351212
rect 119338 351160 119344 351212
rect 119396 351200 119402 351212
rect 153470 351200 153476 351212
rect 119396 351172 153476 351200
rect 119396 351160 119402 351172
rect 153470 351160 153476 351172
rect 153528 351160 153534 351212
rect 193214 351160 193220 351212
rect 193272 351200 193278 351212
rect 195238 351200 195244 351212
rect 193272 351172 195244 351200
rect 193272 351160 193278 351172
rect 195238 351160 195244 351172
rect 195296 351160 195302 351212
rect 228174 351160 228180 351212
rect 228232 351200 228238 351212
rect 229830 351200 229836 351212
rect 228232 351172 229836 351200
rect 228232 351160 228238 351172
rect 229830 351160 229836 351172
rect 229888 351160 229894 351212
rect 57146 351092 57152 351144
rect 57204 351132 57210 351144
rect 59446 351132 59452 351144
rect 57204 351104 59452 351132
rect 57204 351092 57210 351104
rect 59446 351092 59452 351104
rect 59504 351092 59510 351144
rect 77202 351092 77208 351144
rect 77260 351132 77266 351144
rect 80054 351132 80060 351144
rect 77260 351104 80060 351132
rect 77260 351092 77266 351104
rect 80054 351092 80060 351104
rect 80112 351092 80118 351144
rect 80146 351092 80152 351144
rect 80204 351132 80210 351144
rect 92934 351132 92940 351144
rect 80204 351104 92940 351132
rect 80204 351092 80210 351104
rect 92934 351092 92940 351104
rect 92992 351092 92998 351144
rect 62114 351024 62120 351076
rect 62172 351064 62178 351076
rect 66346 351064 66352 351076
rect 62172 351036 66352 351064
rect 62172 351024 62178 351036
rect 66346 351024 66352 351036
rect 66404 351024 66410 351076
rect 78582 351024 78588 351076
rect 78640 351064 78646 351076
rect 84378 351064 84384 351076
rect 78640 351036 84384 351064
rect 78640 351024 78646 351036
rect 84378 351024 84384 351036
rect 84436 351024 84442 351076
rect 187602 351024 187608 351076
rect 187660 351064 187666 351076
rect 193214 351064 193220 351076
rect 187660 351036 193220 351064
rect 187660 351024 187666 351036
rect 193214 351024 193220 351036
rect 193272 351024 193278 351076
rect 79318 350956 79324 351008
rect 79376 350996 79382 351008
rect 88518 350996 88524 351008
rect 79376 350968 88524 350996
rect 79376 350956 79382 350968
rect 88518 350956 88524 350968
rect 88576 350956 88582 351008
rect 173894 350956 173900 351008
rect 173952 350996 173958 351008
rect 174814 350996 174820 351008
rect 173952 350968 174820 350996
rect 173952 350956 173958 350968
rect 174814 350956 174820 350968
rect 174872 350956 174878 351008
rect 124674 350888 124680 350940
rect 124732 350928 124738 350940
rect 125502 350928 125508 350940
rect 124732 350900 125508 350928
rect 124732 350888 124738 350900
rect 125502 350888 125508 350900
rect 125560 350888 125566 350940
rect 134426 350888 134432 350940
rect 134484 350928 134490 350940
rect 135162 350928 135168 350940
rect 134484 350900 135168 350928
rect 134484 350888 134490 350900
rect 135162 350888 135168 350900
rect 135220 350888 135226 350940
rect 183646 350888 183652 350940
rect 183704 350928 183710 350940
rect 184566 350928 184572 350940
rect 183704 350900 184572 350928
rect 183704 350888 183710 350900
rect 184566 350888 184572 350900
rect 184624 350888 184630 350940
rect 201494 350888 201500 350940
rect 201552 350928 201558 350940
rect 202874 350928 202880 350940
rect 201552 350900 202880 350928
rect 201552 350888 201558 350900
rect 202874 350888 202880 350900
rect 202932 350888 202938 350940
rect 226978 350888 226984 350940
rect 227036 350928 227042 350940
rect 228726 350928 228732 350940
rect 227036 350900 228732 350928
rect 227036 350888 227042 350900
rect 228726 350888 228732 350900
rect 228784 350888 228790 350940
rect 230474 350888 230480 350940
rect 230532 350928 230538 350940
rect 231854 350928 231860 350940
rect 230532 350900 231860 350928
rect 230532 350888 230538 350900
rect 231854 350888 231860 350900
rect 231912 350888 231918 350940
rect 233694 350888 233700 350940
rect 233752 350928 233758 350940
rect 235166 350928 235172 350940
rect 233752 350900 235172 350928
rect 233752 350888 233758 350900
rect 235166 350888 235172 350900
rect 235224 350888 235230 350940
rect 272426 350888 272432 350940
rect 272484 350928 272490 350940
rect 274726 350928 274732 350940
rect 272484 350900 274732 350928
rect 272484 350888 272490 350900
rect 274726 350888 274732 350900
rect 274784 350888 274790 350940
rect 37090 350752 37096 350804
rect 37148 350792 37154 350804
rect 37918 350792 37924 350804
rect 37148 350764 37924 350792
rect 37148 350752 37154 350764
rect 37918 350752 37924 350764
rect 37976 350752 37982 350804
rect 222838 350752 222844 350804
rect 222896 350792 222902 350804
rect 224310 350792 224316 350804
rect 222896 350764 224316 350792
rect 222896 350752 222902 350764
rect 224310 350752 224316 350764
rect 224368 350752 224374 350804
rect 115750 350684 115756 350736
rect 115808 350724 115814 350736
rect 149054 350724 149060 350736
rect 115808 350696 149060 350724
rect 115808 350684 115814 350696
rect 149054 350684 149060 350696
rect 149112 350684 149118 350736
rect 112898 350616 112904 350668
rect 112956 350656 112962 350668
rect 146294 350656 146300 350668
rect 112956 350628 146300 350656
rect 112956 350616 112962 350628
rect 146294 350616 146300 350628
rect 146352 350616 146358 350668
rect 106182 350548 106188 350600
rect 106240 350588 106246 350600
rect 153194 350588 153200 350600
rect 106240 350560 153200 350588
rect 106240 350548 106246 350560
rect 153194 350548 153200 350560
rect 153252 350548 153258 350600
rect 3142 336744 3148 336796
rect 3200 336784 3206 336796
rect 6178 336784 6184 336796
rect 3200 336756 6184 336784
rect 3200 336744 3206 336756
rect 6178 336744 6184 336756
rect 6236 336744 6242 336796
rect 303614 327020 303620 327072
rect 303672 327060 303678 327072
rect 417418 327060 417424 327072
rect 303672 327032 417424 327060
rect 303672 327020 303678 327032
rect 417418 327020 417424 327032
rect 417476 327020 417482 327072
rect 303614 325592 303620 325644
rect 303672 325632 303678 325644
rect 563698 325632 563704 325644
rect 303672 325604 563704 325632
rect 303672 325592 303678 325604
rect 563698 325592 563704 325604
rect 563756 325592 563762 325644
rect 21358 323484 21364 323536
rect 21416 323524 21422 323536
rect 22186 323524 22192 323536
rect 21416 323496 22192 323524
rect 21416 323484 21422 323496
rect 22186 323484 22192 323496
rect 22244 323484 22250 323536
rect 22186 321580 22192 321632
rect 22244 321620 22250 321632
rect 22244 321592 23520 321620
rect 22244 321580 22250 321592
rect 23492 321552 23520 321592
rect 303614 321580 303620 321632
rect 303672 321620 303678 321632
rect 580166 321620 580172 321632
rect 303672 321592 580172 321620
rect 303672 321580 303678 321592
rect 580166 321580 580172 321592
rect 580224 321580 580230 321632
rect 26878 321552 26884 321564
rect 23492 321524 26884 321552
rect 26878 321512 26884 321524
rect 26936 321512 26942 321564
rect 100754 321172 100760 321224
rect 100812 321212 100818 321224
rect 106274 321212 106280 321224
rect 100812 321184 106280 321212
rect 100812 321172 100818 321184
rect 106274 321172 106280 321184
rect 106332 321172 106338 321224
rect 111518 321104 111524 321156
rect 111576 321144 111582 321156
rect 117958 321144 117964 321156
rect 111576 321116 117964 321144
rect 111576 321104 111582 321116
rect 117958 321104 117964 321116
rect 118016 321104 118022 321156
rect 231762 321104 231768 321156
rect 231820 321144 231826 321156
rect 235442 321144 235448 321156
rect 231820 321116 235448 321144
rect 231820 321104 231826 321116
rect 235442 321104 235448 321116
rect 235500 321104 235506 321156
rect 92106 321036 92112 321088
rect 92164 321076 92170 321088
rect 96614 321076 96620 321088
rect 92164 321048 96620 321076
rect 92164 321036 92170 321048
rect 96614 321036 96620 321048
rect 96672 321036 96678 321088
rect 108298 321036 108304 321088
rect 108356 321076 108362 321088
rect 115198 321076 115204 321088
rect 108356 321048 115204 321076
rect 108356 321036 108362 321048
rect 115198 321036 115204 321048
rect 115256 321036 115262 321088
rect 228266 321036 228272 321088
rect 228324 321076 228330 321088
rect 232222 321076 232228 321088
rect 228324 321048 232228 321076
rect 228324 321036 228330 321048
rect 232222 321036 232228 321048
rect 232280 321036 232286 321088
rect 101766 320968 101772 321020
rect 101824 321008 101830 321020
rect 106366 321008 106372 321020
rect 101824 320980 106372 321008
rect 101824 320968 101830 320980
rect 106366 320968 106372 320980
rect 106424 320968 106430 321020
rect 109310 320968 109316 321020
rect 109368 321008 109374 321020
rect 119338 321008 119344 321020
rect 109368 320980 119344 321008
rect 109368 320968 109374 320980
rect 119338 320968 119344 320980
rect 119396 320968 119402 321020
rect 75914 320900 75920 320952
rect 75972 320940 75978 320952
rect 78674 320940 78680 320952
rect 75972 320912 78680 320940
rect 75972 320900 75978 320912
rect 78674 320900 78680 320912
rect 78732 320900 78738 320952
rect 93210 320900 93216 320952
rect 93268 320940 93274 320952
rect 97994 320940 98000 320952
rect 93268 320912 98000 320940
rect 93268 320900 93274 320912
rect 97994 320900 98000 320912
rect 98052 320900 98058 320952
rect 102870 320900 102876 320952
rect 102928 320940 102934 320952
rect 108942 320940 108948 320952
rect 102928 320912 108948 320940
rect 102928 320900 102934 320912
rect 108942 320900 108948 320912
rect 109000 320900 109006 320952
rect 115842 320900 115848 320952
rect 115900 320940 115906 320952
rect 126238 320940 126244 320952
rect 115900 320912 126244 320940
rect 115900 320900 115906 320912
rect 126238 320900 126244 320912
rect 126296 320900 126302 320952
rect 24762 320832 24768 320884
rect 24820 320872 24826 320884
rect 26326 320872 26332 320884
rect 24820 320844 26332 320872
rect 24820 320832 24826 320844
rect 26326 320832 26332 320844
rect 26384 320832 26390 320884
rect 34882 320832 34888 320884
rect 34940 320872 34946 320884
rect 35802 320872 35808 320884
rect 34940 320844 35808 320872
rect 34940 320832 34946 320844
rect 35802 320832 35808 320844
rect 35860 320832 35866 320884
rect 54386 320832 54392 320884
rect 54444 320872 54450 320884
rect 55306 320872 55312 320884
rect 54444 320844 55312 320872
rect 54444 320832 54450 320844
rect 55306 320832 55312 320844
rect 55364 320832 55370 320884
rect 64046 320832 64052 320884
rect 64104 320872 64110 320884
rect 64874 320872 64880 320884
rect 64104 320844 64880 320872
rect 64104 320832 64110 320844
rect 64874 320832 64880 320844
rect 64932 320832 64938 320884
rect 72694 320832 72700 320884
rect 72752 320872 72758 320884
rect 74534 320872 74540 320884
rect 72752 320844 74540 320872
rect 72752 320832 72758 320844
rect 74534 320832 74540 320844
rect 74592 320832 74598 320884
rect 82446 320832 82452 320884
rect 82504 320872 82510 320884
rect 85114 320872 85120 320884
rect 82504 320844 85120 320872
rect 82504 320832 82510 320844
rect 85114 320832 85120 320844
rect 85172 320832 85178 320884
rect 85666 320832 85672 320884
rect 85724 320872 85730 320884
rect 89622 320872 89628 320884
rect 85724 320844 89628 320872
rect 85724 320832 85730 320844
rect 89622 320832 89628 320844
rect 89680 320832 89686 320884
rect 106090 320832 106096 320884
rect 106148 320872 106154 320884
rect 121546 320872 121552 320884
rect 106148 320844 121552 320872
rect 106148 320832 106154 320844
rect 121546 320832 121552 320844
rect 121604 320832 121610 320884
rect 198734 320832 198740 320884
rect 198792 320872 198798 320884
rect 202046 320872 202052 320884
rect 198792 320844 202052 320872
rect 198792 320832 198798 320844
rect 202046 320832 202052 320844
rect 202104 320832 202110 320884
rect 247402 320832 247408 320884
rect 247460 320872 247466 320884
rect 249426 320872 249432 320884
rect 247460 320844 249432 320872
rect 247460 320832 247466 320844
rect 249426 320832 249432 320844
rect 249484 320832 249490 320884
rect 73798 320764 73804 320816
rect 73856 320804 73862 320816
rect 75914 320804 75920 320816
rect 73856 320776 75920 320804
rect 73856 320764 73862 320776
rect 75914 320764 75920 320776
rect 75972 320764 75978 320816
rect 110414 320764 110420 320816
rect 110472 320804 110478 320816
rect 113818 320804 113824 320816
rect 110472 320776 113824 320804
rect 110472 320764 110478 320776
rect 113818 320764 113824 320776
rect 113876 320764 113882 320816
rect 146018 320764 146024 320816
rect 146076 320804 146082 320816
rect 152458 320804 152464 320816
rect 146076 320776 152464 320804
rect 146076 320764 146082 320776
rect 152458 320764 152464 320776
rect 152516 320764 152522 320816
rect 227070 320764 227076 320816
rect 227128 320804 227134 320816
rect 231118 320804 231124 320816
rect 227128 320776 231124 320804
rect 227128 320764 227134 320776
rect 231118 320764 231124 320776
rect 231176 320764 231182 320816
rect 246114 320764 246120 320816
rect 246172 320804 246178 320816
rect 248414 320804 248420 320816
rect 246172 320776 248420 320804
rect 246172 320764 246178 320776
rect 248414 320764 248420 320776
rect 248472 320764 248478 320816
rect 256510 320764 256516 320816
rect 256568 320804 256574 320816
rect 258074 320804 258080 320816
rect 256568 320776 258080 320804
rect 256568 320764 256574 320776
rect 258074 320764 258080 320776
rect 258132 320764 258138 320816
rect 83458 320696 83464 320748
rect 83516 320736 83522 320748
rect 85666 320736 85672 320748
rect 83516 320708 85672 320736
rect 83516 320696 83522 320708
rect 85666 320696 85672 320708
rect 85724 320696 85730 320748
rect 248322 320696 248328 320748
rect 248380 320736 248386 320748
rect 250530 320736 250536 320748
rect 248380 320708 250536 320736
rect 248380 320696 248386 320708
rect 250530 320696 250536 320708
rect 250588 320696 250594 320748
rect 226242 320628 226248 320680
rect 226300 320668 226306 320680
rect 230106 320668 230112 320680
rect 226300 320640 230112 320668
rect 226300 320628 226306 320640
rect 230106 320628 230112 320640
rect 230164 320628 230170 320680
rect 98546 320560 98552 320612
rect 98604 320600 98610 320612
rect 103514 320600 103520 320612
rect 98604 320572 103520 320600
rect 98604 320560 98610 320572
rect 103514 320560 103520 320572
rect 103572 320560 103578 320612
rect 204254 320560 204260 320612
rect 204312 320600 204318 320612
rect 206370 320600 206376 320612
rect 204312 320572 206376 320600
rect 204312 320560 204318 320572
rect 206370 320560 206376 320572
rect 206428 320560 206434 320612
rect 208394 320560 208400 320612
rect 208452 320600 208458 320612
rect 210694 320600 210700 320612
rect 208452 320572 210700 320600
rect 208452 320560 208458 320572
rect 210694 320560 210700 320572
rect 210752 320560 210758 320612
rect 202874 320492 202880 320544
rect 202932 320532 202938 320544
rect 205266 320532 205272 320544
rect 202932 320504 205272 320532
rect 202932 320492 202938 320504
rect 205266 320492 205272 320504
rect 205324 320492 205330 320544
rect 23290 320424 23296 320476
rect 23348 320464 23354 320476
rect 25314 320464 25320 320476
rect 23348 320436 25320 320464
rect 23348 320424 23354 320436
rect 25314 320424 25320 320436
rect 25372 320424 25378 320476
rect 91002 320424 91008 320476
rect 91060 320464 91066 320476
rect 95234 320464 95240 320476
rect 91060 320436 95240 320464
rect 91060 320424 91066 320436
rect 95234 320424 95240 320436
rect 95292 320424 95298 320476
rect 99650 320424 99656 320476
rect 99708 320464 99714 320476
rect 104894 320464 104900 320476
rect 99708 320436 104900 320464
rect 99708 320424 99714 320436
rect 104894 320424 104900 320436
rect 104952 320424 104958 320476
rect 195974 320424 195980 320476
rect 196032 320464 196038 320476
rect 198826 320464 198832 320476
rect 196032 320436 198832 320464
rect 196032 320424 196038 320436
rect 198826 320424 198832 320436
rect 198884 320424 198890 320476
rect 235442 320424 235448 320476
rect 235500 320464 235506 320476
rect 238662 320464 238668 320476
rect 235500 320436 238668 320464
rect 235500 320424 235506 320436
rect 238662 320424 238668 320436
rect 238720 320424 238726 320476
rect 78122 320356 78128 320408
rect 78180 320396 78186 320408
rect 81250 320396 81256 320408
rect 78180 320368 81256 320396
rect 78180 320356 78186 320368
rect 81250 320356 81256 320368
rect 81308 320356 81314 320408
rect 88886 320356 88892 320408
rect 88944 320396 88950 320408
rect 92382 320396 92388 320408
rect 88944 320368 92388 320396
rect 88944 320356 88950 320368
rect 92382 320356 92388 320368
rect 92440 320356 92446 320408
rect 94222 320356 94228 320408
rect 94280 320396 94286 320408
rect 99558 320396 99564 320408
rect 94280 320368 99564 320396
rect 94280 320356 94286 320368
rect 99558 320356 99564 320368
rect 99616 320356 99622 320408
rect 236638 320356 236644 320408
rect 236696 320396 236702 320408
rect 239766 320396 239772 320408
rect 236696 320368 239772 320396
rect 236696 320356 236702 320368
rect 239766 320356 239772 320368
rect 239824 320356 239830 320408
rect 25314 320288 25320 320340
rect 25372 320328 25378 320340
rect 27430 320328 27436 320340
rect 25372 320300 27436 320328
rect 25372 320288 25378 320300
rect 27430 320288 27436 320300
rect 27488 320288 27494 320340
rect 66254 320288 66260 320340
rect 66312 320328 66318 320340
rect 67634 320328 67640 320340
rect 66312 320300 67640 320328
rect 66312 320288 66318 320300
rect 67634 320288 67640 320300
rect 67692 320288 67698 320340
rect 71590 320288 71596 320340
rect 71648 320328 71654 320340
rect 73890 320328 73896 320340
rect 71648 320300 73896 320328
rect 71648 320288 71654 320300
rect 73890 320288 73896 320300
rect 73948 320288 73954 320340
rect 80238 320288 80244 320340
rect 80296 320328 80302 320340
rect 82998 320328 83004 320340
rect 80296 320300 83004 320328
rect 80296 320288 80302 320300
rect 82998 320288 83004 320300
rect 83056 320288 83062 320340
rect 86678 320288 86684 320340
rect 86736 320328 86742 320340
rect 91094 320328 91100 320340
rect 86736 320300 91100 320328
rect 86736 320288 86742 320300
rect 91094 320288 91100 320300
rect 91152 320288 91158 320340
rect 97534 320288 97540 320340
rect 97592 320328 97598 320340
rect 102134 320328 102140 320340
rect 97592 320300 102140 320328
rect 97592 320288 97598 320300
rect 102134 320288 102140 320300
rect 102192 320288 102198 320340
rect 103974 320288 103980 320340
rect 104032 320328 104038 320340
rect 109770 320328 109776 320340
rect 104032 320300 109776 320328
rect 104032 320288 104038 320300
rect 109770 320288 109776 320300
rect 109828 320288 109834 320340
rect 184842 320288 184848 320340
rect 184900 320328 184906 320340
rect 186958 320328 186964 320340
rect 184900 320300 186964 320328
rect 184900 320288 184906 320300
rect 186958 320288 186964 320300
rect 187016 320288 187022 320340
rect 198826 320288 198832 320340
rect 198884 320328 198890 320340
rect 200942 320328 200948 320340
rect 198884 320300 200948 320328
rect 198884 320288 198890 320300
rect 200942 320288 200948 320300
rect 201000 320288 201006 320340
rect 229278 320288 229284 320340
rect 229336 320328 229342 320340
rect 233326 320328 233332 320340
rect 229336 320300 233332 320328
rect 229336 320288 229342 320300
rect 233326 320288 233332 320300
rect 233384 320288 233390 320340
rect 238662 320288 238668 320340
rect 238720 320328 238726 320340
rect 241882 320328 241888 320340
rect 238720 320300 241888 320328
rect 238720 320288 238726 320300
rect 241882 320288 241888 320300
rect 241940 320288 241946 320340
rect 242618 320288 242624 320340
rect 242676 320328 242682 320340
rect 245194 320328 245200 320340
rect 242676 320300 245200 320328
rect 242676 320288 242682 320300
rect 245194 320288 245200 320300
rect 245252 320288 245258 320340
rect 253382 320288 253388 320340
rect 253440 320328 253446 320340
rect 254854 320328 254860 320340
rect 253440 320300 254860 320328
rect 253440 320288 253446 320300
rect 254854 320288 254860 320300
rect 254912 320288 254918 320340
rect 27706 320220 27712 320272
rect 27764 320260 27770 320272
rect 29638 320260 29644 320272
rect 27764 320232 29644 320260
rect 27764 320220 27770 320232
rect 29638 320220 29644 320232
rect 29696 320220 29702 320272
rect 30282 320220 30288 320272
rect 30340 320260 30346 320272
rect 31754 320260 31760 320272
rect 30340 320232 31760 320260
rect 30340 320220 30346 320232
rect 31754 320220 31760 320232
rect 31812 320220 31818 320272
rect 33686 320220 33692 320272
rect 33744 320260 33750 320272
rect 34974 320260 34980 320272
rect 33744 320232 34980 320260
rect 33744 320220 33750 320232
rect 34974 320220 34980 320232
rect 35032 320220 35038 320272
rect 61930 320220 61936 320272
rect 61988 320260 61994 320272
rect 63494 320260 63500 320272
rect 61988 320232 63500 320260
rect 61988 320220 61994 320232
rect 63494 320220 63500 320232
rect 63552 320220 63558 320272
rect 68370 320220 68376 320272
rect 68428 320260 68434 320272
rect 70394 320260 70400 320272
rect 68428 320232 70400 320260
rect 68428 320220 68434 320232
rect 70394 320220 70400 320232
rect 70452 320220 70458 320272
rect 70578 320220 70584 320272
rect 70636 320260 70642 320272
rect 73246 320260 73252 320272
rect 70636 320232 73252 320260
rect 70636 320220 70642 320232
rect 73246 320220 73252 320232
rect 73304 320220 73310 320272
rect 77018 320220 77024 320272
rect 77076 320260 77082 320272
rect 79962 320260 79968 320272
rect 77076 320232 79968 320260
rect 77076 320220 77082 320232
rect 79962 320220 79968 320232
rect 80020 320220 80026 320272
rect 81342 320220 81348 320272
rect 81400 320260 81406 320272
rect 82814 320260 82820 320272
rect 81400 320232 82820 320260
rect 81400 320220 81406 320232
rect 82814 320220 82820 320232
rect 82872 320220 82878 320272
rect 89990 320220 89996 320272
rect 90048 320260 90054 320272
rect 92750 320260 92756 320272
rect 90048 320232 92756 320260
rect 90048 320220 90054 320232
rect 92750 320220 92756 320232
rect 92808 320220 92814 320272
rect 96430 320220 96436 320272
rect 96488 320260 96494 320272
rect 100754 320260 100760 320272
rect 96488 320232 100760 320260
rect 96488 320220 96494 320232
rect 100754 320220 100760 320232
rect 100812 320220 100818 320272
rect 105078 320220 105084 320272
rect 105136 320260 105142 320272
rect 110414 320260 110420 320272
rect 105136 320232 110420 320260
rect 105136 320220 105142 320232
rect 110414 320220 110420 320232
rect 110472 320220 110478 320272
rect 163222 320220 163228 320272
rect 163280 320260 163286 320272
rect 167638 320260 167644 320272
rect 163280 320232 167644 320260
rect 163280 320220 163286 320232
rect 167638 320220 167644 320232
rect 167696 320220 167702 320272
rect 181530 320220 181536 320272
rect 181588 320260 181594 320272
rect 184198 320260 184204 320272
rect 181588 320232 184204 320260
rect 181588 320220 181594 320232
rect 184198 320220 184204 320232
rect 184256 320220 184262 320272
rect 192478 320220 192484 320272
rect 192536 320260 192542 320272
rect 196618 320260 196624 320272
rect 192536 320232 196624 320260
rect 192536 320220 192542 320232
rect 196618 320220 196624 320232
rect 196676 320220 196682 320272
rect 202138 320220 202144 320272
rect 202196 320260 202202 320272
rect 204162 320260 204168 320272
rect 202196 320232 204168 320260
rect 202196 320220 202202 320232
rect 204162 320220 204168 320232
rect 204220 320220 204226 320272
rect 233142 320220 233148 320272
rect 233200 320260 233206 320272
rect 236546 320260 236552 320272
rect 233200 320232 236552 320260
rect 233200 320220 233206 320232
rect 236546 320220 236552 320232
rect 236604 320220 236610 320272
rect 237834 320220 237840 320272
rect 237892 320260 237898 320272
rect 240870 320260 240876 320272
rect 237892 320232 240876 320260
rect 237892 320220 237898 320232
rect 240870 320220 240876 320232
rect 240928 320220 240934 320272
rect 241422 320220 241428 320272
rect 241480 320260 241486 320272
rect 244090 320260 244096 320272
rect 241480 320232 244096 320260
rect 241480 320220 241486 320232
rect 244090 320220 244096 320232
rect 244148 320220 244154 320272
rect 245010 320220 245016 320272
rect 245068 320260 245074 320272
rect 247310 320260 247316 320272
rect 245068 320232 247316 320260
rect 245068 320220 245074 320232
rect 247310 320220 247316 320232
rect 247368 320220 247374 320272
rect 251082 320220 251088 320272
rect 251140 320260 251146 320272
rect 252738 320260 252744 320272
rect 251140 320232 252744 320260
rect 251140 320220 251146 320232
rect 252738 320220 252744 320232
rect 252796 320220 252802 320272
rect 254578 320220 254584 320272
rect 254636 320260 254642 320272
rect 255958 320260 255964 320272
rect 254636 320232 255964 320260
rect 254636 320220 254642 320232
rect 255958 320220 255964 320232
rect 256016 320220 256022 320272
rect 257982 320220 257988 320272
rect 258040 320260 258046 320272
rect 259178 320260 259184 320272
rect 258040 320232 259184 320260
rect 258040 320220 258046 320232
rect 259178 320220 259184 320232
rect 259236 320220 259242 320272
rect 22002 320152 22008 320204
rect 22060 320192 22066 320204
rect 24210 320192 24216 320204
rect 22060 320164 24216 320192
rect 22060 320152 22066 320164
rect 24210 320152 24216 320164
rect 24268 320152 24274 320204
rect 26510 320152 26516 320204
rect 26568 320192 26574 320204
rect 28534 320192 28540 320204
rect 26568 320164 28540 320192
rect 26568 320152 26574 320164
rect 28534 320152 28540 320164
rect 28592 320152 28598 320204
rect 28902 320152 28908 320204
rect 28960 320192 28966 320204
rect 30650 320192 30656 320204
rect 28960 320164 30656 320192
rect 28960 320152 28966 320164
rect 30650 320152 30656 320164
rect 30708 320152 30714 320204
rect 31662 320152 31668 320204
rect 31720 320192 31726 320204
rect 32858 320192 32864 320204
rect 31720 320164 32864 320192
rect 31720 320152 31726 320164
rect 32858 320152 32864 320164
rect 32916 320152 32922 320204
rect 33042 320152 33048 320204
rect 33100 320192 33106 320204
rect 33870 320192 33876 320204
rect 33100 320164 33876 320192
rect 33100 320152 33106 320164
rect 33870 320152 33876 320164
rect 33928 320152 33934 320204
rect 35894 320152 35900 320204
rect 35952 320192 35958 320204
rect 37182 320192 37188 320204
rect 35952 320164 37188 320192
rect 35952 320152 35958 320164
rect 37182 320152 37188 320164
rect 37240 320152 37246 320204
rect 37274 320152 37280 320204
rect 37332 320192 37338 320204
rect 38194 320192 38200 320204
rect 37332 320164 38200 320192
rect 37332 320152 37338 320164
rect 38194 320152 38200 320164
rect 38252 320152 38258 320204
rect 38562 320152 38568 320204
rect 38620 320192 38626 320204
rect 39298 320192 39304 320204
rect 38620 320164 39304 320192
rect 38620 320152 38626 320164
rect 39298 320152 39304 320164
rect 39356 320152 39362 320204
rect 42518 320192 42524 320204
rect 41432 320164 42524 320192
rect 41432 320136 41460 320164
rect 42518 320152 42524 320164
rect 42576 320152 42582 320204
rect 42794 320152 42800 320204
rect 42852 320192 42858 320204
rect 43622 320192 43628 320204
rect 42852 320164 43628 320192
rect 42852 320152 42858 320164
rect 43622 320152 43628 320164
rect 43680 320152 43686 320204
rect 46934 320152 46940 320204
rect 46992 320192 46998 320204
rect 47946 320192 47952 320204
rect 46992 320164 47952 320192
rect 46992 320152 46998 320164
rect 47946 320152 47952 320164
rect 48004 320152 48010 320204
rect 59814 320152 59820 320204
rect 59872 320192 59878 320204
rect 60734 320192 60740 320204
rect 59872 320164 60740 320192
rect 59872 320152 59878 320164
rect 60734 320152 60740 320164
rect 60792 320152 60798 320204
rect 60826 320152 60832 320204
rect 60884 320192 60890 320204
rect 62114 320192 62120 320204
rect 60884 320164 62120 320192
rect 60884 320152 60890 320164
rect 62114 320152 62120 320164
rect 62172 320152 62178 320204
rect 63034 320152 63040 320204
rect 63092 320192 63098 320204
rect 64322 320192 64328 320204
rect 63092 320164 64328 320192
rect 63092 320152 63098 320164
rect 64322 320152 64328 320164
rect 64380 320152 64386 320204
rect 65150 320152 65156 320204
rect 65208 320192 65214 320204
rect 66254 320192 66260 320204
rect 65208 320164 66260 320192
rect 65208 320152 65214 320164
rect 66254 320152 66260 320164
rect 66312 320152 66318 320204
rect 67358 320152 67364 320204
rect 67416 320192 67422 320204
rect 69014 320192 69020 320204
rect 67416 320164 69020 320192
rect 67416 320152 67422 320164
rect 69014 320152 69020 320164
rect 69072 320152 69078 320204
rect 69474 320152 69480 320204
rect 69532 320192 69538 320204
rect 71774 320192 71780 320204
rect 69532 320164 71780 320192
rect 69532 320152 69538 320164
rect 71774 320152 71780 320164
rect 71832 320152 71838 320204
rect 74902 320152 74908 320204
rect 74960 320192 74966 320204
rect 77294 320192 77300 320204
rect 74960 320164 77300 320192
rect 74960 320152 74966 320164
rect 77294 320152 77300 320164
rect 77352 320152 77358 320204
rect 79134 320152 79140 320204
rect 79192 320192 79198 320204
rect 81618 320192 81624 320204
rect 79192 320164 81624 320192
rect 79192 320152 79198 320164
rect 81618 320152 81624 320164
rect 81676 320152 81682 320204
rect 84562 320152 84568 320204
rect 84620 320192 84626 320204
rect 87690 320192 87696 320204
rect 84620 320164 87696 320192
rect 84620 320152 84626 320164
rect 87690 320152 87696 320164
rect 87748 320152 87754 320204
rect 87782 320152 87788 320204
rect 87840 320192 87846 320204
rect 90174 320192 90180 320204
rect 87840 320164 90180 320192
rect 87840 320152 87846 320164
rect 90174 320152 90180 320164
rect 90232 320152 90238 320204
rect 95326 320152 95332 320204
rect 95384 320192 95390 320204
rect 98730 320192 98736 320204
rect 95384 320164 98736 320192
rect 95384 320152 95390 320164
rect 98730 320152 98736 320164
rect 98788 320152 98794 320204
rect 107194 320152 107200 320204
rect 107252 320192 107258 320204
rect 112438 320192 112444 320204
rect 107252 320164 112444 320192
rect 107252 320152 107258 320164
rect 112438 320152 112444 320164
rect 112496 320152 112502 320204
rect 114738 320152 114744 320204
rect 114796 320192 114802 320204
rect 115842 320192 115848 320204
rect 114796 320164 115848 320192
rect 114796 320152 114802 320164
rect 115842 320152 115848 320164
rect 115900 320152 115906 320204
rect 119062 320152 119068 320204
rect 119120 320192 119126 320204
rect 119982 320192 119988 320204
rect 119120 320164 119988 320192
rect 119120 320152 119126 320164
rect 119982 320152 119988 320164
rect 120040 320152 120046 320204
rect 120166 320152 120172 320204
rect 120224 320192 120230 320204
rect 121270 320192 121276 320204
rect 120224 320164 121276 320192
rect 120224 320152 120230 320164
rect 121270 320152 121276 320164
rect 121328 320152 121334 320204
rect 124398 320152 124404 320204
rect 124456 320192 124462 320204
rect 125502 320192 125508 320204
rect 124456 320164 125508 320192
rect 124456 320152 124462 320164
rect 125502 320152 125508 320164
rect 125560 320152 125566 320204
rect 128722 320152 128728 320204
rect 128780 320192 128786 320204
rect 129642 320192 129648 320204
rect 128780 320164 129648 320192
rect 128780 320152 128786 320164
rect 129642 320152 129648 320164
rect 129700 320152 129706 320204
rect 129826 320152 129832 320204
rect 129884 320192 129890 320204
rect 130930 320192 130936 320204
rect 129884 320164 130936 320192
rect 129884 320152 129890 320164
rect 130930 320152 130936 320164
rect 130988 320152 130994 320204
rect 133046 320152 133052 320204
rect 133104 320192 133110 320204
rect 133782 320192 133788 320204
rect 133104 320164 133788 320192
rect 133104 320152 133110 320164
rect 133782 320152 133788 320164
rect 133840 320152 133846 320204
rect 134150 320152 134156 320204
rect 134208 320192 134214 320204
rect 135162 320192 135168 320204
rect 134208 320164 135168 320192
rect 134208 320152 134214 320164
rect 135162 320152 135168 320164
rect 135220 320152 135226 320204
rect 135254 320152 135260 320204
rect 135312 320192 135318 320204
rect 136450 320192 136456 320204
rect 135312 320164 136456 320192
rect 135312 320152 135318 320164
rect 136450 320152 136456 320164
rect 136508 320152 136514 320204
rect 138474 320152 138480 320204
rect 138532 320192 138538 320204
rect 139302 320192 139308 320204
rect 138532 320164 139308 320192
rect 138532 320152 138538 320164
rect 139302 320152 139308 320164
rect 139360 320152 139366 320204
rect 139486 320152 139492 320204
rect 139544 320192 139550 320204
rect 141418 320192 141424 320204
rect 139544 320164 141424 320192
rect 139544 320152 139550 320164
rect 141418 320152 141424 320164
rect 141476 320152 141482 320204
rect 143810 320152 143816 320204
rect 143868 320192 143874 320204
rect 144822 320192 144828 320204
rect 143868 320164 144828 320192
rect 143868 320152 143874 320164
rect 144822 320152 144828 320164
rect 144880 320152 144886 320204
rect 144914 320152 144920 320204
rect 144972 320192 144978 320204
rect 146202 320192 146208 320204
rect 144972 320164 146208 320192
rect 144972 320152 144978 320164
rect 146202 320152 146208 320164
rect 146260 320152 146266 320204
rect 148134 320152 148140 320204
rect 148192 320192 148198 320204
rect 148962 320192 148968 320204
rect 148192 320164 148968 320192
rect 148192 320152 148198 320164
rect 148962 320152 148968 320164
rect 149020 320152 149026 320204
rect 149238 320152 149244 320204
rect 149296 320192 149302 320204
rect 150250 320192 150256 320204
rect 149296 320164 150256 320192
rect 149296 320152 149302 320164
rect 150250 320152 150256 320164
rect 150308 320152 150314 320204
rect 153562 320152 153568 320204
rect 153620 320192 153626 320204
rect 154482 320192 154488 320204
rect 153620 320164 154488 320192
rect 153620 320152 153626 320164
rect 154482 320152 154488 320164
rect 154540 320152 154546 320204
rect 154666 320152 154672 320204
rect 154724 320192 154730 320204
rect 155862 320192 155868 320204
rect 154724 320164 155868 320192
rect 154724 320152 154730 320164
rect 155862 320152 155868 320164
rect 155920 320152 155926 320204
rect 157886 320152 157892 320204
rect 157944 320192 157950 320204
rect 158622 320192 158628 320204
rect 157944 320164 158628 320192
rect 157944 320152 157950 320164
rect 158622 320152 158628 320164
rect 158680 320152 158686 320204
rect 158898 320152 158904 320204
rect 158956 320192 158962 320204
rect 160002 320192 160008 320204
rect 158956 320164 160008 320192
rect 158956 320152 158962 320164
rect 160002 320152 160008 320164
rect 160060 320152 160066 320204
rect 164326 320152 164332 320204
rect 164384 320192 164390 320204
rect 165430 320192 165436 320204
rect 164384 320164 165436 320192
rect 164384 320152 164390 320164
rect 165430 320152 165436 320164
rect 165488 320152 165494 320204
rect 168650 320152 168656 320204
rect 168708 320192 168714 320204
rect 169662 320192 169668 320204
rect 168708 320164 169668 320192
rect 168708 320152 168714 320164
rect 169662 320152 169668 320164
rect 169720 320152 169726 320204
rect 169754 320152 169760 320204
rect 169812 320192 169818 320204
rect 170950 320192 170956 320204
rect 169812 320164 170956 320192
rect 169812 320152 169818 320164
rect 170950 320152 170956 320164
rect 171008 320152 171014 320204
rect 172974 320152 172980 320204
rect 173032 320192 173038 320204
rect 173802 320192 173808 320204
rect 173032 320164 173808 320192
rect 173032 320152 173038 320164
rect 173802 320152 173808 320164
rect 173860 320152 173866 320204
rect 173986 320152 173992 320204
rect 174044 320192 174050 320204
rect 175182 320192 175188 320204
rect 174044 320164 175188 320192
rect 174044 320152 174050 320164
rect 175182 320152 175188 320164
rect 175240 320152 175246 320204
rect 178310 320152 178316 320204
rect 178368 320192 178374 320204
rect 179322 320192 179328 320204
rect 178368 320164 179328 320192
rect 178368 320152 178374 320164
rect 179322 320152 179328 320164
rect 179380 320152 179386 320204
rect 179414 320152 179420 320204
rect 179472 320192 179478 320204
rect 180610 320192 180616 320204
rect 179472 320164 180616 320192
rect 179472 320152 179478 320164
rect 180610 320152 180616 320164
rect 180668 320152 180674 320204
rect 182634 320152 182640 320204
rect 182692 320192 182698 320204
rect 183462 320192 183468 320204
rect 182692 320164 183468 320192
rect 182692 320152 182698 320164
rect 183462 320152 183468 320164
rect 183520 320152 183526 320204
rect 183738 320152 183744 320204
rect 183796 320192 183802 320204
rect 184842 320192 184848 320204
rect 183796 320164 184848 320192
rect 183796 320152 183802 320164
rect 184842 320152 184848 320164
rect 184900 320152 184906 320204
rect 197446 320152 197452 320204
rect 197504 320192 197510 320204
rect 199930 320192 199936 320204
rect 197504 320164 199936 320192
rect 197504 320152 197510 320164
rect 199930 320152 199936 320164
rect 199988 320152 199994 320204
rect 201126 320152 201132 320204
rect 201184 320192 201190 320204
rect 203150 320192 203156 320204
rect 201184 320164 203156 320192
rect 201184 320152 201190 320164
rect 203150 320152 203156 320164
rect 203208 320152 203214 320204
rect 207106 320152 207112 320204
rect 207164 320192 207170 320204
rect 209590 320192 209596 320204
rect 207164 320164 209596 320192
rect 207164 320152 207170 320164
rect 209590 320152 209596 320164
rect 209648 320152 209654 320204
rect 219894 320152 219900 320204
rect 219952 320192 219958 320204
rect 224678 320192 224684 320204
rect 219952 320164 224684 320192
rect 219952 320152 219958 320164
rect 224678 320152 224684 320164
rect 224736 320152 224742 320204
rect 224862 320152 224868 320204
rect 224920 320192 224926 320204
rect 229002 320192 229008 320204
rect 224920 320164 229008 320192
rect 224920 320152 224926 320164
rect 229002 320152 229008 320164
rect 229060 320152 229066 320204
rect 230290 320152 230296 320204
rect 230348 320192 230354 320204
rect 234338 320192 234344 320204
rect 230348 320164 234344 320192
rect 230348 320152 230354 320164
rect 234338 320152 234344 320164
rect 234396 320152 234402 320204
rect 234522 320152 234528 320204
rect 234580 320192 234586 320204
rect 237650 320192 237656 320204
rect 234580 320164 237656 320192
rect 234580 320152 234586 320164
rect 237650 320152 237656 320164
rect 237708 320152 237714 320204
rect 240042 320152 240048 320204
rect 240100 320192 240106 320204
rect 242986 320192 242992 320204
rect 240100 320164 242992 320192
rect 240100 320152 240106 320164
rect 242986 320152 242992 320164
rect 243044 320152 243050 320204
rect 243814 320152 243820 320204
rect 243872 320192 243878 320204
rect 246206 320192 246212 320204
rect 243872 320164 246212 320192
rect 243872 320152 243878 320164
rect 246206 320152 246212 320164
rect 246264 320152 246270 320204
rect 249702 320152 249708 320204
rect 249760 320192 249766 320204
rect 251634 320192 251640 320204
rect 249760 320164 251640 320192
rect 249760 320152 249766 320164
rect 251634 320152 251640 320164
rect 251692 320152 251698 320204
rect 252462 320152 252468 320204
rect 252520 320192 252526 320204
rect 253750 320192 253756 320204
rect 252520 320164 253756 320192
rect 252520 320152 252526 320164
rect 253750 320152 253756 320164
rect 253808 320152 253814 320204
rect 255774 320152 255780 320204
rect 255832 320192 255838 320204
rect 256970 320192 256976 320204
rect 255832 320164 256976 320192
rect 255832 320152 255838 320164
rect 256970 320152 256976 320164
rect 257028 320152 257034 320204
rect 259362 320152 259368 320204
rect 259420 320192 259426 320204
rect 260282 320192 260288 320204
rect 259420 320164 260288 320192
rect 259420 320152 259426 320164
rect 260282 320152 260288 320164
rect 260340 320152 260346 320204
rect 263502 320192 263508 320204
rect 262232 320164 263508 320192
rect 41414 320084 41420 320136
rect 41472 320084 41478 320136
rect 262232 320068 262260 320164
rect 263502 320152 263508 320164
rect 263560 320152 263566 320204
rect 263594 320152 263600 320204
rect 263652 320192 263658 320204
rect 264514 320192 264520 320204
rect 263652 320164 264520 320192
rect 263652 320152 263658 320164
rect 264514 320152 264520 320164
rect 264572 320152 264578 320204
rect 267734 320152 267740 320204
rect 267792 320192 267798 320204
rect 268838 320192 268844 320204
rect 267792 320164 268844 320192
rect 267792 320152 267798 320164
rect 268838 320152 268844 320164
rect 268896 320152 268902 320204
rect 269114 320152 269120 320204
rect 269172 320192 269178 320204
rect 269942 320192 269948 320204
rect 269172 320164 269948 320192
rect 269172 320152 269178 320164
rect 269942 320152 269948 320164
rect 270000 320152 270006 320204
rect 262214 320016 262220 320068
rect 262272 320016 262278 320068
rect 22094 319404 22100 319456
rect 22152 319444 22158 319456
rect 113174 319444 113180 319456
rect 22152 319416 113180 319444
rect 22152 319404 22158 319416
rect 113174 319404 113180 319416
rect 113232 319404 113238 319456
rect 113634 319404 113640 319456
rect 113692 319444 113698 319456
rect 128446 319444 128452 319456
rect 113692 319416 128452 319444
rect 113692 319404 113698 319416
rect 128446 319404 128452 319416
rect 128504 319404 128510 319456
rect 195606 319404 195612 319456
rect 195664 319444 195670 319456
rect 280154 319444 280160 319456
rect 195664 319416 280160 319444
rect 195664 319404 195670 319416
rect 280154 319404 280160 319416
rect 280212 319404 280218 319456
rect 20622 318724 20628 318776
rect 20680 318764 20686 318776
rect 23106 318764 23112 318776
rect 20680 318736 23112 318764
rect 20680 318724 20686 318736
rect 23106 318724 23112 318736
rect 23164 318724 23170 318776
rect 90174 318724 90180 318776
rect 90232 318764 90238 318776
rect 92290 318764 92296 318776
rect 90232 318736 92296 318764
rect 90232 318724 90238 318736
rect 92290 318724 92296 318736
rect 92348 318724 92354 318776
rect 192386 318724 192392 318776
rect 192444 318764 192450 318776
rect 197446 318764 197452 318776
rect 192444 318736 197452 318764
rect 192444 318724 192450 318736
rect 197446 318724 197452 318736
rect 197504 318724 197510 318776
rect 201954 318724 201960 318776
rect 202012 318764 202018 318776
rect 208302 318764 208308 318776
rect 202012 318736 208308 318764
rect 202012 318724 202018 318736
rect 208302 318724 208308 318736
rect 208360 318724 208366 318776
rect 211522 318724 211528 318776
rect 211580 318764 211586 318776
rect 217134 318764 217140 318776
rect 211580 318736 217140 318764
rect 211580 318724 211586 318736
rect 217134 318724 217140 318736
rect 217192 318724 217198 318776
rect 223482 318724 223488 318776
rect 223540 318764 223546 318776
rect 227898 318764 227904 318776
rect 223540 318736 227904 318764
rect 223540 318724 223546 318736
rect 227898 318724 227904 318736
rect 227956 318724 227962 318776
rect 200758 318656 200764 318708
rect 200816 318696 200822 318708
rect 206922 318696 206928 318708
rect 200816 318668 206928 318696
rect 200816 318656 200822 318668
rect 206922 318656 206928 318668
rect 206980 318656 206986 318708
rect 220630 318656 220636 318708
rect 220688 318696 220694 318708
rect 225782 318696 225788 318708
rect 220688 318668 225788 318696
rect 220688 318656 220694 318668
rect 225782 318656 225788 318668
rect 225840 318656 225846 318708
rect 202782 318588 202788 318640
rect 202840 318628 202846 318640
rect 207106 318628 207112 318640
rect 202840 318600 207112 318628
rect 202840 318588 202846 318600
rect 207106 318588 207112 318600
rect 207164 318588 207170 318640
rect 92382 318520 92388 318572
rect 92440 318560 92446 318572
rect 93486 318560 93492 318572
rect 92440 318532 93492 318560
rect 92440 318520 92446 318532
rect 93486 318520 93492 318532
rect 93544 318520 93550 318572
rect 98730 318520 98736 318572
rect 98788 318560 98794 318572
rect 100662 318560 100668 318572
rect 98788 318532 100668 318560
rect 98788 318520 98794 318532
rect 100662 318520 100668 318532
rect 100720 318520 100726 318572
rect 106366 318520 106372 318572
rect 106424 318560 106430 318572
rect 107838 318560 107844 318572
rect 106424 318532 107844 318560
rect 106424 318520 106430 318532
rect 107838 318520 107844 318532
rect 107896 318520 107902 318572
rect 194502 318452 194508 318504
rect 194560 318492 194566 318504
rect 198734 318492 198740 318504
rect 194560 318464 198740 318492
rect 194560 318452 194566 318464
rect 198734 318452 198740 318464
rect 198792 318452 198798 318504
rect 209130 318452 209136 318504
rect 209188 318492 209194 318504
rect 215018 318492 215024 318504
rect 209188 318464 215024 318492
rect 209188 318452 209194 318464
rect 215018 318452 215024 318464
rect 215076 318452 215082 318504
rect 85114 318384 85120 318436
rect 85172 318424 85178 318436
rect 86310 318424 86316 318436
rect 85172 318396 86316 318424
rect 85172 318384 85178 318396
rect 86310 318384 86316 318396
rect 86368 318384 86374 318436
rect 85666 318316 85672 318368
rect 85724 318356 85730 318368
rect 87506 318356 87512 318368
rect 85724 318328 87512 318356
rect 85724 318316 85730 318328
rect 87506 318316 87512 318328
rect 87564 318316 87570 318368
rect 195882 318316 195888 318368
rect 195940 318356 195946 318368
rect 201126 318356 201132 318368
rect 195940 318328 201132 318356
rect 195940 318316 195946 318328
rect 201126 318316 201132 318328
rect 201184 318316 201190 318368
rect 204162 318316 204168 318368
rect 204220 318356 204226 318368
rect 208394 318356 208400 318368
rect 204220 318328 208400 318356
rect 204220 318316 204226 318328
rect 208394 318316 208400 318328
rect 208452 318316 208458 318368
rect 191190 318248 191196 318300
rect 191248 318288 191254 318300
rect 195974 318288 195980 318300
rect 191248 318260 195980 318288
rect 191248 318248 191254 318260
rect 195974 318248 195980 318260
rect 196032 318248 196038 318300
rect 199562 318248 199568 318300
rect 199620 318288 199626 318300
rect 204254 318288 204260 318300
rect 199620 318260 204260 318288
rect 199620 318248 199626 318260
rect 204254 318248 204260 318260
rect 204312 318248 204318 318300
rect 217502 318248 217508 318300
rect 217560 318288 217566 318300
rect 222562 318288 222568 318300
rect 217560 318260 222568 318288
rect 217560 318248 217566 318260
rect 222562 318248 222568 318260
rect 222620 318248 222626 318300
rect 87690 318180 87696 318232
rect 87748 318220 87754 318232
rect 88702 318220 88708 318232
rect 87748 318192 88708 318220
rect 87748 318180 87754 318192
rect 88702 318180 88708 318192
rect 88760 318180 88766 318232
rect 207934 318180 207940 318232
rect 207992 318220 207998 318232
rect 213822 318220 213828 318232
rect 207992 318192 213828 318220
rect 207992 318180 207998 318192
rect 213822 318180 213828 318192
rect 213880 318180 213886 318232
rect 198366 318112 198372 318164
rect 198424 318152 198430 318164
rect 202874 318152 202880 318164
rect 198424 318124 202880 318152
rect 198424 318112 198430 318124
rect 202874 318112 202880 318124
rect 202932 318112 202938 318164
rect 189994 318044 190000 318096
rect 190052 318084 190058 318096
rect 197262 318084 197268 318096
rect 190052 318056 197268 318084
rect 190052 318044 190058 318056
rect 197262 318044 197268 318056
rect 197320 318044 197326 318096
rect 218698 318044 218704 318096
rect 218756 318084 218762 318096
rect 223574 318084 223580 318096
rect 218756 318056 223580 318084
rect 218756 318044 218762 318056
rect 223574 318044 223580 318056
rect 223632 318044 223638 318096
rect 213822 317908 213828 317960
rect 213880 317948 213886 317960
rect 219250 317948 219256 317960
rect 213880 317920 219256 317948
rect 213880 317908 213886 317920
rect 219250 317908 219256 317920
rect 219308 317908 219314 317960
rect 222010 317908 222016 317960
rect 222068 317948 222074 317960
rect 226794 317948 226800 317960
rect 222068 317920 226800 317948
rect 222068 317908 222074 317920
rect 226794 317908 226800 317920
rect 226852 317908 226858 317960
rect 193582 317840 193588 317892
rect 193640 317880 193646 317892
rect 198826 317880 198832 317892
rect 193640 317852 198832 317880
rect 193640 317840 193646 317852
rect 198826 317840 198832 317852
rect 198884 317840 198890 317892
rect 210326 317704 210332 317756
rect 210384 317744 210390 317756
rect 216030 317744 216036 317756
rect 210384 317716 216036 317744
rect 210384 317704 210390 317716
rect 216030 317704 216036 317716
rect 216088 317704 216094 317756
rect 206738 317568 206744 317620
rect 206796 317608 206802 317620
rect 212442 317608 212448 317620
rect 206796 317580 212448 317608
rect 206796 317568 206802 317580
rect 212442 317568 212448 317580
rect 212500 317568 212506 317620
rect 216306 317568 216312 317620
rect 216364 317608 216370 317620
rect 221458 317608 221464 317620
rect 216364 317580 221464 317608
rect 216364 317568 216370 317580
rect 221458 317568 221464 317580
rect 221516 317568 221522 317620
rect 82814 317500 82820 317552
rect 82872 317540 82878 317552
rect 85114 317540 85120 317552
rect 82872 317512 85120 317540
rect 82872 317500 82878 317512
rect 85114 317500 85120 317512
rect 85172 317500 85178 317552
rect 197170 317500 197176 317552
rect 197228 317540 197234 317552
rect 202138 317540 202144 317552
rect 197228 317512 202144 317540
rect 197228 317500 197234 317512
rect 202138 317500 202144 317512
rect 202196 317500 202202 317552
rect 205542 317500 205548 317552
rect 205600 317540 205606 317552
rect 211062 317540 211068 317552
rect 205600 317512 211068 317540
rect 205600 317500 205606 317512
rect 211062 317500 211068 317512
rect 211120 317500 211126 317552
rect 217962 317540 217968 317552
rect 212460 317512 217968 317540
rect 212460 317484 212488 317512
rect 217962 317500 217968 317512
rect 218020 317500 218026 317552
rect 92750 317432 92756 317484
rect 92808 317472 92814 317484
rect 94682 317472 94688 317484
rect 92808 317444 94688 317472
rect 92808 317432 92814 317444
rect 94682 317432 94688 317444
rect 94740 317432 94746 317484
rect 188614 317432 188620 317484
rect 188672 317472 188678 317484
rect 192478 317472 192484 317484
rect 188672 317444 192484 317472
rect 188672 317432 188678 317444
rect 192478 317432 192484 317444
rect 192536 317432 192542 317484
rect 212442 317432 212448 317484
rect 212500 317432 212506 317484
rect 215110 317432 215116 317484
rect 215168 317472 215174 317484
rect 220354 317472 220360 317484
rect 215168 317444 220360 317472
rect 215168 317432 215174 317444
rect 220354 317432 220360 317444
rect 220412 317432 220418 317484
rect 2774 316684 2780 316736
rect 2832 316724 2838 316736
rect 3418 316724 3424 316736
rect 2832 316696 3424 316724
rect 2832 316684 2838 316696
rect 3418 316684 3424 316696
rect 3476 316724 3482 316736
rect 288894 316724 288900 316736
rect 3476 316696 288900 316724
rect 3476 316684 3482 316696
rect 288894 316684 288900 316696
rect 288952 316684 288958 316736
rect 26878 315324 26884 315376
rect 26936 315364 26942 315376
rect 111794 315364 111800 315376
rect 26936 315336 111800 315364
rect 26936 315324 26942 315336
rect 111794 315324 111800 315336
rect 111852 315324 111858 315376
rect 15838 315256 15844 315308
rect 15896 315296 15902 315308
rect 185578 315296 185584 315308
rect 15896 315268 185584 315296
rect 15896 315256 15902 315268
rect 185578 315256 185584 315268
rect 185636 315256 185642 315308
rect 111794 313624 111800 313676
rect 111852 313664 111858 313676
rect 113542 313664 113548 313676
rect 111852 313636 113548 313664
rect 111852 313624 111858 313636
rect 113542 313624 113548 313636
rect 113600 313624 113606 313676
rect 303614 311856 303620 311908
rect 303672 311896 303678 311908
rect 335998 311896 336004 311908
rect 303672 311868 336004 311896
rect 303672 311856 303678 311868
rect 335998 311856 336004 311868
rect 336056 311856 336062 311908
rect 113542 311584 113548 311636
rect 113600 311624 113606 311636
rect 116578 311624 116584 311636
rect 113600 311596 116584 311624
rect 113600 311584 113606 311596
rect 116578 311584 116584 311596
rect 116636 311584 116642 311636
rect 303614 310496 303620 310548
rect 303672 310536 303678 310548
rect 341518 310536 341524 310548
rect 303672 310508 341524 310536
rect 303672 310496 303678 310508
rect 341518 310496 341524 310508
rect 341576 310496 341582 310548
rect 303614 309136 303620 309188
rect 303672 309176 303678 309188
rect 340138 309176 340144 309188
rect 303672 309148 340144 309176
rect 303672 309136 303678 309148
rect 340138 309136 340144 309148
rect 340196 309136 340202 309188
rect 303614 306348 303620 306400
rect 303672 306388 303678 306400
rect 560938 306388 560944 306400
rect 303672 306360 560944 306388
rect 303672 306348 303678 306360
rect 560938 306348 560944 306360
rect 560996 306348 561002 306400
rect 282178 305600 282184 305652
rect 282236 305640 282242 305652
rect 300854 305640 300860 305652
rect 282236 305612 300860 305640
rect 282236 305600 282242 305612
rect 300854 305600 300860 305612
rect 300912 305600 300918 305652
rect 296162 303560 296168 303612
rect 296220 303600 296226 303612
rect 580350 303600 580356 303612
rect 296220 303572 580356 303600
rect 296220 303560 296226 303572
rect 580350 303560 580356 303572
rect 580408 303560 580414 303612
rect 3418 293972 3424 294024
rect 3476 294012 3482 294024
rect 15838 294012 15844 294024
rect 3476 293984 15844 294012
rect 3476 293972 3482 293984
rect 15838 293972 15844 293984
rect 15896 293972 15902 294024
rect 11790 275952 11796 276004
rect 11848 275992 11854 276004
rect 17126 275992 17132 276004
rect 11848 275964 17132 275992
rect 11848 275952 11854 275964
rect 17126 275952 17132 275964
rect 17184 275952 17190 276004
rect 304350 275952 304356 276004
rect 304408 275992 304414 276004
rect 580166 275992 580172 276004
rect 304408 275964 580172 275992
rect 304408 275952 304414 275964
rect 580166 275952 580172 275964
rect 580224 275952 580230 276004
rect 117222 236648 117228 236700
rect 117280 236688 117286 236700
rect 132494 236688 132500 236700
rect 117280 236660 132500 236688
rect 117280 236648 117286 236660
rect 132494 236648 132500 236660
rect 132552 236648 132558 236700
rect 113910 235900 113916 235952
rect 113968 235940 113974 235952
rect 281534 235940 281540 235952
rect 113968 235912 281540 235940
rect 113968 235900 113974 235912
rect 281534 235900 281540 235912
rect 281592 235900 281598 235952
rect 180610 235220 180616 235272
rect 180668 235260 180674 235272
rect 194594 235260 194600 235272
rect 180668 235232 194600 235260
rect 180668 235220 180674 235232
rect 194594 235220 194600 235232
rect 194652 235220 194658 235272
rect 10502 233860 10508 233912
rect 10560 233900 10566 233912
rect 299474 233900 299480 233912
rect 10560 233872 299480 233900
rect 10560 233860 10566 233872
rect 299474 233860 299480 233872
rect 299532 233860 299538 233912
rect 146202 232500 146208 232552
rect 146260 232540 146266 232552
rect 160094 232540 160100 232552
rect 146260 232512 160100 232540
rect 146260 232500 146266 232512
rect 160094 232500 160100 232512
rect 160152 232500 160158 232552
rect 227622 232500 227628 232552
rect 227680 232540 227686 232552
rect 313918 232540 313924 232552
rect 227680 232512 313924 232540
rect 227680 232500 227686 232512
rect 313918 232500 313924 232512
rect 313976 232500 313982 232552
rect 143442 231072 143448 231124
rect 143500 231112 143506 231124
rect 157518 231112 157524 231124
rect 143500 231084 157524 231112
rect 143500 231072 143506 231084
rect 157518 231072 157524 231084
rect 157576 231072 157582 231124
rect 166902 231072 166908 231124
rect 166960 231112 166966 231124
rect 180886 231112 180892 231124
rect 166960 231084 180892 231112
rect 166960 231072 166966 231084
rect 180886 231072 180892 231084
rect 180944 231072 180950 231124
rect 214742 231072 214748 231124
rect 214800 231112 214806 231124
rect 305638 231112 305644 231124
rect 214800 231084 305644 231112
rect 214800 231072 214806 231084
rect 305638 231072 305644 231084
rect 305696 231072 305702 231124
rect 140682 229712 140688 229764
rect 140740 229752 140746 229764
rect 155954 229752 155960 229764
rect 140740 229724 155960 229752
rect 140740 229712 140746 229724
rect 155954 229712 155960 229724
rect 156012 229712 156018 229764
rect 159910 229712 159916 229764
rect 159968 229752 159974 229764
rect 175274 229752 175280 229764
rect 159968 229724 175280 229752
rect 159968 229712 159974 229724
rect 175274 229712 175280 229724
rect 175332 229712 175338 229764
rect 214558 229712 214564 229764
rect 214616 229752 214622 229764
rect 308398 229752 308404 229764
rect 214616 229724 308404 229752
rect 214616 229712 214622 229724
rect 308398 229712 308404 229724
rect 308456 229712 308462 229764
rect 304258 229032 304264 229084
rect 304316 229072 304322 229084
rect 579982 229072 579988 229084
rect 304316 229044 579988 229072
rect 304316 229032 304322 229044
rect 579982 229032 579988 229044
rect 580040 229032 580046 229084
rect 139302 228352 139308 228404
rect 139360 228392 139366 228404
rect 154298 228392 154304 228404
rect 139360 228364 154304 228392
rect 139360 228352 139366 228364
rect 154298 228352 154304 228364
rect 154356 228352 154362 228404
rect 155770 228352 155776 228404
rect 155828 228392 155834 228404
rect 171410 228392 171416 228404
rect 155828 228364 171416 228392
rect 155828 228352 155834 228364
rect 171410 228352 171416 228364
rect 171468 228352 171474 228404
rect 175090 228352 175096 228404
rect 175148 228392 175154 228404
rect 190638 228392 190644 228404
rect 175148 228364 190644 228392
rect 175148 228352 175154 228364
rect 190638 228352 190644 228364
rect 190696 228352 190702 228404
rect 214926 228352 214932 228404
rect 214984 228392 214990 228404
rect 287698 228392 287704 228404
rect 214984 228364 287704 228392
rect 214984 228352 214990 228364
rect 287698 228352 287704 228364
rect 287756 228352 287762 228404
rect 135162 227060 135168 227112
rect 135220 227100 135226 227112
rect 149974 227100 149980 227112
rect 135220 227072 149980 227100
rect 135220 227060 135226 227072
rect 149974 227060 149980 227072
rect 150032 227060 150038 227112
rect 162762 227060 162768 227112
rect 162820 227100 162826 227112
rect 177758 227100 177764 227112
rect 162820 227072 177764 227100
rect 162820 227060 162826 227072
rect 177758 227060 177764 227072
rect 177816 227060 177822 227112
rect 15838 226992 15844 227044
rect 15896 227032 15902 227044
rect 120074 227032 120080 227044
rect 15896 227004 120080 227032
rect 15896 226992 15902 227004
rect 120074 226992 120080 227004
rect 120132 226992 120138 227044
rect 121270 226992 121276 227044
rect 121328 227032 121334 227044
rect 136082 227032 136088 227044
rect 121328 227004 136088 227032
rect 121328 226992 121334 227004
rect 136082 226992 136088 227004
rect 136140 226992 136146 227044
rect 147582 226992 147588 227044
rect 147640 227032 147646 227044
rect 162854 227032 162860 227044
rect 147640 227004 162860 227032
rect 147640 226992 147646 227004
rect 162854 226992 162860 227004
rect 162912 226992 162918 227044
rect 214650 226992 214656 227044
rect 214708 227032 214714 227044
rect 309778 227032 309784 227044
rect 214708 227004 309784 227032
rect 214708 226992 214714 227004
rect 309778 226992 309784 227004
rect 309836 226992 309842 227044
rect 14458 225564 14464 225616
rect 14516 225604 14522 225616
rect 411990 225604 411996 225616
rect 14516 225576 411996 225604
rect 14516 225564 14522 225576
rect 411990 225564 411996 225576
rect 412048 225564 412054 225616
rect 119338 224884 119344 224936
rect 119396 224924 119402 224936
rect 125410 224924 125416 224936
rect 119396 224896 125416 224924
rect 119396 224884 119402 224896
rect 125410 224884 125416 224896
rect 125468 224884 125474 224936
rect 125502 224884 125508 224936
rect 125560 224924 125566 224936
rect 133690 224924 133696 224936
rect 125560 224896 133696 224924
rect 125560 224884 125566 224896
rect 133690 224884 133696 224896
rect 133748 224884 133754 224936
rect 133782 224884 133788 224936
rect 133840 224924 133846 224936
rect 139394 224924 139400 224936
rect 133840 224896 139400 224924
rect 133840 224884 133846 224896
rect 139394 224884 139400 224896
rect 139452 224884 139458 224936
rect 144822 224884 144828 224936
rect 144880 224924 144886 224936
rect 159634 224924 159640 224936
rect 144880 224896 159640 224924
rect 144880 224884 144886 224896
rect 159634 224884 159640 224896
rect 159692 224884 159698 224936
rect 160002 224884 160008 224936
rect 160060 224924 160066 224936
rect 174630 224924 174636 224936
rect 160060 224896 174636 224924
rect 160060 224884 160066 224896
rect 174630 224884 174636 224896
rect 174688 224884 174694 224936
rect 176562 224884 176568 224936
rect 176620 224924 176626 224936
rect 191742 224924 191748 224936
rect 176620 224896 191748 224924
rect 176620 224884 176626 224896
rect 191742 224884 191748 224896
rect 191800 224884 191806 224936
rect 115198 224816 115204 224868
rect 115256 224856 115262 224868
rect 124306 224856 124312 224868
rect 115256 224828 124312 224856
rect 115256 224816 115262 224828
rect 124306 224816 124312 224828
rect 124364 224816 124370 224868
rect 130930 224816 130936 224868
rect 130988 224856 130994 224868
rect 145742 224856 145748 224868
rect 130988 224828 145748 224856
rect 130988 224816 130994 224828
rect 145742 224816 145748 224828
rect 145800 224816 145806 224868
rect 152458 224816 152464 224868
rect 152516 224856 152522 224868
rect 161750 224856 161756 224868
rect 152516 224828 161756 224856
rect 152516 224816 152522 224828
rect 161750 224816 161756 224828
rect 161808 224816 161814 224868
rect 169662 224816 169668 224868
rect 169720 224856 169726 224868
rect 183830 224856 183836 224868
rect 169720 224828 183836 224856
rect 169720 224816 169726 224828
rect 183830 224816 183836 224828
rect 183888 224816 183894 224868
rect 184198 224816 184204 224868
rect 184256 224856 184262 224868
rect 197078 224856 197084 224868
rect 184256 224828 197084 224856
rect 184256 224816 184262 224828
rect 197078 224816 197084 224828
rect 197136 224816 197142 224868
rect 119982 224748 119988 224800
rect 120040 224788 120046 224800
rect 126146 224788 126152 224800
rect 120040 224760 126152 224788
rect 120040 224748 120046 224760
rect 126146 224748 126152 224760
rect 126204 224748 126210 224800
rect 126238 224748 126244 224800
rect 126296 224788 126302 224800
rect 131758 224788 131764 224800
rect 126296 224760 131764 224788
rect 126296 224748 126302 224760
rect 131758 224748 131764 224760
rect 131816 224748 131822 224800
rect 136450 224748 136456 224800
rect 136508 224788 136514 224800
rect 151078 224788 151084 224800
rect 136508 224760 151084 224788
rect 136508 224748 136514 224760
rect 151078 224748 151084 224760
rect 151136 224748 151142 224800
rect 154482 224748 154488 224800
rect 154540 224788 154546 224800
rect 169202 224788 169208 224800
rect 154540 224760 169208 224788
rect 154540 224748 154546 224760
rect 169202 224748 169208 224760
rect 169260 224748 169266 224800
rect 172422 224748 172428 224800
rect 172480 224788 172486 224800
rect 172480 224760 184152 224788
rect 172480 224748 172486 224760
rect 117958 224680 117964 224732
rect 118016 224720 118022 224732
rect 127526 224720 127532 224732
rect 118016 224692 127532 224720
rect 118016 224680 118022 224692
rect 127526 224680 127532 224692
rect 127584 224680 127590 224732
rect 128262 224680 128268 224732
rect 128320 224720 128326 224732
rect 143534 224720 143540 224732
rect 128320 224692 143540 224720
rect 128320 224680 128326 224692
rect 143534 224680 143540 224692
rect 143592 224680 143598 224732
rect 153102 224680 153108 224732
rect 153160 224720 153166 224732
rect 168190 224720 168196 224732
rect 153160 224692 168196 224720
rect 153160 224680 153166 224692
rect 168190 224680 168196 224692
rect 168248 224680 168254 224732
rect 175182 224680 175188 224732
rect 175240 224720 175246 224732
rect 184014 224720 184020 224732
rect 175240 224692 184020 224720
rect 175240 224680 175246 224692
rect 184014 224680 184020 224692
rect 184072 224680 184078 224732
rect 184124 224720 184152 224760
rect 186958 224748 186964 224800
rect 187016 224788 187022 224800
rect 200298 224788 200304 224800
rect 187016 224760 200304 224788
rect 187016 224748 187022 224760
rect 200298 224748 200304 224760
rect 200356 224748 200362 224800
rect 187418 224720 187424 224732
rect 184124 224692 187424 224720
rect 187418 224680 187424 224692
rect 187476 224680 187482 224732
rect 115842 224612 115848 224664
rect 115900 224652 115906 224664
rect 130746 224652 130752 224664
rect 115900 224624 130752 224652
rect 115900 224612 115906 224624
rect 130746 224612 130752 224624
rect 130804 224612 130810 224664
rect 132402 224612 132408 224664
rect 132460 224652 132466 224664
rect 147858 224652 147864 224664
rect 132460 224624 147864 224652
rect 132460 224612 132466 224624
rect 147858 224612 147864 224624
rect 147916 224612 147922 224664
rect 148962 224612 148968 224664
rect 149020 224652 149026 224664
rect 163866 224652 163872 224664
rect 149020 224624 163872 224652
rect 149020 224612 149026 224624
rect 163866 224612 163872 224624
rect 163924 224612 163930 224664
rect 177942 224612 177948 224664
rect 178000 224652 178006 224664
rect 192754 224652 192760 224664
rect 178000 224624 192760 224652
rect 178000 224612 178006 224624
rect 192754 224612 192760 224624
rect 192812 224612 192818 224664
rect 113818 224544 113824 224596
rect 113876 224584 113882 224596
rect 126422 224584 126428 224596
rect 113876 224556 126428 224584
rect 113876 224544 113882 224556
rect 126422 224544 126428 224556
rect 126480 224544 126486 224596
rect 126882 224544 126888 224596
rect 126940 224584 126946 224596
rect 142522 224584 142528 224596
rect 126940 224556 142528 224584
rect 126940 224544 126946 224556
rect 142522 224544 142528 224556
rect 142580 224544 142586 224596
rect 150250 224544 150256 224596
rect 150308 224584 150314 224596
rect 164970 224584 164976 224596
rect 150308 224556 164976 224584
rect 150308 224544 150314 224556
rect 164970 224544 164976 224556
rect 165028 224544 165034 224596
rect 165430 224544 165436 224596
rect 165488 224584 165494 224596
rect 179966 224584 179972 224596
rect 165488 224556 179972 224584
rect 165488 224544 165494 224556
rect 179966 224544 179972 224556
rect 180024 224544 180030 224596
rect 184842 224544 184848 224596
rect 184900 224584 184906 224596
rect 199194 224584 199200 224596
rect 184900 224556 199200 224584
rect 184900 224544 184906 224556
rect 199194 224544 199200 224556
rect 199252 224544 199258 224596
rect 113082 224476 113088 224528
rect 113140 224516 113146 224528
rect 128630 224516 128636 224528
rect 113140 224488 128636 224516
rect 113140 224476 113146 224488
rect 128630 224476 128636 224488
rect 128688 224476 128694 224528
rect 131022 224476 131028 224528
rect 131080 224516 131086 224528
rect 146754 224516 146760 224528
rect 131080 224488 146760 224516
rect 131080 224476 131086 224488
rect 146754 224476 146760 224488
rect 146812 224476 146818 224528
rect 151722 224476 151728 224528
rect 151780 224516 151786 224528
rect 167086 224516 167092 224528
rect 151780 224488 167092 224516
rect 151780 224476 151786 224488
rect 167086 224476 167092 224488
rect 167144 224476 167150 224528
rect 168282 224476 168288 224528
rect 168340 224516 168346 224528
rect 183186 224516 183192 224528
rect 168340 224488 183192 224516
rect 168340 224476 168346 224488
rect 183186 224476 183192 224488
rect 183244 224476 183250 224528
rect 183462 224476 183468 224528
rect 183520 224516 183526 224528
rect 198090 224516 198096 224528
rect 183520 224488 198096 224516
rect 183520 224476 183526 224488
rect 198090 224476 198096 224488
rect 198148 224476 198154 224528
rect 118602 224408 118608 224460
rect 118660 224448 118666 224460
rect 133966 224448 133972 224460
rect 118660 224420 133972 224448
rect 118660 224408 118666 224420
rect 133966 224408 133972 224420
rect 134024 224408 134030 224460
rect 136542 224408 136548 224460
rect 136600 224448 136606 224460
rect 152090 224448 152096 224460
rect 136600 224420 152096 224448
rect 136600 224408 136606 224420
rect 152090 224408 152096 224420
rect 152148 224408 152154 224460
rect 155862 224408 155868 224460
rect 155920 224448 155926 224460
rect 170306 224448 170312 224460
rect 155920 224420 170312 224448
rect 155920 224408 155926 224420
rect 170306 224408 170312 224420
rect 170364 224408 170370 224460
rect 170950 224408 170956 224460
rect 171008 224448 171014 224460
rect 185302 224448 185308 224460
rect 171008 224420 185308 224448
rect 171008 224408 171014 224420
rect 185302 224408 185308 224420
rect 185360 224408 185366 224460
rect 186222 224408 186228 224460
rect 186280 224448 186286 224460
rect 201310 224448 201316 224460
rect 186280 224420 201316 224448
rect 186280 224408 186286 224420
rect 201310 224408 201316 224420
rect 201368 224408 201374 224460
rect 121362 224340 121368 224392
rect 121420 224380 121426 224392
rect 137186 224380 137192 224392
rect 121420 224352 137192 224380
rect 121420 224340 121426 224352
rect 137186 224340 137192 224352
rect 137244 224340 137250 224392
rect 137922 224340 137928 224392
rect 137980 224380 137986 224392
rect 153194 224380 153200 224392
rect 137980 224352 153200 224380
rect 137980 224340 137986 224352
rect 153194 224340 153200 224352
rect 153252 224340 153258 224392
rect 165522 224340 165528 224392
rect 165580 224380 165586 224392
rect 180978 224380 180984 224392
rect 165580 224352 180984 224380
rect 165580 224340 165586 224352
rect 180978 224340 180984 224352
rect 181036 224340 181042 224392
rect 187602 224340 187608 224392
rect 187660 224380 187666 224392
rect 202414 224380 202420 224392
rect 187660 224352 202420 224380
rect 187660 224340 187666 224352
rect 202414 224340 202420 224352
rect 202472 224340 202478 224392
rect 122742 224272 122748 224324
rect 122800 224312 122806 224324
rect 138198 224312 138204 224324
rect 122800 224284 138204 224312
rect 122800 224272 122806 224284
rect 138198 224272 138204 224284
rect 138256 224272 138262 224324
rect 142062 224272 142068 224324
rect 142120 224312 142126 224324
rect 157426 224312 157432 224324
rect 142120 224284 157432 224312
rect 142120 224272 142126 224284
rect 157426 224272 157432 224284
rect 157484 224272 157490 224324
rect 161382 224272 161388 224324
rect 161440 224312 161446 224324
rect 176746 224312 176752 224324
rect 161440 224284 176752 224312
rect 161440 224272 161446 224284
rect 176746 224272 176752 224284
rect 176804 224272 176810 224324
rect 180702 224272 180708 224324
rect 180760 224312 180766 224324
rect 195974 224312 195980 224324
rect 180760 224284 195980 224312
rect 180760 224272 180766 224284
rect 195974 224272 195980 224284
rect 196032 224272 196038 224324
rect 112438 224204 112444 224256
rect 112496 224244 112502 224256
rect 123202 224244 123208 224256
rect 112496 224216 123208 224244
rect 112496 224204 112502 224216
rect 123202 224204 123208 224216
rect 123260 224204 123266 224256
rect 125226 224204 125232 224256
rect 125284 224244 125290 224256
rect 141418 224244 141424 224256
rect 125284 224216 141424 224244
rect 125284 224204 125290 224216
rect 141418 224204 141424 224216
rect 141476 224204 141482 224256
rect 150342 224204 150348 224256
rect 150400 224244 150406 224256
rect 166074 224244 166080 224256
rect 150400 224216 166080 224244
rect 150400 224204 150406 224216
rect 166074 224204 166080 224216
rect 166132 224204 166138 224256
rect 171042 224204 171048 224256
rect 171100 224244 171106 224256
rect 186314 224244 186320 224256
rect 171100 224216 186320 224244
rect 171100 224204 171106 224216
rect 186314 224204 186320 224216
rect 186372 224204 186378 224256
rect 188430 224204 188436 224256
rect 188488 224244 188494 224256
rect 203426 224244 203432 224256
rect 188488 224216 203432 224244
rect 188488 224204 188494 224216
rect 203426 224204 203432 224216
rect 203484 224204 203490 224256
rect 210970 224204 210976 224256
rect 211028 224244 211034 224256
rect 286318 224244 286324 224256
rect 211028 224216 286324 224244
rect 211028 224204 211034 224216
rect 286318 224204 286324 224216
rect 286376 224204 286382 224256
rect 139302 224176 139308 224188
rect 135916 224148 139308 224176
rect 126146 224068 126152 224120
rect 126204 224108 126210 224120
rect 134978 224108 134984 224120
rect 126204 224080 134984 224108
rect 126204 224068 126210 224080
rect 134978 224068 134984 224080
rect 135036 224068 135042 224120
rect 124122 224000 124128 224052
rect 124180 224040 124186 224052
rect 135916 224040 135944 224148
rect 139302 224136 139308 224148
rect 139360 224136 139366 224188
rect 139394 224136 139400 224188
rect 139452 224176 139458 224188
rect 148870 224176 148876 224188
rect 139452 224148 148876 224176
rect 139452 224136 139458 224148
rect 148870 224136 148876 224148
rect 148928 224136 148934 224188
rect 158622 224136 158628 224188
rect 158680 224176 158686 224188
rect 173526 224176 173532 224188
rect 158680 224148 173532 224176
rect 158680 224136 158686 224148
rect 173526 224136 173532 224148
rect 173584 224136 173590 224188
rect 173802 224136 173808 224188
rect 173860 224176 173866 224188
rect 188522 224176 188528 224188
rect 173860 224148 188528 224176
rect 173860 224136 173866 224148
rect 188522 224136 188528 224148
rect 188580 224136 188586 224188
rect 144638 224108 144644 224120
rect 124180 224012 135944 224040
rect 137296 224080 144644 224108
rect 124180 224000 124186 224012
rect 129642 223932 129648 223984
rect 129700 223972 129706 223984
rect 137296 223972 137324 224080
rect 144638 224068 144644 224080
rect 144696 224068 144702 224120
rect 157242 224068 157248 224120
rect 157300 224108 157306 224120
rect 172422 224108 172428 224120
rect 157300 224080 172428 224108
rect 157300 224068 157306 224080
rect 172422 224068 172428 224080
rect 172480 224068 172486 224120
rect 179322 224068 179328 224120
rect 179380 224108 179386 224120
rect 193858 224108 193864 224120
rect 179380 224080 193864 224108
rect 179380 224068 179386 224080
rect 193858 224068 193864 224080
rect 193916 224068 193922 224120
rect 141326 224000 141332 224052
rect 141384 224040 141390 224052
rect 155310 224040 155316 224052
rect 141384 224012 155316 224040
rect 141384 224000 141390 224012
rect 155310 224000 155316 224012
rect 155368 224000 155374 224052
rect 167638 224000 167644 224052
rect 167696 224040 167702 224052
rect 178862 224040 178868 224052
rect 167696 224012 178868 224040
rect 167696 224000 167702 224012
rect 178862 224000 178868 224012
rect 178920 224000 178926 224052
rect 184014 224000 184020 224052
rect 184072 224040 184078 224052
rect 189534 224040 189540 224052
rect 184072 224012 189540 224040
rect 184072 224000 184078 224012
rect 189534 224000 189540 224012
rect 189592 224000 189598 224052
rect 129700 223944 137324 223972
rect 129700 223932 129706 223944
rect 133690 223864 133696 223916
rect 133748 223904 133754 223916
rect 140314 223904 140320 223916
rect 133748 223876 140320 223904
rect 133748 223864 133754 223876
rect 140314 223864 140320 223876
rect 140372 223864 140378 223916
rect 229738 223592 229744 223644
rect 229796 223632 229802 223644
rect 283374 223632 283380 223644
rect 229796 223604 283380 223632
rect 229796 223592 229802 223604
rect 283374 223592 283380 223604
rect 283432 223592 283438 223644
rect 13078 222844 13084 222896
rect 13136 222884 13142 222896
rect 411898 222884 411904 222896
rect 13136 222856 411904 222884
rect 13136 222844 13142 222856
rect 411898 222844 411904 222856
rect 411956 222844 411962 222896
rect 231118 222436 231124 222488
rect 231176 222476 231182 222488
rect 235258 222476 235264 222488
rect 231176 222448 235264 222476
rect 231176 222436 231182 222448
rect 235258 222436 235264 222448
rect 235316 222436 235322 222488
rect 120718 221484 120724 221536
rect 120776 221484 120782 221536
rect 55214 220872 55220 220924
rect 55272 220912 55278 220924
rect 116394 220912 116400 220924
rect 55272 220884 116400 220912
rect 55272 220872 55278 220884
rect 116394 220872 116400 220884
rect 116452 220872 116458 220924
rect 9122 220804 9128 220856
rect 9180 220844 9186 220856
rect 120736 220844 120764 221484
rect 9180 220816 120764 220844
rect 9180 220804 9186 220816
rect 215110 220804 215116 220856
rect 215168 220844 215174 220856
rect 226334 220844 226340 220856
rect 215168 220816 226340 220844
rect 215168 220804 215174 220816
rect 226334 220804 226340 220816
rect 226392 220804 226398 220856
rect 215110 220124 215116 220176
rect 215168 220164 215174 220176
rect 226426 220164 226432 220176
rect 215168 220136 226432 220164
rect 215168 220124 215174 220136
rect 226426 220124 226432 220136
rect 226484 220124 226490 220176
rect 11698 220056 11704 220108
rect 11756 220096 11762 220108
rect 116670 220096 116676 220108
rect 11756 220068 116676 220096
rect 11756 220056 11762 220068
rect 116670 220056 116676 220068
rect 116728 220056 116734 220108
rect 215202 220056 215208 220108
rect 215260 220096 215266 220108
rect 226334 220096 226340 220108
rect 215260 220068 226340 220096
rect 215260 220056 215266 220068
rect 226334 220056 226340 220068
rect 226392 220056 226398 220108
rect 116118 219484 116124 219496
rect 114572 219456 116124 219484
rect 104802 219376 104808 219428
rect 104860 219416 104866 219428
rect 114572 219416 114600 219456
rect 116118 219444 116124 219456
rect 116176 219444 116182 219496
rect 104860 219388 114600 219416
rect 104860 219376 104866 219388
rect 215110 218764 215116 218816
rect 215168 218804 215174 218816
rect 226334 218804 226340 218816
rect 215168 218776 226340 218804
rect 215168 218764 215174 218776
rect 226334 218764 226340 218776
rect 226392 218764 226398 218816
rect 215202 218696 215208 218748
rect 215260 218736 215266 218748
rect 226426 218736 226432 218748
rect 215260 218708 226432 218736
rect 215260 218696 215266 218708
rect 226426 218696 226432 218708
rect 226484 218696 226490 218748
rect 116394 218056 116400 218068
rect 114480 218028 116400 218056
rect 104802 217948 104808 218000
rect 104860 217988 104866 218000
rect 114480 217988 114508 218028
rect 116394 218016 116400 218028
rect 116452 218016 116458 218068
rect 104860 217960 114508 217988
rect 104860 217948 104866 217960
rect 215110 217268 215116 217320
rect 215168 217308 215174 217320
rect 226334 217308 226340 217320
rect 215168 217280 226340 217308
rect 215168 217268 215174 217280
rect 226334 217268 226340 217280
rect 226392 217268 226398 217320
rect 116394 216696 116400 216708
rect 107672 216668 116400 216696
rect 104802 216588 104808 216640
rect 104860 216628 104866 216640
rect 107672 216628 107700 216668
rect 116394 216656 116400 216668
rect 116452 216656 116458 216708
rect 104860 216600 107700 216628
rect 104860 216588 104866 216600
rect 215110 216588 215116 216640
rect 215168 216628 215174 216640
rect 226426 216628 226432 216640
rect 215168 216600 226432 216628
rect 215168 216588 215174 216600
rect 226426 216588 226432 216600
rect 226484 216588 226490 216640
rect 104802 215908 104808 215960
rect 104860 215948 104866 215960
rect 115934 215948 115940 215960
rect 104860 215920 115940 215948
rect 104860 215908 104866 215920
rect 115934 215908 115940 215920
rect 115992 215908 115998 215960
rect 215110 215908 215116 215960
rect 215168 215948 215174 215960
rect 226334 215948 226340 215960
rect 215168 215920 226340 215948
rect 215168 215908 215174 215920
rect 226334 215908 226340 215920
rect 226392 215908 226398 215960
rect 116394 215336 116400 215348
rect 114480 215308 116400 215336
rect 104802 215228 104808 215280
rect 104860 215268 104866 215280
rect 114480 215268 114508 215308
rect 116394 215296 116400 215308
rect 116452 215296 116458 215348
rect 104860 215240 114508 215268
rect 104860 215228 104866 215240
rect 215110 215228 215116 215280
rect 215168 215268 215174 215280
rect 226426 215268 226432 215280
rect 215168 215240 226432 215268
rect 215168 215228 215174 215240
rect 226426 215228 226432 215240
rect 226484 215228 226490 215280
rect 215202 215160 215208 215212
rect 215260 215200 215266 215212
rect 226334 215200 226340 215212
rect 215260 215172 226340 215200
rect 215260 215160 215266 215172
rect 226334 215160 226340 215172
rect 226392 215160 226398 215212
rect 116394 213976 116400 213988
rect 113928 213948 116400 213976
rect 104802 213868 104808 213920
rect 104860 213908 104866 213920
rect 113928 213908 113956 213948
rect 116394 213936 116400 213948
rect 116452 213936 116458 213988
rect 104860 213880 113956 213908
rect 104860 213868 104866 213880
rect 215110 213868 215116 213920
rect 215168 213908 215174 213920
rect 226426 213908 226432 213920
rect 215168 213880 226432 213908
rect 215168 213868 215174 213880
rect 226426 213868 226432 213880
rect 226484 213868 226490 213920
rect 214374 213800 214380 213852
rect 214432 213840 214438 213852
rect 226334 213840 226340 213852
rect 214432 213812 226340 213840
rect 214432 213800 214438 213812
rect 226334 213800 226340 213812
rect 226392 213800 226398 213852
rect 115934 212548 115940 212560
rect 114480 212520 115940 212548
rect 104434 212440 104440 212492
rect 104492 212480 104498 212492
rect 114480 212480 114508 212520
rect 115934 212508 115940 212520
rect 115992 212508 115998 212560
rect 104492 212452 114508 212480
rect 104492 212440 104498 212452
rect 215110 212440 215116 212492
rect 215168 212480 215174 212492
rect 226426 212480 226432 212492
rect 215168 212452 226432 212480
rect 215168 212440 215174 212452
rect 226426 212440 226432 212452
rect 226484 212440 226490 212492
rect 215202 212372 215208 212424
rect 215260 212412 215266 212424
rect 226334 212412 226340 212424
rect 215260 212384 226340 212412
rect 215260 212372 215266 212384
rect 226334 212372 226340 212384
rect 226392 212372 226398 212424
rect 116302 211188 116308 211200
rect 114480 211160 116308 211188
rect 104802 211080 104808 211132
rect 104860 211120 104866 211132
rect 114480 211120 114508 211160
rect 116302 211148 116308 211160
rect 116360 211148 116366 211200
rect 104860 211092 114508 211120
rect 104860 211080 104866 211092
rect 214190 211080 214196 211132
rect 214248 211120 214254 211132
rect 226518 211120 226524 211132
rect 214248 211092 226524 211120
rect 214248 211080 214254 211092
rect 226518 211080 226524 211092
rect 226576 211080 226582 211132
rect 116302 209828 116308 209840
rect 113192 209800 116308 209828
rect 104802 209720 104808 209772
rect 104860 209760 104866 209772
rect 113192 209760 113220 209800
rect 116302 209788 116308 209800
rect 116360 209788 116366 209840
rect 104860 209732 113220 209760
rect 104860 209720 104866 209732
rect 215110 209720 215116 209772
rect 215168 209760 215174 209772
rect 226150 209760 226156 209772
rect 215168 209732 226156 209760
rect 215168 209720 215174 209732
rect 226150 209720 226156 209732
rect 226208 209720 226214 209772
rect 214190 209652 214196 209704
rect 214248 209692 214254 209704
rect 226242 209692 226248 209704
rect 214248 209664 226248 209692
rect 214248 209652 214254 209664
rect 226242 209652 226248 209664
rect 226300 209652 226306 209704
rect 116026 208400 116032 208412
rect 114480 208372 116032 208400
rect 104802 208292 104808 208344
rect 104860 208332 104866 208344
rect 114480 208332 114508 208372
rect 116026 208360 116032 208372
rect 116084 208360 116090 208412
rect 104860 208304 114508 208332
rect 104860 208292 104866 208304
rect 215110 208292 215116 208344
rect 215168 208332 215174 208344
rect 226058 208332 226064 208344
rect 215168 208304 226064 208332
rect 215168 208292 215174 208304
rect 226058 208292 226064 208304
rect 226116 208292 226122 208344
rect 214282 208224 214288 208276
rect 214340 208264 214346 208276
rect 225966 208264 225972 208276
rect 214340 208236 225972 208264
rect 214340 208224 214346 208236
rect 225966 208224 225972 208236
rect 226024 208224 226030 208276
rect 113082 207068 113088 207120
rect 113140 207108 113146 207120
rect 116026 207108 116032 207120
rect 113140 207080 116032 207108
rect 113140 207068 113146 207080
rect 116026 207068 116032 207080
rect 116084 207068 116090 207120
rect 115934 207040 115940 207052
rect 114480 207012 115940 207040
rect 104802 206864 104808 206916
rect 104860 206904 104866 206916
rect 114480 206904 114508 207012
rect 115934 207000 115940 207012
rect 115992 207000 115998 207052
rect 215110 206932 215116 206984
rect 215168 206972 215174 206984
rect 226058 206972 226064 206984
rect 215168 206944 226064 206972
rect 215168 206932 215174 206944
rect 226058 206932 226064 206944
rect 226116 206932 226122 206984
rect 104860 206876 114508 206904
rect 104860 206864 104866 206876
rect 214374 206864 214380 206916
rect 214432 206904 214438 206916
rect 226242 206904 226248 206916
rect 214432 206876 226248 206904
rect 214432 206864 214438 206876
rect 226242 206864 226248 206876
rect 226300 206864 226306 206916
rect 104710 206796 104716 206848
rect 104768 206836 104774 206848
rect 113082 206836 113088 206848
rect 104768 206808 113088 206836
rect 104768 206796 104774 206808
rect 113082 206796 113088 206808
rect 113140 206796 113146 206848
rect 115934 205680 115940 205692
rect 114480 205652 115940 205680
rect 104802 205572 104808 205624
rect 104860 205612 104866 205624
rect 114480 205612 114508 205652
rect 115934 205640 115940 205652
rect 115992 205640 115998 205692
rect 104860 205584 114508 205612
rect 104860 205572 104866 205584
rect 215110 205572 215116 205624
rect 215168 205612 215174 205624
rect 226150 205612 226156 205624
rect 215168 205584 226156 205612
rect 215168 205572 215174 205584
rect 226150 205572 226156 205584
rect 226208 205572 226214 205624
rect 116394 204320 116400 204332
rect 114480 204292 116400 204320
rect 104802 204212 104808 204264
rect 104860 204252 104866 204264
rect 114480 204252 114508 204292
rect 116394 204280 116400 204292
rect 116452 204280 116458 204332
rect 104860 204224 114508 204252
rect 104860 204212 104866 204224
rect 215202 204212 215208 204264
rect 215260 204252 215266 204264
rect 225966 204252 225972 204264
rect 215260 204224 225972 204252
rect 215260 204212 215266 204224
rect 225966 204212 225972 204224
rect 226024 204212 226030 204264
rect 215110 204144 215116 204196
rect 215168 204184 215174 204196
rect 225874 204184 225880 204196
rect 215168 204156 225880 204184
rect 215168 204144 215174 204156
rect 225874 204144 225880 204156
rect 225932 204144 225938 204196
rect 116302 202892 116308 202904
rect 114480 202864 116308 202892
rect 104802 202784 104808 202836
rect 104860 202824 104866 202836
rect 114480 202824 114508 202864
rect 116302 202852 116308 202864
rect 116360 202852 116366 202904
rect 104860 202796 114508 202824
rect 104860 202784 104866 202796
rect 214282 202784 214288 202836
rect 214340 202824 214346 202836
rect 226058 202824 226064 202836
rect 214340 202796 226064 202824
rect 214340 202784 214346 202796
rect 226058 202784 226064 202796
rect 226116 202784 226122 202836
rect 215110 202716 215116 202768
rect 215168 202756 215174 202768
rect 225782 202756 225788 202768
rect 215168 202728 225788 202756
rect 215168 202716 215174 202728
rect 225782 202716 225788 202728
rect 225840 202716 225846 202768
rect 116118 201532 116124 201544
rect 114480 201504 116124 201532
rect 104802 201424 104808 201476
rect 104860 201464 104866 201476
rect 114480 201464 114508 201504
rect 116118 201492 116124 201504
rect 116176 201492 116182 201544
rect 104860 201436 114508 201464
rect 104860 201424 104866 201436
rect 214374 201424 214380 201476
rect 214432 201464 214438 201476
rect 225598 201464 225604 201476
rect 214432 201436 225604 201464
rect 214432 201424 214438 201436
rect 225598 201424 225604 201436
rect 225656 201424 225662 201476
rect 215110 201356 215116 201408
rect 215168 201396 215174 201408
rect 226058 201396 226064 201408
rect 215168 201368 226064 201396
rect 215168 201356 215174 201368
rect 226058 201356 226064 201368
rect 226116 201356 226122 201408
rect 116118 200240 116124 200252
rect 113192 200212 116124 200240
rect 104802 200064 104808 200116
rect 104860 200104 104866 200116
rect 113192 200104 113220 200212
rect 116118 200200 116124 200212
rect 116176 200200 116182 200252
rect 113266 200132 113272 200184
rect 113324 200172 113330 200184
rect 115934 200172 115940 200184
rect 113324 200144 115940 200172
rect 113324 200132 113330 200144
rect 115934 200132 115940 200144
rect 115992 200132 115998 200184
rect 104860 200076 113220 200104
rect 104860 200064 104866 200076
rect 214098 200064 214104 200116
rect 214156 200104 214162 200116
rect 226242 200104 226248 200116
rect 214156 200076 226248 200104
rect 214156 200064 214162 200076
rect 226242 200064 226248 200076
rect 226300 200064 226306 200116
rect 224034 198772 224040 198824
rect 224092 198812 224098 198824
rect 226426 198812 226432 198824
rect 224092 198784 226432 198812
rect 224092 198772 224098 198784
rect 226426 198772 226432 198784
rect 226484 198772 226490 198824
rect 113174 198704 113180 198756
rect 113232 198744 113238 198756
rect 116394 198744 116400 198756
rect 113232 198716 116400 198744
rect 113232 198704 113238 198716
rect 116394 198704 116400 198716
rect 116452 198704 116458 198756
rect 224126 198704 224132 198756
rect 224184 198744 224190 198756
rect 226334 198744 226340 198756
rect 224184 198716 226340 198744
rect 224184 198704 224190 198716
rect 226334 198704 226340 198716
rect 226392 198704 226398 198756
rect 104802 198636 104808 198688
rect 104860 198676 104866 198688
rect 113266 198676 113272 198688
rect 104860 198648 113272 198676
rect 104860 198636 104866 198648
rect 113266 198636 113272 198648
rect 113324 198636 113330 198688
rect 215110 198636 215116 198688
rect 215168 198676 215174 198688
rect 225966 198676 225972 198688
rect 215168 198648 225972 198676
rect 215168 198636 215174 198648
rect 225966 198636 225972 198648
rect 226024 198636 226030 198688
rect 214098 198568 214104 198620
rect 214156 198608 214162 198620
rect 225690 198608 225696 198620
rect 214156 198580 225696 198608
rect 214156 198568 214162 198580
rect 225690 198568 225696 198580
rect 225748 198568 225754 198620
rect 223942 197412 223948 197464
rect 224000 197452 224006 197464
rect 226426 197452 226432 197464
rect 224000 197424 226432 197452
rect 224000 197412 224006 197424
rect 226426 197412 226432 197424
rect 226484 197412 226490 197464
rect 116394 197384 116400 197396
rect 114480 197356 116400 197384
rect 104802 197276 104808 197328
rect 104860 197316 104866 197328
rect 113082 197316 113088 197328
rect 104860 197288 113088 197316
rect 104860 197276 104866 197288
rect 113082 197276 113088 197288
rect 113140 197276 113146 197328
rect 104526 197208 104532 197260
rect 104584 197248 104590 197260
rect 114480 197248 114508 197356
rect 116394 197344 116400 197356
rect 116452 197344 116458 197396
rect 224310 197344 224316 197396
rect 224368 197384 224374 197396
rect 226334 197384 226340 197396
rect 224368 197356 226340 197384
rect 224368 197344 224374 197356
rect 226334 197344 226340 197356
rect 226392 197344 226398 197396
rect 214374 197276 214380 197328
rect 214432 197316 214438 197328
rect 226150 197316 226156 197328
rect 214432 197288 226156 197316
rect 214432 197276 214438 197288
rect 226150 197276 226156 197288
rect 226208 197276 226214 197328
rect 104584 197220 114508 197248
rect 104584 197208 104590 197220
rect 215110 197208 215116 197260
rect 215168 197248 215174 197260
rect 225874 197248 225880 197260
rect 215168 197220 225880 197248
rect 215168 197208 215174 197220
rect 225874 197208 225880 197220
rect 225932 197208 225938 197260
rect 224218 196052 224224 196104
rect 224276 196092 224282 196104
rect 226610 196092 226616 196104
rect 224276 196064 226616 196092
rect 224276 196052 224282 196064
rect 226610 196052 226616 196064
rect 226668 196052 226674 196104
rect 116394 196024 116400 196036
rect 114296 195996 116400 196024
rect 104802 195916 104808 195968
rect 104860 195956 104866 195968
rect 114296 195956 114324 195996
rect 116394 195984 116400 195996
rect 116452 195984 116458 196036
rect 224586 195984 224592 196036
rect 224644 196024 224650 196036
rect 226702 196024 226708 196036
rect 224644 195996 226708 196024
rect 224644 195984 224650 195996
rect 226702 195984 226708 195996
rect 226760 195984 226766 196036
rect 104860 195928 114324 195956
rect 104860 195916 104866 195928
rect 215202 195916 215208 195968
rect 215260 195956 215266 195968
rect 226058 195956 226064 195968
rect 215260 195928 226064 195956
rect 215260 195916 215266 195928
rect 226058 195916 226064 195928
rect 226116 195916 226122 195968
rect 215110 195848 215116 195900
rect 215168 195888 215174 195900
rect 226242 195888 226248 195900
rect 215168 195860 226248 195888
rect 215168 195848 215174 195860
rect 226242 195848 226248 195860
rect 226300 195848 226306 195900
rect 115934 194596 115940 194608
rect 114480 194568 115940 194596
rect 104802 194488 104808 194540
rect 104860 194528 104866 194540
rect 114480 194528 114508 194568
rect 115934 194556 115940 194568
rect 115992 194556 115998 194608
rect 224402 194556 224408 194608
rect 224460 194596 224466 194608
rect 226334 194596 226340 194608
rect 224460 194568 226340 194596
rect 224460 194556 224466 194568
rect 226334 194556 226340 194568
rect 226392 194556 226398 194608
rect 104860 194500 114508 194528
rect 104860 194488 104866 194500
rect 215110 194488 215116 194540
rect 215168 194528 215174 194540
rect 225782 194528 225788 194540
rect 215168 194500 225788 194528
rect 215168 194488 215174 194500
rect 225782 194488 225788 194500
rect 225840 194488 225846 194540
rect 220262 193264 220268 193316
rect 220320 193304 220326 193316
rect 226426 193304 226432 193316
rect 220320 193276 226432 193304
rect 220320 193264 220326 193276
rect 226426 193264 226432 193276
rect 226484 193264 226490 193316
rect 116118 193236 116124 193248
rect 114480 193208 116124 193236
rect 104434 193128 104440 193180
rect 104492 193168 104498 193180
rect 114480 193168 114508 193208
rect 116118 193196 116124 193208
rect 116176 193196 116182 193248
rect 215938 193196 215944 193248
rect 215996 193236 216002 193248
rect 226334 193236 226340 193248
rect 215996 193208 226340 193236
rect 215996 193196 216002 193208
rect 226334 193196 226340 193208
rect 226392 193196 226398 193248
rect 104492 193140 114508 193168
rect 104492 193128 104498 193140
rect 215110 193128 215116 193180
rect 215168 193168 215174 193180
rect 224034 193168 224040 193180
rect 215168 193140 224040 193168
rect 215168 193128 215174 193140
rect 224034 193128 224040 193140
rect 224092 193128 224098 193180
rect 215202 193060 215208 193112
rect 215260 193100 215266 193112
rect 224126 193100 224132 193112
rect 215260 193072 224132 193100
rect 215260 193060 215266 193072
rect 224126 193060 224132 193072
rect 224184 193060 224190 193112
rect 113174 191972 113180 192024
rect 113232 192012 113238 192024
rect 116394 192012 116400 192024
rect 113232 191984 116400 192012
rect 113232 191972 113238 191984
rect 116394 191972 116400 191984
rect 116452 191972 116458 192024
rect 113266 191904 113272 191956
rect 113324 191944 113330 191956
rect 116026 191944 116032 191956
rect 113324 191916 116032 191944
rect 113324 191904 113330 191916
rect 116026 191904 116032 191916
rect 116084 191904 116090 191956
rect 224862 191904 224868 191956
rect 224920 191944 224926 191956
rect 226426 191944 226432 191956
rect 224920 191916 226432 191944
rect 224920 191904 224926 191916
rect 226426 191904 226432 191916
rect 226484 191904 226490 191956
rect 218146 191836 218152 191888
rect 218204 191876 218210 191888
rect 226334 191876 226340 191888
rect 218204 191848 226340 191876
rect 218204 191836 218210 191848
rect 226334 191836 226340 191848
rect 226392 191836 226398 191888
rect 104802 191768 104808 191820
rect 104860 191808 104866 191820
rect 113174 191808 113180 191820
rect 104860 191780 113180 191808
rect 104860 191768 104866 191780
rect 113174 191768 113180 191780
rect 113232 191768 113238 191820
rect 214282 191768 214288 191820
rect 214340 191808 214346 191820
rect 224310 191808 224316 191820
rect 214340 191780 224316 191808
rect 214340 191768 214346 191780
rect 224310 191768 224316 191780
rect 224368 191768 224374 191820
rect 215110 191700 215116 191752
rect 215168 191740 215174 191752
rect 223942 191740 223948 191752
rect 215168 191712 223948 191740
rect 215168 191700 215174 191712
rect 223942 191700 223948 191712
rect 224000 191700 224006 191752
rect 215294 191088 215300 191140
rect 215352 191128 215358 191140
rect 226610 191128 226616 191140
rect 215352 191100 226616 191128
rect 215352 191088 215358 191100
rect 226610 191088 226616 191100
rect 226668 191088 226674 191140
rect 221458 190884 221464 190936
rect 221516 190924 221522 190936
rect 226334 190924 226340 190936
rect 221516 190896 226340 190924
rect 221516 190884 221522 190896
rect 226334 190884 226340 190896
rect 226392 190884 226398 190936
rect 113358 190612 113364 190664
rect 113416 190652 113422 190664
rect 116486 190652 116492 190664
rect 113416 190624 116492 190652
rect 113416 190612 113422 190624
rect 116486 190612 116492 190624
rect 116544 190612 116550 190664
rect 222838 190476 222844 190528
rect 222896 190516 222902 190528
rect 226334 190516 226340 190528
rect 222896 190488 226340 190516
rect 222896 190476 222902 190488
rect 226334 190476 226340 190488
rect 226392 190476 226398 190528
rect 104710 190408 104716 190460
rect 104768 190448 104774 190460
rect 113266 190448 113272 190460
rect 104768 190420 113272 190448
rect 104768 190408 104774 190420
rect 113266 190408 113272 190420
rect 113324 190408 113330 190460
rect 214374 190408 214380 190460
rect 214432 190448 214438 190460
rect 224586 190448 224592 190460
rect 214432 190420 224592 190448
rect 214432 190408 214438 190420
rect 224586 190408 224592 190420
rect 224644 190408 224650 190460
rect 215110 190340 215116 190392
rect 215168 190380 215174 190392
rect 224218 190380 224224 190392
rect 215168 190352 224224 190380
rect 215168 190340 215174 190352
rect 224218 190340 224224 190352
rect 224276 190340 224282 190392
rect 218054 189728 218060 189780
rect 218112 189768 218118 189780
rect 226978 189768 226984 189780
rect 218112 189740 226984 189768
rect 218112 189728 218118 189740
rect 226978 189728 226984 189740
rect 227036 189728 227042 189780
rect 114186 189048 114192 189100
rect 114244 189088 114250 189100
rect 116394 189088 116400 189100
rect 114244 189060 116400 189088
rect 114244 189048 114250 189060
rect 116394 189048 116400 189060
rect 116452 189048 116458 189100
rect 220078 189048 220084 189100
rect 220136 189088 220142 189100
rect 226334 189088 226340 189100
rect 220136 189060 226340 189088
rect 220136 189048 220142 189060
rect 226334 189048 226340 189060
rect 226392 189048 226398 189100
rect 104802 188980 104808 189032
rect 104860 189020 104866 189032
rect 113358 189020 113364 189032
rect 104860 188992 113364 189020
rect 104860 188980 104866 188992
rect 113358 188980 113364 188992
rect 113416 188980 113422 189032
rect 214006 188980 214012 189032
rect 214064 189020 214070 189032
rect 224402 189020 224408 189032
rect 214064 188992 224408 189020
rect 214064 188980 214070 188992
rect 224402 188980 224408 188992
rect 224460 188980 224466 189032
rect 221642 187756 221648 187808
rect 221700 187796 221706 187808
rect 226426 187796 226432 187808
rect 221700 187768 226432 187796
rect 221700 187756 221706 187768
rect 226426 187756 226432 187768
rect 226484 187756 226490 187808
rect 113174 187688 113180 187740
rect 113232 187728 113238 187740
rect 116210 187728 116216 187740
rect 113232 187700 116216 187728
rect 113232 187688 113238 187700
rect 116210 187688 116216 187700
rect 116268 187688 116274 187740
rect 216030 187688 216036 187740
rect 216088 187728 216094 187740
rect 226334 187728 226340 187740
rect 216088 187700 226340 187728
rect 216088 187688 216094 187700
rect 226334 187688 226340 187700
rect 226392 187688 226398 187740
rect 104802 187620 104808 187672
rect 104860 187660 104866 187672
rect 114186 187660 114192 187672
rect 104860 187632 114192 187660
rect 104860 187620 104866 187632
rect 114186 187620 114192 187632
rect 114244 187620 114250 187672
rect 215110 187552 215116 187604
rect 215168 187592 215174 187604
rect 220262 187592 220268 187604
rect 215168 187564 220268 187592
rect 215168 187552 215174 187564
rect 220262 187552 220268 187564
rect 220320 187552 220326 187604
rect 215202 187144 215208 187196
rect 215260 187184 215266 187196
rect 218054 187184 218060 187196
rect 215260 187156 218060 187184
rect 215260 187144 215266 187156
rect 218054 187144 218060 187156
rect 218112 187144 218118 187196
rect 218790 186464 218796 186516
rect 218848 186504 218854 186516
rect 226334 186504 226340 186516
rect 218848 186476 226340 186504
rect 218848 186464 218854 186476
rect 226334 186464 226340 186476
rect 226392 186464 226398 186516
rect 116302 186368 116308 186380
rect 114480 186340 116308 186368
rect 104802 186260 104808 186312
rect 104860 186300 104866 186312
rect 113082 186300 113088 186312
rect 104860 186272 113088 186300
rect 104860 186260 104866 186272
rect 113082 186260 113088 186272
rect 113140 186260 113146 186312
rect 104526 186192 104532 186244
rect 104584 186232 104590 186244
rect 114480 186232 114508 186340
rect 116302 186328 116308 186340
rect 116360 186328 116366 186380
rect 220170 186328 220176 186380
rect 220228 186368 220234 186380
rect 226334 186368 226340 186380
rect 220228 186340 226340 186368
rect 220228 186328 220234 186340
rect 226334 186328 226340 186340
rect 226392 186328 226398 186380
rect 104584 186204 114508 186232
rect 104584 186192 104590 186204
rect 214466 185648 214472 185700
rect 214524 185688 214530 185700
rect 224862 185688 224868 185700
rect 214524 185660 224868 185688
rect 214524 185648 214530 185660
rect 224862 185648 224868 185660
rect 224920 185648 224926 185700
rect 215294 185580 215300 185632
rect 215352 185620 215358 185632
rect 226518 185620 226524 185632
rect 215352 185592 226524 185620
rect 215352 185580 215358 185592
rect 226518 185580 226524 185592
rect 226576 185580 226582 185632
rect 213914 185512 213920 185564
rect 213972 185552 213978 185564
rect 215938 185552 215944 185564
rect 213972 185524 215944 185552
rect 213972 185512 213978 185524
rect 215938 185512 215944 185524
rect 215996 185512 216002 185564
rect 114462 184968 114468 185020
rect 114520 185008 114526 185020
rect 116394 185008 116400 185020
rect 114520 184980 116400 185008
rect 114520 184968 114526 184980
rect 116394 184968 116400 184980
rect 116452 184968 116458 185020
rect 116026 184940 116032 184952
rect 114480 184912 116032 184940
rect 104802 184832 104808 184884
rect 104860 184872 104866 184884
rect 114480 184872 114508 184912
rect 116026 184900 116032 184912
rect 116084 184900 116090 184952
rect 224218 184900 224224 184952
rect 224276 184940 224282 184952
rect 226334 184940 226340 184952
rect 224276 184912 226340 184940
rect 224276 184900 224282 184912
rect 226334 184900 226340 184912
rect 226392 184900 226398 184952
rect 104860 184844 114508 184872
rect 104860 184832 104866 184844
rect 227162 184832 227168 184884
rect 227220 184872 227226 184884
rect 230842 184872 230848 184884
rect 227220 184844 230848 184872
rect 227220 184832 227226 184844
rect 230842 184832 230848 184844
rect 230900 184832 230906 184884
rect 214190 184764 214196 184816
rect 214248 184804 214254 184816
rect 218146 184804 218152 184816
rect 214248 184776 218152 184804
rect 214248 184764 214254 184776
rect 218146 184764 218152 184776
rect 218204 184764 218210 184816
rect 224310 183608 224316 183660
rect 224368 183648 224374 183660
rect 226518 183648 226524 183660
rect 224368 183620 226524 183648
rect 224368 183608 224374 183620
rect 226518 183608 226524 183620
rect 226576 183608 226582 183660
rect 114370 183540 114376 183592
rect 114428 183580 114434 183592
rect 116394 183580 116400 183592
rect 114428 183552 116400 183580
rect 114428 183540 114434 183552
rect 116394 183540 116400 183552
rect 116452 183540 116458 183592
rect 215018 183540 215024 183592
rect 215076 183580 215082 183592
rect 226334 183580 226340 183592
rect 215076 183552 226340 183580
rect 215076 183540 215082 183552
rect 226334 183540 226340 183552
rect 226392 183540 226398 183592
rect 104802 183472 104808 183524
rect 104860 183512 104866 183524
rect 114462 183512 114468 183524
rect 104860 183484 114468 183512
rect 104860 183472 104866 183484
rect 114462 183472 114468 183484
rect 114520 183472 114526 183524
rect 215110 182520 215116 182572
rect 215168 182560 215174 182572
rect 221458 182560 221464 182572
rect 215168 182532 221464 182560
rect 215168 182520 215174 182532
rect 221458 182520 221464 182532
rect 221516 182520 221522 182572
rect 222930 182248 222936 182300
rect 222988 182288 222994 182300
rect 226518 182288 226524 182300
rect 222988 182260 226524 182288
rect 222988 182248 222994 182260
rect 226518 182248 226524 182260
rect 226576 182248 226582 182300
rect 113174 182180 113180 182232
rect 113232 182220 113238 182232
rect 115934 182220 115940 182232
rect 113232 182192 115940 182220
rect 113232 182180 113238 182192
rect 115934 182180 115940 182192
rect 115992 182180 115998 182232
rect 214834 182180 214840 182232
rect 214892 182220 214898 182232
rect 226334 182220 226340 182232
rect 214892 182192 226340 182220
rect 214892 182180 214898 182192
rect 226334 182180 226340 182192
rect 226392 182180 226398 182232
rect 104802 182112 104808 182164
rect 104860 182152 104866 182164
rect 114370 182152 114376 182164
rect 104860 182124 114376 182152
rect 104860 182112 104866 182124
rect 114370 182112 114376 182124
rect 114428 182112 114434 182164
rect 214190 182112 214196 182164
rect 214248 182152 214254 182164
rect 222838 182152 222844 182164
rect 214248 182124 222844 182152
rect 214248 182112 214254 182124
rect 222838 182112 222844 182124
rect 222896 182112 222902 182164
rect 335998 182112 336004 182164
rect 336056 182152 336062 182164
rect 579982 182152 579988 182164
rect 336056 182124 579988 182152
rect 336056 182112 336062 182124
rect 579982 182112 579988 182124
rect 580040 182112 580046 182164
rect 218882 181432 218888 181484
rect 218940 181472 218946 181484
rect 226426 181472 226432 181484
rect 218940 181444 226432 181472
rect 218940 181432 218946 181444
rect 226426 181432 226432 181444
rect 226484 181432 226490 181484
rect 113266 181092 113272 181144
rect 113324 181132 113330 181144
rect 115934 181132 115940 181144
rect 113324 181104 115940 181132
rect 113324 181092 113330 181104
rect 115934 181092 115940 181104
rect 115992 181092 115998 181144
rect 221550 180888 221556 180940
rect 221608 180928 221614 180940
rect 226334 180928 226340 180940
rect 221608 180900 226340 180928
rect 221608 180888 221614 180900
rect 226334 180888 226340 180900
rect 226392 180888 226398 180940
rect 104802 180752 104808 180804
rect 104860 180792 104866 180804
rect 113174 180792 113180 180804
rect 104860 180764 113180 180792
rect 104860 180752 104866 180764
rect 113174 180752 113180 180764
rect 113232 180752 113238 180804
rect 214006 180752 214012 180804
rect 214064 180792 214070 180804
rect 225782 180792 225788 180804
rect 214064 180764 225788 180792
rect 214064 180752 214070 180764
rect 225782 180752 225788 180764
rect 225840 180752 225846 180804
rect 214098 179732 214104 179784
rect 214156 179772 214162 179784
rect 220078 179772 220084 179784
rect 214156 179744 220084 179772
rect 214156 179732 214162 179744
rect 220078 179732 220084 179744
rect 220136 179732 220142 179784
rect 221458 179460 221464 179512
rect 221516 179500 221522 179512
rect 226426 179500 226432 179512
rect 221516 179472 226432 179500
rect 221516 179460 221522 179472
rect 226426 179460 226432 179472
rect 226484 179460 226490 179512
rect 113910 179392 113916 179444
rect 113968 179432 113974 179444
rect 116394 179432 116400 179444
rect 113968 179404 116400 179432
rect 113968 179392 113974 179404
rect 116394 179392 116400 179404
rect 116452 179392 116458 179444
rect 225690 179392 225696 179444
rect 225748 179432 225754 179444
rect 227622 179432 227628 179444
rect 225748 179404 227628 179432
rect 225748 179392 225754 179404
rect 227622 179392 227628 179404
rect 227680 179392 227686 179444
rect 104802 179324 104808 179376
rect 104860 179364 104866 179376
rect 113266 179364 113272 179376
rect 104860 179336 113272 179364
rect 104860 179324 104866 179336
rect 113266 179324 113272 179336
rect 113324 179324 113330 179376
rect 213914 179188 213920 179240
rect 213972 179228 213978 179240
rect 216030 179228 216036 179240
rect 213972 179200 216036 179228
rect 213972 179188 213978 179200
rect 216030 179188 216036 179200
rect 216088 179188 216094 179240
rect 215938 178644 215944 178696
rect 215996 178684 216002 178696
rect 226334 178684 226340 178696
rect 215996 178656 226340 178684
rect 215996 178644 216002 178656
rect 226334 178644 226340 178656
rect 226392 178644 226398 178696
rect 214098 178576 214104 178628
rect 214156 178616 214162 178628
rect 221642 178616 221648 178628
rect 214156 178588 221648 178616
rect 214156 178576 214162 178588
rect 221642 178576 221648 178588
rect 221700 178576 221706 178628
rect 114186 178032 114192 178084
rect 114244 178072 114250 178084
rect 115934 178072 115940 178084
rect 114244 178044 115940 178072
rect 114244 178032 114250 178044
rect 115934 178032 115940 178044
rect 115992 178032 115998 178084
rect 220078 178032 220084 178084
rect 220136 178072 220142 178084
rect 226426 178072 226432 178084
rect 220136 178044 226432 178072
rect 220136 178032 220142 178044
rect 226426 178032 226432 178044
rect 226484 178032 226490 178084
rect 104158 177964 104164 178016
rect 104216 178004 104222 178016
rect 113910 178004 113916 178016
rect 104216 177976 113916 178004
rect 104216 177964 104222 177976
rect 113910 177964 113916 177976
rect 113968 177964 113974 178016
rect 224954 177964 224960 178016
rect 225012 178004 225018 178016
rect 226978 178004 226984 178016
rect 225012 177976 226984 178004
rect 225012 177964 225018 177976
rect 226978 177964 226984 177976
rect 227036 177964 227042 178016
rect 215018 177488 215024 177540
rect 215076 177528 215082 177540
rect 218790 177528 218796 177540
rect 215076 177500 218796 177528
rect 215076 177488 215082 177500
rect 218790 177488 218796 177500
rect 218848 177488 218854 177540
rect 113910 176740 113916 176792
rect 113968 176780 113974 176792
rect 115934 176780 115940 176792
rect 113968 176752 115940 176780
rect 113968 176740 113974 176752
rect 115934 176740 115940 176752
rect 115992 176740 115998 176792
rect 114462 176672 114468 176724
rect 114520 176712 114526 176724
rect 116394 176712 116400 176724
rect 114520 176684 116400 176712
rect 114520 176672 114526 176684
rect 116394 176672 116400 176684
rect 116452 176672 116458 176724
rect 218698 176672 218704 176724
rect 218756 176712 218762 176724
rect 226334 176712 226340 176724
rect 218756 176684 226340 176712
rect 218756 176672 218762 176684
rect 226334 176672 226340 176684
rect 226392 176672 226398 176724
rect 104158 176604 104164 176656
rect 104216 176644 104222 176656
rect 114186 176644 114192 176656
rect 104216 176616 114192 176644
rect 104216 176604 104222 176616
rect 114186 176604 114192 176616
rect 114244 176604 114250 176656
rect 215110 176604 215116 176656
rect 215168 176644 215174 176656
rect 225598 176644 225604 176656
rect 215168 176616 225604 176644
rect 215168 176604 215174 176616
rect 225598 176604 225604 176616
rect 225656 176604 225662 176656
rect 215110 176128 215116 176180
rect 215168 176168 215174 176180
rect 220170 176168 220176 176180
rect 215168 176140 220176 176168
rect 215168 176128 215174 176140
rect 220170 176128 220176 176140
rect 220228 176128 220234 176180
rect 220262 175584 220268 175636
rect 220320 175624 220326 175636
rect 227162 175624 227168 175636
rect 220320 175596 227168 175624
rect 220320 175584 220326 175596
rect 227162 175584 227168 175596
rect 227220 175584 227226 175636
rect 114278 175244 114284 175296
rect 114336 175284 114342 175296
rect 116394 175284 116400 175296
rect 114336 175256 116400 175284
rect 114336 175244 114342 175256
rect 116394 175244 116400 175256
rect 116452 175244 116458 175296
rect 222838 175244 222844 175296
rect 222896 175284 222902 175296
rect 227438 175284 227444 175296
rect 222896 175256 227444 175284
rect 222896 175244 222902 175256
rect 227438 175244 227444 175256
rect 227496 175244 227502 175296
rect 104434 175176 104440 175228
rect 104492 175216 104498 175228
rect 114462 175216 114468 175228
rect 104492 175188 114468 175216
rect 104492 175176 104498 175188
rect 114462 175176 114468 175188
rect 114520 175176 114526 175228
rect 214098 175176 214104 175228
rect 214156 175216 214162 175228
rect 224954 175216 224960 175228
rect 214156 175188 224960 175216
rect 214156 175176 214162 175188
rect 224954 175176 224960 175188
rect 225012 175176 225018 175228
rect 104802 175108 104808 175160
rect 104860 175148 104866 175160
rect 113910 175148 113916 175160
rect 104860 175120 113916 175148
rect 104860 175108 104866 175120
rect 113910 175108 113916 175120
rect 113968 175108 113974 175160
rect 215110 175108 215116 175160
rect 215168 175148 215174 175160
rect 224218 175148 224224 175160
rect 215168 175120 224224 175148
rect 215168 175108 215174 175120
rect 224218 175108 224224 175120
rect 224276 175108 224282 175160
rect 114370 173884 114376 173936
rect 114428 173924 114434 173936
rect 115934 173924 115940 173936
rect 114428 173896 115940 173924
rect 114428 173884 114434 173896
rect 115934 173884 115940 173896
rect 115992 173884 115998 173936
rect 225598 173884 225604 173936
rect 225656 173924 225662 173936
rect 227346 173924 227352 173936
rect 225656 173896 227352 173924
rect 225656 173884 225662 173896
rect 227346 173884 227352 173896
rect 227404 173884 227410 173936
rect 104802 173816 104808 173868
rect 104860 173856 104866 173868
rect 114278 173856 114284 173868
rect 104860 173828 114284 173856
rect 104860 173816 104866 173828
rect 114278 173816 114284 173828
rect 114336 173816 114342 173868
rect 214282 173816 214288 173868
rect 214340 173856 214346 173868
rect 224310 173856 224316 173868
rect 214340 173828 224316 173856
rect 214340 173816 214346 173828
rect 224310 173816 224316 173828
rect 224368 173816 224374 173868
rect 224310 173272 224316 173324
rect 224368 173312 224374 173324
rect 226702 173312 226708 173324
rect 224368 173284 226708 173312
rect 224368 173272 224374 173284
rect 226702 173272 226708 173284
rect 226760 173272 226766 173324
rect 113174 172524 113180 172576
rect 113232 172564 113238 172576
rect 116394 172564 116400 172576
rect 113232 172536 116400 172564
rect 113232 172524 113238 172536
rect 116394 172524 116400 172536
rect 116452 172524 116458 172576
rect 104434 172456 104440 172508
rect 104492 172496 104498 172508
rect 114370 172496 114376 172508
rect 104492 172468 114376 172496
rect 104492 172456 104498 172468
rect 114370 172456 114376 172468
rect 114428 172456 114434 172508
rect 214282 172456 214288 172508
rect 214340 172496 214346 172508
rect 222930 172496 222936 172508
rect 214340 172468 222936 172496
rect 214340 172456 214346 172468
rect 222930 172456 222936 172468
rect 222988 172456 222994 172508
rect 215018 171980 215024 172032
rect 215076 172020 215082 172032
rect 218882 172020 218888 172032
rect 215076 171992 218888 172020
rect 215076 171980 215082 171992
rect 218882 171980 218888 171992
rect 218940 171980 218946 172032
rect 113266 171572 113272 171624
rect 113324 171612 113330 171624
rect 116118 171612 116124 171624
rect 113324 171584 116124 171612
rect 113324 171572 113330 171584
rect 116118 171572 116124 171584
rect 116176 171572 116182 171624
rect 104802 171028 104808 171080
rect 104860 171068 104866 171080
rect 113174 171068 113180 171080
rect 104860 171040 113180 171068
rect 104860 171028 104866 171040
rect 113174 171028 113180 171040
rect 113232 171028 113238 171080
rect 113910 169804 113916 169856
rect 113968 169844 113974 169856
rect 116302 169844 116308 169856
rect 113968 169816 116308 169844
rect 113968 169804 113974 169816
rect 116302 169804 116308 169816
rect 116360 169804 116366 169856
rect 104250 169736 104256 169788
rect 104308 169776 104314 169788
rect 116394 169776 116400 169788
rect 104308 169748 116400 169776
rect 104308 169736 104314 169748
rect 116394 169736 116400 169748
rect 116452 169736 116458 169788
rect 104802 169668 104808 169720
rect 104860 169708 104866 169720
rect 113266 169708 113272 169720
rect 104860 169680 113272 169708
rect 104860 169668 104866 169680
rect 113266 169668 113272 169680
rect 113324 169668 113330 169720
rect 215110 169668 215116 169720
rect 215168 169708 215174 169720
rect 225690 169708 225696 169720
rect 215168 169680 225696 169708
rect 215168 169668 215174 169680
rect 225690 169668 225696 169680
rect 225748 169668 225754 169720
rect 215110 168580 215116 168632
rect 215168 168620 215174 168632
rect 221550 168620 221556 168632
rect 215168 168592 221556 168620
rect 215168 168580 215174 168592
rect 221550 168580 221556 168592
rect 221608 168580 221614 168632
rect 104802 168376 104808 168428
rect 104860 168416 104866 168428
rect 116394 168416 116400 168428
rect 104860 168388 116400 168416
rect 104860 168376 104866 168388
rect 116394 168376 116400 168388
rect 116452 168376 116458 168428
rect 104158 168308 104164 168360
rect 104216 168348 104222 168360
rect 113910 168348 113916 168360
rect 104216 168320 113916 168348
rect 104216 168308 104222 168320
rect 113910 168308 113916 168320
rect 113968 168308 113974 168360
rect 213914 168036 213920 168088
rect 213972 168076 213978 168088
rect 215938 168076 215944 168088
rect 213972 168048 215944 168076
rect 213972 168036 213978 168048
rect 215938 168036 215944 168048
rect 215996 168036 216002 168088
rect 215294 167628 215300 167680
rect 215352 167668 215358 167680
rect 227070 167668 227076 167680
rect 215352 167640 227076 167668
rect 215352 167628 215358 167640
rect 227070 167628 227076 167640
rect 227128 167628 227134 167680
rect 214282 167560 214288 167612
rect 214340 167600 214346 167612
rect 221458 167600 221464 167612
rect 214340 167572 221464 167600
rect 214340 167560 214346 167572
rect 221458 167560 221464 167572
rect 221516 167560 221522 167612
rect 114462 167016 114468 167068
rect 114520 167056 114526 167068
rect 115934 167056 115940 167068
rect 114520 167028 115940 167056
rect 114520 167016 114526 167028
rect 115934 167016 115940 167028
rect 115992 167016 115998 167068
rect 232222 166948 232228 167000
rect 232280 166988 232286 167000
rect 232590 166988 232596 167000
rect 232280 166960 232596 166988
rect 232280 166948 232286 166960
rect 232590 166948 232596 166960
rect 232648 166948 232654 167000
rect 214374 166812 214380 166864
rect 214432 166852 214438 166864
rect 220078 166852 220084 166864
rect 214432 166824 220084 166852
rect 214432 166812 214438 166824
rect 220078 166812 220084 166824
rect 220136 166812 220142 166864
rect 217226 165792 217232 165844
rect 217284 165832 217290 165844
rect 220262 165832 220268 165844
rect 217284 165804 220268 165832
rect 217284 165792 217290 165804
rect 220262 165792 220268 165804
rect 220320 165792 220326 165844
rect 113818 165588 113824 165640
rect 113876 165628 113882 165640
rect 115934 165628 115940 165640
rect 113876 165600 115940 165628
rect 113876 165588 113882 165600
rect 115934 165588 115940 165600
rect 115992 165588 115998 165640
rect 104618 165520 104624 165572
rect 104676 165560 104682 165572
rect 114462 165560 114468 165572
rect 104676 165532 114468 165560
rect 104676 165520 104682 165532
rect 114462 165520 114468 165532
rect 114520 165520 114526 165572
rect 214098 165520 214104 165572
rect 214156 165560 214162 165572
rect 224310 165560 224316 165572
rect 214156 165532 224316 165560
rect 214156 165520 214162 165532
rect 224310 165520 224316 165532
rect 224368 165520 224374 165572
rect 114462 164228 114468 164280
rect 114520 164268 114526 164280
rect 116118 164268 116124 164280
rect 114520 164240 116124 164268
rect 114520 164228 114526 164240
rect 116118 164228 116124 164240
rect 116176 164228 116182 164280
rect 104802 164160 104808 164212
rect 104860 164200 104866 164212
rect 113818 164200 113824 164212
rect 104860 164172 113824 164200
rect 104860 164160 104866 164172
rect 113818 164160 113824 164172
rect 113876 164160 113882 164212
rect 214374 164160 214380 164212
rect 214432 164200 214438 164212
rect 225598 164200 225604 164212
rect 214432 164172 225604 164200
rect 214432 164160 214438 164172
rect 225598 164160 225604 164172
rect 225656 164160 225662 164212
rect 232314 164160 232320 164212
rect 232372 164200 232378 164212
rect 232590 164200 232596 164212
rect 232372 164172 232596 164200
rect 232372 164160 232378 164172
rect 232590 164160 232596 164172
rect 232648 164160 232654 164212
rect 214926 164092 214932 164144
rect 214984 164132 214990 164144
rect 218698 164132 218704 164144
rect 214984 164104 218704 164132
rect 214984 164092 214990 164104
rect 218698 164092 218704 164104
rect 218756 164092 218762 164144
rect 214926 163344 214932 163396
rect 214984 163384 214990 163396
rect 217226 163384 217232 163396
rect 214984 163356 217232 163384
rect 214984 163344 214990 163356
rect 217226 163344 217232 163356
rect 217284 163344 217290 163396
rect 113174 162868 113180 162920
rect 113232 162908 113238 162920
rect 116394 162908 116400 162920
rect 113232 162880 116400 162908
rect 113232 162868 113238 162880
rect 116394 162868 116400 162880
rect 116452 162868 116458 162920
rect 104802 162800 104808 162852
rect 104860 162840 104866 162852
rect 114462 162840 114468 162852
rect 104860 162812 114468 162840
rect 104860 162800 104866 162812
rect 114462 162800 114468 162812
rect 114520 162800 114526 162852
rect 214282 162800 214288 162852
rect 214340 162840 214346 162852
rect 226978 162840 226984 162852
rect 214340 162812 226984 162840
rect 214340 162800 214346 162812
rect 226978 162800 226984 162812
rect 227036 162800 227042 162852
rect 215110 162732 215116 162784
rect 215168 162772 215174 162784
rect 222838 162772 222844 162784
rect 215168 162744 222844 162772
rect 215168 162732 215174 162744
rect 222838 162732 222844 162744
rect 222896 162732 222902 162784
rect 113266 161984 113272 162036
rect 113324 162024 113330 162036
rect 116210 162024 116216 162036
rect 113324 161996 116216 162024
rect 113324 161984 113330 161996
rect 116210 161984 116216 161996
rect 116268 161984 116274 162036
rect 103698 161440 103704 161492
rect 103756 161480 103762 161492
rect 116394 161480 116400 161492
rect 103756 161452 116400 161480
rect 103756 161440 103762 161452
rect 116394 161440 116400 161452
rect 116452 161440 116458 161492
rect 104802 161372 104808 161424
rect 104860 161412 104866 161424
rect 113174 161412 113180 161424
rect 104860 161384 113180 161412
rect 104860 161372 104866 161384
rect 113174 161372 113180 161384
rect 113232 161372 113238 161424
rect 215110 161372 215116 161424
rect 215168 161412 215174 161424
rect 229738 161412 229744 161424
rect 215168 161384 229744 161412
rect 215168 161372 215174 161384
rect 229738 161372 229744 161384
rect 229796 161372 229802 161424
rect 104250 160080 104256 160132
rect 104308 160120 104314 160132
rect 116394 160120 116400 160132
rect 104308 160092 116400 160120
rect 104308 160080 104314 160092
rect 116394 160080 116400 160092
rect 116452 160080 116458 160132
rect 104802 160012 104808 160064
rect 104860 160052 104866 160064
rect 113266 160052 113272 160064
rect 104860 160024 113272 160052
rect 104860 160012 104866 160024
rect 113266 160012 113272 160024
rect 113324 160012 113330 160064
rect 104802 158720 104808 158772
rect 104860 158760 104866 158772
rect 116394 158760 116400 158772
rect 104860 158732 116400 158760
rect 104860 158720 104866 158732
rect 116394 158720 116400 158732
rect 116452 158720 116458 158772
rect 104342 157360 104348 157412
rect 104400 157400 104406 157412
rect 116394 157400 116400 157412
rect 104400 157372 116400 157400
rect 104400 157360 104406 157372
rect 116394 157360 116400 157372
rect 116452 157360 116458 157412
rect 114278 155932 114284 155984
rect 114336 155972 114342 155984
rect 116026 155972 116032 155984
rect 114336 155944 116032 155972
rect 114336 155932 114342 155944
rect 116026 155932 116032 155944
rect 116084 155932 116090 155984
rect 215110 155932 215116 155984
rect 215168 155972 215174 155984
rect 224678 155972 224684 155984
rect 215168 155944 224684 155972
rect 215168 155932 215174 155944
rect 224678 155932 224684 155944
rect 224736 155932 224742 155984
rect 113450 154640 113456 154692
rect 113508 154680 113514 154692
rect 116026 154680 116032 154692
rect 113508 154652 116032 154680
rect 113508 154640 113514 154652
rect 116026 154640 116032 154652
rect 116084 154640 116090 154692
rect 214374 154640 214380 154692
rect 214432 154680 214438 154692
rect 224586 154680 224592 154692
rect 214432 154652 224592 154680
rect 214432 154640 214438 154652
rect 224586 154640 224592 154652
rect 224644 154640 224650 154692
rect 104158 154572 104164 154624
rect 104216 154612 104222 154624
rect 116394 154612 116400 154624
rect 104216 154584 116400 154612
rect 104216 154572 104222 154584
rect 116394 154572 116400 154584
rect 116452 154572 116458 154624
rect 215110 154572 215116 154624
rect 215168 154612 215174 154624
rect 225598 154612 225604 154624
rect 215168 154584 225604 154612
rect 215168 154572 215174 154584
rect 225598 154572 225604 154584
rect 225656 154572 225662 154624
rect 104618 154504 104624 154556
rect 104676 154544 104682 154556
rect 114278 154544 114284 154556
rect 104676 154516 114284 154544
rect 104676 154504 104682 154516
rect 114278 154504 114284 154516
rect 114336 154504 114342 154556
rect 215202 153280 215208 153332
rect 215260 153320 215266 153332
rect 224862 153320 224868 153332
rect 215260 153292 224868 153320
rect 215260 153280 215266 153292
rect 224862 153280 224868 153292
rect 224920 153280 224926 153332
rect 103790 153212 103796 153264
rect 103848 153252 103854 153264
rect 115934 153252 115940 153264
rect 103848 153224 115940 153252
rect 103848 153212 103854 153224
rect 115934 153212 115940 153224
rect 115992 153212 115998 153264
rect 215110 153212 215116 153264
rect 215168 153252 215174 153264
rect 224770 153252 224776 153264
rect 215168 153224 224776 153252
rect 215168 153212 215174 153224
rect 224770 153212 224776 153224
rect 224828 153212 224834 153264
rect 104802 153144 104808 153196
rect 104860 153184 104866 153196
rect 113450 153184 113456 153196
rect 104860 153156 113456 153184
rect 104860 153144 104866 153156
rect 113450 153144 113456 153156
rect 113508 153144 113514 153196
rect 214006 151852 214012 151904
rect 214064 151892 214070 151904
rect 224494 151892 224500 151904
rect 214064 151864 224500 151892
rect 214064 151852 214070 151864
rect 224494 151852 224500 151864
rect 224552 151852 224558 151904
rect 103698 151784 103704 151836
rect 103756 151824 103762 151836
rect 116394 151824 116400 151836
rect 103756 151796 116400 151824
rect 103756 151784 103762 151796
rect 116394 151784 116400 151796
rect 116452 151784 116458 151836
rect 218698 151784 218704 151836
rect 218756 151824 218762 151836
rect 286134 151824 286140 151836
rect 218756 151796 286140 151824
rect 218756 151784 218762 151796
rect 286134 151784 286140 151796
rect 286192 151784 286198 151836
rect 214374 150492 214380 150544
rect 214432 150532 214438 150544
rect 216674 150532 216680 150544
rect 214432 150504 216680 150532
rect 214432 150492 214438 150504
rect 216674 150492 216680 150504
rect 216732 150492 216738 150544
rect 104342 150424 104348 150476
rect 104400 150464 104406 150476
rect 116394 150464 116400 150476
rect 104400 150436 116400 150464
rect 104400 150424 104406 150436
rect 116394 150424 116400 150436
rect 116452 150424 116458 150476
rect 215110 150424 215116 150476
rect 215168 150464 215174 150476
rect 224034 150464 224040 150476
rect 215168 150436 224040 150464
rect 215168 150424 215174 150436
rect 224034 150424 224040 150436
rect 224092 150424 224098 150476
rect 224678 150356 224684 150408
rect 224736 150396 224742 150408
rect 227438 150396 227444 150408
rect 224736 150368 227444 150396
rect 224736 150356 224742 150368
rect 227438 150356 227444 150368
rect 227496 150356 227502 150408
rect 232130 149676 232136 149728
rect 232188 149716 232194 149728
rect 232498 149716 232504 149728
rect 232188 149688 232504 149716
rect 232188 149676 232194 149688
rect 232498 149676 232504 149688
rect 232556 149676 232562 149728
rect 214374 149200 214380 149252
rect 214432 149240 214438 149252
rect 216858 149240 216864 149252
rect 214432 149212 216864 149240
rect 214432 149200 214438 149212
rect 216858 149200 216864 149212
rect 216916 149200 216922 149252
rect 104434 149064 104440 149116
rect 104492 149104 104498 149116
rect 116394 149104 116400 149116
rect 104492 149076 116400 149104
rect 104492 149064 104498 149076
rect 116394 149064 116400 149076
rect 116452 149064 116458 149116
rect 215110 149064 215116 149116
rect 215168 149104 215174 149116
rect 224218 149104 224224 149116
rect 215168 149076 224224 149104
rect 215168 149064 215174 149076
rect 224218 149064 224224 149076
rect 224276 149064 224282 149116
rect 214742 148996 214748 149048
rect 214800 149036 214806 149048
rect 227438 149036 227444 149048
rect 214800 149008 227444 149036
rect 214800 148996 214806 149008
rect 227438 148996 227444 149008
rect 227496 148996 227502 149048
rect 224586 148928 224592 148980
rect 224644 148968 224650 148980
rect 227530 148968 227536 148980
rect 224644 148940 227536 148968
rect 224644 148928 224650 148940
rect 227530 148928 227536 148940
rect 227588 148928 227594 148980
rect 104802 147636 104808 147688
rect 104860 147676 104866 147688
rect 116394 147676 116400 147688
rect 104860 147648 116400 147676
rect 104860 147636 104866 147648
rect 116394 147636 116400 147648
rect 116452 147636 116458 147688
rect 215110 147636 215116 147688
rect 215168 147676 215174 147688
rect 216766 147676 216772 147688
rect 215168 147648 216772 147676
rect 215168 147636 215174 147648
rect 216766 147636 216772 147648
rect 216824 147636 216830 147688
rect 224862 147568 224868 147620
rect 224920 147608 224926 147620
rect 226702 147608 226708 147620
rect 224920 147580 226708 147608
rect 224920 147568 224926 147580
rect 226702 147568 226708 147580
rect 226760 147568 226766 147620
rect 224770 147500 224776 147552
rect 224828 147540 224834 147552
rect 226518 147540 226524 147552
rect 224828 147512 226524 147540
rect 224828 147500 224834 147512
rect 226518 147500 226524 147512
rect 226576 147500 226582 147552
rect 113634 146344 113640 146396
rect 113692 146384 113698 146396
rect 115934 146384 115940 146396
rect 113692 146356 115940 146384
rect 113692 146344 113698 146356
rect 115934 146344 115940 146356
rect 115992 146344 115998 146396
rect 215202 146344 215208 146396
rect 215260 146384 215266 146396
rect 217686 146384 217692 146396
rect 215260 146356 217692 146384
rect 215260 146344 215266 146356
rect 217686 146344 217692 146356
rect 217744 146344 217750 146396
rect 104158 146276 104164 146328
rect 104216 146316 104222 146328
rect 116394 146316 116400 146328
rect 104216 146288 116400 146316
rect 104216 146276 104222 146288
rect 116394 146276 116400 146288
rect 116452 146276 116458 146328
rect 214834 146276 214840 146328
rect 214892 146316 214898 146328
rect 227622 146316 227628 146328
rect 214892 146288 227628 146316
rect 214892 146276 214898 146288
rect 227622 146276 227628 146288
rect 227680 146276 227686 146328
rect 216674 146208 216680 146260
rect 216732 146248 216738 146260
rect 226702 146248 226708 146260
rect 216732 146220 226708 146248
rect 216732 146208 216738 146220
rect 226702 146208 226708 146220
rect 226760 146208 226766 146260
rect 224494 146140 224500 146192
rect 224552 146180 224558 146192
rect 227438 146180 227444 146192
rect 224552 146152 227444 146180
rect 224552 146140 224558 146152
rect 227438 146140 227444 146152
rect 227496 146140 227502 146192
rect 215202 144984 215208 145036
rect 215260 145024 215266 145036
rect 217410 145024 217416 145036
rect 215260 144996 217416 145024
rect 215260 144984 215266 144996
rect 217410 144984 217416 144996
rect 217468 144984 217474 145036
rect 104526 144916 104532 144968
rect 104584 144956 104590 144968
rect 116026 144956 116032 144968
rect 104584 144928 116032 144956
rect 104584 144916 104590 144928
rect 116026 144916 116032 144928
rect 116084 144916 116090 144968
rect 215018 144916 215024 144968
rect 215076 144956 215082 144968
rect 227254 144956 227260 144968
rect 215076 144928 227260 144956
rect 215076 144916 215082 144928
rect 227254 144916 227260 144928
rect 227312 144916 227318 144968
rect 104618 144848 104624 144900
rect 104676 144888 104682 144900
rect 113634 144888 113640 144900
rect 104676 144860 113640 144888
rect 104676 144848 104682 144860
rect 113634 144848 113640 144860
rect 113692 144848 113698 144900
rect 216858 144848 216864 144900
rect 216916 144888 216922 144900
rect 226518 144888 226524 144900
rect 216916 144860 226524 144888
rect 216916 144848 216922 144860
rect 226518 144848 226524 144860
rect 226576 144848 226582 144900
rect 224034 144780 224040 144832
rect 224092 144820 224098 144832
rect 227438 144820 227444 144832
rect 224092 144792 227444 144820
rect 224092 144780 224098 144792
rect 227438 144780 227444 144792
rect 227496 144780 227502 144832
rect 215202 143624 215208 143676
rect 215260 143664 215266 143676
rect 216674 143664 216680 143676
rect 215260 143636 216680 143664
rect 215260 143624 215266 143636
rect 216674 143624 216680 143636
rect 216732 143624 216738 143676
rect 103514 143556 103520 143608
rect 103572 143596 103578 143608
rect 116394 143596 116400 143608
rect 103572 143568 116400 143596
rect 103572 143556 103578 143568
rect 116394 143556 116400 143568
rect 116452 143556 116458 143608
rect 214466 143556 214472 143608
rect 214524 143596 214530 143608
rect 227530 143596 227536 143608
rect 214524 143568 227536 143596
rect 214524 143556 214530 143568
rect 227530 143556 227536 143568
rect 227588 143556 227594 143608
rect 216766 143488 216772 143540
rect 216824 143528 216830 143540
rect 226886 143528 226892 143540
rect 216824 143500 226892 143528
rect 216824 143488 216830 143500
rect 226886 143488 226892 143500
rect 226944 143488 226950 143540
rect 224218 143420 224224 143472
rect 224276 143460 224282 143472
rect 227438 143460 227444 143472
rect 224276 143432 227444 143460
rect 224276 143420 224282 143432
rect 227438 143420 227444 143432
rect 227496 143420 227502 143472
rect 215202 142196 215208 142248
rect 215260 142236 215266 142248
rect 216766 142236 216772 142248
rect 215260 142208 216772 142236
rect 215260 142196 215266 142208
rect 216766 142196 216772 142208
rect 216824 142196 216830 142248
rect 103698 142128 103704 142180
rect 103756 142168 103762 142180
rect 116394 142168 116400 142180
rect 103756 142140 116400 142168
rect 103756 142128 103762 142140
rect 116394 142128 116400 142140
rect 116452 142128 116458 142180
rect 215110 142128 215116 142180
rect 215168 142168 215174 142180
rect 227346 142168 227352 142180
rect 215168 142140 227352 142168
rect 215168 142128 215174 142140
rect 227346 142128 227352 142140
rect 227404 142128 227410 142180
rect 217686 142060 217692 142112
rect 217744 142100 217750 142112
rect 226702 142100 226708 142112
rect 217744 142072 226708 142100
rect 217744 142060 217750 142072
rect 226702 142060 226708 142072
rect 226760 142060 226766 142112
rect 104342 140768 104348 140820
rect 104400 140808 104406 140820
rect 116394 140808 116400 140820
rect 104400 140780 116400 140808
rect 104400 140768 104406 140780
rect 116394 140768 116400 140780
rect 116452 140768 116458 140820
rect 215110 140768 215116 140820
rect 215168 140808 215174 140820
rect 226702 140808 226708 140820
rect 215168 140780 226708 140808
rect 215168 140768 215174 140780
rect 226702 140768 226708 140780
rect 226760 140768 226766 140820
rect 217410 140700 217416 140752
rect 217468 140740 217474 140752
rect 227070 140740 227076 140752
rect 217468 140712 227076 140740
rect 217468 140700 217474 140712
rect 227070 140700 227076 140712
rect 227128 140700 227134 140752
rect 113542 139476 113548 139528
rect 113600 139516 113606 139528
rect 116302 139516 116308 139528
rect 113600 139488 116308 139516
rect 113600 139476 113606 139488
rect 116302 139476 116308 139488
rect 116360 139476 116366 139528
rect 214374 139476 214380 139528
rect 214432 139516 214438 139528
rect 226610 139516 226616 139528
rect 214432 139488 226616 139516
rect 214432 139476 214438 139488
rect 226610 139476 226616 139488
rect 226668 139476 226674 139528
rect 104802 139408 104808 139460
rect 104860 139448 104866 139460
rect 116394 139448 116400 139460
rect 104860 139420 116400 139448
rect 104860 139408 104866 139420
rect 116394 139408 116400 139420
rect 116452 139408 116458 139460
rect 215110 139408 215116 139460
rect 215168 139448 215174 139460
rect 226518 139448 226524 139460
rect 215168 139420 226524 139448
rect 215168 139408 215174 139420
rect 226518 139408 226524 139420
rect 226576 139408 226582 139460
rect 216674 139340 216680 139392
rect 216732 139380 216738 139392
rect 227438 139380 227444 139392
rect 216732 139352 227444 139380
rect 216732 139340 216738 139352
rect 227438 139340 227444 139352
rect 227496 139340 227502 139392
rect 215110 138048 215116 138100
rect 215168 138088 215174 138100
rect 226794 138088 226800 138100
rect 215168 138060 226800 138088
rect 215168 138048 215174 138060
rect 226794 138048 226800 138060
rect 226852 138048 226858 138100
rect 214466 137980 214472 138032
rect 214524 138020 214530 138032
rect 226426 138020 226432 138032
rect 214524 137992 226432 138020
rect 214524 137980 214530 137992
rect 226426 137980 226432 137992
rect 226484 137980 226490 138032
rect 216766 137912 216772 137964
rect 216824 137952 216830 137964
rect 227438 137952 227444 137964
rect 216824 137924 227444 137952
rect 216824 137912 216830 137924
rect 227438 137912 227444 137924
rect 227496 137912 227502 137964
rect 215110 136688 215116 136740
rect 215168 136728 215174 136740
rect 227254 136728 227260 136740
rect 215168 136700 227260 136728
rect 215168 136688 215174 136700
rect 227254 136688 227260 136700
rect 227312 136688 227318 136740
rect 104710 136620 104716 136672
rect 104768 136660 104774 136672
rect 116394 136660 116400 136672
rect 104768 136632 116400 136660
rect 104768 136620 104774 136632
rect 116394 136620 116400 136632
rect 116452 136620 116458 136672
rect 214282 136620 214288 136672
rect 214340 136660 214346 136672
rect 227438 136660 227444 136672
rect 214340 136632 227444 136660
rect 214340 136620 214346 136632
rect 227438 136620 227444 136632
rect 227496 136620 227502 136672
rect 104342 135260 104348 135312
rect 104400 135300 104406 135312
rect 115934 135300 115940 135312
rect 104400 135272 115940 135300
rect 104400 135260 104406 135272
rect 115934 135260 115940 135272
rect 115992 135260 115998 135312
rect 214190 135260 214196 135312
rect 214248 135300 214254 135312
rect 226518 135300 226524 135312
rect 214248 135272 226524 135300
rect 214248 135260 214254 135272
rect 226518 135260 226524 135272
rect 226576 135260 226582 135312
rect 104802 135192 104808 135244
rect 104860 135232 104866 135244
rect 113542 135232 113548 135244
rect 104860 135204 113548 135232
rect 104860 135192 104866 135204
rect 113542 135192 113548 135204
rect 113600 135192 113606 135244
rect 341518 135192 341524 135244
rect 341576 135232 341582 135244
rect 580166 135232 580172 135244
rect 341576 135204 580172 135232
rect 341576 135192 341582 135204
rect 580166 135192 580172 135204
rect 580224 135192 580230 135244
rect 215110 133968 215116 134020
rect 215168 134008 215174 134020
rect 226702 134008 226708 134020
rect 215168 133980 226708 134008
rect 215168 133968 215174 133980
rect 226702 133968 226708 133980
rect 226760 133968 226766 134020
rect 109862 133900 109868 133952
rect 109920 133940 109926 133952
rect 116394 133940 116400 133952
rect 109920 133912 116400 133940
rect 109920 133900 109926 133912
rect 116394 133900 116400 133912
rect 116452 133900 116458 133952
rect 215202 133900 215208 133952
rect 215260 133940 215266 133952
rect 227530 133940 227536 133952
rect 215260 133912 227536 133940
rect 215260 133900 215266 133912
rect 227530 133900 227536 133912
rect 227588 133900 227594 133952
rect 104802 133832 104808 133884
rect 104860 133872 104866 133884
rect 115842 133872 115848 133884
rect 104860 133844 115848 133872
rect 104860 133832 104866 133844
rect 115842 133832 115848 133844
rect 115900 133832 115906 133884
rect 114554 132880 114560 132932
rect 114612 132920 114618 132932
rect 117130 132920 117136 132932
rect 114612 132892 117136 132920
rect 114612 132880 114618 132892
rect 117130 132880 117136 132892
rect 117188 132880 117194 132932
rect 214006 132540 214012 132592
rect 214064 132580 214070 132592
rect 227346 132580 227352 132592
rect 214064 132552 227352 132580
rect 214064 132540 214070 132552
rect 227346 132540 227352 132552
rect 227404 132540 227410 132592
rect 215110 132472 215116 132524
rect 215168 132512 215174 132524
rect 227438 132512 227444 132524
rect 215168 132484 227444 132512
rect 215168 132472 215174 132484
rect 227438 132472 227444 132484
rect 227496 132472 227502 132524
rect 215110 131180 215116 131232
rect 215168 131220 215174 131232
rect 226518 131220 226524 131232
rect 215168 131192 226524 131220
rect 215168 131180 215174 131192
rect 226518 131180 226524 131192
rect 226576 131180 226582 131232
rect 113726 131112 113732 131164
rect 113784 131152 113790 131164
rect 116118 131152 116124 131164
rect 113784 131124 116124 131152
rect 113784 131112 113790 131124
rect 116118 131112 116124 131124
rect 116176 131112 116182 131164
rect 214374 131112 214380 131164
rect 214432 131152 214438 131164
rect 227070 131152 227076 131164
rect 214432 131124 227076 131152
rect 214432 131112 214438 131124
rect 227070 131112 227076 131124
rect 227128 131112 227134 131164
rect 103974 130704 103980 130756
rect 104032 130744 104038 130756
rect 109862 130744 109868 130756
rect 104032 130716 109868 130744
rect 104032 130704 104038 130716
rect 109862 130704 109868 130716
rect 109920 130704 109926 130756
rect 100754 130364 100760 130416
rect 100812 130404 100818 130416
rect 116394 130404 116400 130416
rect 100812 130376 116400 130404
rect 100812 130364 100818 130376
rect 116394 130364 116400 130376
rect 116452 130364 116458 130416
rect 214190 129752 214196 129804
rect 214248 129792 214254 129804
rect 227530 129792 227536 129804
rect 214248 129764 227536 129792
rect 214248 129752 214254 129764
rect 227530 129752 227536 129764
rect 227588 129752 227594 129804
rect 104802 129684 104808 129736
rect 104860 129724 104866 129736
rect 114554 129724 114560 129736
rect 104860 129696 114560 129724
rect 104860 129684 104866 129696
rect 114554 129684 114560 129696
rect 114612 129684 114618 129736
rect 116394 129316 116400 129328
rect 10428 129288 116400 129316
rect 10428 129260 10456 129288
rect 116394 129276 116400 129288
rect 116452 129276 116458 129328
rect 10410 129208 10416 129260
rect 10468 129208 10474 129260
rect 214190 129004 214196 129056
rect 214248 129044 214254 129056
rect 227438 129044 227444 129056
rect 214248 129016 227444 129044
rect 214248 129004 214254 129016
rect 227438 129004 227444 129016
rect 227496 129004 227502 129056
rect 214006 128324 214012 128376
rect 214064 128364 214070 128376
rect 226334 128364 226340 128376
rect 214064 128336 226340 128364
rect 214064 128324 214070 128336
rect 226334 128324 226340 128336
rect 226392 128324 226398 128376
rect 9030 128256 9036 128308
rect 9088 128296 9094 128308
rect 116394 128296 116400 128308
rect 9088 128268 116400 128296
rect 9088 128256 9094 128268
rect 116394 128256 116400 128268
rect 116452 128256 116458 128308
rect 104802 128188 104808 128240
rect 104860 128228 104866 128240
rect 113726 128228 113732 128240
rect 104860 128200 113732 128228
rect 104860 128188 104866 128200
rect 113726 128188 113732 128200
rect 113784 128188 113790 128240
rect 215110 127576 215116 127628
rect 215168 127616 215174 127628
rect 227438 127616 227444 127628
rect 215168 127588 227444 127616
rect 215168 127576 215174 127588
rect 227438 127576 227444 127588
rect 227496 127576 227502 127628
rect 215110 126964 215116 127016
rect 215168 127004 215174 127016
rect 227438 127004 227444 127016
rect 215168 126976 227444 127004
rect 215168 126964 215174 126976
rect 227438 126964 227444 126976
rect 227496 126964 227502 127016
rect 10318 126896 10324 126948
rect 10376 126936 10382 126948
rect 116394 126936 116400 126948
rect 10376 126908 116400 126936
rect 10376 126896 10382 126908
rect 116394 126896 116400 126908
rect 116452 126896 116458 126948
rect 215110 126216 215116 126268
rect 215168 126256 215174 126268
rect 227438 126256 227444 126268
rect 215168 126228 227444 126256
rect 215168 126216 215174 126228
rect 227438 126216 227444 126228
rect 227496 126216 227502 126268
rect 215110 125604 215116 125656
rect 215168 125644 215174 125656
rect 227438 125644 227444 125656
rect 215168 125616 227444 125644
rect 215168 125604 215174 125616
rect 227438 125604 227444 125616
rect 227496 125604 227502 125656
rect 8938 125536 8944 125588
rect 8996 125576 9002 125588
rect 116394 125576 116400 125588
rect 8996 125548 116400 125576
rect 8996 125536 9002 125548
rect 116394 125536 116400 125548
rect 116452 125536 116458 125588
rect 78214 125468 78220 125520
rect 78272 125508 78278 125520
rect 100754 125508 100760 125520
rect 78272 125480 100760 125508
rect 78272 125468 78278 125480
rect 100754 125468 100760 125480
rect 100812 125468 100818 125520
rect 215110 124856 215116 124908
rect 215168 124896 215174 124908
rect 227254 124896 227260 124908
rect 215168 124868 227260 124896
rect 215168 124856 215174 124868
rect 227254 124856 227260 124868
rect 227312 124856 227318 124908
rect 215110 124108 215116 124160
rect 215168 124148 215174 124160
rect 227254 124148 227260 124160
rect 215168 124120 227260 124148
rect 215168 124108 215174 124120
rect 227254 124108 227260 124120
rect 227312 124108 227318 124160
rect 215110 123428 215116 123480
rect 215168 123468 215174 123480
rect 227254 123468 227260 123480
rect 215168 123440 227260 123468
rect 215168 123428 215174 123440
rect 227254 123428 227260 123440
rect 227312 123428 227318 123480
rect 215110 122748 215116 122800
rect 215168 122788 215174 122800
rect 227438 122788 227444 122800
rect 215168 122760 227444 122788
rect 215168 122748 215174 122760
rect 227438 122748 227444 122760
rect 227496 122748 227502 122800
rect 215110 122068 215116 122120
rect 215168 122108 215174 122120
rect 227438 122108 227444 122120
rect 215168 122080 227444 122108
rect 215168 122068 215174 122080
rect 227438 122068 227444 122080
rect 227496 122068 227502 122120
rect 50982 121456 50988 121508
rect 51040 121496 51046 121508
rect 116394 121496 116400 121508
rect 51040 121468 116400 121496
rect 51040 121456 51046 121468
rect 116394 121456 116400 121468
rect 116452 121456 116458 121508
rect 215110 121388 215116 121440
rect 215168 121428 215174 121440
rect 227438 121428 227444 121440
rect 215168 121400 227444 121428
rect 215168 121388 215174 121400
rect 227438 121388 227444 121400
rect 227496 121388 227502 121440
rect 215110 120708 215116 120760
rect 215168 120748 215174 120760
rect 227438 120748 227444 120760
rect 215168 120720 227444 120748
rect 215168 120708 215174 120720
rect 227438 120708 227444 120720
rect 227496 120708 227502 120760
rect 100018 120096 100024 120148
rect 100076 120136 100082 120148
rect 116394 120136 116400 120148
rect 100076 120108 116400 120136
rect 100076 120096 100082 120108
rect 116394 120096 116400 120108
rect 116452 120096 116458 120148
rect 214190 120028 214196 120080
rect 214248 120068 214254 120080
rect 227438 120068 227444 120080
rect 214248 120040 227444 120068
rect 214248 120028 214254 120040
rect 227438 120028 227444 120040
rect 227496 120028 227502 120080
rect 94774 118668 94780 118720
rect 94832 118708 94838 118720
rect 116394 118708 116400 118720
rect 94832 118680 116400 118708
rect 94832 118668 94838 118680
rect 116394 118668 116400 118680
rect 116452 118668 116458 118720
rect 214282 118600 214288 118652
rect 214340 118640 214346 118652
rect 226334 118640 226340 118652
rect 214340 118612 226340 118640
rect 214340 118600 214346 118612
rect 226334 118600 226340 118612
rect 226392 118600 226398 118652
rect 215110 118532 215116 118584
rect 215168 118572 215174 118584
rect 226426 118572 226432 118584
rect 215168 118544 226432 118572
rect 215168 118532 215174 118544
rect 226426 118532 226432 118544
rect 226484 118532 226490 118584
rect 94682 117308 94688 117360
rect 94740 117348 94746 117360
rect 116394 117348 116400 117360
rect 94740 117320 116400 117348
rect 94740 117308 94746 117320
rect 116394 117308 116400 117320
rect 116452 117308 116458 117360
rect 215202 117240 215208 117292
rect 215260 117280 215266 117292
rect 227438 117280 227444 117292
rect 215260 117252 227444 117280
rect 215260 117240 215266 117252
rect 227438 117240 227444 117252
rect 227496 117240 227502 117292
rect 215110 117172 215116 117224
rect 215168 117212 215174 117224
rect 226242 117212 226248 117224
rect 215168 117184 226248 117212
rect 215168 117172 215174 117184
rect 226242 117172 226248 117184
rect 226300 117172 226306 117224
rect 94866 116016 94872 116068
rect 94924 116056 94930 116068
rect 116302 116056 116308 116068
rect 94924 116028 116308 116056
rect 94924 116016 94930 116028
rect 116302 116016 116308 116028
rect 116360 116016 116366 116068
rect 94590 115948 94596 116000
rect 94648 115988 94654 116000
rect 116394 115988 116400 116000
rect 94648 115960 116400 115988
rect 94648 115948 94654 115960
rect 116394 115948 116400 115960
rect 116452 115948 116458 116000
rect 215202 115880 215208 115932
rect 215260 115920 215266 115932
rect 227438 115920 227444 115932
rect 215260 115892 227444 115920
rect 215260 115880 215266 115892
rect 227438 115880 227444 115892
rect 227496 115880 227502 115932
rect 215110 115812 215116 115864
rect 215168 115852 215174 115864
rect 226150 115852 226156 115864
rect 215168 115824 226156 115852
rect 215168 115812 215174 115824
rect 226150 115812 226156 115824
rect 226208 115812 226214 115864
rect 94498 114520 94504 114572
rect 94556 114560 94562 114572
rect 116394 114560 116400 114572
rect 94556 114532 116400 114560
rect 94556 114520 94562 114532
rect 116394 114520 116400 114532
rect 116452 114520 116458 114572
rect 215110 114452 215116 114504
rect 215168 114492 215174 114504
rect 227070 114492 227076 114504
rect 215168 114464 227076 114492
rect 215168 114452 215174 114464
rect 227070 114452 227076 114464
rect 227128 114452 227134 114504
rect 214006 114384 214012 114436
rect 214064 114424 214070 114436
rect 226242 114424 226248 114436
rect 214064 114396 226248 114424
rect 214064 114384 214070 114396
rect 226242 114384 226248 114396
rect 226300 114384 226306 114436
rect 95878 113160 95884 113212
rect 95936 113200 95942 113212
rect 116394 113200 116400 113212
rect 95936 113172 116400 113200
rect 95936 113160 95942 113172
rect 116394 113160 116400 113172
rect 116452 113160 116458 113212
rect 214374 113092 214380 113144
rect 214432 113132 214438 113144
rect 226150 113132 226156 113144
rect 214432 113104 226156 113132
rect 214432 113092 214438 113104
rect 226150 113092 226156 113104
rect 226208 113092 226214 113144
rect 98638 111800 98644 111852
rect 98696 111840 98702 111852
rect 116394 111840 116400 111852
rect 98696 111812 116400 111840
rect 98696 111800 98702 111812
rect 116394 111800 116400 111812
rect 116452 111800 116458 111852
rect 215202 111732 215208 111784
rect 215260 111772 215266 111784
rect 226242 111772 226248 111784
rect 215260 111744 226248 111772
rect 215260 111732 215266 111744
rect 226242 111732 226248 111744
rect 226300 111732 226306 111784
rect 215110 111664 215116 111716
rect 215168 111704 215174 111716
rect 226058 111704 226064 111716
rect 215168 111676 226064 111704
rect 215168 111664 215174 111676
rect 226058 111664 226064 111676
rect 226116 111664 226122 111716
rect 104158 110440 104164 110492
rect 104216 110480 104222 110492
rect 116394 110480 116400 110492
rect 104216 110452 116400 110480
rect 104216 110440 104222 110452
rect 116394 110440 116400 110452
rect 116452 110440 116458 110492
rect 215110 110372 215116 110424
rect 215168 110412 215174 110424
rect 225966 110412 225972 110424
rect 215168 110384 225972 110412
rect 215168 110372 215174 110384
rect 225966 110372 225972 110384
rect 226024 110372 226030 110424
rect 214466 110304 214472 110356
rect 214524 110344 214530 110356
rect 226150 110344 226156 110356
rect 214524 110316 226156 110344
rect 214524 110304 214530 110316
rect 226150 110304 226156 110316
rect 226208 110304 226214 110356
rect 94958 109012 94964 109064
rect 95016 109052 95022 109064
rect 116394 109052 116400 109064
rect 95016 109024 116400 109052
rect 95016 109012 95022 109024
rect 116394 109012 116400 109024
rect 116452 109012 116458 109064
rect 215202 108944 215208 108996
rect 215260 108984 215266 108996
rect 226242 108984 226248 108996
rect 215260 108956 226248 108984
rect 215260 108944 215266 108956
rect 226242 108944 226248 108956
rect 226300 108944 226306 108996
rect 215110 108876 215116 108928
rect 215168 108916 215174 108928
rect 225782 108916 225788 108928
rect 215168 108888 225788 108916
rect 215168 108876 215174 108888
rect 225782 108876 225788 108888
rect 225840 108876 225846 108928
rect 105538 107720 105544 107772
rect 105596 107760 105602 107772
rect 116302 107760 116308 107772
rect 105596 107732 116308 107760
rect 105596 107720 105602 107732
rect 116302 107720 116308 107732
rect 116360 107720 116366 107772
rect 97258 107652 97264 107704
rect 97316 107692 97322 107704
rect 116394 107692 116400 107704
rect 97316 107664 116400 107692
rect 97316 107652 97322 107664
rect 116394 107652 116400 107664
rect 116452 107652 116458 107704
rect 214190 107584 214196 107636
rect 214248 107624 214254 107636
rect 226058 107624 226064 107636
rect 214248 107596 226064 107624
rect 214248 107584 214254 107596
rect 226058 107584 226064 107596
rect 226116 107584 226122 107636
rect 101398 106292 101404 106344
rect 101456 106332 101462 106344
rect 116394 106332 116400 106344
rect 101456 106304 116400 106332
rect 101456 106292 101462 106304
rect 116394 106292 116400 106304
rect 116452 106292 116458 106344
rect 215110 106224 215116 106276
rect 215168 106264 215174 106276
rect 225690 106264 225696 106276
rect 215168 106236 225696 106264
rect 215168 106224 215174 106236
rect 225690 106224 225696 106236
rect 225748 106224 225754 106276
rect 214374 106156 214380 106208
rect 214432 106196 214438 106208
rect 226150 106196 226156 106208
rect 214432 106168 226156 106196
rect 214432 106156 214438 106168
rect 226150 106156 226156 106168
rect 226208 106156 226214 106208
rect 97350 104864 97356 104916
rect 97408 104904 97414 104916
rect 116394 104904 116400 104916
rect 97408 104876 116400 104904
rect 97408 104864 97414 104876
rect 116394 104864 116400 104876
rect 116452 104864 116458 104916
rect 224770 104864 224776 104916
rect 224828 104904 224834 104916
rect 227438 104904 227444 104916
rect 224828 104876 227444 104904
rect 224828 104864 224834 104876
rect 227438 104864 227444 104876
rect 227496 104864 227502 104916
rect 215110 104796 215116 104848
rect 215168 104836 215174 104848
rect 225598 104836 225604 104848
rect 215168 104808 225604 104836
rect 215168 104796 215174 104808
rect 225598 104796 225604 104808
rect 225656 104796 225662 104848
rect 214374 104728 214380 104780
rect 214432 104768 214438 104780
rect 226242 104768 226248 104780
rect 214432 104740 226248 104768
rect 214432 104728 214438 104740
rect 226242 104728 226248 104740
rect 226300 104728 226306 104780
rect 224862 103640 224868 103692
rect 224920 103680 224926 103692
rect 227438 103680 227444 103692
rect 224920 103652 227444 103680
rect 224920 103640 224926 103652
rect 227438 103640 227444 103652
rect 227496 103640 227502 103692
rect 102778 103504 102784 103556
rect 102836 103544 102842 103556
rect 116394 103544 116400 103556
rect 102836 103516 116400 103544
rect 102836 103504 102842 103516
rect 116394 103504 116400 103516
rect 116452 103504 116458 103556
rect 215110 103436 215116 103488
rect 215168 103476 215174 103488
rect 226058 103476 226064 103488
rect 215168 103448 226064 103476
rect 215168 103436 215174 103448
rect 226058 103436 226064 103448
rect 226116 103436 226122 103488
rect 215202 103368 215208 103420
rect 215260 103408 215266 103420
rect 225782 103408 225788 103420
rect 215260 103380 225788 103408
rect 215260 103368 215266 103380
rect 225782 103368 225788 103380
rect 225840 103368 225846 103420
rect 95970 102144 95976 102196
rect 96028 102184 96034 102196
rect 116302 102184 116308 102196
rect 96028 102156 116308 102184
rect 96028 102144 96034 102156
rect 116302 102144 116308 102156
rect 116360 102144 116366 102196
rect 215110 102076 215116 102128
rect 215168 102116 215174 102128
rect 225874 102116 225880 102128
rect 215168 102088 225880 102116
rect 215168 102076 215174 102088
rect 225874 102076 225880 102088
rect 225932 102076 225938 102128
rect 314194 102076 314200 102128
rect 314252 102116 314258 102128
rect 338390 102116 338396 102128
rect 314252 102088 338396 102116
rect 314252 102076 314258 102088
rect 338390 102076 338396 102088
rect 338448 102076 338454 102128
rect 98730 100716 98736 100768
rect 98788 100756 98794 100768
rect 116394 100756 116400 100768
rect 98788 100728 116400 100756
rect 98788 100716 98794 100728
rect 116394 100716 116400 100728
rect 116452 100716 116458 100768
rect 214466 100648 214472 100700
rect 214524 100688 214530 100700
rect 226150 100688 226156 100700
rect 214524 100660 226156 100688
rect 214524 100648 214530 100660
rect 226150 100648 226156 100660
rect 226208 100648 226214 100700
rect 232130 100648 232136 100700
rect 232188 100688 232194 100700
rect 258074 100688 258080 100700
rect 232188 100660 258080 100688
rect 232188 100648 232194 100660
rect 258074 100648 258080 100660
rect 258132 100648 258138 100700
rect 215110 100580 215116 100632
rect 215168 100620 215174 100632
rect 225966 100620 225972 100632
rect 215168 100592 225972 100620
rect 215168 100580 215174 100592
rect 225966 100580 225972 100592
rect 226024 100580 226030 100632
rect 100110 99356 100116 99408
rect 100168 99396 100174 99408
rect 116394 99396 116400 99408
rect 100168 99368 116400 99396
rect 100168 99356 100174 99368
rect 116394 99356 116400 99368
rect 116452 99356 116458 99408
rect 214650 99288 214656 99340
rect 214708 99328 214714 99340
rect 226242 99328 226248 99340
rect 214708 99300 226248 99328
rect 214708 99288 214714 99300
rect 226242 99288 226248 99300
rect 226300 99288 226306 99340
rect 232130 99288 232136 99340
rect 232188 99328 232194 99340
rect 232498 99328 232504 99340
rect 232188 99300 232504 99328
rect 232188 99288 232194 99300
rect 232498 99288 232504 99300
rect 232556 99288 232562 99340
rect 215110 99220 215116 99272
rect 215168 99260 215174 99272
rect 224770 99260 224776 99272
rect 215168 99232 224776 99260
rect 215168 99220 215174 99232
rect 224770 99220 224776 99232
rect 224828 99220 224834 99272
rect 95142 98948 95148 99000
rect 95200 98988 95206 99000
rect 100018 98988 100024 99000
rect 95200 98960 100024 98988
rect 95200 98948 95206 98960
rect 100018 98948 100024 98960
rect 100076 98948 100082 99000
rect 106918 97996 106924 98048
rect 106976 98036 106982 98048
rect 116394 98036 116400 98048
rect 106976 98008 116400 98036
rect 106976 97996 106982 98008
rect 116394 97996 116400 98008
rect 116452 97996 116458 98048
rect 214098 97928 214104 97980
rect 214156 97968 214162 97980
rect 224862 97968 224868 97980
rect 214156 97940 224868 97968
rect 214156 97928 214162 97940
rect 224862 97928 224868 97940
rect 224920 97928 224926 97980
rect 214558 96976 214564 97028
rect 214616 97016 214622 97028
rect 218698 97016 218704 97028
rect 214616 96988 218704 97016
rect 214616 96976 214622 96988
rect 218698 96976 218704 96988
rect 218756 96976 218762 97028
rect 96062 96636 96068 96688
rect 96120 96676 96126 96688
rect 116394 96676 116400 96688
rect 96120 96648 116400 96676
rect 96120 96636 96126 96648
rect 116394 96636 116400 96648
rect 116452 96636 116458 96688
rect 94682 95208 94688 95260
rect 94740 95248 94746 95260
rect 116302 95248 116308 95260
rect 94740 95220 116308 95248
rect 94740 95208 94746 95220
rect 116302 95208 116308 95220
rect 116360 95208 116366 95260
rect 215110 95140 215116 95192
rect 215168 95180 215174 95192
rect 576118 95180 576124 95192
rect 215168 95152 576124 95180
rect 215168 95140 215174 95152
rect 576118 95140 576124 95152
rect 576176 95140 576182 95192
rect 94590 93848 94596 93900
rect 94648 93888 94654 93900
rect 116394 93888 116400 93900
rect 94648 93860 116400 93888
rect 94648 93848 94654 93860
rect 116394 93848 116400 93860
rect 116452 93848 116458 93900
rect 215202 93780 215208 93832
rect 215260 93820 215266 93832
rect 578878 93820 578884 93832
rect 215260 93792 578884 93820
rect 215260 93780 215266 93792
rect 578878 93780 578884 93792
rect 578936 93780 578942 93832
rect 215110 93712 215116 93764
rect 215168 93752 215174 93764
rect 577498 93752 577504 93764
rect 215168 93724 577504 93752
rect 215168 93712 215174 93724
rect 577498 93712 577504 93724
rect 577556 93712 577562 93764
rect 94866 93644 94872 93696
rect 94924 93684 94930 93696
rect 95878 93684 95884 93696
rect 94924 93656 95884 93684
rect 94924 93644 94930 93656
rect 95878 93644 95884 93656
rect 95936 93644 95942 93696
rect 94406 93304 94412 93356
rect 94464 93344 94470 93356
rect 98638 93344 98644 93356
rect 94464 93316 98644 93344
rect 94464 93304 94470 93316
rect 98638 93304 98644 93316
rect 98696 93304 98702 93356
rect 98822 93100 98828 93152
rect 98880 93140 98886 93152
rect 116670 93140 116676 93152
rect 98880 93112 116676 93140
rect 98880 93100 98886 93112
rect 116670 93100 116676 93112
rect 116728 93100 116734 93152
rect 101490 92488 101496 92540
rect 101548 92528 101554 92540
rect 116394 92528 116400 92540
rect 101548 92500 116400 92528
rect 101548 92488 101554 92500
rect 116394 92488 116400 92500
rect 116452 92488 116458 92540
rect 95142 92420 95148 92472
rect 95200 92460 95206 92472
rect 104158 92460 104164 92472
rect 95200 92432 104164 92460
rect 95200 92420 95206 92432
rect 104158 92420 104164 92432
rect 104216 92420 104222 92472
rect 104250 91060 104256 91112
rect 104308 91100 104314 91112
rect 116394 91100 116400 91112
rect 104308 91072 116400 91100
rect 104308 91060 104314 91072
rect 116394 91060 116400 91072
rect 116452 91060 116458 91112
rect 95050 90992 95056 91044
rect 95108 91032 95114 91044
rect 105538 91032 105544 91044
rect 95108 91004 105544 91032
rect 95108 90992 95114 91004
rect 105538 90992 105544 91004
rect 105596 90992 105602 91044
rect 97442 89700 97448 89752
rect 97500 89740 97506 89752
rect 116394 89740 116400 89752
rect 97500 89712 116400 89740
rect 97500 89700 97506 89712
rect 116394 89700 116400 89712
rect 116452 89700 116458 89752
rect 214466 89700 214472 89752
rect 214524 89740 214530 89752
rect 227346 89740 227352 89752
rect 214524 89712 227352 89740
rect 214524 89700 214530 89712
rect 227346 89700 227352 89712
rect 227404 89700 227410 89752
rect 95142 89292 95148 89344
rect 95200 89332 95206 89344
rect 97258 89332 97264 89344
rect 95200 89304 97264 89332
rect 95200 89292 95206 89304
rect 97258 89292 97264 89304
rect 97316 89292 97322 89344
rect 215110 88408 215116 88460
rect 215168 88448 215174 88460
rect 221458 88448 221464 88460
rect 215168 88420 221464 88448
rect 215168 88408 215174 88420
rect 221458 88408 221464 88420
rect 221516 88408 221522 88460
rect 97534 88340 97540 88392
rect 97592 88380 97598 88392
rect 115934 88380 115940 88392
rect 97592 88352 115940 88380
rect 97592 88340 97598 88352
rect 115934 88340 115940 88352
rect 115992 88340 115998 88392
rect 214098 88340 214104 88392
rect 214156 88380 214162 88392
rect 222838 88380 222844 88392
rect 214156 88352 222844 88380
rect 214156 88340 214162 88352
rect 222838 88340 222844 88352
rect 222896 88340 222902 88392
rect 340138 88272 340144 88324
rect 340196 88312 340202 88324
rect 580166 88312 580172 88324
rect 340196 88284 580172 88312
rect 340196 88272 340202 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 95142 88204 95148 88256
rect 95200 88244 95206 88256
rect 101398 88244 101404 88256
rect 95200 88216 101404 88244
rect 95200 88204 95206 88216
rect 101398 88204 101404 88216
rect 101456 88204 101462 88256
rect 94406 87864 94412 87916
rect 94464 87904 94470 87916
rect 97350 87904 97356 87916
rect 94464 87876 97356 87904
rect 94464 87864 94470 87876
rect 97350 87864 97356 87876
rect 97408 87864 97414 87916
rect 215018 87048 215024 87100
rect 215076 87088 215082 87100
rect 218698 87088 218704 87100
rect 215076 87060 218704 87088
rect 215076 87048 215082 87060
rect 218698 87048 218704 87060
rect 218756 87048 218762 87100
rect 98638 86980 98644 87032
rect 98696 87020 98702 87032
rect 116394 87020 116400 87032
rect 98696 86992 116400 87020
rect 98696 86980 98702 86992
rect 116394 86980 116400 86992
rect 116452 86980 116458 87032
rect 215110 86980 215116 87032
rect 215168 87020 215174 87032
rect 224218 87020 224224 87032
rect 215168 86992 224224 87020
rect 215168 86980 215174 86992
rect 224218 86980 224224 86992
rect 224276 86980 224282 87032
rect 232314 86912 232320 86964
rect 232372 86952 232378 86964
rect 232498 86952 232504 86964
rect 232372 86924 232504 86952
rect 232372 86912 232378 86924
rect 232498 86912 232504 86924
rect 232556 86912 232562 86964
rect 94498 86708 94504 86760
rect 94556 86748 94562 86760
rect 102778 86748 102784 86760
rect 94556 86720 102784 86748
rect 94556 86708 94562 86720
rect 102778 86708 102784 86720
rect 102836 86708 102842 86760
rect 94038 86164 94044 86216
rect 94096 86204 94102 86216
rect 98730 86204 98736 86216
rect 94096 86176 98736 86204
rect 94096 86164 94102 86176
rect 98730 86164 98736 86176
rect 98788 86164 98794 86216
rect 102870 85552 102876 85604
rect 102928 85592 102934 85604
rect 116118 85592 116124 85604
rect 102928 85564 116124 85592
rect 102928 85552 102934 85564
rect 116118 85552 116124 85564
rect 116176 85552 116182 85604
rect 215110 85552 215116 85604
rect 215168 85592 215174 85604
rect 225598 85592 225604 85604
rect 215168 85564 225604 85592
rect 215168 85552 215174 85564
rect 225598 85552 225604 85564
rect 225656 85552 225662 85604
rect 94866 85484 94872 85536
rect 94924 85524 94930 85536
rect 95970 85524 95976 85536
rect 94924 85496 95976 85524
rect 94924 85484 94930 85496
rect 95970 85484 95976 85496
rect 96028 85484 96034 85536
rect 95142 84804 95148 84856
rect 95200 84844 95206 84856
rect 98822 84844 98828 84856
rect 95200 84816 98828 84844
rect 95200 84804 95206 84816
rect 98822 84804 98828 84816
rect 98880 84804 98886 84856
rect 100018 84804 100024 84856
rect 100076 84844 100082 84856
rect 116394 84844 116400 84856
rect 100076 84816 116400 84844
rect 100076 84804 100082 84816
rect 116394 84804 116400 84816
rect 116452 84804 116458 84856
rect 215202 84192 215208 84244
rect 215260 84232 215266 84244
rect 227070 84232 227076 84244
rect 215260 84204 227076 84232
rect 215260 84192 215266 84204
rect 227070 84192 227076 84204
rect 227128 84192 227134 84244
rect 320818 83512 320824 83564
rect 320876 83552 320882 83564
rect 412082 83552 412088 83564
rect 320876 83524 412088 83552
rect 320876 83512 320882 83524
rect 412082 83512 412088 83524
rect 412140 83512 412146 83564
rect 284478 83444 284484 83496
rect 284536 83484 284542 83496
rect 580258 83484 580264 83496
rect 284536 83456 580264 83484
rect 284536 83444 284542 83456
rect 580258 83444 580264 83456
rect 580316 83444 580322 83496
rect 94222 83376 94228 83428
rect 94280 83416 94286 83428
rect 100110 83416 100116 83428
rect 94280 83388 100116 83416
rect 94280 83376 94286 83388
rect 100110 83376 100116 83388
rect 100168 83376 100174 83428
rect 95878 82832 95884 82884
rect 95936 82872 95942 82884
rect 116394 82872 116400 82884
rect 95936 82844 116400 82872
rect 95936 82832 95942 82844
rect 116394 82832 116400 82844
rect 116452 82832 116458 82884
rect 215938 82832 215944 82884
rect 215996 82872 216002 82884
rect 248138 82872 248144 82884
rect 215996 82844 248144 82872
rect 215996 82832 216002 82844
rect 248138 82832 248144 82844
rect 248196 82832 248202 82884
rect 95142 82764 95148 82816
rect 95200 82804 95206 82816
rect 106918 82804 106924 82816
rect 95200 82776 106924 82804
rect 95200 82764 95206 82776
rect 106918 82764 106924 82776
rect 106976 82764 106982 82816
rect 94958 81404 94964 81456
rect 95016 81444 95022 81456
rect 97534 81444 97540 81456
rect 95016 81416 97540 81444
rect 95016 81404 95022 81416
rect 97534 81404 97540 81416
rect 97592 81404 97598 81456
rect 98730 81404 98736 81456
rect 98788 81444 98794 81456
rect 115934 81444 115940 81456
rect 98788 81416 115940 81444
rect 98788 81404 98794 81416
rect 115934 81404 115940 81416
rect 115992 81404 115998 81456
rect 214190 81404 214196 81456
rect 214248 81444 214254 81456
rect 227162 81444 227168 81456
rect 214248 81416 227168 81444
rect 214248 81404 214254 81416
rect 227162 81404 227168 81416
rect 227220 81404 227226 81456
rect 94406 81336 94412 81388
rect 94464 81376 94470 81388
rect 96062 81376 96068 81388
rect 94464 81348 96068 81376
rect 94464 81336 94470 81348
rect 96062 81336 96068 81348
rect 96120 81336 96126 81388
rect 214558 81336 214564 81388
rect 214616 81376 214622 81388
rect 227438 81376 227444 81388
rect 214616 81348 227444 81376
rect 214616 81336 214622 81348
rect 227438 81336 227444 81348
rect 227496 81336 227502 81388
rect 214742 81268 214748 81320
rect 214800 81308 214806 81320
rect 227530 81308 227536 81320
rect 214800 81280 227536 81308
rect 214800 81268 214806 81280
rect 227530 81268 227536 81280
rect 227588 81268 227594 81320
rect 95234 80656 95240 80708
rect 95292 80696 95298 80708
rect 116578 80696 116584 80708
rect 95292 80668 116584 80696
rect 95292 80656 95298 80668
rect 116578 80656 116584 80668
rect 116636 80656 116642 80708
rect 97258 80044 97264 80096
rect 97316 80084 97322 80096
rect 116394 80084 116400 80096
rect 97316 80056 116400 80084
rect 97316 80044 97322 80056
rect 116394 80044 116400 80056
rect 116452 80044 116458 80096
rect 214006 80044 214012 80096
rect 214064 80084 214070 80096
rect 216122 80084 216128 80096
rect 214064 80056 216128 80084
rect 214064 80044 214070 80056
rect 216122 80044 216128 80056
rect 216180 80044 216186 80096
rect 232314 80044 232320 80096
rect 232372 80044 232378 80096
rect 221458 79976 221464 80028
rect 221516 80016 221522 80028
rect 227438 80016 227444 80028
rect 221516 79988 227444 80016
rect 221516 79976 221522 79988
rect 227438 79976 227444 79988
rect 227496 79976 227502 80028
rect 232332 79960 232360 80044
rect 232314 79908 232320 79960
rect 232372 79908 232378 79960
rect 96062 79296 96068 79348
rect 96120 79336 96126 79348
rect 117038 79336 117044 79348
rect 96120 79308 117044 79336
rect 96120 79296 96126 79308
rect 117038 79296 117044 79308
rect 117096 79296 117102 79348
rect 215110 78752 215116 78804
rect 215168 78792 215174 78804
rect 221550 78792 221556 78804
rect 215168 78764 221556 78792
rect 215168 78752 215174 78764
rect 221550 78752 221556 78764
rect 221608 78752 221614 78804
rect 102778 78684 102784 78736
rect 102836 78724 102842 78736
rect 116394 78724 116400 78736
rect 102836 78696 116400 78724
rect 102836 78684 102842 78696
rect 116394 78684 116400 78696
rect 116452 78684 116458 78736
rect 94406 78616 94412 78668
rect 94464 78656 94470 78668
rect 101490 78656 101496 78668
rect 94464 78628 101496 78656
rect 94464 78616 94470 78628
rect 101490 78616 101496 78628
rect 101548 78616 101554 78668
rect 218698 78616 218704 78668
rect 218756 78656 218762 78668
rect 227530 78656 227536 78668
rect 218756 78628 227536 78656
rect 218756 78616 218762 78628
rect 227530 78616 227536 78628
rect 227588 78616 227594 78668
rect 222838 78548 222844 78600
rect 222896 78588 222902 78600
rect 227438 78588 227444 78600
rect 222896 78560 227444 78588
rect 222896 78548 222902 78560
rect 227438 78548 227444 78560
rect 227496 78548 227502 78600
rect 94222 77936 94228 77988
rect 94280 77976 94286 77988
rect 104250 77976 104256 77988
rect 94280 77948 104256 77976
rect 94280 77936 94286 77948
rect 104250 77936 104256 77948
rect 104308 77936 104314 77988
rect 101398 77256 101404 77308
rect 101456 77296 101462 77308
rect 116394 77296 116400 77308
rect 101456 77268 116400 77296
rect 101456 77256 101462 77268
rect 116394 77256 116400 77268
rect 116452 77256 116458 77308
rect 214742 77256 214748 77308
rect 214800 77296 214806 77308
rect 218790 77296 218796 77308
rect 214800 77268 218796 77296
rect 214800 77256 214806 77268
rect 218790 77256 218796 77268
rect 218848 77256 218854 77308
rect 215202 77188 215208 77240
rect 215260 77228 215266 77240
rect 227530 77228 227536 77240
rect 215260 77200 227536 77228
rect 215260 77188 215266 77200
rect 227530 77188 227536 77200
rect 227588 77188 227594 77240
rect 224218 77120 224224 77172
rect 224276 77160 224282 77172
rect 227438 77160 227444 77172
rect 224276 77132 227444 77160
rect 224276 77120 224282 77132
rect 227438 77120 227444 77132
rect 227496 77120 227502 77172
rect 94038 76848 94044 76900
rect 94096 76888 94102 76900
rect 102870 76888 102876 76900
rect 94096 76860 102876 76888
rect 94096 76848 94102 76860
rect 102870 76848 102876 76860
rect 102928 76848 102934 76900
rect 95970 75896 95976 75948
rect 96028 75936 96034 75948
rect 116394 75936 116400 75948
rect 96028 75908 116400 75936
rect 96028 75896 96034 75908
rect 116394 75896 116400 75908
rect 116452 75896 116458 75948
rect 215202 75896 215208 75948
rect 215260 75936 215266 75948
rect 218054 75936 218060 75948
rect 215260 75908 218060 75936
rect 215260 75896 215266 75908
rect 218054 75896 218060 75908
rect 218112 75896 218118 75948
rect 214650 75828 214656 75880
rect 214708 75868 214714 75880
rect 227438 75868 227444 75880
rect 214708 75840 227444 75868
rect 214708 75828 214714 75840
rect 227438 75828 227444 75840
rect 227496 75828 227502 75880
rect 94590 75692 94596 75744
rect 94648 75732 94654 75744
rect 97442 75732 97448 75744
rect 94648 75704 97448 75732
rect 94648 75692 94654 75704
rect 97442 75692 97448 75704
rect 97500 75692 97506 75744
rect 215202 74604 215208 74656
rect 215260 74644 215266 74656
rect 216030 74644 216036 74656
rect 215260 74616 216036 74644
rect 215260 74604 215266 74616
rect 216030 74604 216036 74616
rect 216088 74604 216094 74656
rect 94590 74536 94596 74588
rect 94648 74576 94654 74588
rect 116394 74576 116400 74588
rect 94648 74548 116400 74576
rect 94648 74536 94654 74548
rect 116394 74536 116400 74548
rect 116452 74536 116458 74588
rect 214834 74468 214840 74520
rect 214892 74508 214898 74520
rect 227438 74508 227444 74520
rect 214892 74480 227444 74508
rect 214892 74468 214898 74480
rect 227438 74468 227444 74480
rect 227496 74468 227502 74520
rect 95142 74196 95148 74248
rect 95200 74236 95206 74248
rect 98638 74236 98644 74248
rect 95200 74208 98644 74236
rect 95200 74196 95206 74208
rect 98638 74196 98644 74208
rect 98696 74196 98702 74248
rect 96614 73788 96620 73840
rect 96672 73828 96678 73840
rect 116578 73828 116584 73840
rect 96672 73800 116584 73828
rect 96672 73788 96678 73800
rect 116578 73788 116584 73800
rect 116636 73788 116642 73840
rect 214834 73448 214840 73500
rect 214892 73488 214898 73500
rect 215110 73488 215116 73500
rect 214892 73460 215116 73488
rect 214892 73448 214898 73460
rect 215110 73448 215116 73460
rect 215168 73448 215174 73500
rect 215110 73312 215116 73364
rect 215168 73352 215174 73364
rect 220722 73352 220728 73364
rect 215168 73324 220728 73352
rect 215168 73312 215174 73324
rect 220722 73312 220728 73324
rect 220780 73312 220786 73364
rect 98822 73176 98828 73228
rect 98880 73216 98886 73228
rect 116394 73216 116400 73228
rect 98880 73188 116400 73216
rect 98880 73176 98886 73188
rect 116394 73176 116400 73188
rect 116452 73176 116458 73228
rect 214926 73108 214932 73160
rect 214984 73148 214990 73160
rect 227438 73148 227444 73160
rect 214984 73120 227444 73148
rect 214984 73108 214990 73120
rect 227438 73108 227444 73120
rect 227496 73108 227502 73160
rect 216122 73040 216128 73092
rect 216180 73080 216186 73092
rect 227530 73080 227536 73092
rect 216180 73052 227536 73080
rect 216180 73040 216186 73052
rect 227530 73040 227536 73052
rect 227588 73040 227594 73092
rect 94406 72632 94412 72684
rect 94464 72672 94470 72684
rect 100018 72672 100024 72684
rect 94464 72644 100024 72672
rect 94464 72632 94470 72644
rect 100018 72632 100024 72644
rect 100076 72632 100082 72684
rect 94774 71748 94780 71800
rect 94832 71788 94838 71800
rect 116394 71788 116400 71800
rect 94832 71760 116400 71788
rect 94832 71748 94838 71760
rect 116394 71748 116400 71760
rect 116452 71748 116458 71800
rect 94222 71680 94228 71732
rect 94280 71720 94286 71732
rect 96062 71720 96068 71732
rect 94280 71692 96068 71720
rect 94280 71680 94286 71692
rect 96062 71680 96068 71692
rect 96120 71680 96126 71732
rect 215018 71680 215024 71732
rect 215076 71720 215082 71732
rect 227438 71720 227444 71732
rect 215076 71692 227444 71720
rect 215076 71680 215082 71692
rect 227438 71680 227444 71692
rect 227496 71680 227502 71732
rect 221550 71612 221556 71664
rect 221608 71652 221614 71664
rect 227530 71652 227536 71664
rect 221608 71624 227536 71652
rect 221608 71612 221614 71624
rect 227530 71612 227536 71624
rect 227588 71612 227594 71664
rect 95050 70456 95056 70508
rect 95108 70496 95114 70508
rect 98730 70496 98736 70508
rect 95108 70468 98736 70496
rect 95108 70456 95114 70468
rect 98730 70456 98736 70468
rect 98788 70456 98794 70508
rect 100018 70456 100024 70508
rect 100076 70496 100082 70508
rect 116302 70496 116308 70508
rect 100076 70468 116308 70496
rect 100076 70456 100082 70468
rect 116302 70456 116308 70468
rect 116360 70456 116366 70508
rect 215110 70456 215116 70508
rect 215168 70496 215174 70508
rect 224126 70496 224132 70508
rect 215168 70468 224132 70496
rect 215168 70456 215174 70468
rect 224126 70456 224132 70468
rect 224184 70456 224190 70508
rect 94498 70388 94504 70440
rect 94556 70428 94562 70440
rect 116394 70428 116400 70440
rect 94556 70400 116400 70428
rect 94556 70388 94562 70400
rect 116394 70388 116400 70400
rect 116452 70388 116458 70440
rect 214098 70388 214104 70440
rect 214156 70428 214162 70440
rect 224862 70428 224868 70440
rect 214156 70400 224868 70428
rect 214156 70388 214162 70400
rect 224862 70388 224868 70400
rect 224920 70388 224926 70440
rect 214558 70320 214564 70372
rect 214616 70360 214622 70372
rect 227438 70360 227444 70372
rect 214616 70332 227444 70360
rect 214616 70320 214622 70332
rect 227438 70320 227444 70332
rect 227496 70320 227502 70372
rect 94866 70252 94872 70304
rect 94924 70292 94930 70304
rect 95878 70292 95884 70304
rect 94924 70264 95884 70292
rect 94924 70252 94930 70264
rect 95878 70252 95884 70264
rect 95936 70252 95942 70304
rect 218790 70252 218796 70304
rect 218848 70292 218854 70304
rect 226518 70292 226524 70304
rect 218848 70264 226524 70292
rect 218848 70252 218854 70264
rect 226518 70252 226524 70264
rect 226576 70252 226582 70304
rect 95142 69844 95148 69896
rect 95200 69884 95206 69896
rect 102778 69884 102784 69896
rect 95200 69856 102784 69884
rect 95200 69844 95206 69856
rect 102778 69844 102784 69856
rect 102836 69844 102842 69896
rect 214926 69096 214932 69148
rect 214984 69136 214990 69148
rect 224402 69136 224408 69148
rect 214984 69108 224408 69136
rect 214984 69096 214990 69108
rect 224402 69096 224408 69108
rect 224460 69096 224466 69148
rect 96062 69028 96068 69080
rect 96120 69068 96126 69080
rect 116394 69068 116400 69080
rect 96120 69040 116400 69068
rect 96120 69028 96126 69040
rect 116394 69028 116400 69040
rect 116452 69028 116458 69080
rect 215110 69028 215116 69080
rect 215168 69068 215174 69080
rect 224586 69068 224592 69080
rect 215168 69040 224592 69068
rect 215168 69028 215174 69040
rect 224586 69028 224592 69040
rect 224644 69028 224650 69080
rect 214466 68960 214472 69012
rect 214524 69000 214530 69012
rect 227438 69000 227444 69012
rect 214524 68972 227444 69000
rect 214524 68960 214530 68972
rect 227438 68960 227444 68972
rect 227496 68960 227502 69012
rect 218054 68892 218060 68944
rect 218112 68932 218118 68944
rect 227530 68932 227536 68944
rect 218112 68904 227536 68932
rect 218112 68892 218118 68904
rect 227530 68892 227536 68904
rect 227588 68892 227594 68944
rect 94038 68552 94044 68604
rect 94096 68592 94102 68604
rect 97258 68592 97264 68604
rect 94096 68564 97264 68592
rect 94096 68552 94102 68564
rect 97258 68552 97264 68564
rect 97316 68552 97322 68604
rect 215202 67668 215208 67720
rect 215260 67708 215266 67720
rect 224218 67708 224224 67720
rect 215260 67680 224224 67708
rect 215260 67668 215266 67680
rect 224218 67668 224224 67680
rect 224276 67668 224282 67720
rect 94682 67600 94688 67652
rect 94740 67640 94746 67652
rect 116394 67640 116400 67652
rect 94740 67612 116400 67640
rect 94740 67600 94746 67612
rect 116394 67600 116400 67612
rect 116452 67600 116458 67652
rect 215110 67600 215116 67652
rect 215168 67640 215174 67652
rect 224770 67640 224776 67652
rect 215168 67612 224776 67640
rect 215168 67600 215174 67612
rect 224770 67600 224776 67612
rect 224828 67600 224834 67652
rect 214834 67532 214840 67584
rect 214892 67572 214898 67584
rect 227438 67572 227444 67584
rect 214892 67544 227444 67572
rect 214892 67532 214898 67544
rect 227438 67532 227444 67544
rect 227496 67532 227502 67584
rect 95142 67464 95148 67516
rect 95200 67504 95206 67516
rect 96614 67504 96620 67516
rect 95200 67476 96620 67504
rect 95200 67464 95206 67476
rect 96614 67464 96620 67476
rect 96672 67464 96678 67516
rect 216030 67464 216036 67516
rect 216088 67504 216094 67516
rect 227530 67504 227536 67516
rect 216088 67476 227536 67504
rect 216088 67464 216094 67476
rect 227530 67464 227536 67476
rect 227588 67464 227594 67516
rect 97258 66240 97264 66292
rect 97316 66280 97322 66292
rect 116394 66280 116400 66292
rect 97316 66252 116400 66280
rect 97316 66240 97322 66252
rect 116394 66240 116400 66252
rect 116452 66240 116458 66292
rect 215110 66240 215116 66292
rect 215168 66280 215174 66292
rect 224678 66280 224684 66292
rect 215168 66252 224684 66280
rect 215168 66240 215174 66252
rect 224678 66240 224684 66252
rect 224736 66240 224742 66292
rect 214282 66172 214288 66224
rect 214340 66212 214346 66224
rect 227438 66212 227444 66224
rect 214340 66184 227444 66212
rect 214340 66172 214346 66184
rect 227438 66172 227444 66184
rect 227496 66172 227502 66224
rect 220722 66104 220728 66156
rect 220780 66144 220786 66156
rect 227530 66144 227536 66156
rect 220780 66116 227536 66144
rect 220780 66104 220786 66116
rect 227530 66104 227536 66116
rect 227588 66104 227594 66156
rect 94406 65968 94412 66020
rect 94464 66008 94470 66020
rect 95970 66008 95976 66020
rect 94464 65980 95976 66008
rect 94464 65968 94470 65980
rect 95970 65968 95976 65980
rect 96028 65968 96034 66020
rect 94130 65900 94136 65952
rect 94188 65940 94194 65952
rect 101398 65940 101404 65952
rect 94188 65912 101404 65940
rect 94188 65900 94194 65912
rect 101398 65900 101404 65912
rect 101456 65900 101462 65952
rect 213914 65152 213920 65204
rect 213972 65192 213978 65204
rect 216858 65192 216864 65204
rect 213972 65164 216864 65192
rect 213972 65152 213978 65164
rect 216858 65152 216864 65164
rect 216916 65152 216922 65204
rect 94866 64880 94872 64932
rect 94924 64920 94930 64932
rect 116394 64920 116400 64932
rect 94924 64892 116400 64920
rect 94924 64880 94930 64892
rect 116394 64880 116400 64892
rect 116452 64880 116458 64932
rect 214006 64880 214012 64932
rect 214064 64920 214070 64932
rect 224494 64920 224500 64932
rect 214064 64892 224500 64920
rect 214064 64880 214070 64892
rect 224494 64880 224500 64892
rect 224552 64880 224558 64932
rect 214650 64676 214656 64728
rect 214708 64716 214714 64728
rect 227254 64716 227260 64728
rect 214708 64688 227260 64716
rect 214708 64676 214714 64688
rect 227254 64676 227260 64688
rect 227312 64676 227318 64728
rect 224862 64472 224868 64524
rect 224920 64512 224926 64524
rect 227438 64512 227444 64524
rect 224920 64484 227444 64512
rect 224920 64472 224926 64484
rect 227438 64472 227444 64484
rect 227496 64472 227502 64524
rect 224126 64200 224132 64252
rect 224184 64240 224190 64252
rect 227530 64240 227536 64252
rect 224184 64212 227536 64240
rect 224184 64200 224190 64212
rect 227530 64200 227536 64212
rect 227588 64200 227594 64252
rect 214098 63588 214104 63640
rect 214156 63628 214162 63640
rect 216950 63628 216956 63640
rect 214156 63600 216956 63628
rect 214156 63588 214162 63600
rect 216950 63588 216956 63600
rect 217008 63588 217014 63640
rect 95234 63520 95240 63572
rect 95292 63560 95298 63572
rect 115934 63560 115940 63572
rect 95292 63532 115940 63560
rect 95292 63520 95298 63532
rect 115934 63520 115940 63532
rect 115992 63520 115998 63572
rect 215110 63520 215116 63572
rect 215168 63560 215174 63572
rect 224310 63560 224316 63572
rect 215168 63532 224316 63560
rect 215168 63520 215174 63532
rect 224310 63520 224316 63532
rect 224368 63520 224374 63572
rect 224586 63452 224592 63504
rect 224644 63492 224650 63504
rect 227070 63492 227076 63504
rect 224644 63464 227076 63492
rect 224644 63452 224650 63464
rect 227070 63452 227076 63464
rect 227128 63452 227134 63504
rect 224402 63384 224408 63436
rect 224460 63424 224466 63436
rect 227438 63424 227444 63436
rect 224460 63396 227444 63424
rect 224460 63384 224466 63396
rect 227438 63384 227444 63396
rect 227496 63384 227502 63436
rect 95142 63180 95148 63232
rect 95200 63220 95206 63232
rect 98822 63220 98828 63232
rect 95200 63192 98828 63220
rect 95200 63180 95206 63192
rect 98822 63180 98828 63192
rect 98880 63180 98886 63232
rect 487614 62772 487620 62824
rect 487672 62812 487678 62824
rect 573358 62812 573364 62824
rect 487672 62784 573364 62812
rect 487672 62772 487678 62784
rect 573358 62772 573364 62784
rect 573416 62772 573422 62824
rect 214374 62160 214380 62212
rect 214432 62200 214438 62212
rect 216674 62200 216680 62212
rect 214432 62172 216680 62200
rect 214432 62160 214438 62172
rect 216674 62160 216680 62172
rect 216732 62160 216738 62212
rect 94590 62092 94596 62144
rect 94648 62132 94654 62144
rect 116394 62132 116400 62144
rect 94648 62104 116400 62132
rect 94648 62092 94654 62104
rect 116394 62092 116400 62104
rect 116452 62092 116458 62144
rect 215110 62092 215116 62144
rect 215168 62132 215174 62144
rect 224126 62132 224132 62144
rect 215168 62104 224132 62132
rect 215168 62092 215174 62104
rect 224126 62092 224132 62104
rect 224184 62092 224190 62144
rect 224770 62024 224776 62076
rect 224828 62064 224834 62076
rect 226702 62064 226708 62076
rect 224828 62036 226708 62064
rect 224828 62024 224834 62036
rect 226702 62024 226708 62036
rect 226760 62024 226766 62076
rect 224218 61956 224224 62008
rect 224276 61996 224282 62008
rect 227438 61996 227444 62008
rect 224276 61968 227444 61996
rect 224276 61956 224282 61968
rect 227438 61956 227444 61968
rect 227496 61956 227502 62008
rect 94314 61752 94320 61804
rect 94372 61792 94378 61804
rect 100018 61792 100024 61804
rect 94372 61764 100024 61792
rect 94372 61752 94378 61764
rect 100018 61752 100024 61764
rect 100076 61752 100082 61804
rect 214742 60800 214748 60852
rect 214800 60840 214806 60852
rect 216766 60840 216772 60852
rect 214800 60812 216772 60840
rect 214800 60800 214806 60812
rect 216766 60800 216772 60812
rect 216824 60800 216830 60852
rect 94774 60732 94780 60784
rect 94832 60772 94838 60784
rect 116394 60772 116400 60784
rect 94832 60744 116400 60772
rect 94832 60732 94838 60744
rect 116394 60732 116400 60744
rect 116452 60732 116458 60784
rect 215110 60732 215116 60784
rect 215168 60772 215174 60784
rect 224402 60772 224408 60784
rect 215168 60744 224408 60772
rect 215168 60732 215174 60744
rect 224402 60732 224408 60744
rect 224460 60732 224466 60784
rect 216858 60664 216864 60716
rect 216916 60704 216922 60716
rect 227530 60704 227536 60716
rect 216916 60676 227536 60704
rect 216916 60664 216922 60676
rect 227530 60664 227536 60676
rect 227588 60664 227594 60716
rect 224678 60596 224684 60648
rect 224736 60636 224742 60648
rect 227438 60636 227444 60648
rect 224736 60608 227444 60636
rect 224736 60596 224742 60608
rect 227438 60596 227444 60608
rect 227496 60596 227502 60648
rect 96154 59984 96160 60036
rect 96212 60024 96218 60036
rect 116486 60024 116492 60036
rect 96212 59996 116492 60024
rect 96212 59984 96218 59996
rect 116486 59984 116492 59996
rect 116544 59984 116550 60036
rect 94314 59848 94320 59900
rect 94372 59888 94378 59900
rect 96062 59888 96068 59900
rect 94372 59860 96068 59888
rect 94372 59848 94378 59860
rect 96062 59848 96068 59860
rect 96120 59848 96126 59900
rect 97350 59372 97356 59424
rect 97408 59412 97414 59424
rect 116394 59412 116400 59424
rect 97408 59384 116400 59412
rect 97408 59372 97414 59384
rect 116394 59372 116400 59384
rect 116452 59372 116458 59424
rect 214374 59372 214380 59424
rect 214432 59412 214438 59424
rect 217318 59412 217324 59424
rect 214432 59384 217324 59412
rect 214432 59372 214438 59384
rect 217318 59372 217324 59384
rect 217376 59372 217382 59424
rect 216950 59304 216956 59356
rect 217008 59344 217014 59356
rect 227530 59344 227536 59356
rect 217008 59316 227536 59344
rect 217008 59304 217014 59316
rect 227530 59304 227536 59316
rect 227588 59304 227594 59356
rect 224494 59236 224500 59288
rect 224552 59276 224558 59288
rect 227438 59276 227444 59288
rect 224552 59248 227444 59276
rect 224552 59236 224558 59248
rect 227438 59236 227444 59248
rect 227496 59236 227502 59288
rect 214282 58012 214288 58064
rect 214340 58052 214346 58064
rect 217686 58052 217692 58064
rect 214340 58024 217692 58052
rect 214340 58012 214346 58024
rect 217686 58012 217692 58024
rect 217744 58012 217750 58064
rect 94958 57944 94964 57996
rect 95016 57984 95022 57996
rect 116394 57984 116400 57996
rect 95016 57956 116400 57984
rect 95016 57944 95022 57956
rect 116394 57944 116400 57956
rect 116452 57944 116458 57996
rect 214374 57944 214380 57996
rect 214432 57984 214438 57996
rect 217778 57984 217784 57996
rect 214432 57956 217784 57984
rect 214432 57944 214438 57956
rect 217778 57944 217784 57956
rect 217836 57944 217842 57996
rect 94406 57876 94412 57928
rect 94464 57916 94470 57928
rect 97258 57916 97264 57928
rect 94464 57888 97264 57916
rect 94464 57876 94470 57888
rect 97258 57876 97264 57888
rect 97316 57876 97322 57928
rect 216674 57876 216680 57928
rect 216732 57916 216738 57928
rect 227438 57916 227444 57928
rect 216732 57888 227444 57916
rect 216732 57876 216738 57888
rect 227438 57876 227444 57888
rect 227496 57876 227502 57928
rect 224310 57808 224316 57860
rect 224368 57848 224374 57860
rect 227254 57848 227260 57860
rect 224368 57820 227260 57848
rect 224368 57808 224374 57820
rect 227254 57808 227260 57820
rect 227312 57808 227318 57860
rect 213914 56652 213920 56704
rect 213972 56692 213978 56704
rect 216858 56692 216864 56704
rect 213972 56664 216864 56692
rect 213972 56652 213978 56664
rect 216858 56652 216864 56664
rect 216916 56652 216922 56704
rect 95234 56584 95240 56636
rect 95292 56624 95298 56636
rect 116302 56624 116308 56636
rect 95292 56596 116308 56624
rect 95292 56584 95298 56596
rect 116302 56584 116308 56596
rect 116360 56584 116366 56636
rect 214006 56584 214012 56636
rect 214064 56624 214070 56636
rect 216674 56624 216680 56636
rect 214064 56596 216680 56624
rect 214064 56584 214070 56596
rect 216674 56584 216680 56596
rect 216732 56584 216738 56636
rect 216766 56516 216772 56568
rect 216824 56556 216830 56568
rect 227438 56556 227444 56568
rect 216824 56528 227444 56556
rect 216824 56516 216830 56528
rect 227438 56516 227444 56528
rect 227496 56516 227502 56568
rect 224126 56448 224132 56500
rect 224184 56488 224190 56500
rect 227254 56488 227260 56500
rect 224184 56460 227260 56488
rect 224184 56448 224190 56460
rect 227254 56448 227260 56460
rect 227312 56448 227318 56500
rect 94038 55292 94044 55344
rect 94096 55332 94102 55344
rect 116302 55332 116308 55344
rect 94096 55304 116308 55332
rect 94096 55292 94102 55304
rect 116302 55292 116308 55304
rect 116360 55292 116366 55344
rect 94130 55224 94136 55276
rect 94188 55264 94194 55276
rect 116394 55264 116400 55276
rect 94188 55236 116400 55264
rect 94188 55224 94194 55236
rect 116394 55224 116400 55236
rect 116452 55224 116458 55276
rect 215110 55224 215116 55276
rect 215168 55264 215174 55276
rect 227530 55264 227536 55276
rect 215168 55236 227536 55264
rect 215168 55224 215174 55236
rect 227530 55224 227536 55236
rect 227588 55224 227594 55276
rect 217318 55156 217324 55208
rect 217376 55196 217382 55208
rect 217376 55168 224264 55196
rect 217376 55156 217382 55168
rect 224236 55060 224264 55168
rect 224402 55156 224408 55208
rect 224460 55196 224466 55208
rect 227438 55196 227444 55208
rect 224460 55168 227444 55196
rect 224460 55156 224466 55168
rect 227438 55156 227444 55168
rect 227496 55156 227502 55208
rect 226518 55060 226524 55072
rect 224236 55032 226524 55060
rect 226518 55020 226524 55032
rect 226576 55020 226582 55072
rect 94590 54680 94596 54732
rect 94648 54720 94654 54732
rect 96154 54720 96160 54732
rect 94648 54692 96160 54720
rect 94648 54680 94654 54692
rect 96154 54680 96160 54692
rect 96212 54680 96218 54732
rect 214742 53864 214748 53916
rect 214800 53904 214806 53916
rect 226518 53904 226524 53916
rect 214800 53876 226524 53904
rect 214800 53864 214806 53876
rect 226518 53864 226524 53876
rect 226576 53864 226582 53916
rect 94866 53796 94872 53848
rect 94924 53836 94930 53848
rect 116394 53836 116400 53848
rect 94924 53808 116400 53836
rect 94924 53796 94930 53808
rect 116394 53796 116400 53808
rect 116452 53796 116458 53848
rect 215110 53796 215116 53848
rect 215168 53836 215174 53848
rect 226978 53836 226984 53848
rect 215168 53808 226984 53836
rect 215168 53796 215174 53808
rect 226978 53796 226984 53808
rect 227036 53796 227042 53848
rect 217778 53728 217784 53780
rect 217836 53768 217842 53780
rect 227438 53768 227444 53780
rect 217836 53740 227444 53768
rect 217836 53728 217842 53740
rect 227438 53728 227444 53740
rect 227496 53728 227502 53780
rect 217686 53660 217692 53712
rect 217744 53700 217750 53712
rect 227254 53700 227260 53712
rect 217744 53672 227260 53700
rect 217744 53660 217750 53672
rect 227254 53660 227260 53672
rect 227312 53660 227318 53712
rect 215110 52504 215116 52556
rect 215168 52544 215174 52556
rect 226794 52544 226800 52556
rect 215168 52516 226800 52544
rect 215168 52504 215174 52516
rect 226794 52504 226800 52516
rect 226852 52504 226858 52556
rect 94774 52436 94780 52488
rect 94832 52476 94838 52488
rect 116394 52476 116400 52488
rect 94832 52448 116400 52476
rect 94832 52436 94838 52448
rect 116394 52436 116400 52448
rect 116452 52436 116458 52488
rect 214742 52436 214748 52488
rect 214800 52476 214806 52488
rect 226702 52476 226708 52488
rect 214800 52448 226708 52476
rect 214800 52436 214806 52448
rect 226702 52436 226708 52448
rect 226760 52436 226766 52488
rect 95142 52368 95148 52420
rect 95200 52408 95206 52420
rect 97350 52408 97356 52420
rect 95200 52380 97356 52408
rect 95200 52368 95206 52380
rect 97350 52368 97356 52380
rect 97408 52368 97414 52420
rect 216674 52368 216680 52420
rect 216732 52408 216738 52420
rect 227438 52408 227444 52420
rect 216732 52380 227444 52408
rect 216732 52368 216738 52380
rect 227438 52368 227444 52380
rect 227496 52368 227502 52420
rect 216858 52300 216864 52352
rect 216916 52340 216922 52352
rect 227254 52340 227260 52352
rect 216916 52312 227260 52340
rect 216916 52300 216922 52312
rect 227254 52300 227260 52312
rect 227312 52300 227318 52352
rect 215110 51144 215116 51196
rect 215168 51184 215174 51196
rect 226610 51184 226616 51196
rect 215168 51156 226616 51184
rect 215168 51144 215174 51156
rect 226610 51144 226616 51156
rect 226668 51144 226674 51196
rect 95050 51076 95056 51128
rect 95108 51116 95114 51128
rect 115934 51116 115940 51128
rect 95108 51088 115940 51116
rect 95108 51076 95114 51088
rect 115934 51076 115940 51088
rect 115992 51076 115998 51128
rect 214558 51076 214564 51128
rect 214616 51116 214622 51128
rect 226334 51116 226340 51128
rect 214616 51088 226340 51116
rect 214616 51076 214622 51088
rect 226334 51076 226340 51088
rect 226392 51076 226398 51128
rect 214374 49784 214380 49836
rect 214432 49824 214438 49836
rect 227346 49824 227352 49836
rect 214432 49796 227352 49824
rect 214432 49784 214438 49796
rect 227346 49784 227352 49796
rect 227404 49784 227410 49836
rect 95142 49716 95148 49768
rect 95200 49756 95206 49768
rect 116394 49756 116400 49768
rect 95200 49728 116400 49756
rect 95200 49716 95206 49728
rect 116394 49716 116400 49728
rect 116452 49716 116458 49768
rect 215110 49716 215116 49768
rect 215168 49756 215174 49768
rect 227070 49756 227076 49768
rect 215168 49728 227076 49756
rect 215168 49716 215174 49728
rect 227070 49716 227076 49728
rect 227128 49716 227134 49768
rect 94958 48356 94964 48408
rect 95016 48396 95022 48408
rect 116118 48396 116124 48408
rect 95016 48368 116124 48396
rect 95016 48356 95022 48368
rect 116118 48356 116124 48368
rect 116176 48356 116182 48408
rect 94406 48288 94412 48340
rect 94464 48328 94470 48340
rect 116394 48328 116400 48340
rect 94464 48300 116400 48328
rect 94464 48288 94470 48300
rect 116394 48288 116400 48300
rect 116452 48288 116458 48340
rect 215110 48288 215116 48340
rect 215168 48328 215174 48340
rect 227530 48328 227536 48340
rect 215168 48300 227536 48328
rect 215168 48288 215174 48300
rect 227530 48288 227536 48300
rect 227588 48288 227594 48340
rect 214742 46996 214748 47048
rect 214800 47036 214806 47048
rect 227438 47036 227444 47048
rect 214800 47008 227444 47036
rect 214800 46996 214806 47008
rect 227438 46996 227444 47008
rect 227496 46996 227502 47048
rect 94130 46928 94136 46980
rect 94188 46968 94194 46980
rect 116394 46968 116400 46980
rect 94188 46940 116400 46968
rect 94188 46928 94194 46940
rect 116394 46928 116400 46940
rect 116452 46928 116458 46980
rect 214006 46928 214012 46980
rect 214064 46968 214070 46980
rect 227622 46968 227628 46980
rect 214064 46940 227628 46968
rect 214064 46928 214070 46940
rect 227622 46928 227628 46940
rect 227680 46928 227686 46980
rect 215110 45636 215116 45688
rect 215168 45676 215174 45688
rect 226702 45676 226708 45688
rect 215168 45648 226708 45676
rect 215168 45636 215174 45648
rect 226702 45636 226708 45648
rect 226760 45636 226766 45688
rect 93946 45568 93952 45620
rect 94004 45608 94010 45620
rect 116394 45608 116400 45620
rect 94004 45580 116400 45608
rect 94004 45568 94010 45580
rect 116394 45568 116400 45580
rect 116452 45568 116458 45620
rect 215202 45568 215208 45620
rect 215260 45608 215266 45620
rect 227070 45608 227076 45620
rect 215260 45580 227076 45608
rect 215260 45568 215266 45580
rect 227070 45568 227076 45580
rect 227128 45568 227134 45620
rect 215110 44208 215116 44260
rect 215168 44248 215174 44260
rect 227346 44248 227352 44260
rect 215168 44220 227352 44248
rect 215168 44208 215174 44220
rect 227346 44208 227352 44220
rect 227404 44208 227410 44260
rect 95050 44140 95056 44192
rect 95108 44180 95114 44192
rect 116394 44180 116400 44192
rect 95108 44152 116400 44180
rect 95108 44140 95114 44152
rect 116394 44140 116400 44152
rect 116452 44140 116458 44192
rect 214466 44140 214472 44192
rect 214524 44180 214530 44192
rect 227438 44180 227444 44192
rect 214524 44152 227444 44180
rect 214524 44140 214530 44152
rect 227438 44140 227444 44152
rect 227496 44140 227502 44192
rect 94590 42780 94596 42832
rect 94648 42820 94654 42832
rect 115934 42820 115940 42832
rect 94648 42792 115940 42820
rect 94648 42780 94654 42792
rect 115934 42780 115940 42792
rect 115992 42780 115998 42832
rect 214374 42780 214380 42832
rect 214432 42820 214438 42832
rect 226426 42820 226432 42832
rect 214432 42792 226432 42820
rect 214432 42780 214438 42792
rect 226426 42780 226432 42792
rect 226484 42780 226490 42832
rect 215110 41488 215116 41540
rect 215168 41528 215174 41540
rect 226610 41528 226616 41540
rect 215168 41500 226616 41528
rect 215168 41488 215174 41500
rect 226610 41488 226616 41500
rect 226668 41488 226674 41540
rect 95142 41420 95148 41472
rect 95200 41460 95206 41472
rect 116394 41460 116400 41472
rect 95200 41432 116400 41460
rect 95200 41420 95206 41432
rect 116394 41420 116400 41432
rect 116452 41420 116458 41472
rect 214098 41420 214104 41472
rect 214156 41460 214162 41472
rect 226334 41460 226340 41472
rect 214156 41432 226340 41460
rect 214156 41420 214162 41432
rect 226334 41420 226340 41432
rect 226392 41420 226398 41472
rect 560938 41352 560944 41404
rect 560996 41392 561002 41404
rect 580166 41392 580172 41404
rect 560996 41364 580172 41392
rect 560996 41352 561002 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 94498 40128 94504 40180
rect 94556 40168 94562 40180
rect 116302 40168 116308 40180
rect 94556 40140 116308 40168
rect 94556 40128 94562 40140
rect 116302 40128 116308 40140
rect 116360 40128 116366 40180
rect 215110 40128 215116 40180
rect 215168 40168 215174 40180
rect 226886 40168 226892 40180
rect 215168 40140 226892 40168
rect 215168 40128 215174 40140
rect 226886 40128 226892 40140
rect 226944 40128 226950 40180
rect 95050 40060 95056 40112
rect 95108 40100 95114 40112
rect 116394 40100 116400 40112
rect 95108 40072 116400 40100
rect 95108 40060 95114 40072
rect 116394 40060 116400 40072
rect 116452 40060 116458 40112
rect 214650 40060 214656 40112
rect 214708 40100 214714 40112
rect 227070 40100 227076 40112
rect 214708 40072 227076 40100
rect 214708 40060 214714 40072
rect 227070 40060 227076 40072
rect 227128 40060 227134 40112
rect 214466 38700 214472 38752
rect 214524 38740 214530 38752
rect 227438 38740 227444 38752
rect 214524 38712 227444 38740
rect 214524 38700 214530 38712
rect 227438 38700 227444 38712
rect 227496 38700 227502 38752
rect 94590 38632 94596 38684
rect 94648 38672 94654 38684
rect 116394 38672 116400 38684
rect 94648 38644 116400 38672
rect 94648 38632 94654 38644
rect 116394 38632 116400 38644
rect 116452 38632 116458 38684
rect 215110 38632 215116 38684
rect 215168 38672 215174 38684
rect 227530 38672 227536 38684
rect 215168 38644 227536 38672
rect 215168 38632 215174 38644
rect 227530 38632 227536 38644
rect 227588 38632 227594 38684
rect 93854 37272 93860 37324
rect 93912 37312 93918 37324
rect 116394 37312 116400 37324
rect 93912 37284 116400 37312
rect 93912 37272 93918 37284
rect 116394 37272 116400 37284
rect 116452 37272 116458 37324
rect 215110 37272 215116 37324
rect 215168 37312 215174 37324
rect 227438 37312 227444 37324
rect 215168 37284 227444 37312
rect 215168 37272 215174 37284
rect 227438 37272 227444 37284
rect 227496 37272 227502 37324
rect 214558 35980 214564 36032
rect 214616 36020 214622 36032
rect 227530 36020 227536 36032
rect 214616 35992 227536 36020
rect 214616 35980 214622 35992
rect 227530 35980 227536 35992
rect 227588 35980 227594 36032
rect 93946 35912 93952 35964
rect 94004 35952 94010 35964
rect 116394 35952 116400 35964
rect 94004 35924 116400 35952
rect 94004 35912 94010 35924
rect 116394 35912 116400 35924
rect 116452 35912 116458 35964
rect 215110 35912 215116 35964
rect 215168 35952 215174 35964
rect 227438 35952 227444 35964
rect 215168 35924 227444 35952
rect 215168 35912 215174 35924
rect 227438 35912 227444 35924
rect 227496 35912 227502 35964
rect 3418 35844 3424 35896
rect 3476 35884 3482 35896
rect 9122 35884 9128 35896
rect 3476 35856 9128 35884
rect 3476 35844 3482 35856
rect 9122 35844 9128 35856
rect 9180 35844 9186 35896
rect 215110 34552 215116 34604
rect 215168 34592 215174 34604
rect 227346 34592 227352 34604
rect 215168 34564 227352 34592
rect 215168 34552 215174 34564
rect 227346 34552 227352 34564
rect 227404 34552 227410 34604
rect 95142 34484 95148 34536
rect 95200 34524 95206 34536
rect 116394 34524 116400 34536
rect 95200 34496 116400 34524
rect 95200 34484 95206 34496
rect 116394 34484 116400 34496
rect 116452 34484 116458 34536
rect 214650 34484 214656 34536
rect 214708 34524 214714 34536
rect 227438 34524 227444 34536
rect 214708 34496 227444 34524
rect 214708 34484 214714 34496
rect 227438 34484 227444 34496
rect 227496 34484 227502 34536
rect 215110 33192 215116 33244
rect 215168 33232 215174 33244
rect 227530 33232 227536 33244
rect 215168 33204 227536 33232
rect 215168 33192 215174 33204
rect 227530 33192 227536 33204
rect 227588 33192 227594 33244
rect 95142 33124 95148 33176
rect 95200 33164 95206 33176
rect 116302 33164 116308 33176
rect 95200 33136 116308 33164
rect 95200 33124 95206 33136
rect 116302 33124 116308 33136
rect 116360 33124 116366 33176
rect 214558 33124 214564 33176
rect 214616 33164 214622 33176
rect 227438 33164 227444 33176
rect 214616 33136 227444 33164
rect 214616 33124 214622 33136
rect 227438 33124 227444 33136
rect 227496 33124 227502 33176
rect 213914 32512 213920 32564
rect 213972 32552 213978 32564
rect 215938 32552 215944 32564
rect 213972 32524 215944 32552
rect 213972 32512 213978 32524
rect 215938 32512 215944 32524
rect 215996 32512 216002 32564
rect 95142 32376 95148 32428
rect 95200 32416 95206 32428
rect 116394 32416 116400 32428
rect 95200 32388 116400 32416
rect 95200 32376 95206 32388
rect 116394 32376 116400 32388
rect 116452 32376 116458 32428
rect 215110 32376 215116 32428
rect 215168 32416 215174 32428
rect 227438 32416 227444 32428
rect 215168 32388 227444 32416
rect 215168 32376 215174 32388
rect 227438 32376 227444 32388
rect 227496 32376 227502 32428
rect 71682 31764 71688 31816
rect 71740 31804 71746 31816
rect 116394 31804 116400 31816
rect 71740 31776 116400 31804
rect 71740 31764 71746 31776
rect 116394 31764 116400 31776
rect 116452 31764 116458 31816
rect 29914 30268 29920 30320
rect 29972 30308 29978 30320
rect 32306 30308 32312 30320
rect 29972 30280 32312 30308
rect 29972 30268 29978 30280
rect 32306 30268 32312 30280
rect 32364 30308 32370 30320
rect 119982 30308 119988 30320
rect 32364 30280 119988 30308
rect 32364 30268 32370 30280
rect 119982 30268 119988 30280
rect 120040 30308 120046 30320
rect 231946 30308 231952 30320
rect 120040 30280 231952 30308
rect 120040 30268 120046 30280
rect 231946 30268 231952 30280
rect 232004 30308 232010 30320
rect 284570 30308 284576 30320
rect 232004 30280 284576 30308
rect 232004 30268 232010 30280
rect 284570 30268 284576 30280
rect 284628 30268 284634 30320
rect 115842 30200 115848 30252
rect 115900 30240 115906 30252
rect 203242 30240 203248 30252
rect 115900 30212 203248 30240
rect 115900 30200 115906 30212
rect 203242 30200 203248 30212
rect 203300 30200 203306 30252
rect 107562 30132 107568 30184
rect 107620 30172 107626 30184
rect 198090 30172 198096 30184
rect 107620 30144 198096 30172
rect 107620 30132 107626 30144
rect 198090 30132 198096 30144
rect 198148 30132 198154 30184
rect 51718 30064 51724 30116
rect 51776 30104 51782 30116
rect 143350 30104 143356 30116
rect 51776 30076 143356 30104
rect 51776 30064 51782 30076
rect 143350 30064 143356 30076
rect 143408 30064 143414 30116
rect 57238 29996 57244 30048
rect 57296 30036 57302 30048
rect 148594 30036 148600 30048
rect 57296 30008 148600 30036
rect 57296 29996 57302 30008
rect 148594 29996 148600 30008
rect 148652 29996 148658 30048
rect 32398 29928 32404 29980
rect 32456 29968 32462 29980
rect 134702 29968 134708 29980
rect 32456 29940 134708 29968
rect 32456 29928 32462 29940
rect 134702 29928 134708 29940
rect 134760 29928 134766 29980
rect 28258 29860 28264 29912
rect 28316 29900 28322 29912
rect 131206 29900 131212 29912
rect 28316 29872 131212 29900
rect 28316 29860 28322 29872
rect 131206 29860 131212 29872
rect 131264 29860 131270 29912
rect 164878 29860 164884 29912
rect 164936 29900 164942 29912
rect 185026 29900 185032 29912
rect 164936 29872 185032 29900
rect 164936 29860 164942 29872
rect 185026 29860 185032 29872
rect 185084 29860 185090 29912
rect 24118 29792 24124 29844
rect 24176 29832 24182 29844
rect 127710 29832 127716 29844
rect 24176 29804 127716 29832
rect 24176 29792 24182 29804
rect 127710 29792 127716 29804
rect 127768 29792 127774 29844
rect 159358 29792 159364 29844
rect 159416 29832 159422 29844
rect 179782 29832 179788 29844
rect 159416 29804 179788 29832
rect 159416 29792 159422 29804
rect 179782 29792 179788 29804
rect 179840 29792 179846 29844
rect 31018 29724 31024 29776
rect 31076 29764 31082 29776
rect 140774 29764 140780 29776
rect 31076 29736 140780 29764
rect 31076 29724 31082 29736
rect 140774 29724 140780 29736
rect 140832 29724 140838 29776
rect 166258 29724 166264 29776
rect 166316 29764 166322 29776
rect 190270 29764 190276 29776
rect 166316 29736 190276 29764
rect 166316 29724 166322 29736
rect 190270 29724 190276 29736
rect 190328 29724 190334 29776
rect 22738 29656 22744 29708
rect 22796 29696 22802 29708
rect 133782 29696 133788 29708
rect 22796 29668 133788 29696
rect 22796 29656 22802 29668
rect 133782 29656 133788 29668
rect 133840 29656 133846 29708
rect 169018 29656 169024 29708
rect 169076 29696 169082 29708
rect 195422 29696 195428 29708
rect 169076 29668 195428 29696
rect 169076 29656 169082 29668
rect 195422 29656 195428 29668
rect 195480 29656 195486 29708
rect 25498 29588 25504 29640
rect 25556 29628 25562 29640
rect 137278 29628 137284 29640
rect 25556 29600 137284 29628
rect 25556 29588 25562 29600
rect 137278 29588 137284 29600
rect 137336 29588 137342 29640
rect 171778 29588 171784 29640
rect 171836 29628 171842 29640
rect 200666 29628 200672 29640
rect 171836 29600 200672 29628
rect 171836 29588 171842 29600
rect 200666 29588 200672 29600
rect 200724 29588 200730 29640
rect 118602 29520 118608 29572
rect 118660 29560 118666 29572
rect 205818 29560 205824 29572
rect 118660 29532 205824 29560
rect 118660 29520 118666 29532
rect 205818 29520 205824 29532
rect 205876 29520 205882 29572
rect 61378 29452 61384 29504
rect 61436 29492 61442 29504
rect 123386 29492 123392 29504
rect 61436 29464 123392 29492
rect 61436 29452 61442 29464
rect 123386 29452 123392 29464
rect 123444 29452 123450 29504
rect 123478 29452 123484 29504
rect 123536 29492 123542 29504
rect 208486 29492 208492 29504
rect 123536 29464 208492 29492
rect 123536 29452 123542 29464
rect 208486 29452 208492 29464
rect 208544 29452 208550 29504
rect 69658 29384 69664 29436
rect 69716 29424 69722 29436
rect 124306 29424 124312 29436
rect 69716 29396 124312 29424
rect 69716 29384 69722 29396
rect 124306 29384 124312 29396
rect 124364 29384 124370 29436
rect 126238 29384 126244 29436
rect 126296 29424 126302 29436
rect 211062 29424 211068 29436
rect 126296 29396 211068 29424
rect 126296 29384 126302 29396
rect 211062 29384 211068 29396
rect 211120 29384 211126 29436
rect 142798 28976 142804 29028
rect 142856 29016 142862 29028
rect 146018 29016 146024 29028
rect 142856 28988 146024 29016
rect 142856 28976 142862 28988
rect 146018 28976 146024 28988
rect 146076 28976 146082 29028
rect 199010 28908 199016 28960
rect 199068 28948 199074 28960
rect 199102 28948 199108 28960
rect 199068 28920 199108 28948
rect 199068 28908 199074 28920
rect 199102 28908 199108 28920
rect 199160 28908 199166 28960
rect 135254 28840 135260 28892
rect 135312 28880 135318 28892
rect 136174 28880 136180 28892
rect 135312 28852 136180 28880
rect 135312 28840 135318 28852
rect 136174 28840 136180 28852
rect 136232 28840 136238 28892
rect 138106 28840 138112 28892
rect 138164 28880 138170 28892
rect 138750 28880 138756 28892
rect 138164 28852 138756 28880
rect 138164 28840 138170 28852
rect 138750 28840 138756 28852
rect 138808 28840 138814 28892
rect 113082 28364 113088 28416
rect 113140 28404 113146 28416
rect 201494 28404 201500 28416
rect 113140 28376 201500 28404
rect 113140 28364 113146 28376
rect 201494 28364 201500 28376
rect 201552 28364 201558 28416
rect 50982 28296 50988 28348
rect 51040 28336 51046 28348
rect 156414 28336 156420 28348
rect 51040 28308 156420 28336
rect 51040 28296 51046 28308
rect 156414 28296 156420 28308
rect 156472 28296 156478 28348
rect 8938 28228 8944 28280
rect 8996 28268 9002 28280
rect 121638 28268 121644 28280
rect 8996 28240 121644 28268
rect 8996 28228 9002 28240
rect 121638 28228 121644 28240
rect 121696 28228 121702 28280
rect 125502 28228 125508 28280
rect 125560 28268 125566 28280
rect 210234 28268 210240 28280
rect 125560 28240 210240 28268
rect 125560 28228 125566 28240
rect 210234 28228 210240 28240
rect 210292 28228 210298 28280
rect 117222 27072 117228 27124
rect 117280 27112 117286 27124
rect 204162 27112 204168 27124
rect 117280 27084 204168 27112
rect 117280 27072 117286 27084
rect 204162 27072 204168 27084
rect 204220 27072 204226 27124
rect 107470 27004 107476 27056
rect 107528 27044 107534 27056
rect 197170 27044 197176 27056
rect 107528 27016 197176 27044
rect 107528 27004 107534 27016
rect 197170 27004 197176 27016
rect 197228 27004 197234 27056
rect 62022 26936 62028 26988
rect 62080 26976 62086 26988
rect 164234 26976 164240 26988
rect 62080 26948 164240 26976
rect 62080 26936 62086 26948
rect 164234 26936 164240 26948
rect 164292 26936 164298 26988
rect 11698 26868 11704 26920
rect 11756 26908 11762 26920
rect 125134 26908 125140 26920
rect 11756 26880 125140 26908
rect 11756 26868 11762 26880
rect 125134 26868 125140 26880
rect 125192 26868 125198 26920
rect 125870 26732 125876 26784
rect 125928 26772 125934 26784
rect 126606 26772 126612 26784
rect 125928 26744 126612 26772
rect 125928 26732 125934 26744
rect 126606 26732 126612 26744
rect 126664 26732 126670 26784
rect 154574 26732 154580 26784
rect 154632 26772 154638 26784
rect 155126 26772 155132 26784
rect 154632 26744 155132 26772
rect 154632 26732 154638 26744
rect 155126 26732 155132 26744
rect 155184 26732 155190 26784
rect 186498 26256 186504 26308
rect 186556 26296 186562 26308
rect 187326 26296 187332 26308
rect 186556 26268 187332 26296
rect 186556 26256 186562 26268
rect 187326 26256 187332 26268
rect 187384 26256 187390 26308
rect 85482 25644 85488 25696
rect 85540 25684 85546 25696
rect 181530 25684 181536 25696
rect 85540 25656 181536 25684
rect 85540 25644 85546 25656
rect 181530 25644 181536 25656
rect 181588 25644 181594 25696
rect 68922 25576 68928 25628
rect 68980 25616 68986 25628
rect 169386 25616 169392 25628
rect 68980 25588 169392 25616
rect 68980 25576 68986 25588
rect 169386 25576 169392 25588
rect 169444 25576 169450 25628
rect 59262 25508 59268 25560
rect 59320 25548 59326 25560
rect 161566 25548 161572 25560
rect 59320 25520 161572 25548
rect 59320 25508 59326 25520
rect 161566 25508 161572 25520
rect 161624 25508 161630 25560
rect 96522 24216 96528 24268
rect 96580 24256 96586 24268
rect 189166 24256 189172 24268
rect 96580 24228 189172 24256
rect 96580 24216 96586 24228
rect 189166 24216 189172 24228
rect 189224 24216 189230 24268
rect 63402 24148 63408 24200
rect 63460 24188 63466 24200
rect 164234 24188 164240 24200
rect 63460 24160 164240 24188
rect 63460 24148 63466 24160
rect 164234 24148 164240 24160
rect 164292 24148 164298 24200
rect 57882 24080 57888 24132
rect 57940 24120 57946 24132
rect 161474 24120 161480 24132
rect 57940 24092 161480 24120
rect 57940 24080 57946 24092
rect 161474 24080 161480 24092
rect 161532 24080 161538 24132
rect 182174 23740 182180 23792
rect 182232 23780 182238 23792
rect 182910 23780 182916 23792
rect 182232 23752 182916 23780
rect 182232 23740 182238 23752
rect 182910 23740 182916 23752
rect 182968 23740 182974 23792
rect 89622 22856 89628 22908
rect 89680 22896 89686 22908
rect 184198 22896 184204 22908
rect 89680 22868 184204 22896
rect 89680 22856 89686 22868
rect 184198 22856 184204 22868
rect 184256 22856 184262 22908
rect 64782 22788 64788 22840
rect 64840 22828 64846 22840
rect 165890 22828 165896 22840
rect 64840 22800 165896 22828
rect 64840 22788 64846 22800
rect 165890 22788 165896 22800
rect 165948 22788 165954 22840
rect 56502 22720 56508 22772
rect 56560 22760 56566 22772
rect 158806 22760 158812 22772
rect 56560 22732 158812 22760
rect 56560 22720 56566 22732
rect 158806 22720 158812 22732
rect 158864 22720 158870 22772
rect 175458 22040 175464 22092
rect 175516 22040 175522 22092
rect 175476 22012 175504 22040
rect 175550 22012 175556 22024
rect 175476 21984 175556 22012
rect 175550 21972 175556 21984
rect 175608 21972 175614 22024
rect 100662 21564 100668 21616
rect 100720 21604 100726 21616
rect 192110 21604 192116 21616
rect 100720 21576 192116 21604
rect 100720 21564 100726 21576
rect 192110 21564 192116 21576
rect 192168 21564 192174 21616
rect 82722 21496 82728 21548
rect 82780 21536 82786 21548
rect 178126 21536 178132 21548
rect 82780 21508 178132 21536
rect 82780 21496 82786 21508
rect 178126 21496 178132 21508
rect 178184 21496 178190 21548
rect 72970 21428 72976 21480
rect 73028 21468 73034 21480
rect 171226 21468 171232 21480
rect 73028 21440 171232 21468
rect 73028 21428 73034 21440
rect 171226 21428 171232 21440
rect 171284 21428 171290 21480
rect 52362 21360 52368 21412
rect 52420 21400 52426 21412
rect 156046 21400 156052 21412
rect 52420 21372 156052 21400
rect 52420 21360 52426 21372
rect 156046 21360 156052 21372
rect 156104 21360 156110 21412
rect 119982 20136 119988 20188
rect 120040 20176 120046 20188
rect 205818 20176 205824 20188
rect 120040 20148 205824 20176
rect 120040 20136 120046 20148
rect 205818 20136 205824 20148
rect 205876 20136 205882 20188
rect 75822 20068 75828 20120
rect 75880 20108 75886 20120
rect 173894 20108 173900 20120
rect 75880 20080 173900 20108
rect 75880 20068 75886 20080
rect 173894 20068 173900 20080
rect 173952 20068 173958 20120
rect 48222 20000 48228 20052
rect 48280 20040 48286 20052
rect 154666 20040 154672 20052
rect 48280 20012 154672 20040
rect 48280 20000 48286 20012
rect 154666 20000 154672 20012
rect 154724 20000 154730 20052
rect 10962 19932 10968 19984
rect 11020 19972 11026 19984
rect 125870 19972 125876 19984
rect 11020 19944 125876 19972
rect 11020 19932 11026 19944
rect 125870 19932 125876 19944
rect 125928 19932 125934 19984
rect 199102 19320 199108 19372
rect 199160 19360 199166 19372
rect 199194 19360 199200 19372
rect 199160 19332 199200 19360
rect 199160 19320 199166 19332
rect 199194 19320 199200 19332
rect 199252 19320 199258 19372
rect 148042 19252 148048 19304
rect 148100 19292 148106 19304
rect 151998 19292 152004 19304
rect 148100 19264 152004 19292
rect 148100 19252 148106 19264
rect 151998 19252 152004 19264
rect 152056 19252 152062 19304
rect 208486 19252 208492 19304
rect 208544 19292 208550 19304
rect 208670 19292 208676 19304
rect 208544 19264 208676 19292
rect 208544 19252 208550 19264
rect 208670 19252 208676 19264
rect 208728 19252 208734 19304
rect 79962 18640 79968 18692
rect 80020 18680 80026 18692
rect 176654 18680 176660 18692
rect 80020 18652 176660 18680
rect 80020 18640 80026 18652
rect 176654 18640 176660 18652
rect 176712 18640 176718 18692
rect 30282 18572 30288 18624
rect 30340 18612 30346 18624
rect 140866 18612 140872 18624
rect 30340 18584 140872 18612
rect 30340 18572 30346 18584
rect 140866 18572 140872 18584
rect 140924 18572 140930 18624
rect 129642 17960 129648 18012
rect 129700 18000 129706 18012
rect 406470 18000 406476 18012
rect 129700 17972 406476 18000
rect 129700 17960 129706 17972
rect 406470 17960 406476 17972
rect 406528 17960 406534 18012
rect 414382 17620 414388 17672
rect 414440 17660 414446 17672
rect 414440 17632 440556 17660
rect 414440 17620 414446 17632
rect 440528 17524 440556 17632
rect 440528 17496 449940 17524
rect 414290 17416 414296 17468
rect 414348 17456 414354 17468
rect 449912 17456 449940 17496
rect 414348 17428 430712 17456
rect 449912 17428 459508 17456
rect 414348 17416 414354 17428
rect 287054 17348 287060 17400
rect 287112 17388 287118 17400
rect 296530 17388 296536 17400
rect 287112 17360 296536 17388
rect 287112 17348 287118 17360
rect 296530 17348 296536 17360
rect 296588 17348 296594 17400
rect 393958 17348 393964 17400
rect 394016 17388 394022 17400
rect 410518 17388 410524 17400
rect 394016 17360 410524 17388
rect 394016 17348 394022 17360
rect 410518 17348 410524 17360
rect 410576 17348 410582 17400
rect 410610 17348 410616 17400
rect 410668 17388 410674 17400
rect 410668 17360 418844 17388
rect 410668 17348 410674 17360
rect 38562 17280 38568 17332
rect 38620 17320 38626 17332
rect 147766 17320 147772 17332
rect 38620 17292 147772 17320
rect 38620 17280 38626 17292
rect 147766 17280 147772 17292
rect 147824 17280 147830 17332
rect 246942 17280 246948 17332
rect 247000 17320 247006 17332
rect 270494 17320 270500 17332
rect 247000 17292 270500 17320
rect 247000 17280 247006 17292
rect 270494 17280 270500 17292
rect 270552 17280 270558 17332
rect 300762 17280 300768 17332
rect 300820 17320 300826 17332
rect 414382 17320 414388 17332
rect 300820 17292 414388 17320
rect 300820 17280 300826 17292
rect 414382 17280 414388 17292
rect 414440 17280 414446 17332
rect 17862 17212 17868 17264
rect 17920 17252 17926 17264
rect 131298 17252 131304 17264
rect 17920 17224 131304 17252
rect 17920 17212 17926 17224
rect 131298 17212 131304 17224
rect 131356 17212 131362 17264
rect 278682 17212 278688 17264
rect 278740 17252 278746 17264
rect 414290 17252 414296 17264
rect 278740 17224 414296 17252
rect 278740 17212 278746 17224
rect 414290 17212 414296 17224
rect 414348 17212 414354 17264
rect 418816 17252 418844 17360
rect 430684 17252 430712 17428
rect 459480 17388 459508 17428
rect 459480 17360 462912 17388
rect 462884 17320 462912 17360
rect 462884 17292 468984 17320
rect 468956 17252 468984 17292
rect 418816 17224 427400 17252
rect 430684 17224 439636 17252
rect 267642 17144 267648 17196
rect 267700 17184 267706 17196
rect 393958 17184 393964 17196
rect 267700 17156 393964 17184
rect 267700 17144 267706 17156
rect 393958 17144 393964 17156
rect 394016 17144 394022 17196
rect 427372 17184 427400 17224
rect 439608 17184 439636 17224
rect 440252 17224 449940 17252
rect 468956 17224 470088 17252
rect 440252 17184 440280 17224
rect 427372 17156 439544 17184
rect 439608 17156 440280 17184
rect 449912 17184 449940 17224
rect 449912 17156 459508 17184
rect 270586 17076 270592 17128
rect 270644 17116 270650 17128
rect 287054 17116 287060 17128
rect 270644 17088 287060 17116
rect 270644 17076 270650 17088
rect 287054 17076 287060 17088
rect 287112 17076 287118 17128
rect 296530 17076 296536 17128
rect 296588 17116 296594 17128
rect 296588 17088 439452 17116
rect 296588 17076 296594 17088
rect 439424 17060 439452 17088
rect 217962 17008 217968 17060
rect 218020 17048 218026 17060
rect 424594 17048 424600 17060
rect 218020 17020 424600 17048
rect 218020 17008 218026 17020
rect 424594 17008 424600 17020
rect 424652 17008 424658 17060
rect 439406 17008 439412 17060
rect 439464 17008 439470 17060
rect 439516 17048 439544 17156
rect 459480 17116 459508 17156
rect 459480 17088 462636 17116
rect 462608 17060 462636 17088
rect 470060 17060 470088 17224
rect 459094 17048 459100 17060
rect 439516 17020 459100 17048
rect 459094 17008 459100 17020
rect 459152 17008 459158 17060
rect 462590 17008 462596 17060
rect 462648 17008 462654 17060
rect 470042 17008 470048 17060
rect 470100 17008 470106 17060
rect 202782 16940 202788 16992
rect 202840 16980 202846 16992
rect 418706 16980 418712 16992
rect 202840 16952 418712 16980
rect 202840 16940 202846 16952
rect 418706 16940 418712 16952
rect 418764 16940 418770 16992
rect 425606 16940 425612 16992
rect 425664 16980 425670 16992
rect 425664 16952 430160 16980
rect 425664 16940 425670 16952
rect 193122 16872 193128 16924
rect 193180 16912 193186 16924
rect 430022 16912 430028 16924
rect 193180 16884 430028 16912
rect 193180 16872 193186 16884
rect 430022 16872 430028 16884
rect 430080 16872 430086 16924
rect 184842 16804 184848 16856
rect 184900 16844 184906 16856
rect 429930 16844 429936 16856
rect 184900 16816 429936 16844
rect 184900 16804 184906 16816
rect 429930 16804 429936 16816
rect 429988 16804 429994 16856
rect 164142 16736 164148 16788
rect 164200 16776 164206 16788
rect 425790 16776 425796 16788
rect 164200 16748 425796 16776
rect 164200 16736 164206 16748
rect 425790 16736 425796 16748
rect 425848 16736 425854 16788
rect 430132 16776 430160 16952
rect 430132 16748 430896 16776
rect 160002 16668 160008 16720
rect 160060 16708 160066 16720
rect 424226 16708 424232 16720
rect 160060 16680 424232 16708
rect 160060 16668 160066 16680
rect 424226 16668 424232 16680
rect 424284 16668 424290 16720
rect 430868 16708 430896 16748
rect 435358 16736 435364 16788
rect 435416 16776 435422 16788
rect 442994 16776 443000 16788
rect 435416 16748 443000 16776
rect 435416 16736 435422 16748
rect 442994 16736 443000 16748
rect 443052 16736 443058 16788
rect 438394 16708 438400 16720
rect 430868 16680 438400 16708
rect 438394 16668 438400 16680
rect 438452 16668 438458 16720
rect 132402 16600 132408 16652
rect 132460 16640 132466 16652
rect 415394 16640 415400 16652
rect 132460 16612 415400 16640
rect 132460 16600 132466 16612
rect 415394 16600 415400 16612
rect 415452 16600 415458 16652
rect 418706 16600 418712 16652
rect 418764 16640 418770 16652
rect 425606 16640 425612 16652
rect 418764 16612 425612 16640
rect 418764 16600 418770 16612
rect 425606 16600 425612 16612
rect 425664 16600 425670 16652
rect 429930 16600 429936 16652
rect 429988 16640 429994 16652
rect 432690 16640 432696 16652
rect 429988 16612 432696 16640
rect 429988 16600 429994 16612
rect 432690 16600 432696 16612
rect 432748 16600 432754 16652
rect 430022 16532 430028 16584
rect 430080 16572 430086 16584
rect 434990 16572 434996 16584
rect 430080 16544 434996 16572
rect 430080 16532 430086 16544
rect 434990 16532 434996 16544
rect 435048 16532 435054 16584
rect 479058 16396 479064 16448
rect 479116 16436 479122 16448
rect 479794 16436 479800 16448
rect 479116 16408 479800 16436
rect 479116 16396 479122 16408
rect 479794 16396 479800 16408
rect 479852 16396 479858 16448
rect 534350 16396 534356 16448
rect 534408 16436 534414 16448
rect 534994 16436 535000 16448
rect 534408 16408 535000 16436
rect 534408 16396 534414 16408
rect 534994 16396 535000 16408
rect 535052 16396 535058 16448
rect 187602 16192 187608 16244
rect 187660 16232 187666 16244
rect 433702 16232 433708 16244
rect 187660 16204 433708 16232
rect 187660 16192 187666 16204
rect 433702 16192 433708 16204
rect 433760 16192 433766 16244
rect 180702 16124 180708 16176
rect 180760 16164 180766 16176
rect 431402 16164 431408 16176
rect 180760 16136 431408 16164
rect 180760 16124 180766 16136
rect 431402 16124 431408 16136
rect 431460 16124 431466 16176
rect 387702 16056 387708 16108
rect 387760 16096 387766 16108
rect 498102 16096 498108 16108
rect 387760 16068 498108 16096
rect 387760 16056 387766 16068
rect 498102 16056 498108 16068
rect 498160 16056 498166 16108
rect 376202 15988 376208 16040
rect 376260 16028 376266 16040
rect 494698 16028 494704 16040
rect 376260 16000 494704 16028
rect 376260 15988 376266 16000
rect 494698 15988 494704 16000
rect 494756 15988 494762 16040
rect 55122 15920 55128 15972
rect 55180 15960 55186 15972
rect 158714 15960 158720 15972
rect 55180 15932 158720 15960
rect 55180 15920 55186 15932
rect 158714 15920 158720 15932
rect 158772 15920 158778 15972
rect 311158 15920 311164 15972
rect 311216 15960 311222 15972
rect 450998 15960 451004 15972
rect 311216 15932 451004 15960
rect 311216 15920 311222 15932
rect 450998 15920 451004 15932
rect 451056 15920 451062 15972
rect 34422 15852 34428 15904
rect 34480 15892 34486 15904
rect 143534 15892 143540 15904
rect 34480 15864 143540 15892
rect 34480 15852 34486 15864
rect 143534 15852 143540 15864
rect 143592 15852 143598 15904
rect 339402 15852 339408 15904
rect 339460 15892 339466 15904
rect 482370 15892 482376 15904
rect 339460 15864 482376 15892
rect 339460 15852 339466 15864
rect 482370 15852 482376 15864
rect 482428 15852 482434 15904
rect 326338 15784 326344 15836
rect 326396 15824 326402 15836
rect 471698 15824 471704 15836
rect 326396 15796 471704 15824
rect 326396 15784 326402 15796
rect 471698 15784 471704 15796
rect 471756 15784 471762 15836
rect 333238 15716 333244 15768
rect 333296 15756 333302 15768
rect 479702 15756 479708 15768
rect 333296 15728 479708 15756
rect 333296 15716 333302 15728
rect 479702 15716 479708 15728
rect 479760 15716 479766 15768
rect 282178 15648 282184 15700
rect 282236 15688 282242 15700
rect 439498 15688 439504 15700
rect 282236 15660 439504 15688
rect 282236 15648 282242 15660
rect 439498 15648 439504 15660
rect 439556 15648 439562 15700
rect 275278 15580 275284 15632
rect 275336 15620 275342 15632
rect 437198 15620 437204 15632
rect 275336 15592 437204 15620
rect 275336 15580 275342 15592
rect 437198 15580 437204 15592
rect 437256 15580 437262 15632
rect 280062 15512 280068 15564
rect 280120 15552 280126 15564
rect 463234 15552 463240 15564
rect 280120 15524 463240 15552
rect 280120 15512 280126 15524
rect 463234 15512 463240 15524
rect 463292 15512 463298 15564
rect 259362 15444 259368 15496
rect 259420 15484 259426 15496
rect 456702 15484 456708 15496
rect 259420 15456 456708 15484
rect 259420 15444 259426 15456
rect 456702 15444 456708 15456
rect 456760 15444 456766 15496
rect 248322 15376 248328 15428
rect 248380 15416 248386 15428
rect 453298 15416 453304 15428
rect 248380 15388 453304 15416
rect 248380 15376 248386 15388
rect 453298 15376 453304 15388
rect 453356 15376 453362 15428
rect 234522 15308 234528 15360
rect 234580 15348 234586 15360
rect 448698 15348 448704 15360
rect 234580 15320 448704 15348
rect 234580 15308 234586 15320
rect 448698 15308 448704 15320
rect 448756 15308 448762 15360
rect 405642 15240 405648 15292
rect 405700 15280 405706 15292
rect 503898 15280 503904 15292
rect 405700 15252 503904 15280
rect 405700 15240 405706 15252
rect 503898 15240 503904 15252
rect 503956 15240 503962 15292
rect 398742 15172 398748 15224
rect 398800 15212 398806 15224
rect 501598 15212 501604 15224
rect 398800 15184 501604 15212
rect 398800 15172 398806 15184
rect 501598 15172 501604 15184
rect 501656 15172 501662 15224
rect 368658 15104 368664 15156
rect 368716 15144 368722 15156
rect 476298 15144 476304 15156
rect 368716 15116 476304 15144
rect 368716 15104 368722 15116
rect 476298 15104 476304 15116
rect 476356 15104 476362 15156
rect 525058 15104 525064 15156
rect 525116 15144 525122 15156
rect 534534 15144 534540 15156
rect 525116 15116 534540 15144
rect 525116 15104 525122 15116
rect 534534 15104 534540 15116
rect 534592 15104 534598 15156
rect 535362 15104 535368 15156
rect 535420 15144 535426 15156
rect 545666 15144 545672 15156
rect 535420 15116 545672 15144
rect 535420 15104 535426 15116
rect 545666 15104 545672 15116
rect 545724 15104 545730 15156
rect 390462 15036 390468 15088
rect 390520 15076 390526 15088
rect 498838 15076 498844 15088
rect 390520 15048 498844 15076
rect 390520 15036 390526 15048
rect 498838 15036 498844 15048
rect 498896 15036 498902 15088
rect 527910 15036 527916 15088
rect 527968 15076 527974 15088
rect 539134 15076 539140 15088
rect 527968 15048 539140 15076
rect 527968 15036 527974 15048
rect 539134 15036 539140 15048
rect 539192 15036 539198 15088
rect 368382 14968 368388 15020
rect 368440 15008 368446 15020
rect 491938 15008 491944 15020
rect 368440 14980 491944 15008
rect 368440 14968 368446 14980
rect 491938 14968 491944 14980
rect 491996 14968 492002 15020
rect 530578 14968 530584 15020
rect 530636 15008 530642 15020
rect 541434 15008 541440 15020
rect 530636 14980 541440 15008
rect 530636 14968 530642 14980
rect 541434 14968 541440 14980
rect 541492 14968 541498 15020
rect 357342 14900 357348 14952
rect 357400 14940 357406 14952
rect 488534 14940 488540 14952
rect 357400 14912 488540 14940
rect 357400 14900 357406 14912
rect 488534 14900 488540 14912
rect 488592 14900 488598 14952
rect 511902 14900 511908 14952
rect 511960 14940 511966 14952
rect 537938 14940 537944 14952
rect 511960 14912 537944 14940
rect 511960 14900 511966 14912
rect 537938 14900 537944 14912
rect 537996 14900 538002 14952
rect 350166 14832 350172 14884
rect 350224 14872 350230 14884
rect 486234 14872 486240 14884
rect 350224 14844 486240 14872
rect 350224 14832 350230 14844
rect 486234 14832 486240 14844
rect 486292 14832 486298 14884
rect 491938 14832 491944 14884
rect 491996 14872 492002 14884
rect 520734 14872 520740 14884
rect 491996 14844 520740 14872
rect 491996 14832 492002 14844
rect 520734 14832 520740 14844
rect 520792 14832 520798 14884
rect 527818 14832 527824 14884
rect 527876 14872 527882 14884
rect 540238 14872 540244 14884
rect 527876 14844 540244 14872
rect 527876 14832 527882 14844
rect 540238 14832 540244 14844
rect 540296 14832 540302 14884
rect 329742 14764 329748 14816
rect 329800 14804 329806 14816
rect 479334 14804 479340 14816
rect 329800 14776 479340 14804
rect 329800 14764 329806 14776
rect 479334 14764 479340 14776
rect 479392 14764 479398 14816
rect 482922 14764 482928 14816
rect 482980 14804 482986 14816
rect 528738 14804 528744 14816
rect 482980 14776 528744 14804
rect 482980 14764 482986 14776
rect 528738 14764 528744 14776
rect 528796 14764 528802 14816
rect 531958 14764 531964 14816
rect 532016 14804 532022 14816
rect 543734 14804 543740 14816
rect 532016 14776 543740 14804
rect 532016 14764 532022 14776
rect 543734 14764 543740 14776
rect 543792 14764 543798 14816
rect 93762 14696 93768 14748
rect 93820 14736 93826 14748
rect 186498 14736 186504 14748
rect 93820 14708 186504 14736
rect 93820 14696 93826 14708
rect 186498 14696 186504 14708
rect 186556 14696 186562 14748
rect 314562 14696 314568 14748
rect 314620 14736 314626 14748
rect 474734 14736 474740 14748
rect 314620 14708 474740 14736
rect 314620 14696 314626 14708
rect 474734 14696 474740 14708
rect 474792 14696 474798 14748
rect 478782 14696 478788 14748
rect 478840 14736 478846 14748
rect 527634 14736 527640 14748
rect 478840 14708 527640 14736
rect 478840 14696 478846 14708
rect 527634 14696 527640 14708
rect 527692 14696 527698 14748
rect 531222 14696 531228 14748
rect 531280 14736 531286 14748
rect 544470 14736 544476 14748
rect 531280 14708 544476 14736
rect 531280 14696 531286 14708
rect 544470 14696 544476 14708
rect 544528 14696 544534 14748
rect 66162 14628 66168 14680
rect 66220 14668 66226 14680
rect 166994 14668 167000 14680
rect 66220 14640 167000 14668
rect 66220 14628 66226 14640
rect 166994 14628 167000 14640
rect 167052 14628 167058 14680
rect 250530 14628 250536 14680
rect 250588 14668 250594 14680
rect 419442 14668 419448 14680
rect 250588 14640 419448 14668
rect 250588 14628 250594 14640
rect 419442 14628 419448 14640
rect 419500 14628 419506 14680
rect 420638 14668 420644 14680
rect 419552 14640 420644 14668
rect 147582 14560 147588 14612
rect 147640 14600 147646 14612
rect 419552 14600 419580 14640
rect 420638 14628 420644 14640
rect 420696 14628 420702 14680
rect 426986 14628 426992 14680
rect 427044 14668 427050 14680
rect 435634 14668 435640 14680
rect 427044 14640 435640 14668
rect 427044 14628 427050 14640
rect 435634 14628 435640 14640
rect 435692 14628 435698 14680
rect 440418 14628 440424 14680
rect 440476 14668 440482 14680
rect 444466 14668 444472 14680
rect 440476 14640 444472 14668
rect 440476 14628 440482 14640
rect 444466 14628 444472 14640
rect 444524 14628 444530 14680
rect 464982 14628 464988 14680
rect 465040 14668 465046 14680
rect 523034 14668 523040 14680
rect 465040 14640 523040 14668
rect 465040 14628 465046 14640
rect 523034 14628 523040 14640
rect 523092 14628 523098 14680
rect 528462 14628 528468 14680
rect 528520 14668 528526 14680
rect 543366 14668 543372 14680
rect 528520 14640 543372 14668
rect 528520 14628 528526 14640
rect 543366 14628 543372 14640
rect 543424 14628 543430 14680
rect 555602 14628 555608 14680
rect 555660 14668 555666 14680
rect 561674 14668 561680 14680
rect 555660 14640 561680 14668
rect 555660 14628 555666 14640
rect 561674 14628 561680 14640
rect 561732 14628 561738 14680
rect 147640 14572 419580 14600
rect 147640 14560 147646 14572
rect 419626 14560 419632 14612
rect 419684 14600 419690 14612
rect 483198 14600 483204 14612
rect 419684 14572 483204 14600
rect 419684 14560 419690 14572
rect 483198 14560 483204 14572
rect 483256 14560 483262 14612
rect 503622 14560 503628 14612
rect 503680 14600 503686 14612
rect 535638 14600 535644 14612
rect 503680 14572 535644 14600
rect 503680 14560 503686 14572
rect 535638 14560 535644 14572
rect 535696 14560 535702 14612
rect 536742 14560 536748 14612
rect 536800 14600 536806 14612
rect 546034 14600 546040 14612
rect 536800 14572 546040 14600
rect 536800 14560 536806 14572
rect 546034 14560 546040 14572
rect 546092 14560 546098 14612
rect 554866 14560 554872 14612
rect 554924 14600 554930 14612
rect 563146 14600 563152 14612
rect 554924 14572 563152 14600
rect 554924 14560 554930 14572
rect 563146 14560 563152 14572
rect 563204 14560 563210 14612
rect 154482 14492 154488 14544
rect 154540 14532 154546 14544
rect 154540 14504 419672 14532
rect 154540 14492 154546 14504
rect 28902 14424 28908 14476
rect 28960 14464 28966 14476
rect 139394 14464 139400 14476
rect 28960 14436 139400 14464
rect 28960 14424 28966 14436
rect 139394 14424 139400 14436
rect 139452 14424 139458 14476
rect 143442 14424 143448 14476
rect 143500 14464 143506 14476
rect 419534 14464 419540 14476
rect 143500 14436 419540 14464
rect 143500 14424 143506 14436
rect 419534 14424 419540 14436
rect 419592 14424 419598 14476
rect 419644 14464 419672 14504
rect 420914 14492 420920 14544
rect 420972 14532 420978 14544
rect 420972 14504 426572 14532
rect 420972 14492 420978 14504
rect 422938 14464 422944 14476
rect 419644 14436 422944 14464
rect 422938 14424 422944 14436
rect 422996 14424 423002 14476
rect 423122 14424 423128 14476
rect 423180 14464 423186 14476
rect 426434 14464 426440 14476
rect 423180 14436 426440 14464
rect 423180 14424 423186 14436
rect 426434 14424 426440 14436
rect 426492 14424 426498 14476
rect 426544 14464 426572 14504
rect 428458 14492 428464 14544
rect 428516 14532 428522 14544
rect 431034 14532 431040 14544
rect 428516 14504 431040 14532
rect 428516 14492 428522 14504
rect 431034 14492 431040 14504
rect 431092 14492 431098 14544
rect 433242 14492 433248 14544
rect 433300 14532 433306 14544
rect 512638 14532 512644 14544
rect 433300 14504 512644 14532
rect 433300 14492 433306 14504
rect 512638 14492 512644 14504
rect 512696 14492 512702 14544
rect 525702 14492 525708 14544
rect 525760 14532 525766 14544
rect 542538 14532 542544 14544
rect 525760 14504 542544 14532
rect 525760 14492 525766 14504
rect 542538 14492 542544 14504
rect 542596 14492 542602 14544
rect 555234 14492 555240 14544
rect 555292 14532 555298 14544
rect 563054 14532 563060 14544
rect 555292 14504 563060 14532
rect 555292 14492 555298 14504
rect 563054 14492 563060 14504
rect 563112 14492 563118 14544
rect 506198 14464 506204 14476
rect 426544 14436 506204 14464
rect 506198 14424 506204 14436
rect 506256 14424 506262 14476
rect 507762 14424 507768 14476
rect 507820 14464 507826 14476
rect 536834 14464 536840 14476
rect 507820 14436 536840 14464
rect 507820 14424 507826 14436
rect 536834 14424 536840 14436
rect 536892 14424 536898 14476
rect 538122 14424 538128 14476
rect 538180 14464 538186 14476
rect 546770 14464 546776 14476
rect 538180 14436 546776 14464
rect 538180 14424 538186 14436
rect 546770 14424 546776 14436
rect 546828 14424 546834 14476
rect 557902 14424 557908 14476
rect 557960 14464 557966 14476
rect 570598 14464 570604 14476
rect 557960 14436 570604 14464
rect 557960 14424 557966 14436
rect 570598 14424 570604 14436
rect 570656 14424 570662 14476
rect 397362 14356 397368 14408
rect 397420 14396 397426 14408
rect 501138 14396 501144 14408
rect 397420 14368 501144 14396
rect 397420 14356 397426 14368
rect 501138 14356 501144 14368
rect 501196 14356 501202 14408
rect 523954 14356 523960 14408
rect 524012 14396 524018 14408
rect 524012 14368 528324 14396
rect 524012 14356 524018 14368
rect 408402 14288 408408 14340
rect 408460 14328 408466 14340
rect 504634 14328 504640 14340
rect 408460 14300 504640 14328
rect 408460 14288 408466 14300
rect 504634 14288 504640 14300
rect 504692 14288 504698 14340
rect 528296 14328 528324 14368
rect 528646 14356 528652 14408
rect 528704 14396 528710 14408
rect 529290 14396 529296 14408
rect 528704 14368 529296 14396
rect 528704 14356 528710 14368
rect 529290 14356 529296 14368
rect 529348 14356 529354 14408
rect 536098 14356 536104 14408
rect 536156 14396 536162 14408
rect 544838 14396 544844 14408
rect 536156 14368 544844 14396
rect 536156 14356 536162 14368
rect 544838 14356 544844 14368
rect 544896 14356 544902 14408
rect 532234 14328 532240 14340
rect 528296 14300 532240 14328
rect 532234 14288 532240 14300
rect 532292 14288 532298 14340
rect 553670 14288 553676 14340
rect 553728 14328 553734 14340
rect 556982 14328 556988 14340
rect 553728 14300 556988 14328
rect 553728 14288 553734 14300
rect 556982 14288 556988 14300
rect 557040 14288 557046 14340
rect 378042 14220 378048 14272
rect 378100 14260 378106 14272
rect 467834 14260 467840 14272
rect 378100 14232 467840 14260
rect 378100 14220 378106 14232
rect 467834 14220 467840 14232
rect 467892 14220 467898 14272
rect 471974 14220 471980 14272
rect 472032 14260 472038 14272
rect 525334 14260 525340 14272
rect 472032 14232 525340 14260
rect 472032 14220 472038 14232
rect 525334 14220 525340 14232
rect 525392 14220 525398 14272
rect 554038 14220 554044 14272
rect 554096 14260 554102 14272
rect 556614 14260 556620 14272
rect 554096 14232 556620 14260
rect 554096 14220 554102 14232
rect 556614 14220 556620 14232
rect 556672 14220 556678 14272
rect 384114 14152 384120 14204
rect 384172 14192 384178 14204
rect 418338 14192 418344 14204
rect 384172 14164 418344 14192
rect 384172 14152 384178 14164
rect 418338 14152 418344 14164
rect 418396 14152 418402 14204
rect 418522 14152 418528 14204
rect 418580 14192 418586 14204
rect 506934 14192 506940 14204
rect 418580 14164 506940 14192
rect 418580 14152 418586 14164
rect 506934 14152 506940 14164
rect 506992 14152 506998 14204
rect 543642 14152 543648 14204
rect 543700 14192 543706 14204
rect 548334 14192 548340 14204
rect 543700 14164 548340 14192
rect 543700 14152 543706 14164
rect 548334 14152 548340 14164
rect 548392 14152 548398 14204
rect 554498 14152 554504 14204
rect 554556 14192 554562 14204
rect 556890 14192 556896 14204
rect 554556 14164 556896 14192
rect 554556 14152 554562 14164
rect 556890 14152 556896 14164
rect 556948 14152 556954 14204
rect 419534 14084 419540 14136
rect 419592 14124 419598 14136
rect 482002 14124 482008 14136
rect 419592 14096 482008 14124
rect 419592 14084 419598 14096
rect 482002 14084 482008 14096
rect 482060 14084 482066 14136
rect 545022 14084 545028 14136
rect 545080 14124 545086 14136
rect 548702 14124 548708 14136
rect 545080 14096 548708 14124
rect 545080 14084 545086 14096
rect 548702 14084 548708 14096
rect 548760 14084 548766 14136
rect 552198 14084 552204 14136
rect 552256 14124 552262 14136
rect 555234 14124 555240 14136
rect 552256 14096 555240 14124
rect 552256 14084 552262 14096
rect 555234 14084 555240 14096
rect 555292 14084 555298 14136
rect 411254 14016 411260 14068
rect 411312 14056 411318 14068
rect 411312 14028 419396 14056
rect 411312 14016 411318 14028
rect 419368 13988 419396 14028
rect 419442 14016 419448 14068
rect 419500 14056 419506 14068
rect 425238 14056 425244 14068
rect 419500 14028 425244 14056
rect 419500 14016 419506 14028
rect 425238 14016 425244 14028
rect 425296 14016 425302 14068
rect 546310 14016 546316 14068
rect 546368 14056 546374 14068
rect 549070 14056 549076 14068
rect 546368 14028 549076 14056
rect 546368 14016 546374 14028
rect 549070 14016 549076 14028
rect 549128 14016 549134 14068
rect 552934 14016 552940 14068
rect 552992 14056 552998 14068
rect 555510 14056 555516 14068
rect 552992 14028 555516 14056
rect 552992 14016 552998 14028
rect 555510 14016 555516 14028
rect 555568 14016 555574 14068
rect 422202 13988 422208 14000
rect 419368 13960 422208 13988
rect 422202 13948 422208 13960
rect 422260 13948 422266 14000
rect 547690 13948 547696 14000
rect 547748 13988 547754 14000
rect 549898 13988 549904 14000
rect 547748 13960 549904 13988
rect 547748 13948 547754 13960
rect 549898 13948 549904 13960
rect 549956 13948 549962 14000
rect 553302 13948 553308 14000
rect 553360 13988 553366 14000
rect 555418 13988 555424 14000
rect 553360 13960 555424 13988
rect 553360 13948 553366 13960
rect 555418 13948 555424 13960
rect 555476 13948 555482 14000
rect 559834 13948 559840 14000
rect 559892 13988 559898 14000
rect 560202 13988 560208 14000
rect 559892 13960 560208 13988
rect 559892 13948 559898 13960
rect 560202 13948 560208 13960
rect 560260 13948 560266 14000
rect 425054 13880 425060 13932
rect 425112 13920 425118 13932
rect 428734 13920 428740 13932
rect 425112 13892 428740 13920
rect 425112 13880 425118 13892
rect 428734 13880 428740 13892
rect 428792 13880 428798 13932
rect 544378 13880 544384 13932
rect 544436 13920 544442 13932
rect 546402 13920 546408 13932
rect 544436 13892 546408 13920
rect 544436 13880 544442 13892
rect 546402 13880 546408 13892
rect 546460 13880 546466 13932
rect 547782 13880 547788 13932
rect 547840 13920 547846 13932
rect 549438 13920 549444 13932
rect 547840 13892 549444 13920
rect 547840 13880 547846 13892
rect 549438 13880 549444 13892
rect 549496 13880 549502 13932
rect 551370 13880 551376 13932
rect 551428 13920 551434 13932
rect 551830 13920 551836 13932
rect 551428 13892 551836 13920
rect 551428 13880 551434 13892
rect 551830 13880 551836 13892
rect 551888 13880 551894 13932
rect 552566 13880 552572 13932
rect 552624 13920 552630 13932
rect 554866 13920 554872 13932
rect 552624 13892 554872 13920
rect 552624 13880 552630 13892
rect 554866 13880 554872 13892
rect 554924 13880 554930 13932
rect 557534 13880 557540 13932
rect 557592 13920 557598 13932
rect 558730 13920 558736 13932
rect 557592 13892 558736 13920
rect 557592 13880 557598 13892
rect 558730 13880 558736 13892
rect 558788 13880 558794 13932
rect 559098 13880 559104 13932
rect 559156 13920 559162 13932
rect 560018 13920 560024 13932
rect 559156 13892 560024 13920
rect 559156 13880 559162 13892
rect 560018 13880 560024 13892
rect 560076 13880 560082 13932
rect 377876 13824 378272 13852
rect 375190 13744 375196 13796
rect 375248 13784 375254 13796
rect 377876 13784 377904 13824
rect 375248 13756 377904 13784
rect 378244 13784 378272 13824
rect 545758 13812 545764 13864
rect 545816 13852 545822 13864
rect 547138 13852 547144 13864
rect 545816 13824 547144 13852
rect 545816 13812 545822 13824
rect 547138 13812 547144 13824
rect 547196 13812 547202 13864
rect 549162 13812 549168 13864
rect 549220 13852 549226 13864
rect 550266 13852 550272 13864
rect 549220 13824 550272 13852
rect 549220 13812 549226 13824
rect 550266 13812 550272 13824
rect 550324 13812 550330 13864
rect 551738 13812 551744 13864
rect 551796 13852 551802 13864
rect 553394 13852 553400 13864
rect 551796 13824 553400 13852
rect 551796 13812 551802 13824
rect 553394 13812 553400 13824
rect 553452 13812 553458 13864
rect 556338 13812 556344 13864
rect 556396 13852 556402 13864
rect 557258 13852 557264 13864
rect 556396 13824 557264 13852
rect 556396 13812 556402 13824
rect 557258 13812 557264 13824
rect 557316 13812 557322 13864
rect 558270 13812 558276 13864
rect 558328 13852 558334 13864
rect 558822 13852 558828 13864
rect 558328 13824 558828 13852
rect 558328 13812 558334 13824
rect 558822 13812 558828 13824
rect 558880 13812 558886 13864
rect 559466 13812 559472 13864
rect 559524 13852 559530 13864
rect 560110 13852 560116 13864
rect 559524 13824 560116 13852
rect 559524 13812 559530 13824
rect 560110 13812 560116 13824
rect 560168 13812 560174 13864
rect 560570 13812 560576 13864
rect 560628 13852 560634 13864
rect 561582 13852 561588 13864
rect 560628 13824 561588 13852
rect 560628 13812 560634 13824
rect 561582 13812 561588 13824
rect 561640 13812 561646 13864
rect 493870 13784 493876 13796
rect 378244 13756 493876 13784
rect 375248 13744 375254 13756
rect 493870 13744 493876 13756
rect 493928 13744 493934 13796
rect 293862 13676 293868 13728
rect 293920 13716 293926 13728
rect 378042 13716 378048 13728
rect 293920 13688 378048 13716
rect 293920 13676 293926 13688
rect 378042 13676 378048 13688
rect 378100 13676 378106 13728
rect 378134 13676 378140 13728
rect 378192 13716 378198 13728
rect 495066 13716 495072 13728
rect 378192 13688 495072 13716
rect 378192 13676 378198 13688
rect 495066 13676 495072 13688
rect 495124 13676 495130 13728
rect 320082 13608 320088 13660
rect 320140 13648 320146 13660
rect 368658 13648 368664 13660
rect 320140 13620 368664 13648
rect 320140 13608 320146 13620
rect 368658 13608 368664 13620
rect 368716 13608 368722 13660
rect 371142 13608 371148 13660
rect 371200 13648 371206 13660
rect 492766 13648 492772 13660
rect 371200 13620 492772 13648
rect 371200 13608 371206 13620
rect 492766 13608 492772 13620
rect 492824 13608 492830 13660
rect 364242 13540 364248 13592
rect 364300 13580 364306 13592
rect 490466 13580 490472 13592
rect 364300 13552 490472 13580
rect 364300 13540 364306 13552
rect 490466 13540 490472 13552
rect 490524 13540 490530 13592
rect 360102 13472 360108 13524
rect 360160 13512 360166 13524
rect 489270 13512 489276 13524
rect 360160 13484 489276 13512
rect 360160 13472 360166 13484
rect 489270 13472 489276 13484
rect 489328 13472 489334 13524
rect 504358 13472 504364 13524
rect 504416 13512 504422 13524
rect 516134 13512 516140 13524
rect 504416 13484 516140 13512
rect 504416 13472 504422 13484
rect 516134 13472 516140 13484
rect 516192 13472 516198 13524
rect 269022 13404 269028 13456
rect 269080 13444 269086 13456
rect 459738 13444 459744 13456
rect 269080 13416 459744 13444
rect 269080 13404 269086 13416
rect 459738 13404 459744 13416
rect 459796 13404 459802 13456
rect 499114 13404 499120 13456
rect 499172 13444 499178 13456
rect 511534 13444 511540 13456
rect 499172 13416 511540 13444
rect 499172 13404 499178 13416
rect 511534 13404 511540 13416
rect 511592 13404 511598 13456
rect 226242 13336 226248 13388
rect 226300 13376 226306 13388
rect 445938 13376 445944 13388
rect 226300 13348 445944 13376
rect 226300 13336 226306 13348
rect 445938 13336 445944 13348
rect 445996 13336 446002 13388
rect 500218 13336 500224 13388
rect 500276 13376 500282 13388
rect 513834 13376 513840 13388
rect 500276 13348 513840 13376
rect 500276 13336 500282 13348
rect 513834 13336 513840 13348
rect 513892 13336 513898 13388
rect 190362 13268 190368 13320
rect 190420 13308 190426 13320
rect 434438 13308 434444 13320
rect 190420 13280 434444 13308
rect 190420 13268 190426 13280
rect 434438 13268 434444 13280
rect 434496 13268 434502 13320
rect 456978 13268 456984 13320
rect 457036 13308 457042 13320
rect 457438 13308 457444 13320
rect 457036 13280 457444 13308
rect 457036 13268 457042 13280
rect 457438 13268 457444 13280
rect 457496 13268 457502 13320
rect 496722 13268 496728 13320
rect 496780 13308 496786 13320
rect 533338 13308 533344 13320
rect 496780 13280 533344 13308
rect 496780 13268 496786 13280
rect 533338 13268 533344 13280
rect 533396 13268 533402 13320
rect 140682 13200 140688 13252
rect 140740 13240 140746 13252
rect 384114 13240 384120 13252
rect 140740 13212 384120 13240
rect 140740 13200 140746 13212
rect 384114 13200 384120 13212
rect 384172 13200 384178 13252
rect 384482 13200 384488 13252
rect 384540 13240 384546 13252
rect 497366 13240 497372 13252
rect 384540 13212 497372 13240
rect 384540 13200 384546 13212
rect 497366 13200 497372 13212
rect 497424 13200 497430 13252
rect 498102 13200 498108 13252
rect 498160 13240 498166 13252
rect 533798 13240 533804 13252
rect 498160 13212 533804 13240
rect 498160 13200 498166 13212
rect 533798 13200 533804 13212
rect 533856 13200 533862 13252
rect 42702 13132 42708 13184
rect 42760 13172 42766 13184
rect 149330 13172 149336 13184
rect 42760 13144 149336 13172
rect 42760 13132 42766 13144
rect 149330 13132 149336 13144
rect 149388 13132 149394 13184
rect 153102 13132 153108 13184
rect 153160 13172 153166 13184
rect 409138 13172 409144 13184
rect 153160 13144 409144 13172
rect 153160 13132 153166 13144
rect 409138 13132 409144 13144
rect 409196 13132 409202 13184
rect 436738 13132 436744 13184
rect 436796 13172 436802 13184
rect 466638 13172 466644 13184
rect 436796 13144 466644 13172
rect 436796 13132 436802 13144
rect 466638 13132 466644 13144
rect 466696 13132 466702 13184
rect 495342 13132 495348 13184
rect 495400 13172 495406 13184
rect 532602 13172 532608 13184
rect 495400 13144 532608 13172
rect 495400 13132 495406 13144
rect 532602 13132 532608 13144
rect 532660 13132 532666 13184
rect 533982 13132 533988 13184
rect 534040 13172 534046 13184
rect 545298 13172 545304 13184
rect 534040 13144 545304 13172
rect 534040 13132 534046 13144
rect 545298 13132 545304 13144
rect 545356 13132 545362 13184
rect 22002 13064 22008 13116
rect 22060 13104 22066 13116
rect 135346 13104 135352 13116
rect 22060 13076 135352 13104
rect 22060 13064 22066 13076
rect 135346 13064 135352 13076
rect 135404 13064 135410 13116
rect 150342 13064 150348 13116
rect 150400 13104 150406 13116
rect 421466 13104 421472 13116
rect 150400 13076 421472 13104
rect 150400 13064 150406 13076
rect 421466 13064 421472 13076
rect 421524 13064 421530 13116
rect 424962 13064 424968 13116
rect 425020 13104 425026 13116
rect 509970 13104 509976 13116
rect 425020 13076 509976 13104
rect 425020 13064 425026 13076
rect 509970 13064 509976 13076
rect 510028 13064 510034 13116
rect 517422 13064 517428 13116
rect 517480 13104 517486 13116
rect 539870 13104 539876 13116
rect 517480 13076 539876 13104
rect 517480 13064 517486 13076
rect 539870 13064 539876 13076
rect 539928 13064 539934 13116
rect 382182 12996 382188 13048
rect 382240 13036 382246 13048
rect 496170 13036 496176 13048
rect 382240 13008 496176 13036
rect 382240 12996 382246 13008
rect 496170 12996 496176 13008
rect 496228 12996 496234 13048
rect 389082 12928 389088 12980
rect 389140 12968 389146 12980
rect 498470 12968 498476 12980
rect 389140 12940 498476 12968
rect 389140 12928 389146 12940
rect 498470 12928 498476 12940
rect 498528 12928 498534 12980
rect 391842 12860 391848 12912
rect 391900 12900 391906 12912
rect 391900 12872 490696 12900
rect 391900 12860 391906 12872
rect 407022 12792 407028 12844
rect 407080 12832 407086 12844
rect 490558 12832 490564 12844
rect 407080 12804 490564 12832
rect 407080 12792 407086 12804
rect 490558 12792 490564 12804
rect 490616 12792 490622 12844
rect 415302 12724 415308 12776
rect 415360 12764 415366 12776
rect 422570 12764 422576 12776
rect 415360 12736 422576 12764
rect 415360 12724 415366 12736
rect 422570 12724 422576 12736
rect 422628 12724 422634 12776
rect 422754 12724 422760 12776
rect 422812 12764 422818 12776
rect 447042 12764 447048 12776
rect 422812 12736 447048 12764
rect 422812 12724 422818 12736
rect 447042 12724 447048 12736
rect 447100 12724 447106 12776
rect 476022 12724 476028 12776
rect 476080 12764 476086 12776
rect 490668 12764 490696 12872
rect 490742 12792 490748 12844
rect 490800 12832 490806 12844
rect 504266 12832 504272 12844
rect 490800 12804 504272 12832
rect 490800 12792 490806 12804
rect 504266 12792 504272 12804
rect 504324 12792 504330 12844
rect 561674 12792 561680 12844
rect 561732 12832 561738 12844
rect 564434 12832 564440 12844
rect 561732 12804 564440 12832
rect 561732 12792 561738 12804
rect 564434 12792 564440 12804
rect 564492 12792 564498 12844
rect 499666 12764 499672 12776
rect 476080 12736 490604 12764
rect 490668 12736 499672 12764
rect 476080 12724 476086 12736
rect 395982 12656 395988 12708
rect 396040 12696 396046 12708
rect 396040 12668 418384 12696
rect 396040 12656 396046 12668
rect 409138 12588 409144 12640
rect 409196 12628 409202 12640
rect 415302 12628 415308 12640
rect 409196 12600 415308 12628
rect 409196 12588 409202 12600
rect 415302 12588 415308 12600
rect 415360 12588 415366 12640
rect 418356 12560 418384 12668
rect 421558 12656 421564 12708
rect 421616 12696 421622 12708
rect 427078 12696 427084 12708
rect 421616 12668 427084 12696
rect 421616 12656 421622 12668
rect 427078 12656 427084 12668
rect 427136 12656 427142 12708
rect 427998 12656 428004 12708
rect 428056 12696 428062 12708
rect 444374 12696 444380 12708
rect 428056 12668 444380 12696
rect 428056 12656 428062 12668
rect 444374 12656 444380 12668
rect 444432 12656 444438 12708
rect 489638 12696 489644 12708
rect 447612 12668 489644 12696
rect 422294 12560 422300 12572
rect 418356 12532 422300 12560
rect 422294 12520 422300 12532
rect 422352 12520 422358 12572
rect 444374 12520 444380 12572
rect 444432 12560 444438 12572
rect 447612 12560 447640 12668
rect 489638 12656 489644 12668
rect 489696 12656 489702 12708
rect 490576 12696 490604 12736
rect 499666 12724 499672 12736
rect 499724 12724 499730 12776
rect 500770 12696 500776 12708
rect 490576 12668 500776 12696
rect 500770 12656 500776 12668
rect 500828 12656 500834 12708
rect 466178 12628 466184 12640
rect 444432 12532 447640 12560
rect 453960 12600 466184 12628
rect 444432 12520 444438 12532
rect 427078 12452 427084 12504
rect 427136 12492 427142 12504
rect 427998 12492 428004 12504
rect 427136 12464 428004 12492
rect 427136 12452 427142 12464
rect 427998 12452 428004 12464
rect 428056 12452 428062 12504
rect 447042 12452 447048 12504
rect 447100 12492 447106 12504
rect 453960 12492 453988 12600
rect 466178 12588 466184 12600
rect 466236 12588 466242 12640
rect 471882 12588 471888 12640
rect 471940 12628 471946 12640
rect 476022 12628 476028 12640
rect 471940 12600 476028 12628
rect 471940 12588 471946 12600
rect 476022 12588 476028 12600
rect 476080 12588 476086 12640
rect 447100 12464 453988 12492
rect 447100 12452 447106 12464
rect 320450 12384 320456 12436
rect 320508 12424 320514 12436
rect 476666 12424 476672 12436
rect 320508 12396 476672 12424
rect 320508 12384 320514 12396
rect 476666 12384 476672 12396
rect 476724 12384 476730 12436
rect 313366 12316 313372 12368
rect 313424 12356 313430 12368
rect 313424 12328 316816 12356
rect 313424 12316 313430 12328
rect 316678 12288 316684 12300
rect 302252 12260 316684 12288
rect 299106 12112 299112 12164
rect 299164 12152 299170 12164
rect 302252 12152 302280 12260
rect 316678 12248 316684 12260
rect 316736 12248 316742 12300
rect 316788 12288 316816 12328
rect 316954 12316 316960 12368
rect 317012 12356 317018 12368
rect 475470 12356 475476 12368
rect 317012 12328 475476 12356
rect 317012 12316 317018 12328
rect 475470 12316 475476 12328
rect 475528 12316 475534 12368
rect 474366 12288 474372 12300
rect 316788 12260 474372 12288
rect 474366 12248 474372 12260
rect 474424 12248 474430 12300
rect 484486 12248 484492 12300
rect 484544 12288 484550 12300
rect 485038 12288 485044 12300
rect 484544 12260 485044 12288
rect 484544 12248 484550 12260
rect 485038 12248 485044 12260
rect 485096 12248 485102 12300
rect 306190 12180 306196 12232
rect 306248 12220 306254 12232
rect 472066 12220 472072 12232
rect 306248 12192 472072 12220
rect 306248 12180 306254 12192
rect 472066 12180 472072 12192
rect 472124 12180 472130 12232
rect 473446 12180 473452 12232
rect 473504 12220 473510 12232
rect 473998 12220 474004 12232
rect 473504 12192 474004 12220
rect 473504 12180 473510 12192
rect 473998 12180 474004 12192
rect 474056 12180 474062 12232
rect 501230 12180 501236 12232
rect 501288 12220 501294 12232
rect 534902 12220 534908 12232
rect 501288 12192 534908 12220
rect 501288 12180 501294 12192
rect 534902 12180 534908 12192
rect 534960 12180 534966 12232
rect 299164 12124 302280 12152
rect 299164 12112 299170 12124
rect 302602 12112 302608 12164
rect 302660 12152 302666 12164
rect 470870 12152 470876 12164
rect 302660 12124 470876 12152
rect 302660 12112 302666 12124
rect 470870 12112 470876 12124
rect 470928 12112 470934 12164
rect 484302 12112 484308 12164
rect 484360 12152 484366 12164
rect 529198 12152 529204 12164
rect 484360 12124 529204 12152
rect 484360 12112 484366 12124
rect 529198 12112 529204 12124
rect 529256 12112 529262 12164
rect 325602 12044 325608 12096
rect 325660 12084 325666 12096
rect 335354 12084 335360 12096
rect 325660 12056 335360 12084
rect 325660 12044 325666 12056
rect 335354 12044 335360 12056
rect 335412 12044 335418 12096
rect 342990 12044 342996 12096
rect 343048 12084 343054 12096
rect 355318 12084 355324 12096
rect 343048 12056 355324 12084
rect 343048 12044 343054 12056
rect 355318 12044 355324 12056
rect 355376 12044 355382 12096
rect 364150 12044 364156 12096
rect 364208 12084 364214 12096
rect 374638 12084 374644 12096
rect 364208 12056 374644 12084
rect 364208 12044 364214 12056
rect 374638 12044 374644 12056
rect 374696 12044 374702 12096
rect 384298 12044 384304 12096
rect 384356 12084 384362 12096
rect 393958 12084 393964 12096
rect 384356 12056 393964 12084
rect 384356 12044 384362 12056
rect 393958 12044 393964 12056
rect 394016 12044 394022 12096
rect 403618 12044 403624 12096
rect 403676 12084 403682 12096
rect 413278 12084 413284 12096
rect 403676 12056 413284 12084
rect 403676 12044 403682 12056
rect 413278 12044 413284 12056
rect 413336 12044 413342 12096
rect 422202 12044 422208 12096
rect 422260 12084 422266 12096
rect 431954 12084 431960 12096
rect 422260 12056 431960 12084
rect 422260 12044 422266 12056
rect 431954 12044 431960 12056
rect 432012 12044 432018 12096
rect 442258 12044 442264 12096
rect 442316 12084 442322 12096
rect 461486 12084 461492 12096
rect 442316 12056 461492 12084
rect 442316 12044 442322 12056
rect 461486 12044 461492 12056
rect 461544 12044 461550 12096
rect 468570 12084 468576 12096
rect 461596 12056 468576 12084
rect 295518 11976 295524 12028
rect 295576 12016 295582 12028
rect 461596 12016 461624 12056
rect 468570 12044 468576 12056
rect 468628 12044 468634 12096
rect 478690 12044 478696 12096
rect 478748 12084 478754 12096
rect 527266 12084 527272 12096
rect 478748 12056 527272 12084
rect 478748 12044 478754 12056
rect 527266 12044 527272 12056
rect 527324 12044 527330 12096
rect 467466 12016 467472 12028
rect 295576 11988 461624 12016
rect 461688 11988 467472 12016
rect 295576 11976 295582 11988
rect 291930 11908 291936 11960
rect 291988 11948 291994 11960
rect 461688 11948 461716 11988
rect 467466 11976 467472 11988
rect 467524 11976 467530 12028
rect 473906 11976 473912 12028
rect 473964 12016 473970 12028
rect 526070 12016 526076 12028
rect 473964 11988 526076 12016
rect 473964 11976 473970 11988
rect 526070 11976 526076 11988
rect 526128 11976 526134 12028
rect 291988 11920 461716 11948
rect 291988 11908 291994 11920
rect 472710 11908 472716 11960
rect 472768 11948 472774 11960
rect 525426 11948 525432 11960
rect 472768 11920 525432 11948
rect 472768 11908 472774 11920
rect 525426 11908 525432 11920
rect 525484 11908 525490 11960
rect 46842 11840 46848 11892
rect 46900 11880 46906 11892
rect 148042 11880 148048 11892
rect 46900 11852 148048 11880
rect 46900 11840 46906 11852
rect 148042 11840 148048 11852
rect 148100 11840 148106 11892
rect 288342 11840 288348 11892
rect 288400 11880 288406 11892
rect 466270 11880 466276 11892
rect 288400 11852 466276 11880
rect 288400 11840 288406 11852
rect 466270 11840 466276 11852
rect 466328 11840 466334 11892
rect 470502 11840 470508 11892
rect 470560 11880 470566 11892
rect 524966 11880 524972 11892
rect 470560 11852 524972 11880
rect 470560 11840 470566 11852
rect 524966 11840 524972 11852
rect 525024 11840 525030 11892
rect 27522 11772 27528 11824
rect 27580 11812 27586 11824
rect 138106 11812 138112 11824
rect 27580 11784 138112 11812
rect 27580 11772 27586 11784
rect 138106 11772 138112 11784
rect 138164 11772 138170 11824
rect 284754 11772 284760 11824
rect 284812 11812 284818 11824
rect 465166 11812 465172 11824
rect 284812 11784 465172 11812
rect 284812 11772 284818 11784
rect 465166 11772 465172 11784
rect 465224 11772 465230 11824
rect 466822 11772 466828 11824
rect 466880 11812 466886 11824
rect 523770 11812 523776 11824
rect 466880 11784 523776 11812
rect 466880 11772 466886 11784
rect 523770 11772 523776 11784
rect 523828 11772 523834 11824
rect 529842 11772 529848 11824
rect 529900 11812 529906 11824
rect 544102 11812 544108 11824
rect 529900 11784 544108 11812
rect 529900 11772 529906 11784
rect 544102 11772 544108 11784
rect 544160 11772 544166 11824
rect 133782 11704 133788 11756
rect 133840 11744 133846 11756
rect 416038 11744 416044 11756
rect 133840 11716 416044 11744
rect 133840 11704 133846 11716
rect 416038 11704 416044 11716
rect 416096 11704 416102 11756
rect 416682 11704 416688 11756
rect 416740 11744 416746 11756
rect 507302 11744 507308 11756
rect 416740 11716 507308 11744
rect 416740 11704 416746 11716
rect 507302 11704 507308 11716
rect 507360 11704 507366 11756
rect 526438 11704 526444 11756
rect 526496 11744 526502 11756
rect 542170 11744 542176 11756
rect 526496 11716 542176 11744
rect 526496 11704 526502 11716
rect 542170 11704 542176 11716
rect 542228 11704 542234 11756
rect 556798 11704 556804 11756
rect 556856 11744 556862 11756
rect 568574 11744 568580 11756
rect 556856 11716 568580 11744
rect 556856 11704 556862 11716
rect 568574 11704 568580 11716
rect 568632 11704 568638 11756
rect 324222 11636 324228 11688
rect 324280 11676 324286 11688
rect 477494 11676 477500 11688
rect 324280 11648 477500 11676
rect 324280 11636 324286 11648
rect 477494 11636 477500 11648
rect 477552 11636 477558 11688
rect 483106 11636 483112 11688
rect 483164 11676 483170 11688
rect 483658 11676 483664 11688
rect 483164 11648 483664 11676
rect 483164 11636 483170 11648
rect 483658 11636 483664 11648
rect 483716 11636 483722 11688
rect 512086 11636 512092 11688
rect 512144 11676 512150 11688
rect 512914 11676 512920 11688
rect 512144 11648 512920 11676
rect 512144 11636 512150 11648
rect 512914 11636 512920 11648
rect 512972 11636 512978 11688
rect 316678 11568 316684 11620
rect 316736 11608 316742 11620
rect 325602 11608 325608 11620
rect 316736 11580 325608 11608
rect 316736 11568 316742 11580
rect 325602 11568 325608 11580
rect 325660 11568 325666 11620
rect 335354 11568 335360 11620
rect 335412 11608 335418 11620
rect 342990 11608 342996 11620
rect 335412 11580 342996 11608
rect 335412 11568 335418 11580
rect 342990 11568 342996 11580
rect 343048 11568 343054 11620
rect 349062 11568 349068 11620
rect 349120 11608 349126 11620
rect 485866 11608 485872 11620
rect 349120 11580 485872 11608
rect 349120 11568 349126 11580
rect 485866 11568 485872 11580
rect 485924 11568 485930 11620
rect 335998 11500 336004 11552
rect 336056 11540 336062 11552
rect 473170 11540 473176 11552
rect 336056 11512 473176 11540
rect 336056 11500 336062 11512
rect 473170 11500 473176 11512
rect 473228 11500 473234 11552
rect 355318 11432 355324 11484
rect 355376 11472 355382 11484
rect 364150 11472 364156 11484
rect 355376 11444 364156 11472
rect 355376 11432 355382 11444
rect 364150 11432 364156 11444
rect 364208 11432 364214 11484
rect 374638 11432 374644 11484
rect 374696 11472 374702 11484
rect 384298 11472 384304 11484
rect 374696 11444 384304 11472
rect 374696 11432 374702 11444
rect 384298 11432 384304 11444
rect 384356 11432 384362 11484
rect 400214 11432 400220 11484
rect 400272 11472 400278 11484
rect 502334 11472 502340 11484
rect 400272 11444 502340 11472
rect 400272 11432 400278 11444
rect 502334 11432 502340 11444
rect 502392 11432 502398 11484
rect 393958 11364 393964 11416
rect 394016 11404 394022 11416
rect 403618 11404 403624 11416
rect 394016 11376 403624 11404
rect 394016 11364 394022 11376
rect 403618 11364 403624 11376
rect 403676 11364 403682 11416
rect 409690 11364 409696 11416
rect 409748 11404 409754 11416
rect 505370 11404 505376 11416
rect 409748 11376 505376 11404
rect 409748 11364 409754 11376
rect 505370 11364 505376 11376
rect 505428 11364 505434 11416
rect 413278 11296 413284 11348
rect 413336 11336 413342 11348
rect 422202 11336 422208 11348
rect 413336 11308 422208 11336
rect 413336 11296 413342 11308
rect 422202 11296 422208 11308
rect 422260 11296 422266 11348
rect 425054 11296 425060 11348
rect 425112 11336 425118 11348
rect 425514 11336 425520 11348
rect 425112 11308 425520 11336
rect 425112 11296 425118 11308
rect 425514 11296 425520 11308
rect 425572 11296 425578 11348
rect 434806 11296 434812 11348
rect 434864 11336 434870 11348
rect 435726 11336 435732 11348
rect 434864 11308 435732 11336
rect 434864 11296 434870 11308
rect 435726 11296 435732 11308
rect 435784 11296 435790 11348
rect 468294 11296 468300 11348
rect 468352 11336 468358 11348
rect 518434 11336 518440 11348
rect 468352 11308 518440 11336
rect 468352 11296 468358 11308
rect 518434 11296 518440 11308
rect 518492 11296 518498 11348
rect 431954 11228 431960 11280
rect 432012 11268 432018 11280
rect 442258 11268 442264 11280
rect 432012 11240 442264 11268
rect 432012 11228 432018 11240
rect 442258 11228 442264 11240
rect 442316 11228 442322 11280
rect 461486 11228 461492 11280
rect 461544 11268 461550 11280
rect 469766 11268 469772 11280
rect 461544 11240 469772 11268
rect 461544 11228 461550 11240
rect 469766 11228 469772 11240
rect 469824 11228 469830 11280
rect 441706 11024 441712 11076
rect 441764 11064 441770 11076
rect 441982 11064 441988 11076
rect 441764 11036 441988 11064
rect 441764 11024 441770 11036
rect 441982 11024 441988 11036
rect 442040 11024 442046 11076
rect 281258 10956 281264 11008
rect 281316 10996 281322 11008
rect 463970 10996 463976 11008
rect 281316 10968 463976 10996
rect 281316 10956 281322 10968
rect 463970 10956 463976 10968
rect 464028 10956 464034 11008
rect 489914 10956 489920 11008
rect 489972 10996 489978 11008
rect 509142 10996 509148 11008
rect 489972 10968 509148 10996
rect 489972 10956 489978 10968
rect 509142 10956 509148 10968
rect 509200 10956 509206 11008
rect 263502 10888 263508 10940
rect 263560 10928 263566 10940
rect 458266 10928 458272 10940
rect 263560 10900 458272 10928
rect 263560 10888 263566 10900
rect 458266 10888 458272 10900
rect 458324 10888 458330 10940
rect 506382 10888 506388 10940
rect 506440 10928 506446 10940
rect 536466 10928 536472 10940
rect 506440 10900 536472 10928
rect 506440 10888 506446 10900
rect 536466 10888 536472 10900
rect 536524 10888 536530 10940
rect 253842 10820 253848 10872
rect 253900 10860 253906 10872
rect 454770 10860 454776 10872
rect 253900 10832 454776 10860
rect 253900 10820 253906 10832
rect 454770 10820 454776 10832
rect 454828 10820 454834 10872
rect 474734 10820 474740 10872
rect 474792 10860 474798 10872
rect 509234 10860 509240 10872
rect 474792 10832 509240 10860
rect 474792 10820 474798 10832
rect 509234 10820 509240 10832
rect 509292 10820 509298 10872
rect 530302 10860 530308 10872
rect 509344 10832 530308 10860
rect 249702 10752 249708 10804
rect 249760 10792 249766 10804
rect 453666 10792 453672 10804
rect 249760 10764 453672 10792
rect 249760 10752 249766 10764
rect 453666 10752 453672 10764
rect 453724 10752 453730 10804
rect 487062 10752 487068 10804
rect 487120 10792 487126 10804
rect 489914 10792 489920 10804
rect 487120 10764 489920 10792
rect 487120 10752 487126 10764
rect 489914 10752 489920 10764
rect 489972 10752 489978 10804
rect 509142 10752 509148 10804
rect 509200 10792 509206 10804
rect 509344 10792 509372 10832
rect 530302 10820 530308 10832
rect 530360 10820 530366 10872
rect 509200 10764 509372 10792
rect 509200 10752 509206 10764
rect 245562 10684 245568 10736
rect 245620 10724 245626 10736
rect 452470 10724 452476 10736
rect 245620 10696 452476 10724
rect 245620 10684 245626 10696
rect 452470 10684 452476 10696
rect 452528 10684 452534 10736
rect 452654 10684 452660 10736
rect 452712 10724 452718 10736
rect 480438 10724 480444 10736
rect 452712 10696 480444 10724
rect 452712 10684 452718 10696
rect 480438 10684 480444 10696
rect 480496 10684 480502 10736
rect 481542 10684 481548 10736
rect 481600 10724 481606 10736
rect 528370 10724 528376 10736
rect 481600 10696 528376 10724
rect 481600 10684 481606 10696
rect 528370 10684 528376 10696
rect 528428 10684 528434 10736
rect 240042 10616 240048 10668
rect 240100 10656 240106 10668
rect 450538 10656 450544 10668
rect 240100 10628 450544 10656
rect 240100 10616 240106 10628
rect 450538 10616 450544 10628
rect 450596 10616 450602 10668
rect 456058 10616 456064 10668
rect 456116 10656 456122 10668
rect 520274 10656 520280 10668
rect 456116 10628 520280 10656
rect 456116 10616 456122 10628
rect 520274 10616 520280 10628
rect 520332 10616 520338 10668
rect 235902 10548 235908 10600
rect 235960 10588 235966 10600
rect 448790 10588 448796 10600
rect 235960 10560 448796 10588
rect 235960 10548 235966 10560
rect 448790 10548 448796 10560
rect 448848 10548 448854 10600
rect 452470 10548 452476 10600
rect 452528 10588 452534 10600
rect 518894 10588 518900 10600
rect 452528 10560 518900 10588
rect 452528 10548 452534 10560
rect 518894 10548 518900 10560
rect 518952 10548 518958 10600
rect 231762 10480 231768 10532
rect 231820 10520 231826 10532
rect 447594 10520 447600 10532
rect 231820 10492 447600 10520
rect 231820 10480 231826 10492
rect 447594 10480 447600 10492
rect 447652 10480 447658 10532
rect 448146 10480 448152 10532
rect 448204 10520 448210 10532
rect 514938 10520 514944 10532
rect 448204 10492 514944 10520
rect 448204 10480 448210 10492
rect 514938 10480 514944 10492
rect 514996 10480 515002 10532
rect 86126 10412 86132 10464
rect 86184 10452 86190 10464
rect 182266 10452 182272 10464
rect 86184 10424 182272 10452
rect 86184 10412 86190 10424
rect 182266 10412 182272 10424
rect 182324 10412 182330 10464
rect 229002 10412 229008 10464
rect 229060 10452 229066 10464
rect 446766 10452 446772 10464
rect 229060 10424 446772 10452
rect 229060 10412 229066 10424
rect 446766 10412 446772 10424
rect 446824 10412 446830 10464
rect 448974 10412 448980 10464
rect 449032 10452 449038 10464
rect 518066 10452 518072 10464
rect 449032 10424 518072 10452
rect 449032 10412 449038 10424
rect 518066 10412 518072 10424
rect 518124 10412 518130 10464
rect 31662 10344 31668 10396
rect 31720 10384 31726 10396
rect 142246 10384 142252 10396
rect 31720 10356 142252 10384
rect 31720 10344 31726 10356
rect 142246 10344 142252 10356
rect 142304 10344 142310 10396
rect 220722 10344 220728 10396
rect 220780 10384 220786 10396
rect 440418 10384 440424 10396
rect 220780 10356 440424 10384
rect 220780 10344 220786 10356
rect 440418 10344 440424 10356
rect 440476 10344 440482 10396
rect 440602 10344 440608 10396
rect 440660 10384 440666 10396
rect 515398 10384 515404 10396
rect 440660 10356 515404 10384
rect 440660 10344 440666 10356
rect 515398 10344 515404 10356
rect 515456 10344 515462 10396
rect 9030 10276 9036 10328
rect 9088 10316 9094 10328
rect 120074 10316 120080 10328
rect 9088 10288 120080 10316
rect 9088 10276 9094 10288
rect 120074 10276 120080 10288
rect 120132 10276 120138 10328
rect 135162 10276 135168 10328
rect 135220 10316 135226 10328
rect 416866 10316 416872 10328
rect 135220 10288 416872 10316
rect 135220 10276 135226 10288
rect 416866 10276 416872 10288
rect 416924 10276 416930 10328
rect 417050 10276 417056 10328
rect 417108 10316 417114 10328
rect 507670 10316 507676 10328
rect 417108 10288 507676 10316
rect 417108 10276 417114 10288
rect 507670 10276 507676 10288
rect 507728 10276 507734 10328
rect 522666 10276 522672 10328
rect 522724 10316 522730 10328
rect 541802 10316 541808 10328
rect 522724 10288 541808 10316
rect 522724 10276 522730 10288
rect 541802 10276 541808 10288
rect 541860 10276 541866 10328
rect 322842 10208 322848 10260
rect 322900 10248 322906 10260
rect 477034 10248 477040 10260
rect 322900 10220 477040 10248
rect 322900 10208 322906 10220
rect 477034 10208 477040 10220
rect 477092 10208 477098 10260
rect 352558 10140 352564 10192
rect 352616 10180 352622 10192
rect 486970 10180 486976 10192
rect 352616 10152 486976 10180
rect 352616 10140 352622 10152
rect 486970 10140 486976 10152
rect 487028 10140 487034 10192
rect 364978 10072 364984 10124
rect 365036 10112 365042 10124
rect 456334 10112 456340 10124
rect 365036 10084 456340 10112
rect 365036 10072 365042 10084
rect 456334 10072 456340 10084
rect 456392 10072 456398 10124
rect 418798 10004 418804 10056
rect 418856 10044 418862 10056
rect 503070 10044 503076 10056
rect 418856 10016 503076 10044
rect 418856 10004 418862 10016
rect 503070 10004 503076 10016
rect 503128 10004 503134 10056
rect 338022 9936 338028 9988
rect 338080 9976 338086 9988
rect 419534 9976 419540 9988
rect 338080 9948 419540 9976
rect 338080 9936 338086 9948
rect 419534 9936 419540 9948
rect 419592 9936 419598 9988
rect 442350 9936 442356 9988
rect 442408 9976 442414 9988
rect 515766 9976 515772 9988
rect 442408 9948 515772 9976
rect 442408 9936 442414 9948
rect 515766 9936 515772 9948
rect 515824 9936 515830 9988
rect 445754 9868 445760 9920
rect 445812 9908 445818 9920
rect 473538 9908 473544 9920
rect 445812 9880 473544 9908
rect 445812 9868 445818 9880
rect 473538 9868 473544 9880
rect 473596 9868 473602 9920
rect 450078 9800 450084 9852
rect 450136 9840 450142 9852
rect 475838 9840 475844 9852
rect 450136 9812 475844 9840
rect 450136 9800 450142 9812
rect 475838 9800 475844 9812
rect 475896 9800 475902 9852
rect 208486 9664 208492 9716
rect 208544 9704 208550 9716
rect 208762 9704 208768 9716
rect 208544 9676 208768 9704
rect 208544 9664 208550 9676
rect 208762 9664 208768 9676
rect 208820 9664 208826 9716
rect 376202 9664 376208 9716
rect 376260 9704 376266 9716
rect 376386 9704 376392 9716
rect 376260 9676 376392 9704
rect 376260 9664 376266 9676
rect 376386 9664 376392 9676
rect 376444 9664 376450 9716
rect 451826 9664 451832 9716
rect 451884 9704 451890 9716
rect 452102 9704 452108 9716
rect 451884 9676 452108 9704
rect 451884 9664 451890 9676
rect 452102 9664 452108 9676
rect 452160 9664 452166 9716
rect 458634 9664 458640 9716
rect 458692 9704 458698 9716
rect 459002 9704 459008 9716
rect 458692 9676 459008 9704
rect 458692 9664 458698 9676
rect 459002 9664 459008 9676
rect 459060 9664 459066 9716
rect 459922 9664 459928 9716
rect 459980 9704 459986 9716
rect 460566 9704 460572 9716
rect 459980 9676 460572 9704
rect 459980 9664 459986 9676
rect 460566 9664 460572 9676
rect 460624 9664 460630 9716
rect 470594 9664 470600 9716
rect 470652 9704 470658 9716
rect 471238 9704 471244 9716
rect 470652 9676 471244 9704
rect 470652 9664 470658 9676
rect 471238 9664 471244 9676
rect 471296 9664 471302 9716
rect 471514 9664 471520 9716
rect 471572 9704 471578 9716
rect 471974 9704 471980 9716
rect 471572 9676 471980 9704
rect 471572 9664 471578 9676
rect 471974 9664 471980 9676
rect 472032 9664 472038 9716
rect 472158 9664 472164 9716
rect 472216 9704 472222 9716
rect 472802 9704 472808 9716
rect 472216 9676 472808 9704
rect 472216 9664 472222 9676
rect 472802 9664 472808 9676
rect 472860 9664 472866 9716
rect 497090 9664 497096 9716
rect 497148 9704 497154 9716
rect 497734 9704 497740 9716
rect 497148 9676 497740 9704
rect 497148 9664 497154 9676
rect 497734 9664 497740 9676
rect 497792 9664 497798 9716
rect 530118 9664 530124 9716
rect 530176 9704 530182 9716
rect 530670 9704 530676 9716
rect 530176 9676 530676 9704
rect 530176 9664 530182 9676
rect 530670 9664 530676 9676
rect 530728 9664 530734 9716
rect 202782 9596 202788 9648
rect 202840 9596 202846 9648
rect 253750 9596 253756 9648
rect 253808 9636 253814 9648
rect 455138 9636 455144 9648
rect 253808 9608 455144 9636
rect 253808 9596 253814 9608
rect 455138 9596 455144 9608
rect 455196 9596 455202 9648
rect 509234 9596 509240 9648
rect 509292 9636 509298 9648
rect 517238 9636 517244 9648
rect 509292 9608 517244 9636
rect 509292 9596 509298 9608
rect 517238 9596 517244 9608
rect 517296 9596 517302 9648
rect 202506 9528 202512 9580
rect 202564 9568 202570 9580
rect 202800 9568 202828 9596
rect 202564 9540 202828 9568
rect 202564 9528 202570 9540
rect 228910 9528 228916 9580
rect 228968 9568 228974 9580
rect 447134 9568 447140 9580
rect 228968 9540 447140 9568
rect 228968 9528 228974 9540
rect 447134 9528 447140 9540
rect 447192 9528 447198 9580
rect 218146 9460 218152 9512
rect 218204 9500 218210 9512
rect 443638 9500 443644 9512
rect 218204 9472 443644 9500
rect 218204 9460 218210 9472
rect 443638 9460 443644 9472
rect 443696 9460 443702 9512
rect 454126 9460 454132 9512
rect 454184 9500 454190 9512
rect 493134 9500 493140 9512
rect 454184 9472 493140 9500
rect 454184 9460 454190 9472
rect 493134 9460 493140 9472
rect 493192 9460 493198 9512
rect 204346 9392 204352 9444
rect 204404 9432 204410 9444
rect 436462 9432 436468 9444
rect 204404 9404 436468 9432
rect 204404 9392 204410 9404
rect 436462 9392 436468 9404
rect 436520 9392 436526 9444
rect 439774 9392 439780 9444
rect 439832 9432 439838 9444
rect 490834 9432 490840 9444
rect 439832 9404 490840 9432
rect 439832 9392 439838 9404
rect 490834 9392 490840 9404
rect 490892 9392 490898 9444
rect 510614 9392 510620 9444
rect 510672 9432 510678 9444
rect 521838 9432 521844 9444
rect 510672 9404 521844 9432
rect 510672 9392 510678 9404
rect 521838 9392 521844 9404
rect 521896 9392 521902 9444
rect 203886 9324 203892 9376
rect 203944 9364 203950 9376
rect 439038 9364 439044 9376
rect 203944 9336 439044 9364
rect 203944 9324 203950 9336
rect 439038 9324 439044 9336
rect 439096 9324 439102 9376
rect 445386 9324 445392 9376
rect 445444 9364 445450 9376
rect 516870 9364 516876 9376
rect 445444 9336 516876 9364
rect 445444 9324 445450 9336
rect 516870 9324 516876 9336
rect 516928 9324 516934 9376
rect 186038 9256 186044 9308
rect 186096 9296 186102 9308
rect 433334 9296 433340 9308
rect 186096 9268 433340 9296
rect 186096 9256 186102 9268
rect 433334 9256 433340 9268
rect 433392 9256 433398 9308
rect 438210 9256 438216 9308
rect 438268 9296 438274 9308
rect 514570 9296 514576 9308
rect 438268 9268 514576 9296
rect 438268 9256 438274 9268
rect 514570 9256 514576 9268
rect 514628 9256 514634 9308
rect 514662 9256 514668 9308
rect 514720 9296 514726 9308
rect 519538 9296 519544 9308
rect 514720 9268 519544 9296
rect 514720 9256 514726 9268
rect 519538 9256 519544 9268
rect 519596 9256 519602 9308
rect 531314 9256 531320 9308
rect 531372 9296 531378 9308
rect 540882 9296 540888 9308
rect 531372 9268 540888 9296
rect 531372 9256 531378 9268
rect 540882 9256 540888 9268
rect 540940 9256 540946 9308
rect 541066 9256 541072 9308
rect 541124 9296 541130 9308
rect 541124 9268 541296 9296
rect 541124 9256 541130 9268
rect 181346 9188 181352 9240
rect 181404 9228 181410 9240
rect 431034 9228 431040 9240
rect 181404 9200 431040 9228
rect 181404 9188 181410 9200
rect 431034 9188 431040 9200
rect 431092 9188 431098 9240
rect 431126 9188 431132 9240
rect 431184 9228 431190 9240
rect 512270 9228 512276 9240
rect 431184 9200 512276 9228
rect 431184 9188 431190 9200
rect 512270 9188 512276 9200
rect 512328 9188 512334 9240
rect 69474 9120 69480 9172
rect 69532 9160 69538 9172
rect 169754 9160 169760 9172
rect 69532 9132 169760 9160
rect 69532 9120 69538 9132
rect 169754 9120 169760 9132
rect 169812 9120 169818 9172
rect 182542 9120 182548 9172
rect 182600 9160 182606 9172
rect 432138 9160 432144 9172
rect 182600 9132 432144 9160
rect 182600 9120 182606 9132
rect 432138 9120 432144 9132
rect 432196 9120 432202 9172
rect 434622 9120 434628 9172
rect 434680 9160 434686 9172
rect 513466 9160 513472 9172
rect 434680 9132 513472 9160
rect 434680 9120 434686 9132
rect 513466 9120 513472 9132
rect 513524 9120 513530 9172
rect 520274 9120 520280 9172
rect 520332 9160 520338 9172
rect 531314 9160 531320 9172
rect 520332 9132 531320 9160
rect 520332 9120 520338 9132
rect 531314 9120 531320 9132
rect 531372 9120 531378 9172
rect 168190 9052 168196 9104
rect 168248 9092 168254 9104
rect 427262 9092 427268 9104
rect 168248 9064 427268 9092
rect 168248 9052 168254 9064
rect 427262 9052 427268 9064
rect 427320 9052 427326 9104
rect 427538 9052 427544 9104
rect 427596 9092 427602 9104
rect 511166 9092 511172 9104
rect 427596 9064 511172 9092
rect 427596 9052 427602 9064
rect 511166 9052 511172 9064
rect 511224 9052 511230 9104
rect 540882 9052 540888 9104
rect 540940 9092 540946 9104
rect 541268 9092 541296 9268
rect 540940 9064 541296 9092
rect 540940 9052 540946 9064
rect 151538 8984 151544 9036
rect 151596 9024 151602 9036
rect 411254 9024 411260 9036
rect 151596 8996 411260 9024
rect 151596 8984 151602 8996
rect 411254 8984 411260 8996
rect 411312 8984 411318 9036
rect 414474 8984 414480 9036
rect 414532 9024 414538 9036
rect 418522 9024 418528 9036
rect 414532 8996 418528 9024
rect 414532 8984 414538 8996
rect 418522 8984 418528 8996
rect 418580 8984 418586 9036
rect 419166 8984 419172 9036
rect 419224 9024 419230 9036
rect 508498 9024 508504 9036
rect 419224 8996 508504 9024
rect 419224 8984 419230 8996
rect 508498 8984 508504 8996
rect 508556 8984 508562 9036
rect 519078 8984 519084 9036
rect 519136 9024 519142 9036
rect 540698 9024 540704 9036
rect 519136 8996 540704 9024
rect 519136 8984 519142 8996
rect 540698 8984 540704 8996
rect 540756 8984 540762 9036
rect 23106 8916 23112 8968
rect 23164 8956 23170 8968
rect 135254 8956 135260 8968
rect 23164 8928 135260 8956
rect 23164 8916 23170 8928
rect 135254 8916 135260 8928
rect 135312 8916 135318 8968
rect 156322 8916 156328 8968
rect 156380 8956 156386 8968
rect 423766 8956 423772 8968
rect 156380 8928 423772 8956
rect 156380 8916 156386 8928
rect 423766 8916 423772 8928
rect 423824 8916 423830 8968
rect 426342 8916 426348 8968
rect 426400 8956 426406 8968
rect 510798 8956 510804 8968
rect 426400 8928 510804 8956
rect 426400 8916 426406 8928
rect 510798 8916 510804 8928
rect 510856 8916 510862 8968
rect 513190 8916 513196 8968
rect 513248 8956 513254 8968
rect 538766 8956 538772 8968
rect 513248 8928 538772 8956
rect 513248 8916 513254 8928
rect 538766 8916 538772 8928
rect 538824 8916 538830 8968
rect 334710 8848 334716 8900
rect 334768 8888 334774 8900
rect 481266 8888 481272 8900
rect 334768 8860 481272 8888
rect 334768 8848 334774 8860
rect 481266 8848 481272 8860
rect 481324 8848 481330 8900
rect 345658 8780 345664 8832
rect 345716 8820 345722 8832
rect 481634 8820 481640 8832
rect 345716 8792 481640 8820
rect 345716 8780 345722 8792
rect 481634 8780 481640 8792
rect 481692 8780 481698 8832
rect 510798 8780 510804 8832
rect 510856 8820 510862 8832
rect 511810 8820 511816 8832
rect 510856 8792 511816 8820
rect 510856 8780 510862 8792
rect 511810 8780 511816 8792
rect 511868 8780 511874 8832
rect 399018 8712 399024 8764
rect 399076 8752 399082 8764
rect 501966 8752 501972 8764
rect 399076 8724 501972 8752
rect 399076 8712 399082 8724
rect 501966 8712 501972 8724
rect 502024 8712 502030 8764
rect 412082 8644 412088 8696
rect 412140 8684 412146 8696
rect 420914 8684 420920 8696
rect 412140 8656 420920 8684
rect 412140 8644 412146 8656
rect 420914 8644 420920 8656
rect 420972 8644 420978 8696
rect 422754 8644 422760 8696
rect 422812 8684 422818 8696
rect 509602 8684 509608 8696
rect 422812 8656 509608 8684
rect 422812 8644 422818 8656
rect 509602 8644 509608 8656
rect 509660 8644 509666 8696
rect 371418 8576 371424 8628
rect 371476 8616 371482 8628
rect 454034 8616 454040 8628
rect 371476 8588 454040 8616
rect 371476 8576 371482 8588
rect 454034 8576 454040 8588
rect 454092 8576 454098 8628
rect 433334 8508 433340 8560
rect 433392 8548 433398 8560
rect 464338 8548 464344 8560
rect 433392 8520 464344 8548
rect 433392 8508 433398 8520
rect 464338 8508 464344 8520
rect 464396 8508 464402 8560
rect 307202 8304 307208 8356
rect 307260 8344 307266 8356
rect 307386 8344 307392 8356
rect 307260 8316 307392 8344
rect 307260 8304 307266 8316
rect 307386 8304 307392 8316
rect 307444 8304 307450 8356
rect 384482 8304 384488 8356
rect 384540 8344 384546 8356
rect 384666 8344 384672 8356
rect 384540 8316 384672 8344
rect 384540 8304 384546 8316
rect 384666 8304 384672 8316
rect 384724 8304 384730 8356
rect 372798 8236 372804 8288
rect 372856 8276 372862 8288
rect 493502 8276 493508 8288
rect 372856 8248 493508 8276
rect 372856 8236 372862 8248
rect 493502 8236 493508 8248
rect 493560 8236 493566 8288
rect 369210 8168 369216 8220
rect 369268 8208 369274 8220
rect 492398 8208 492404 8220
rect 369268 8180 492404 8208
rect 369268 8168 369274 8180
rect 492398 8168 492404 8180
rect 492456 8168 492462 8220
rect 113542 8100 113548 8152
rect 113600 8140 113606 8152
rect 201586 8140 201592 8152
rect 113600 8112 201592 8140
rect 113600 8100 113606 8112
rect 201586 8100 201592 8112
rect 201644 8100 201650 8152
rect 365714 8100 365720 8152
rect 365772 8140 365778 8152
rect 491202 8140 491208 8152
rect 365772 8112 491208 8140
rect 365772 8100 365778 8112
rect 491202 8100 491208 8112
rect 491260 8100 491266 8152
rect 117130 8032 117136 8084
rect 117188 8072 117194 8084
rect 204254 8072 204260 8084
rect 117188 8044 204260 8072
rect 117188 8032 117194 8044
rect 204254 8032 204260 8044
rect 204312 8032 204318 8084
rect 362126 8032 362132 8084
rect 362184 8072 362190 8084
rect 490098 8072 490104 8084
rect 362184 8044 490104 8072
rect 362184 8032 362190 8044
rect 490098 8032 490104 8044
rect 490156 8032 490162 8084
rect 109954 7964 109960 8016
rect 110012 8004 110018 8016
rect 199194 8004 199200 8016
rect 110012 7976 199200 8004
rect 110012 7964 110018 7976
rect 199194 7964 199200 7976
rect 199252 7964 199258 8016
rect 358538 7964 358544 8016
rect 358596 8004 358602 8016
rect 488902 8004 488908 8016
rect 358596 7976 488908 8004
rect 358596 7964 358602 7976
rect 488902 7964 488908 7976
rect 488960 7964 488966 8016
rect 510338 8004 510344 8016
rect 509528 7976 510344 8004
rect 102778 7896 102784 7948
rect 102836 7936 102842 7948
rect 194686 7936 194692 7948
rect 102836 7908 194692 7936
rect 102836 7896 102842 7908
rect 194686 7896 194692 7908
rect 194744 7896 194750 7948
rect 354950 7896 354956 7948
rect 355008 7936 355014 7948
rect 487798 7936 487804 7948
rect 355008 7908 487804 7936
rect 355008 7896 355014 7908
rect 487798 7896 487804 7908
rect 487856 7896 487862 7948
rect 99282 7828 99288 7880
rect 99340 7868 99346 7880
rect 191834 7868 191840 7880
rect 99340 7840 191840 7868
rect 99340 7828 99346 7840
rect 191834 7828 191840 7840
rect 191892 7828 191898 7880
rect 351362 7828 351368 7880
rect 351420 7868 351426 7880
rect 486602 7868 486608 7880
rect 351420 7840 486608 7868
rect 351420 7828 351426 7840
rect 486602 7828 486608 7840
rect 486660 7828 486666 7880
rect 493870 7828 493876 7880
rect 493928 7868 493934 7880
rect 509528 7868 509556 7976
rect 510338 7964 510344 7976
rect 510396 7964 510402 8016
rect 493928 7840 509556 7868
rect 493928 7828 493934 7840
rect 509602 7828 509608 7880
rect 509660 7868 509666 7880
rect 537570 7868 537576 7880
rect 509660 7840 537576 7868
rect 509660 7828 509666 7840
rect 537570 7828 537576 7840
rect 537628 7828 537634 7880
rect 92106 7760 92112 7812
rect 92164 7800 92170 7812
rect 186314 7800 186320 7812
rect 92164 7772 186320 7800
rect 92164 7760 92170 7772
rect 186314 7760 186320 7772
rect 186372 7760 186378 7812
rect 347866 7760 347872 7812
rect 347924 7800 347930 7812
rect 485498 7800 485504 7812
rect 347924 7772 485504 7800
rect 347924 7760 347930 7772
rect 485498 7760 485504 7772
rect 485556 7760 485562 7812
rect 490558 7760 490564 7812
rect 490616 7800 490622 7812
rect 531498 7800 531504 7812
rect 490616 7772 531504 7800
rect 490616 7760 490622 7772
rect 531498 7760 531504 7772
rect 531556 7760 531562 7812
rect 34974 7692 34980 7744
rect 35032 7732 35038 7744
rect 145006 7732 145012 7744
rect 35032 7704 145012 7732
rect 35032 7692 35038 7704
rect 145006 7692 145012 7704
rect 145064 7692 145070 7744
rect 344278 7692 344284 7744
rect 344336 7732 344342 7744
rect 484026 7732 484032 7744
rect 344336 7704 484032 7732
rect 344336 7692 344342 7704
rect 484026 7692 484032 7704
rect 484084 7692 484090 7744
rect 489362 7692 489368 7744
rect 489420 7732 489426 7744
rect 531038 7732 531044 7744
rect 489420 7704 531044 7732
rect 489420 7692 489426 7704
rect 531038 7692 531044 7704
rect 531096 7692 531102 7744
rect 18322 7624 18328 7676
rect 18380 7664 18386 7676
rect 132586 7664 132592 7676
rect 18380 7636 132592 7664
rect 18380 7624 18386 7636
rect 132586 7624 132592 7636
rect 132644 7624 132650 7676
rect 285950 7624 285956 7676
rect 286008 7664 286014 7676
rect 456794 7664 456800 7676
rect 286008 7636 456800 7664
rect 286008 7624 286014 7636
rect 456794 7624 456800 7636
rect 456852 7624 456858 7676
rect 456886 7624 456892 7676
rect 456944 7664 456950 7676
rect 457622 7664 457628 7676
rect 456944 7636 457628 7664
rect 456944 7624 456950 7636
rect 457622 7624 457628 7636
rect 457680 7624 457686 7676
rect 485774 7624 485780 7676
rect 485832 7664 485838 7676
rect 529934 7664 529940 7676
rect 485832 7636 529940 7664
rect 485832 7624 485838 7636
rect 529934 7624 529940 7636
rect 529992 7624 529998 7676
rect 13630 7556 13636 7608
rect 13688 7596 13694 7608
rect 128538 7596 128544 7608
rect 13688 7568 128544 7596
rect 13688 7556 13694 7568
rect 128538 7556 128544 7568
rect 128596 7556 128602 7608
rect 159910 7556 159916 7608
rect 159968 7596 159974 7608
rect 424870 7596 424876 7608
rect 159968 7568 424876 7596
rect 159968 7556 159974 7568
rect 424870 7556 424876 7568
rect 424928 7556 424934 7608
rect 426250 7556 426256 7608
rect 426308 7596 426314 7608
rect 496538 7596 496544 7608
rect 426308 7568 496544 7596
rect 426308 7556 426314 7568
rect 496538 7556 496544 7568
rect 496596 7556 496602 7608
rect 504818 7556 504824 7608
rect 504876 7596 504882 7608
rect 535822 7596 535828 7608
rect 504876 7568 535828 7596
rect 504876 7556 504882 7568
rect 535822 7556 535828 7568
rect 535880 7556 535886 7608
rect 383562 7488 383568 7540
rect 383620 7528 383626 7540
rect 496998 7528 497004 7540
rect 383620 7500 497004 7528
rect 383620 7488 383626 7500
rect 496998 7488 497004 7500
rect 497056 7488 497062 7540
rect 408494 7420 408500 7472
rect 408552 7460 408558 7472
rect 504726 7460 504732 7472
rect 408552 7432 504732 7460
rect 408552 7420 408558 7432
rect 504726 7420 504732 7432
rect 504784 7420 504790 7472
rect 413186 7352 413192 7404
rect 413244 7392 413250 7404
rect 506566 7392 506572 7404
rect 413244 7364 506572 7392
rect 413244 7352 413250 7364
rect 506566 7352 506572 7364
rect 506624 7352 506630 7404
rect 340690 7284 340696 7336
rect 340748 7324 340754 7336
rect 419626 7324 419632 7336
rect 340748 7296 419632 7324
rect 340748 7284 340754 7296
rect 419626 7284 419632 7296
rect 419684 7284 419690 7336
rect 420362 7284 420368 7336
rect 420420 7324 420426 7336
rect 508866 7324 508872 7336
rect 420420 7296 508872 7324
rect 420420 7284 420426 7296
rect 508866 7284 508872 7296
rect 508924 7284 508930 7336
rect 385034 7216 385040 7268
rect 385092 7256 385098 7268
rect 461210 7256 461216 7268
rect 385092 7228 461216 7256
rect 385092 7216 385098 7228
rect 461210 7216 461216 7228
rect 461268 7216 461274 7268
rect 437566 7148 437572 7200
rect 437624 7188 437630 7200
rect 438026 7188 438032 7200
rect 437624 7160 438032 7188
rect 437624 7148 437630 7160
rect 438026 7148 438032 7160
rect 438084 7148 438090 7200
rect 448698 7148 448704 7200
rect 448756 7188 448762 7200
rect 449618 7188 449624 7200
rect 448756 7160 449624 7188
rect 448756 7148 448762 7160
rect 449618 7148 449624 7160
rect 449676 7148 449682 7200
rect 456794 7148 456800 7200
rect 456852 7188 456858 7200
rect 465534 7188 465540 7200
rect 456852 7160 465540 7188
rect 456852 7148 456858 7160
rect 465534 7148 465540 7160
rect 465592 7148 465598 7200
rect 429470 6876 429476 6928
rect 429528 6916 429534 6928
rect 430114 6916 430120 6928
rect 429528 6888 430120 6916
rect 429528 6876 429534 6888
rect 430114 6876 430120 6888
rect 430172 6876 430178 6928
rect 476206 6876 476212 6928
rect 476264 6916 476270 6928
rect 477218 6916 477224 6928
rect 476264 6888 477224 6916
rect 476264 6876 476270 6888
rect 477218 6876 477224 6888
rect 477276 6876 477282 6928
rect 67174 6808 67180 6860
rect 67232 6848 67238 6860
rect 168374 6848 168380 6860
rect 67232 6820 168380 6848
rect 67232 6808 67238 6820
rect 168374 6808 168380 6820
rect 168432 6808 168438 6860
rect 297910 6808 297916 6860
rect 297968 6848 297974 6860
rect 469398 6848 469404 6860
rect 297968 6820 469404 6848
rect 297968 6808 297974 6820
rect 469398 6808 469404 6820
rect 469456 6808 469462 6860
rect 493686 6808 493692 6860
rect 493744 6848 493750 6860
rect 498930 6848 498936 6860
rect 493744 6820 498936 6848
rect 493744 6808 493750 6820
rect 498930 6808 498936 6820
rect 498988 6808 498994 6860
rect 63586 6740 63592 6792
rect 63644 6780 63650 6792
rect 165614 6780 165620 6792
rect 63644 6752 165620 6780
rect 63644 6740 63650 6752
rect 165614 6740 165620 6752
rect 165672 6740 165678 6792
rect 294322 6740 294328 6792
rect 294380 6780 294386 6792
rect 467926 6780 467932 6792
rect 294380 6752 467932 6780
rect 294380 6740 294386 6752
rect 467926 6740 467932 6752
rect 467984 6740 467990 6792
rect 502426 6740 502432 6792
rect 502484 6780 502490 6792
rect 534350 6780 534356 6792
rect 502484 6752 534356 6780
rect 502484 6740 502490 6752
rect 534350 6740 534356 6752
rect 534408 6740 534414 6792
rect 59998 6672 60004 6724
rect 60056 6712 60062 6724
rect 162854 6712 162860 6724
rect 60056 6684 162860 6712
rect 60056 6672 60062 6684
rect 162854 6672 162860 6684
rect 162912 6672 162918 6724
rect 290734 6672 290740 6724
rect 290792 6712 290798 6724
rect 466914 6712 466920 6724
rect 290792 6684 466920 6712
rect 290792 6672 290798 6684
rect 466914 6672 466920 6684
rect 466972 6672 466978 6724
rect 498930 6672 498936 6724
rect 498988 6712 498994 6724
rect 534166 6712 534172 6724
rect 498988 6684 534172 6712
rect 498988 6672 498994 6684
rect 534166 6672 534172 6684
rect 534224 6672 534230 6724
rect 52822 6604 52828 6656
rect 52880 6644 52886 6656
rect 157334 6644 157340 6656
rect 52880 6616 157340 6644
rect 52880 6604 52886 6616
rect 157334 6604 157340 6616
rect 157392 6604 157398 6656
rect 287146 6604 287152 6656
rect 287204 6644 287210 6656
rect 465626 6644 465632 6656
rect 287204 6616 465632 6644
rect 287204 6604 287210 6616
rect 465626 6604 465632 6616
rect 465684 6604 465690 6656
rect 495250 6604 495256 6656
rect 495308 6644 495314 6656
rect 532878 6644 532884 6656
rect 495308 6616 532884 6644
rect 495308 6604 495314 6616
rect 532878 6604 532884 6616
rect 532936 6604 532942 6656
rect 56410 6536 56416 6588
rect 56468 6576 56474 6588
rect 160094 6576 160100 6588
rect 56468 6548 160100 6576
rect 56468 6536 56474 6548
rect 160094 6536 160100 6548
rect 160152 6536 160158 6588
rect 283650 6536 283656 6588
rect 283708 6576 283714 6588
rect 464430 6576 464436 6588
rect 283708 6548 464436 6576
rect 283708 6536 283714 6548
rect 464430 6536 464436 6548
rect 464488 6536 464494 6588
rect 491754 6536 491760 6588
rect 491812 6576 491818 6588
rect 531682 6576 531688 6588
rect 491812 6548 531688 6576
rect 491812 6536 491818 6548
rect 531682 6536 531688 6548
rect 531740 6536 531746 6588
rect 49326 6468 49332 6520
rect 49384 6508 49390 6520
rect 154574 6508 154580 6520
rect 49384 6480 154580 6508
rect 49384 6468 49390 6480
rect 154574 6468 154580 6480
rect 154632 6468 154638 6520
rect 279970 6468 279976 6520
rect 280028 6508 280034 6520
rect 463326 6508 463332 6520
rect 280028 6480 463332 6508
rect 280028 6468 280034 6480
rect 463326 6468 463332 6480
rect 463384 6468 463390 6520
rect 488166 6468 488172 6520
rect 488224 6508 488230 6520
rect 530118 6508 530124 6520
rect 488224 6480 530124 6508
rect 488224 6468 488230 6480
rect 530118 6468 530124 6480
rect 530176 6468 530182 6520
rect 44542 6400 44548 6452
rect 44600 6440 44606 6452
rect 151814 6440 151820 6452
rect 44600 6412 151820 6440
rect 44600 6400 44606 6412
rect 151814 6400 151820 6412
rect 151872 6400 151878 6452
rect 276474 6400 276480 6452
rect 276532 6440 276538 6452
rect 276532 6412 459968 6440
rect 276532 6400 276538 6412
rect 40954 6332 40960 6384
rect 41012 6372 41018 6384
rect 149054 6372 149060 6384
rect 41012 6344 149060 6372
rect 41012 6332 41018 6344
rect 149054 6332 149060 6344
rect 149112 6332 149118 6384
rect 269298 6332 269304 6384
rect 269356 6372 269362 6384
rect 459830 6372 459836 6384
rect 269356 6344 459836 6372
rect 269356 6332 269362 6344
rect 459830 6332 459836 6344
rect 459888 6332 459894 6384
rect 459940 6372 459968 6412
rect 462314 6400 462320 6452
rect 462372 6440 462378 6452
rect 484486 6440 484492 6452
rect 462372 6412 484492 6440
rect 462372 6400 462378 6412
rect 484486 6400 484492 6412
rect 484544 6400 484550 6452
rect 484578 6400 484584 6452
rect 484636 6440 484642 6452
rect 528646 6440 528652 6452
rect 484636 6412 528652 6440
rect 484636 6400 484642 6412
rect 528646 6400 528652 6412
rect 528704 6400 528710 6452
rect 462406 6372 462412 6384
rect 459940 6344 462412 6372
rect 462406 6332 462412 6344
rect 462464 6332 462470 6384
rect 479886 6332 479892 6384
rect 479944 6372 479950 6384
rect 527726 6372 527732 6384
rect 479944 6344 527732 6372
rect 479944 6332 479950 6344
rect 527726 6332 527732 6344
rect 527784 6332 527790 6384
rect 37366 6264 37372 6316
rect 37424 6304 37430 6316
rect 146294 6304 146300 6316
rect 37424 6276 146300 6304
rect 37424 6264 37430 6276
rect 146294 6264 146300 6276
rect 146352 6264 146358 6316
rect 161106 6264 161112 6316
rect 161164 6304 161170 6316
rect 250530 6304 250536 6316
rect 161164 6276 250536 6304
rect 161164 6264 161170 6276
rect 250530 6264 250536 6276
rect 250588 6264 250594 6316
rect 261018 6264 261024 6316
rect 261076 6304 261082 6316
rect 456978 6304 456984 6316
rect 261076 6276 456984 6304
rect 261076 6264 261082 6276
rect 456978 6264 456984 6276
rect 457036 6264 457042 6316
rect 476298 6264 476304 6316
rect 476356 6304 476362 6316
rect 526622 6304 526628 6316
rect 476356 6276 526628 6304
rect 476356 6264 476362 6276
rect 526622 6264 526628 6276
rect 526680 6264 526686 6316
rect 8846 6196 8852 6248
rect 8904 6236 8910 6248
rect 125594 6236 125600 6248
rect 8904 6208 125600 6236
rect 8904 6196 8910 6208
rect 125594 6196 125600 6208
rect 125652 6196 125658 6248
rect 221734 6196 221740 6248
rect 221792 6236 221798 6248
rect 444650 6236 444656 6248
rect 221792 6208 444656 6236
rect 221792 6196 221798 6208
rect 444650 6196 444656 6208
rect 444708 6196 444714 6248
rect 463234 6196 463240 6248
rect 463292 6236 463298 6248
rect 522390 6236 522396 6248
rect 463292 6208 522396 6236
rect 463292 6196 463298 6208
rect 522390 6196 522396 6208
rect 522448 6196 522454 6248
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 121638 6168 121644 6180
rect 4120 6140 121644 6168
rect 4120 6128 4126 6140
rect 121638 6128 121644 6140
rect 121696 6128 121702 6180
rect 206278 6128 206284 6180
rect 206336 6168 206342 6180
rect 439590 6168 439596 6180
rect 206336 6140 439596 6168
rect 206336 6128 206342 6140
rect 439590 6128 439596 6140
rect 439648 6128 439654 6180
rect 459646 6128 459652 6180
rect 459704 6168 459710 6180
rect 521194 6168 521200 6180
rect 459704 6140 521200 6168
rect 459704 6128 459710 6140
rect 521194 6128 521200 6140
rect 521252 6128 521258 6180
rect 70670 6060 70676 6112
rect 70728 6100 70734 6112
rect 171134 6100 171140 6112
rect 70728 6072 171140 6100
rect 70728 6060 70734 6072
rect 171134 6060 171140 6072
rect 171192 6060 171198 6112
rect 301406 6060 301412 6112
rect 301464 6100 301470 6112
rect 470226 6100 470232 6112
rect 301464 6072 470232 6100
rect 301464 6060 301470 6072
rect 470226 6060 470232 6072
rect 470284 6060 470290 6112
rect 74258 5992 74264 6044
rect 74316 6032 74322 6044
rect 172606 6032 172612 6044
rect 74316 6004 172612 6032
rect 74316 5992 74322 6004
rect 172606 5992 172612 6004
rect 172664 5992 172670 6044
rect 327626 5992 327632 6044
rect 327684 6032 327690 6044
rect 478966 6032 478972 6044
rect 327684 6004 478972 6032
rect 327684 5992 327690 6004
rect 478966 5992 478972 6004
rect 479024 5992 479030 6044
rect 77846 5924 77852 5976
rect 77904 5964 77910 5976
rect 175550 5964 175556 5976
rect 77904 5936 175556 5964
rect 77904 5924 77910 5936
rect 175550 5924 175556 5936
rect 175608 5924 175614 5976
rect 353754 5924 353760 5976
rect 353812 5964 353818 5976
rect 487154 5964 487160 5976
rect 353812 5936 487160 5964
rect 353812 5924 353818 5936
rect 487154 5924 487160 5936
rect 487212 5924 487218 5976
rect 356146 5856 356152 5908
rect 356204 5896 356210 5908
rect 487246 5896 487252 5908
rect 356204 5868 487252 5896
rect 356204 5856 356210 5868
rect 487246 5856 487252 5868
rect 487304 5856 487310 5908
rect 394234 5788 394240 5840
rect 394292 5828 394298 5840
rect 500126 5828 500132 5840
rect 394292 5800 500132 5828
rect 394292 5788 394298 5800
rect 500126 5788 500132 5800
rect 500184 5788 500190 5840
rect 439038 5720 439044 5772
rect 439096 5760 439102 5772
rect 477586 5760 477592 5772
rect 439096 5732 477592 5760
rect 439096 5720 439102 5732
rect 477586 5720 477592 5732
rect 477644 5720 477650 5772
rect 457254 5652 457260 5704
rect 457312 5692 457318 5704
rect 491938 5692 491944 5704
rect 457312 5664 491944 5692
rect 457312 5652 457318 5664
rect 491938 5652 491944 5664
rect 491996 5652 492002 5704
rect 455966 5584 455972 5636
rect 456024 5624 456030 5636
rect 481726 5624 481732 5636
rect 456024 5596 481732 5624
rect 456024 5584 456030 5596
rect 481726 5584 481732 5596
rect 481784 5584 481790 5636
rect 535270 5584 535276 5636
rect 535328 5624 535334 5636
rect 542722 5624 542728 5636
rect 535328 5596 542728 5624
rect 535328 5584 535334 5596
rect 542722 5584 542728 5596
rect 542780 5584 542786 5636
rect 570598 5516 570604 5568
rect 570656 5556 570662 5568
rect 572622 5556 572628 5568
rect 570656 5528 572628 5556
rect 570656 5516 570662 5528
rect 572622 5516 572628 5528
rect 572680 5516 572686 5568
rect 108758 5448 108764 5500
rect 108816 5488 108822 5500
rect 198734 5488 198740 5500
rect 108816 5460 198740 5488
rect 108816 5448 108822 5460
rect 198734 5448 198740 5460
rect 198792 5448 198798 5500
rect 263594 5448 263600 5500
rect 263652 5488 263658 5500
rect 421098 5488 421104 5500
rect 263652 5460 421104 5488
rect 263652 5448 263658 5460
rect 421098 5448 421104 5460
rect 421156 5448 421162 5500
rect 437014 5448 437020 5500
rect 437072 5488 437078 5500
rect 513558 5488 513564 5500
rect 437072 5460 513564 5488
rect 437072 5448 437078 5460
rect 513558 5448 513564 5460
rect 513616 5448 513622 5500
rect 101582 5380 101588 5432
rect 101640 5420 101646 5432
rect 193214 5420 193220 5432
rect 101640 5392 193220 5420
rect 101640 5380 101646 5392
rect 193214 5380 193220 5392
rect 193272 5380 193278 5432
rect 303798 5380 303804 5432
rect 303856 5420 303862 5432
rect 470594 5420 470600 5432
rect 303856 5392 470600 5420
rect 303856 5380 303862 5392
rect 470594 5380 470600 5392
rect 470652 5380 470658 5432
rect 508406 5380 508412 5432
rect 508464 5420 508470 5432
rect 537018 5420 537024 5432
rect 508464 5392 537024 5420
rect 508464 5380 508470 5392
rect 537018 5380 537024 5392
rect 537076 5380 537082 5432
rect 98086 5312 98092 5364
rect 98144 5352 98150 5364
rect 190454 5352 190460 5364
rect 98144 5324 190460 5352
rect 98144 5312 98150 5324
rect 190454 5312 190460 5324
rect 190512 5312 190518 5364
rect 256234 5312 256240 5364
rect 256292 5352 256298 5364
rect 455782 5352 455788 5364
rect 256292 5324 455788 5352
rect 256292 5312 256298 5324
rect 455782 5312 455788 5324
rect 455840 5312 455846 5364
rect 465626 5312 465632 5364
rect 465684 5352 465690 5364
rect 523126 5352 523132 5364
rect 465684 5324 523132 5352
rect 465684 5312 465690 5324
rect 523126 5312 523132 5324
rect 523184 5312 523190 5364
rect 94498 5244 94504 5296
rect 94556 5284 94562 5296
rect 187694 5284 187700 5296
rect 94556 5256 187700 5284
rect 94556 5244 94562 5256
rect 187694 5244 187700 5256
rect 187752 5244 187758 5296
rect 255038 5244 255044 5296
rect 255096 5284 255102 5296
rect 455506 5284 455512 5296
rect 255096 5256 455512 5284
rect 255096 5244 255102 5256
rect 455506 5244 455512 5256
rect 455564 5244 455570 5296
rect 462038 5244 462044 5296
rect 462096 5284 462102 5296
rect 522022 5284 522028 5296
rect 462096 5256 522028 5284
rect 462096 5244 462102 5256
rect 522022 5244 522028 5256
rect 522080 5244 522086 5296
rect 87322 5176 87328 5228
rect 87380 5216 87386 5228
rect 182174 5216 182180 5228
rect 87380 5188 182180 5216
rect 87380 5176 87386 5188
rect 182174 5176 182180 5188
rect 182232 5176 182238 5228
rect 235994 5176 236000 5228
rect 236052 5216 236058 5228
rect 449158 5216 449164 5228
rect 236052 5188 449164 5216
rect 236052 5176 236058 5188
rect 449158 5176 449164 5188
rect 449216 5176 449222 5228
rect 458450 5176 458456 5228
rect 458508 5216 458514 5228
rect 520918 5216 520924 5228
rect 458508 5188 520924 5216
rect 458508 5176 458514 5188
rect 520918 5176 520924 5188
rect 520976 5176 520982 5228
rect 90910 5108 90916 5160
rect 90968 5148 90974 5160
rect 185118 5148 185124 5160
rect 90968 5120 185124 5148
rect 90968 5108 90974 5120
rect 185118 5108 185124 5120
rect 185176 5108 185182 5160
rect 230106 5108 230112 5160
rect 230164 5148 230170 5160
rect 447410 5148 447416 5160
rect 230164 5120 447416 5148
rect 230164 5108 230170 5120
rect 447410 5108 447416 5120
rect 447468 5108 447474 5160
rect 454862 5108 454868 5160
rect 454920 5148 454926 5160
rect 519630 5148 519636 5160
rect 454920 5120 519636 5148
rect 454920 5108 454926 5120
rect 519630 5108 519636 5120
rect 519688 5108 519694 5160
rect 83826 5040 83832 5092
rect 83884 5080 83890 5092
rect 179506 5080 179512 5092
rect 83884 5052 179512 5080
rect 83884 5040 83890 5052
rect 179506 5040 179512 5052
rect 179564 5040 179570 5092
rect 226518 5040 226524 5092
rect 226576 5080 226582 5092
rect 446122 5080 446128 5092
rect 226576 5052 446128 5080
rect 226576 5040 226582 5052
rect 446122 5040 446128 5052
rect 446180 5040 446186 5092
rect 451274 5040 451280 5092
rect 451332 5080 451338 5092
rect 518618 5080 518624 5092
rect 451332 5052 518624 5080
rect 451332 5040 451338 5052
rect 518618 5040 518624 5052
rect 518676 5040 518682 5092
rect 80238 4972 80244 5024
rect 80296 5012 80302 5024
rect 178034 5012 178040 5024
rect 80296 4984 178040 5012
rect 80296 4972 80302 4984
rect 178034 4972 178040 4984
rect 178092 4972 178098 5024
rect 219342 4972 219348 5024
rect 219400 5012 219406 5024
rect 443822 5012 443828 5024
rect 219400 4984 443828 5012
rect 219400 4972 219406 4984
rect 443822 4972 443828 4984
rect 443880 4972 443886 5024
rect 447778 4972 447784 5024
rect 447836 5012 447842 5024
rect 517606 5012 517612 5024
rect 447836 4984 517612 5012
rect 447836 4972 447842 4984
rect 517606 4972 517612 4984
rect 517664 4972 517670 5024
rect 76650 4904 76656 4956
rect 76708 4944 76714 4956
rect 175274 4944 175280 4956
rect 76708 4916 175280 4944
rect 76708 4904 76714 4916
rect 175274 4904 175280 4916
rect 175332 4904 175338 4956
rect 215846 4904 215852 4956
rect 215904 4944 215910 4956
rect 442718 4944 442724 4956
rect 215904 4916 442724 4944
rect 215904 4904 215910 4916
rect 442718 4904 442724 4916
rect 442776 4904 442782 4956
rect 443914 4904 443920 4956
rect 443972 4944 443978 4956
rect 516318 4944 516324 4956
rect 443972 4916 516324 4944
rect 443972 4904 443978 4916
rect 516318 4904 516324 4916
rect 516376 4904 516382 4956
rect 73062 4836 73068 4888
rect 73120 4876 73126 4888
rect 172514 4876 172520 4888
rect 73120 4848 172520 4876
rect 73120 4836 73126 4848
rect 172514 4836 172520 4848
rect 172572 4836 172578 4888
rect 178954 4836 178960 4888
rect 179012 4876 179018 4888
rect 428458 4876 428464 4888
rect 179012 4848 428464 4876
rect 179012 4836 179018 4848
rect 428458 4836 428464 4848
rect 428516 4836 428522 4888
rect 433518 4836 433524 4888
rect 433576 4876 433582 4888
rect 512086 4876 512092 4888
rect 433576 4848 512092 4876
rect 433576 4836 433582 4848
rect 512086 4836 512092 4848
rect 512144 4836 512150 4888
rect 515582 4836 515588 4888
rect 515640 4876 515646 4888
rect 539226 4876 539232 4888
rect 515640 4848 539232 4876
rect 515640 4836 515646 4848
rect 539226 4836 539232 4848
rect 539284 4836 539290 4888
rect 12434 4768 12440 4820
rect 12492 4808 12498 4820
rect 128354 4808 128360 4820
rect 12492 4780 128360 4808
rect 12492 4768 12498 4780
rect 128354 4768 128360 4780
rect 128412 4768 128418 4820
rect 167086 4768 167092 4820
rect 167144 4808 167150 4820
rect 426526 4808 426532 4820
rect 167144 4780 426532 4808
rect 167144 4768 167150 4780
rect 426526 4768 426532 4780
rect 426584 4768 426590 4820
rect 429930 4768 429936 4820
rect 429988 4808 429994 4820
rect 510798 4808 510804 4820
rect 429988 4780 510804 4808
rect 429988 4768 429994 4780
rect 510798 4768 510804 4780
rect 510856 4768 510862 4820
rect 511994 4768 512000 4820
rect 512052 4808 512058 4820
rect 538398 4808 538404 4820
rect 512052 4780 538404 4808
rect 512052 4768 512058 4780
rect 538398 4768 538404 4780
rect 538456 4768 538462 4820
rect 105170 4700 105176 4752
rect 105228 4740 105234 4752
rect 195974 4740 195980 4752
rect 105228 4712 195980 4740
rect 105228 4700 105234 4712
rect 195974 4700 195980 4712
rect 196032 4700 196038 4752
rect 331214 4700 331220 4752
rect 331272 4740 331278 4752
rect 479058 4740 479064 4752
rect 331272 4712 479064 4740
rect 331272 4700 331278 4712
rect 479058 4700 479064 4712
rect 479116 4700 479122 4752
rect 482278 4700 482284 4752
rect 482336 4740 482342 4752
rect 482922 4740 482928 4752
rect 482336 4712 482928 4740
rect 482336 4700 482342 4712
rect 482922 4700 482928 4712
rect 482980 4700 482986 4752
rect 120626 4632 120632 4684
rect 120684 4672 120690 4684
rect 207014 4672 207020 4684
rect 120684 4644 207020 4672
rect 120684 4632 120690 4644
rect 207014 4632 207020 4644
rect 207072 4632 207078 4684
rect 375282 4632 375288 4684
rect 375340 4672 375346 4684
rect 494146 4672 494152 4684
rect 375340 4644 494152 4672
rect 375340 4632 375346 4644
rect 494146 4632 494152 4644
rect 494204 4632 494210 4684
rect 123018 4564 123024 4616
rect 123076 4604 123082 4616
rect 208762 4604 208768 4616
rect 123076 4576 208768 4604
rect 123076 4564 123082 4576
rect 208762 4564 208768 4576
rect 208820 4564 208826 4616
rect 403710 4564 403716 4616
rect 403768 4604 403774 4616
rect 503162 4604 503168 4616
rect 403768 4576 503168 4604
rect 403768 4564 403774 4576
rect 503162 4564 503168 4576
rect 503220 4564 503226 4616
rect 378134 4496 378140 4548
rect 378192 4536 378198 4548
rect 458358 4536 458364 4548
rect 378192 4508 458364 4536
rect 378192 4496 378198 4508
rect 458358 4496 458364 4508
rect 458416 4496 458422 4548
rect 469122 4496 469128 4548
rect 469180 4536 469186 4548
rect 524598 4536 524604 4548
rect 469180 4508 524604 4536
rect 469180 4496 469186 4508
rect 524598 4496 524604 4508
rect 524656 4496 524662 4548
rect 411162 4428 411168 4480
rect 411220 4468 411226 4480
rect 422294 4468 422300 4480
rect 411220 4440 422300 4468
rect 411220 4428 411226 4440
rect 422294 4428 422300 4440
rect 422352 4428 422358 4480
rect 427078 4428 427084 4480
rect 427136 4468 427142 4480
rect 461762 4468 461768 4480
rect 427136 4440 461768 4468
rect 427136 4428 427142 4440
rect 461762 4428 461768 4440
rect 461820 4428 461826 4480
rect 384850 4360 384856 4412
rect 384908 4400 384914 4412
rect 393222 4400 393228 4412
rect 384908 4372 393228 4400
rect 384908 4360 384914 4372
rect 393222 4360 393228 4372
rect 393280 4360 393286 4412
rect 442994 4360 443000 4412
rect 443052 4400 443058 4412
rect 468662 4400 468668 4412
rect 443052 4372 468668 4400
rect 443052 4360 443058 4372
rect 468662 4360 468668 4372
rect 468720 4360 468726 4412
rect 389266 4264 389272 4276
rect 386892 4236 389272 4264
rect 381096 4168 382320 4196
rect 1670 4088 1676 4140
rect 1728 4128 1734 4140
rect 9030 4128 9036 4140
rect 1728 4100 9036 4128
rect 1728 4088 1734 4100
rect 9030 4088 9036 4100
rect 9088 4088 9094 4140
rect 81434 4088 81440 4140
rect 81492 4128 81498 4140
rect 82722 4128 82728 4140
rect 81492 4100 82728 4128
rect 81492 4088 81498 4100
rect 82722 4088 82728 4100
rect 82780 4088 82786 4140
rect 84930 4088 84936 4140
rect 84988 4128 84994 4140
rect 85482 4128 85488 4140
rect 84988 4100 85488 4128
rect 84988 4088 84994 4100
rect 85482 4088 85488 4100
rect 85540 4088 85546 4140
rect 88518 4088 88524 4140
rect 88576 4128 88582 4140
rect 89622 4128 89628 4140
rect 88576 4100 89628 4128
rect 88576 4088 88582 4100
rect 89622 4088 89628 4100
rect 89680 4088 89686 4140
rect 93302 4088 93308 4140
rect 93360 4128 93366 4140
rect 93762 4128 93768 4140
rect 93360 4100 93768 4128
rect 93360 4088 93366 4100
rect 93762 4088 93768 4100
rect 93820 4088 93826 4140
rect 95694 4088 95700 4140
rect 95752 4128 95758 4140
rect 96522 4128 96528 4140
rect 95752 4100 96528 4128
rect 95752 4088 95758 4100
rect 96522 4088 96528 4100
rect 96580 4088 96586 4140
rect 103514 4088 103520 4140
rect 103572 4128 103578 4140
rect 112990 4128 112996 4140
rect 103572 4100 112996 4128
rect 103572 4088 103578 4100
rect 112990 4088 112996 4100
rect 113048 4088 113054 4140
rect 121822 4088 121828 4140
rect 121880 4128 121886 4140
rect 123478 4128 123484 4140
rect 121880 4100 123484 4128
rect 121880 4088 121886 4100
rect 123478 4088 123484 4100
rect 123536 4088 123542 4140
rect 137278 4088 137284 4140
rect 137336 4128 137342 4140
rect 198182 4128 198188 4140
rect 137336 4100 198188 4128
rect 137336 4088 137342 4100
rect 198182 4088 198188 4100
rect 198240 4088 198246 4140
rect 200390 4088 200396 4140
rect 200448 4128 200454 4140
rect 201402 4128 201408 4140
rect 200448 4100 201408 4128
rect 200448 4088 200454 4100
rect 201402 4088 201408 4100
rect 201460 4088 201466 4140
rect 214650 4088 214656 4140
rect 214708 4128 214714 4140
rect 215202 4128 215208 4140
rect 214708 4100 215208 4128
rect 214708 4088 214714 4100
rect 215202 4088 215208 4100
rect 215260 4088 215266 4140
rect 271690 4088 271696 4140
rect 271748 4128 271754 4140
rect 381096 4128 381124 4168
rect 271748 4100 381124 4128
rect 271748 4088 271754 4100
rect 381170 4088 381176 4140
rect 381228 4128 381234 4140
rect 382182 4128 382188 4140
rect 381228 4100 382188 4128
rect 381228 4088 381234 4100
rect 382182 4088 382188 4100
rect 382240 4088 382246 4140
rect 382292 4128 382320 4168
rect 385034 4128 385040 4140
rect 382292 4100 385040 4128
rect 385034 4088 385040 4100
rect 385092 4088 385098 4140
rect 111150 4020 111156 4072
rect 111208 4060 111214 4072
rect 171594 4060 171600 4072
rect 111208 4032 171600 4060
rect 111208 4020 111214 4032
rect 171594 4020 171600 4032
rect 171652 4020 171658 4072
rect 171778 4020 171784 4072
rect 171836 4060 171842 4072
rect 172422 4060 172428 4072
rect 171836 4032 172428 4060
rect 171836 4020 171842 4032
rect 172422 4020 172428 4032
rect 172480 4020 172486 4072
rect 197998 4020 198004 4072
rect 198056 4060 198062 4072
rect 275278 4060 275284 4072
rect 198056 4032 275284 4060
rect 198056 4020 198062 4032
rect 275278 4020 275284 4032
rect 275336 4020 275342 4072
rect 277670 4020 277676 4072
rect 277728 4060 277734 4072
rect 278682 4060 278688 4072
rect 277728 4032 278688 4060
rect 277728 4020 277734 4032
rect 278682 4020 278688 4032
rect 278740 4020 278746 4072
rect 278866 4020 278872 4072
rect 278924 4060 278930 4072
rect 280062 4060 280068 4072
rect 278924 4032 280068 4060
rect 278924 4020 278930 4032
rect 280062 4020 280068 4032
rect 280120 4020 280126 4072
rect 293126 4020 293132 4072
rect 293184 4060 293190 4072
rect 293862 4060 293868 4072
rect 293184 4032 293868 4060
rect 293184 4020 293190 4032
rect 293862 4020 293868 4032
rect 293920 4020 293926 4072
rect 300302 4020 300308 4072
rect 300360 4060 300366 4072
rect 300762 4060 300768 4072
rect 300360 4032 300768 4060
rect 300360 4020 300366 4032
rect 300762 4020 300768 4032
rect 300820 4020 300826 4072
rect 313918 4020 313924 4072
rect 313976 4060 313982 4072
rect 323026 4060 323032 4072
rect 313976 4032 323032 4060
rect 313976 4020 313982 4032
rect 323026 4020 323032 4032
rect 323084 4020 323090 4072
rect 325234 4020 325240 4072
rect 325292 4060 325298 4072
rect 386892 4060 386920 4236
rect 389266 4224 389272 4236
rect 389324 4224 389330 4276
rect 387058 4088 387064 4140
rect 387116 4128 387122 4140
rect 387702 4128 387708 4140
rect 387116 4100 387708 4128
rect 387116 4088 387122 4100
rect 387702 4088 387708 4100
rect 387760 4088 387766 4140
rect 389450 4088 389456 4140
rect 389508 4128 389514 4140
rect 390462 4128 390468 4140
rect 389508 4100 390468 4128
rect 389508 4088 389514 4100
rect 390462 4088 390468 4100
rect 390520 4088 390526 4140
rect 395430 4088 395436 4140
rect 395488 4128 395494 4140
rect 395982 4128 395988 4140
rect 395488 4100 395988 4128
rect 395488 4088 395494 4100
rect 395982 4088 395988 4100
rect 396040 4088 396046 4140
rect 396626 4088 396632 4140
rect 396684 4128 396690 4140
rect 397362 4128 397368 4140
rect 396684 4100 397368 4128
rect 396684 4088 396690 4100
rect 397362 4088 397368 4100
rect 397420 4088 397426 4140
rect 397454 4088 397460 4140
rect 397512 4128 397518 4140
rect 499758 4128 499764 4140
rect 397512 4100 499764 4128
rect 397512 4088 397518 4100
rect 499758 4088 499764 4100
rect 499816 4088 499822 4140
rect 516778 4088 516784 4140
rect 516836 4128 516842 4140
rect 517422 4128 517428 4140
rect 516836 4100 517428 4128
rect 516836 4088 516842 4100
rect 517422 4088 517428 4100
rect 517480 4088 517486 4140
rect 525058 4088 525064 4140
rect 525116 4128 525122 4140
rect 525702 4128 525708 4140
rect 525116 4100 525708 4128
rect 525116 4088 525122 4100
rect 525702 4088 525708 4100
rect 525760 4088 525766 4140
rect 527450 4088 527456 4140
rect 527508 4128 527514 4140
rect 528462 4128 528468 4140
rect 527508 4100 528468 4128
rect 527508 4088 527514 4100
rect 528462 4088 528468 4100
rect 528520 4088 528526 4140
rect 533430 4088 533436 4140
rect 533488 4128 533494 4140
rect 533982 4128 533988 4140
rect 533488 4100 533988 4128
rect 533488 4088 533494 4100
rect 533982 4088 533988 4100
rect 534040 4088 534046 4140
rect 542906 4088 542912 4140
rect 542964 4128 542970 4140
rect 543642 4128 543648 4140
rect 542964 4100 543648 4128
rect 542964 4088 542970 4100
rect 543642 4088 543648 4100
rect 543700 4088 543706 4140
rect 558730 4088 558736 4140
rect 558788 4128 558794 4140
rect 571426 4128 571432 4140
rect 558788 4100 571432 4128
rect 558788 4088 558794 4100
rect 571426 4088 571432 4100
rect 571484 4088 571490 4140
rect 325292 4032 386920 4060
rect 325292 4020 325298 4032
rect 389266 4020 389272 4072
rect 389324 4060 389330 4072
rect 439038 4060 439044 4072
rect 389324 4032 439044 4060
rect 389324 4020 389330 4032
rect 439038 4020 439044 4032
rect 439096 4020 439102 4072
rect 441798 4020 441804 4072
rect 441856 4060 441862 4072
rect 442350 4060 442356 4072
rect 441856 4032 442356 4060
rect 441856 4020 441862 4032
rect 442350 4020 442356 4032
rect 442408 4020 442414 4072
rect 446582 4020 446588 4072
rect 446640 4060 446646 4072
rect 509234 4060 509240 4072
rect 446640 4032 509240 4060
rect 446640 4020 446646 4032
rect 509234 4020 509240 4032
rect 509292 4020 509298 4072
rect 557350 4020 557356 4072
rect 557408 4060 557414 4072
rect 570230 4060 570236 4072
rect 557408 4032 570236 4060
rect 557408 4020 557414 4032
rect 570230 4020 570236 4032
rect 570288 4020 570294 4072
rect 39758 3952 39764 4004
rect 39816 3992 39822 4004
rect 57238 3992 57244 4004
rect 39816 3964 57244 3992
rect 39816 3952 39822 3964
rect 57238 3952 57244 3964
rect 57296 3952 57302 4004
rect 103974 3952 103980 4004
rect 104032 3992 104038 4004
rect 169018 3992 169024 4004
rect 104032 3964 169024 3992
rect 104032 3952 104038 3964
rect 169018 3952 169024 3964
rect 169076 3952 169082 4004
rect 172974 3952 172980 4004
rect 173032 3992 173038 4004
rect 250438 3992 250444 4004
rect 173032 3964 250444 3992
rect 173032 3952 173038 3964
rect 250438 3952 250444 3964
rect 250496 3952 250502 4004
rect 250530 3952 250536 4004
rect 250588 3992 250594 4004
rect 258442 3992 258448 4004
rect 250588 3964 258448 3992
rect 250588 3952 250594 3964
rect 258442 3952 258448 3964
rect 258500 3952 258506 4004
rect 258534 3952 258540 4004
rect 258592 3992 258598 4004
rect 263594 3992 263600 4004
rect 258592 3964 263600 3992
rect 258592 3952 258598 3964
rect 263594 3952 263600 3964
rect 263652 3952 263658 4004
rect 267734 3952 267740 4004
rect 267792 3992 267798 4004
rect 282730 3992 282736 4004
rect 267792 3964 282736 3992
rect 267792 3952 267798 3964
rect 282730 3952 282736 3964
rect 282788 3952 282794 4004
rect 304994 3952 305000 4004
rect 305052 3992 305058 4004
rect 326338 3992 326344 4004
rect 305052 3964 326344 3992
rect 305052 3952 305058 3964
rect 326338 3952 326344 3964
rect 326396 3952 326402 4004
rect 335998 3992 336004 4004
rect 326816 3964 336004 3992
rect 17126 3884 17132 3936
rect 17184 3924 17190 3936
rect 24118 3924 24124 3936
rect 17184 3896 24124 3924
rect 17184 3884 17190 3896
rect 24118 3884 24124 3896
rect 24176 3884 24182 3936
rect 32674 3884 32680 3936
rect 32732 3924 32738 3936
rect 51718 3924 51724 3936
rect 32732 3896 51724 3924
rect 32732 3884 32738 3896
rect 51718 3884 51724 3896
rect 51776 3884 51782 3936
rect 96890 3884 96896 3936
rect 96948 3924 96954 3936
rect 166258 3924 166264 3936
rect 96948 3896 166264 3924
rect 96948 3884 96954 3896
rect 166258 3884 166264 3896
rect 166316 3884 166322 3936
rect 196802 3884 196808 3936
rect 196860 3924 196866 3936
rect 204346 3924 204352 3936
rect 196860 3896 204352 3924
rect 196860 3884 196866 3896
rect 204346 3884 204352 3896
rect 204404 3884 204410 3936
rect 208670 3884 208676 3936
rect 208728 3924 208734 3936
rect 282822 3924 282828 3936
rect 208728 3896 282828 3924
rect 208728 3884 208734 3896
rect 282822 3884 282828 3896
rect 282880 3884 282886 3936
rect 282914 3884 282920 3936
rect 282972 3924 282978 3936
rect 289814 3924 289820 3936
rect 282972 3896 289820 3924
rect 282972 3884 282978 3896
rect 289814 3884 289820 3896
rect 289872 3884 289878 3936
rect 309778 3884 309784 3936
rect 309836 3924 309842 3936
rect 326816 3924 326844 3964
rect 335998 3952 336004 3964
rect 336056 3952 336062 4004
rect 339494 3952 339500 4004
rect 339552 3992 339558 4004
rect 339552 3964 340276 3992
rect 339552 3952 339558 3964
rect 335262 3924 335268 3936
rect 309836 3896 326844 3924
rect 326908 3896 335268 3924
rect 309836 3884 309842 3896
rect 5258 3816 5264 3868
rect 5316 3856 5322 3868
rect 61378 3856 61384 3868
rect 5316 3828 61384 3856
rect 5316 3816 5322 3828
rect 61378 3816 61384 3828
rect 61436 3816 61442 3868
rect 82630 3816 82636 3868
rect 82688 3856 82694 3868
rect 82688 3828 89760 3856
rect 82688 3816 82694 3828
rect 6454 3748 6460 3800
rect 6512 3788 6518 3800
rect 69658 3788 69664 3800
rect 6512 3760 69664 3788
rect 6512 3748 6518 3760
rect 69658 3748 69664 3760
rect 69716 3748 69722 3800
rect 89732 3788 89760 3828
rect 89806 3816 89812 3868
rect 89864 3856 89870 3868
rect 164878 3856 164884 3868
rect 89864 3828 164884 3856
rect 89864 3816 89870 3828
rect 164878 3816 164884 3828
rect 164936 3816 164942 3868
rect 209866 3816 209872 3868
rect 209924 3856 209930 3868
rect 307754 3856 307760 3868
rect 209924 3828 307760 3856
rect 209924 3816 209930 3828
rect 307754 3816 307760 3828
rect 307812 3816 307818 3868
rect 318058 3816 318064 3868
rect 318116 3856 318122 3868
rect 318116 3828 322980 3856
rect 318116 3816 318122 3828
rect 103514 3788 103520 3800
rect 89732 3760 103520 3788
rect 103514 3748 103520 3760
rect 103572 3748 103578 3800
rect 112990 3748 112996 3800
rect 113048 3788 113054 3800
rect 113174 3788 113180 3800
rect 113048 3760 113180 3788
rect 113048 3748 113054 3760
rect 113174 3748 113180 3760
rect 113232 3748 113238 3800
rect 122742 3748 122748 3800
rect 122800 3788 122806 3800
rect 132494 3788 132500 3800
rect 122800 3760 132500 3788
rect 122800 3748 122806 3760
rect 132494 3748 132500 3760
rect 132552 3748 132558 3800
rect 145834 3748 145840 3800
rect 145892 3788 145898 3800
rect 159358 3788 159364 3800
rect 145892 3760 159364 3788
rect 145892 3748 145898 3760
rect 159358 3748 159364 3760
rect 159416 3748 159422 3800
rect 165890 3748 165896 3800
rect 165948 3788 165954 3800
rect 246298 3788 246304 3800
rect 165948 3760 246304 3788
rect 165948 3748 165954 3760
rect 246298 3748 246304 3760
rect 246356 3748 246362 3800
rect 252646 3748 252652 3800
rect 252704 3788 252710 3800
rect 253842 3788 253848 3800
rect 252704 3760 253848 3788
rect 252704 3748 252710 3760
rect 253842 3748 253848 3760
rect 253900 3748 253906 3800
rect 258442 3748 258448 3800
rect 258500 3788 258506 3800
rect 267734 3788 267740 3800
rect 258500 3760 267740 3788
rect 258500 3748 258506 3760
rect 267734 3748 267740 3760
rect 267792 3748 267798 3800
rect 307662 3748 307668 3800
rect 307720 3788 307726 3800
rect 313918 3788 313924 3800
rect 307720 3760 313924 3788
rect 307720 3748 307726 3760
rect 313918 3748 313924 3760
rect 313976 3748 313982 3800
rect 46934 3680 46940 3732
rect 46992 3720 46998 3732
rect 145926 3720 145932 3732
rect 46992 3692 145932 3720
rect 46992 3680 46998 3692
rect 145926 3680 145932 3692
rect 145984 3680 145990 3732
rect 149238 3680 149244 3732
rect 149296 3720 149302 3732
rect 150342 3720 150348 3732
rect 149296 3692 150348 3720
rect 149296 3680 149302 3692
rect 150342 3680 150348 3692
rect 150400 3680 150406 3732
rect 153930 3680 153936 3732
rect 153988 3720 153994 3732
rect 154482 3720 154488 3732
rect 153988 3692 154488 3720
rect 153988 3680 153994 3692
rect 154482 3680 154488 3692
rect 154540 3680 154546 3732
rect 174170 3680 174176 3732
rect 174228 3720 174234 3732
rect 273162 3720 273168 3732
rect 174228 3692 273168 3720
rect 174228 3680 174234 3692
rect 273162 3680 273168 3692
rect 273220 3680 273226 3732
rect 321646 3680 321652 3732
rect 321704 3720 321710 3732
rect 322842 3720 322848 3732
rect 321704 3692 322848 3720
rect 321704 3680 321710 3692
rect 322842 3680 322848 3692
rect 322900 3680 322906 3732
rect 322952 3720 322980 3828
rect 323026 3816 323032 3868
rect 323084 3856 323090 3868
rect 326908 3856 326936 3896
rect 335262 3884 335268 3896
rect 335320 3884 335326 3936
rect 337746 3884 337752 3936
rect 337804 3924 337810 3936
rect 340138 3924 340144 3936
rect 337804 3896 340144 3924
rect 337804 3884 337810 3896
rect 340138 3884 340144 3896
rect 340196 3884 340202 3936
rect 340248 3924 340276 3964
rect 340322 3952 340328 4004
rect 340380 3992 340386 4004
rect 345658 3992 345664 4004
rect 340380 3964 345664 3992
rect 340380 3952 340386 3964
rect 345658 3952 345664 3964
rect 345716 3952 345722 4004
rect 346670 3952 346676 4004
rect 346728 3992 346734 4004
rect 364334 3992 364340 4004
rect 346728 3964 364340 3992
rect 346728 3952 346734 3964
rect 364334 3952 364340 3964
rect 364392 3952 364398 4004
rect 370406 3952 370412 4004
rect 370464 3992 370470 4004
rect 371142 3992 371148 4004
rect 370464 3964 371148 3992
rect 370464 3952 370470 3964
rect 371142 3952 371148 3964
rect 371200 3952 371206 4004
rect 373994 3952 374000 4004
rect 374052 3992 374058 4004
rect 375190 3992 375196 4004
rect 374052 3964 375196 3992
rect 374052 3952 374058 3964
rect 375190 3952 375196 3964
rect 375248 3952 375254 4004
rect 377582 3952 377588 4004
rect 377640 3992 377646 4004
rect 378042 3992 378048 4004
rect 377640 3964 378048 3992
rect 377640 3952 377646 3964
rect 378042 3952 378048 3964
rect 378100 3952 378106 4004
rect 378226 3952 378232 4004
rect 378284 3992 378290 4004
rect 384298 3992 384304 4004
rect 378284 3964 384304 3992
rect 378284 3952 378290 3964
rect 384298 3952 384304 3964
rect 384356 3952 384362 4004
rect 393958 3952 393964 4004
rect 394016 3992 394022 4004
rect 403618 3992 403624 4004
rect 394016 3964 403624 3992
rect 394016 3952 394022 3964
rect 403618 3952 403624 3964
rect 403676 3952 403682 4004
rect 404906 3952 404912 4004
rect 404964 3992 404970 4004
rect 405642 3992 405648 4004
rect 404964 3964 405648 3992
rect 404964 3952 404970 3964
rect 405642 3952 405648 3964
rect 405700 3952 405706 4004
rect 406102 3952 406108 4004
rect 406160 3992 406166 4004
rect 407022 3992 407028 4004
rect 406160 3964 407028 3992
rect 406160 3952 406166 3964
rect 407022 3952 407028 3964
rect 407080 3952 407086 4004
rect 407298 3952 407304 4004
rect 407356 3992 407362 4004
rect 408402 3992 408408 4004
rect 407356 3964 408408 3992
rect 407356 3952 407362 3964
rect 408402 3952 408408 3964
rect 408460 3952 408466 4004
rect 413278 3952 413284 4004
rect 413336 3992 413342 4004
rect 422294 3992 422300 4004
rect 413336 3964 422300 3992
rect 413336 3952 413342 3964
rect 422294 3952 422300 3964
rect 422352 3952 422358 4004
rect 431862 3952 431868 4004
rect 431920 3992 431926 4004
rect 431954 3992 431960 4004
rect 431920 3964 431960 3992
rect 431920 3952 431926 3964
rect 431954 3952 431960 3964
rect 432012 3952 432018 4004
rect 439314 3952 439320 4004
rect 439372 3992 439378 4004
rect 462314 3992 462320 4004
rect 439372 3964 462320 3992
rect 439372 3952 439378 3964
rect 462314 3952 462320 3964
rect 462372 3952 462378 4004
rect 464430 3952 464436 4004
rect 464488 3992 464494 4004
rect 464982 3992 464988 4004
rect 464488 3964 464988 3992
rect 464488 3952 464494 3964
rect 464982 3952 464988 3964
rect 465040 3952 465046 4004
rect 492950 3952 492956 4004
rect 493008 3992 493014 4004
rect 523954 3992 523960 4004
rect 493008 3964 523960 3992
rect 493008 3952 493014 3964
rect 523954 3952 523960 3964
rect 524012 3952 524018 4004
rect 535730 3952 535736 4004
rect 535788 3992 535794 4004
rect 536742 3992 536748 4004
rect 535788 3964 536748 3992
rect 535788 3952 535794 3964
rect 536742 3952 536748 3964
rect 536800 3952 536806 4004
rect 558822 3952 558828 4004
rect 558880 3992 558886 4004
rect 573818 3992 573824 4004
rect 558880 3964 573824 3992
rect 558880 3952 558886 3964
rect 573818 3952 573824 3964
rect 573876 3952 573882 4004
rect 455966 3924 455972 3936
rect 340248 3896 455972 3924
rect 455966 3884 455972 3896
rect 456024 3884 456030 3936
rect 475102 3884 475108 3936
rect 475160 3924 475166 3936
rect 526254 3924 526260 3936
rect 475160 3896 526260 3924
rect 475160 3884 475166 3896
rect 526254 3884 526260 3896
rect 526312 3884 526318 3936
rect 558638 3884 558644 3936
rect 558696 3924 558702 3936
rect 575014 3924 575020 3936
rect 558696 3896 575020 3924
rect 558696 3884 558702 3896
rect 575014 3884 575020 3896
rect 575072 3884 575078 3936
rect 323084 3828 326936 3856
rect 323084 3816 323090 3828
rect 332410 3816 332416 3868
rect 332468 3856 332474 3868
rect 452654 3856 452660 3868
rect 332468 3828 452660 3856
rect 332468 3816 332474 3828
rect 452654 3816 452660 3828
rect 452712 3816 452718 3868
rect 460842 3816 460848 3868
rect 460900 3856 460906 3868
rect 510614 3856 510620 3868
rect 460900 3828 510620 3856
rect 460900 3816 460906 3828
rect 510614 3816 510620 3828
rect 510672 3816 510678 3868
rect 517882 3816 517888 3868
rect 517940 3856 517946 3868
rect 527818 3856 527824 3868
rect 517940 3828 527824 3856
rect 517940 3816 517946 3828
rect 527818 3816 527824 3828
rect 527876 3816 527882 3868
rect 556982 3816 556988 3868
rect 557040 3856 557046 3868
rect 559558 3856 559564 3868
rect 557040 3828 559564 3856
rect 557040 3816 557046 3828
rect 559558 3816 559564 3828
rect 559616 3816 559622 3868
rect 560018 3816 560024 3868
rect 560076 3856 560082 3868
rect 576210 3856 576216 3868
rect 560076 3828 576216 3856
rect 560076 3816 560082 3828
rect 576210 3816 576216 3828
rect 576268 3816 576274 3868
rect 335262 3748 335268 3800
rect 335320 3788 335326 3800
rect 371418 3788 371424 3800
rect 335320 3760 371424 3788
rect 335320 3748 335326 3760
rect 371418 3748 371424 3760
rect 371476 3748 371482 3800
rect 385862 3748 385868 3800
rect 385920 3788 385926 3800
rect 497090 3788 497096 3800
rect 385920 3760 497096 3788
rect 385920 3748 385926 3760
rect 497090 3748 497096 3760
rect 497148 3748 497154 3800
rect 560110 3748 560116 3800
rect 560168 3788 560174 3800
rect 577406 3788 577412 3800
rect 560168 3760 577412 3788
rect 560168 3748 560174 3760
rect 577406 3748 577412 3760
rect 577464 3748 577470 3800
rect 439590 3720 439596 3732
rect 322952 3692 439596 3720
rect 439590 3680 439596 3692
rect 439648 3680 439654 3732
rect 469030 3680 469036 3732
rect 469088 3720 469094 3732
rect 469088 3692 470732 3720
rect 469088 3680 469094 3692
rect 24302 3612 24308 3664
rect 24360 3652 24366 3664
rect 25498 3652 25504 3664
rect 24360 3624 25504 3652
rect 24360 3612 24366 3624
rect 25498 3612 25504 3624
rect 25556 3612 25562 3664
rect 25590 3612 25596 3664
rect 25648 3652 25654 3664
rect 32398 3652 32404 3664
rect 25648 3624 32404 3652
rect 25648 3612 25654 3624
rect 32398 3612 32404 3624
rect 32456 3612 32462 3664
rect 36170 3612 36176 3664
rect 36228 3652 36234 3664
rect 36228 3624 42840 3652
rect 36228 3612 36234 3624
rect 16022 3544 16028 3596
rect 16080 3584 16086 3596
rect 28258 3584 28264 3596
rect 16080 3556 28264 3584
rect 16080 3544 16086 3556
rect 28258 3544 28264 3556
rect 28316 3544 28322 3596
rect 29086 3544 29092 3596
rect 29144 3584 29150 3596
rect 31018 3584 31024 3596
rect 29144 3556 31024 3584
rect 29144 3544 29150 3556
rect 31018 3544 31024 3556
rect 31076 3544 31082 3596
rect 33870 3544 33876 3596
rect 33928 3584 33934 3596
rect 34422 3584 34428 3596
rect 33928 3556 34428 3584
rect 33928 3544 33934 3556
rect 34422 3544 34428 3556
rect 34480 3544 34486 3596
rect 42150 3544 42156 3596
rect 42208 3584 42214 3596
rect 42702 3584 42708 3596
rect 42208 3556 42708 3584
rect 42208 3544 42214 3556
rect 42702 3544 42708 3556
rect 42760 3544 42766 3596
rect 42812 3584 42840 3624
rect 43346 3612 43352 3664
rect 43404 3652 43410 3664
rect 150434 3652 150440 3664
rect 43404 3624 145972 3652
rect 43404 3612 43410 3624
rect 142798 3584 142804 3596
rect 42812 3556 142804 3584
rect 142798 3544 142804 3556
rect 142856 3544 142862 3596
rect 145944 3584 145972 3624
rect 146220 3624 150440 3652
rect 146220 3584 146248 3624
rect 150434 3612 150440 3624
rect 150492 3612 150498 3664
rect 150526 3612 150532 3664
rect 150584 3652 150590 3664
rect 153194 3652 153200 3664
rect 150584 3624 153200 3652
rect 150584 3612 150590 3624
rect 153194 3612 153200 3624
rect 153252 3612 153258 3664
rect 163498 3612 163504 3664
rect 163556 3652 163562 3664
rect 164142 3652 164148 3664
rect 163556 3624 164148 3652
rect 163556 3612 163562 3624
rect 164142 3612 164148 3624
rect 164200 3612 164206 3664
rect 164694 3612 164700 3664
rect 164752 3652 164758 3664
rect 165522 3652 165528 3664
rect 164752 3624 165528 3652
rect 164752 3612 164758 3624
rect 165522 3612 165528 3624
rect 165580 3612 165586 3664
rect 180150 3612 180156 3664
rect 180208 3652 180214 3664
rect 180702 3652 180708 3664
rect 180208 3624 180708 3652
rect 180208 3612 180214 3624
rect 180702 3612 180708 3624
rect 180760 3612 180766 3664
rect 189626 3612 189632 3664
rect 189684 3652 189690 3664
rect 190362 3652 190368 3664
rect 189684 3624 190368 3652
rect 189684 3612 189690 3624
rect 190362 3612 190368 3624
rect 190420 3612 190426 3664
rect 207474 3612 207480 3664
rect 207532 3652 207538 3664
rect 289722 3652 289728 3664
rect 207532 3624 289728 3652
rect 207532 3612 207538 3624
rect 289722 3612 289728 3624
rect 289780 3612 289786 3664
rect 289906 3612 289912 3664
rect 289964 3652 289970 3664
rect 337746 3652 337752 3664
rect 289964 3624 337752 3652
rect 289964 3612 289970 3624
rect 337746 3612 337752 3624
rect 337804 3612 337810 3664
rect 338298 3612 338304 3664
rect 338356 3652 338362 3664
rect 339402 3652 339408 3664
rect 338356 3624 339408 3652
rect 338356 3612 338362 3624
rect 339402 3612 339408 3624
rect 339460 3612 339466 3664
rect 363322 3612 363328 3664
rect 363380 3652 363386 3664
rect 364242 3652 364248 3664
rect 363380 3624 364248 3652
rect 363380 3612 363386 3624
rect 364242 3612 364248 3624
rect 364300 3612 364306 3664
rect 378870 3612 378876 3664
rect 378928 3652 378934 3664
rect 434714 3652 434720 3664
rect 378928 3624 434720 3652
rect 378928 3612 378934 3624
rect 434714 3612 434720 3624
rect 434772 3612 434778 3664
rect 446398 3612 446404 3664
rect 446456 3652 446462 3664
rect 455966 3652 455972 3664
rect 446456 3624 455972 3652
rect 446456 3612 446462 3624
rect 455966 3612 455972 3624
rect 456024 3612 456030 3664
rect 470704 3652 470732 3692
rect 477494 3680 477500 3732
rect 477552 3720 477558 3732
rect 478690 3720 478696 3732
rect 477552 3692 478696 3720
rect 477552 3680 477558 3692
rect 478690 3680 478696 3692
rect 478748 3680 478754 3732
rect 481082 3680 481088 3732
rect 481140 3720 481146 3732
rect 481542 3720 481548 3732
rect 481140 3692 481548 3720
rect 481140 3680 481146 3692
rect 481542 3680 481548 3692
rect 481600 3680 481606 3732
rect 483014 3680 483020 3732
rect 483072 3680 483078 3732
rect 483124 3692 483428 3720
rect 471882 3652 471888 3664
rect 470704 3624 471888 3652
rect 471882 3612 471888 3624
rect 471940 3612 471946 3664
rect 472066 3612 472072 3664
rect 472124 3652 472130 3664
rect 483032 3652 483060 3680
rect 472124 3624 483060 3652
rect 472124 3612 472130 3624
rect 258534 3584 258540 3596
rect 145944 3556 146248 3584
rect 150636 3556 258540 3584
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 10962 3516 10968 3528
rect 10100 3488 10968 3516
rect 10100 3476 10106 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11238 3476 11244 3528
rect 11296 3516 11302 3528
rect 17126 3516 17132 3528
rect 11296 3488 17132 3516
rect 11296 3476 11302 3488
rect 17126 3476 17132 3488
rect 17184 3476 17190 3528
rect 17218 3476 17224 3528
rect 17276 3516 17282 3528
rect 17862 3516 17868 3528
rect 17276 3488 17868 3516
rect 17276 3476 17282 3488
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 25498 3476 25504 3528
rect 25556 3516 25562 3528
rect 25556 3488 132540 3516
rect 25556 3476 25562 3488
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 10502 3448 10508 3460
rect 624 3420 10508 3448
rect 624 3408 630 3420
rect 10502 3408 10508 3420
rect 10560 3408 10566 3460
rect 14826 3408 14832 3460
rect 14884 3448 14890 3460
rect 14884 3420 124168 3448
rect 14884 3408 14890 3420
rect 20714 3340 20720 3392
rect 20772 3380 20778 3392
rect 25590 3380 25596 3392
rect 20772 3352 25596 3380
rect 20772 3340 20778 3352
rect 25590 3340 25596 3352
rect 25648 3340 25654 3392
rect 45738 3340 45744 3392
rect 45796 3380 45802 3392
rect 46842 3380 46848 3392
rect 45796 3352 46848 3380
rect 45796 3340 45802 3352
rect 46842 3340 46848 3352
rect 46900 3340 46906 3392
rect 50522 3340 50528 3392
rect 50580 3380 50586 3392
rect 50982 3380 50988 3392
rect 50580 3352 50988 3380
rect 50580 3340 50586 3352
rect 50982 3340 50988 3352
rect 51040 3340 51046 3392
rect 51626 3340 51632 3392
rect 51684 3380 51690 3392
rect 52362 3380 52368 3392
rect 51684 3352 52368 3380
rect 51684 3340 51690 3352
rect 52362 3340 52368 3352
rect 52420 3340 52426 3392
rect 54018 3340 54024 3392
rect 54076 3380 54082 3392
rect 55122 3380 55128 3392
rect 54076 3352 55128 3380
rect 54076 3340 54082 3352
rect 55122 3340 55128 3352
rect 55180 3340 55186 3392
rect 55214 3340 55220 3392
rect 55272 3380 55278 3392
rect 56502 3380 56508 3392
rect 55272 3352 56508 3380
rect 55272 3340 55278 3352
rect 56502 3340 56508 3352
rect 56560 3340 56566 3392
rect 58802 3340 58808 3392
rect 58860 3380 58866 3392
rect 59262 3380 59268 3392
rect 58860 3352 59268 3380
rect 58860 3340 58866 3352
rect 59262 3340 59268 3352
rect 59320 3340 59326 3392
rect 61194 3340 61200 3392
rect 61252 3380 61258 3392
rect 62022 3380 62028 3392
rect 61252 3352 62028 3380
rect 61252 3340 61258 3352
rect 62022 3340 62028 3352
rect 62080 3340 62086 3392
rect 62390 3340 62396 3392
rect 62448 3380 62454 3392
rect 63402 3380 63408 3392
rect 62448 3352 63408 3380
rect 62448 3340 62454 3352
rect 63402 3340 63408 3352
rect 63460 3340 63466 3392
rect 68278 3340 68284 3392
rect 68336 3380 68342 3392
rect 68922 3380 68928 3392
rect 68336 3352 68928 3380
rect 68336 3340 68342 3352
rect 68922 3340 68928 3352
rect 68980 3340 68986 3392
rect 71866 3340 71872 3392
rect 71924 3380 71930 3392
rect 72970 3380 72976 3392
rect 71924 3352 72976 3380
rect 71924 3340 71930 3352
rect 72970 3340 72976 3352
rect 73028 3340 73034 3392
rect 79042 3340 79048 3392
rect 79100 3380 79106 3392
rect 79962 3380 79968 3392
rect 79100 3352 79968 3380
rect 79100 3340 79106 3352
rect 79962 3340 79968 3352
rect 80020 3340 80026 3392
rect 106366 3340 106372 3392
rect 106424 3380 106430 3392
rect 107470 3380 107476 3392
rect 106424 3352 107476 3380
rect 106424 3340 106430 3352
rect 107470 3340 107476 3352
rect 107528 3340 107534 3392
rect 112346 3340 112352 3392
rect 112404 3380 112410 3392
rect 113082 3380 113088 3392
rect 112404 3352 113088 3380
rect 112404 3340 112410 3352
rect 113082 3340 113088 3352
rect 113140 3340 113146 3392
rect 114738 3340 114744 3392
rect 114796 3380 114802 3392
rect 115842 3380 115848 3392
rect 114796 3352 115848 3380
rect 114796 3340 114802 3352
rect 115842 3340 115848 3352
rect 115900 3340 115906 3392
rect 119430 3340 119436 3392
rect 119488 3380 119494 3392
rect 119982 3380 119988 3392
rect 119488 3352 119988 3380
rect 119488 3340 119494 3352
rect 119982 3340 119988 3352
rect 120040 3340 120046 3392
rect 113174 3272 113180 3324
rect 113232 3312 113238 3324
rect 122742 3312 122748 3324
rect 113232 3284 122748 3312
rect 113232 3272 113238 3284
rect 122742 3272 122748 3284
rect 122800 3272 122806 3324
rect 124140 3312 124168 3420
rect 124214 3408 124220 3460
rect 124272 3448 124278 3460
rect 125502 3448 125508 3460
rect 124272 3420 125508 3448
rect 124272 3408 124278 3420
rect 125502 3408 125508 3420
rect 125560 3408 125566 3460
rect 128998 3408 129004 3460
rect 129056 3448 129062 3460
rect 129642 3448 129648 3460
rect 129056 3420 129648 3448
rect 129056 3408 129062 3420
rect 129642 3408 129648 3420
rect 129700 3408 129706 3460
rect 130194 3408 130200 3460
rect 130252 3448 130258 3460
rect 131022 3448 131028 3460
rect 130252 3420 131028 3448
rect 130252 3408 130258 3420
rect 131022 3408 131028 3420
rect 131080 3408 131086 3460
rect 131390 3408 131396 3460
rect 131448 3448 131454 3460
rect 132402 3448 132408 3460
rect 131448 3420 132408 3448
rect 131448 3408 131454 3420
rect 132402 3408 132408 3420
rect 132460 3408 132466 3460
rect 125410 3340 125416 3392
rect 125468 3380 125474 3392
rect 126238 3380 126244 3392
rect 125468 3352 126244 3380
rect 125468 3340 125474 3352
rect 126238 3340 126244 3352
rect 126296 3340 126302 3392
rect 132512 3380 132540 3488
rect 132586 3476 132592 3528
rect 132644 3516 132650 3528
rect 133782 3516 133788 3528
rect 132644 3488 133788 3516
rect 132644 3476 132650 3488
rect 133782 3476 133788 3488
rect 133840 3476 133846 3528
rect 136082 3476 136088 3528
rect 136140 3516 136146 3528
rect 136542 3516 136548 3528
rect 136140 3488 136548 3516
rect 136140 3476 136146 3488
rect 136542 3476 136548 3488
rect 136600 3476 136606 3528
rect 139670 3476 139676 3528
rect 139728 3516 139734 3528
rect 140682 3516 140688 3528
rect 139728 3488 140688 3516
rect 139728 3476 139734 3488
rect 140682 3476 140688 3488
rect 140740 3476 140746 3528
rect 150526 3516 150532 3528
rect 147968 3488 150532 3516
rect 145834 3448 145840 3460
rect 138308 3420 145840 3448
rect 138198 3380 138204 3392
rect 132512 3352 138204 3380
rect 138198 3340 138204 3352
rect 138256 3340 138262 3392
rect 129826 3312 129832 3324
rect 124140 3284 129832 3312
rect 129826 3272 129832 3284
rect 129884 3272 129890 3324
rect 132494 3272 132500 3324
rect 132552 3312 132558 3324
rect 138308 3312 138336 3420
rect 145834 3408 145840 3420
rect 145892 3408 145898 3460
rect 146110 3408 146116 3460
rect 146168 3448 146174 3460
rect 147968 3448 147996 3488
rect 150526 3476 150532 3488
rect 150584 3476 150590 3528
rect 146168 3420 147996 3448
rect 146168 3408 146174 3420
rect 148042 3408 148048 3460
rect 148100 3448 148106 3460
rect 150636 3448 150664 3556
rect 258534 3544 258540 3556
rect 258592 3544 258598 3596
rect 258626 3544 258632 3596
rect 258684 3584 258690 3596
rect 259362 3584 259368 3596
rect 258684 3556 259368 3584
rect 258684 3544 258690 3556
rect 259362 3544 259368 3556
rect 259420 3544 259426 3596
rect 266998 3544 267004 3596
rect 267056 3584 267062 3596
rect 267642 3584 267648 3596
rect 267056 3556 267648 3584
rect 267056 3544 267062 3556
rect 267642 3544 267648 3556
rect 267700 3544 267706 3596
rect 268102 3544 268108 3596
rect 268160 3584 268166 3596
rect 269022 3584 269028 3596
rect 268160 3556 269028 3584
rect 268160 3544 268166 3556
rect 269022 3544 269028 3556
rect 269080 3544 269086 3596
rect 282730 3544 282736 3596
rect 282788 3584 282794 3596
rect 289630 3584 289636 3596
rect 282788 3556 289636 3584
rect 282788 3544 282794 3556
rect 289630 3544 289636 3556
rect 289688 3544 289694 3596
rect 298094 3544 298100 3596
rect 298152 3584 298158 3596
rect 307662 3584 307668 3596
rect 298152 3556 307668 3584
rect 298152 3544 298158 3556
rect 307662 3544 307668 3556
rect 307720 3544 307726 3596
rect 316586 3544 316592 3596
rect 316644 3584 316650 3596
rect 445754 3584 445760 3596
rect 316644 3556 445760 3584
rect 316644 3544 316650 3556
rect 445754 3544 445760 3556
rect 445812 3544 445818 3596
rect 461578 3544 461584 3596
rect 461636 3584 461642 3596
rect 483124 3584 483152 3692
rect 483400 3652 483428 3692
rect 483474 3680 483480 3732
rect 483532 3720 483538 3732
rect 484302 3720 484308 3732
rect 483532 3692 484308 3720
rect 483532 3680 483538 3692
rect 484302 3680 484308 3692
rect 484360 3680 484366 3732
rect 484394 3680 484400 3732
rect 484452 3720 484458 3732
rect 527910 3720 527916 3732
rect 484452 3692 492628 3720
rect 484452 3680 484458 3692
rect 492600 3652 492628 3692
rect 519556 3692 527916 3720
rect 495526 3652 495532 3664
rect 483400 3624 483612 3652
rect 492600 3624 495532 3652
rect 461636 3556 483152 3584
rect 483584 3584 483612 3624
rect 495526 3612 495532 3624
rect 495584 3612 495590 3664
rect 500236 3624 505416 3652
rect 500236 3584 500264 3624
rect 483584 3556 500264 3584
rect 461636 3544 461642 3556
rect 500310 3544 500316 3596
rect 500368 3584 500374 3596
rect 505278 3584 505284 3596
rect 500368 3556 505284 3584
rect 500368 3544 500374 3556
rect 505278 3544 505284 3556
rect 505336 3544 505342 3596
rect 505388 3584 505416 3624
rect 505388 3556 512040 3584
rect 150710 3476 150716 3528
rect 150768 3516 150774 3528
rect 384850 3516 384856 3528
rect 150768 3488 384856 3516
rect 150768 3476 150774 3488
rect 384850 3476 384856 3488
rect 384908 3476 384914 3528
rect 393038 3476 393044 3528
rect 393096 3516 393102 3528
rect 397454 3516 397460 3528
rect 393096 3488 397460 3516
rect 393096 3476 393102 3488
rect 397454 3476 397460 3488
rect 397512 3476 397518 3528
rect 397822 3476 397828 3528
rect 397880 3516 397886 3528
rect 398742 3516 398748 3528
rect 397880 3488 398748 3516
rect 397880 3476 397886 3488
rect 398742 3476 398748 3488
rect 398800 3476 398806 3528
rect 410886 3476 410892 3528
rect 410944 3516 410950 3528
rect 483198 3516 483204 3528
rect 410944 3488 483204 3516
rect 410944 3476 410950 3488
rect 483198 3476 483204 3488
rect 483256 3476 483262 3528
rect 483382 3476 483388 3528
rect 483440 3516 483446 3528
rect 483440 3488 495480 3516
rect 483440 3476 483446 3488
rect 148100 3420 150664 3448
rect 148100 3408 148106 3420
rect 155126 3408 155132 3460
rect 155184 3448 155190 3460
rect 411162 3448 411168 3460
rect 155184 3420 411168 3448
rect 155184 3408 155190 3420
rect 411162 3408 411168 3420
rect 411220 3408 411226 3460
rect 415670 3408 415676 3460
rect 415728 3448 415734 3460
rect 416682 3448 416688 3460
rect 415728 3420 416688 3448
rect 415728 3408 415734 3420
rect 416682 3408 416688 3420
rect 416740 3408 416746 3460
rect 423950 3408 423956 3460
rect 424008 3448 424014 3460
rect 424962 3448 424968 3460
rect 424008 3420 424968 3448
rect 424008 3408 424014 3420
rect 424962 3408 424968 3420
rect 425020 3408 425026 3460
rect 428734 3408 428740 3460
rect 428792 3448 428798 3460
rect 439498 3448 439504 3460
rect 428792 3420 439504 3448
rect 428792 3408 428798 3420
rect 439498 3408 439504 3420
rect 439556 3408 439562 3460
rect 439682 3408 439688 3460
rect 439740 3448 439746 3460
rect 439740 3420 444144 3448
rect 439740 3408 439746 3420
rect 140866 3340 140872 3392
rect 140924 3380 140930 3392
rect 191742 3380 191748 3392
rect 140924 3352 151860 3380
rect 140924 3340 140930 3352
rect 132552 3284 138336 3312
rect 132552 3272 132558 3284
rect 146846 3272 146852 3324
rect 146904 3312 146910 3324
rect 147582 3312 147588 3324
rect 146904 3284 147588 3312
rect 146904 3272 146910 3284
rect 147582 3272 147588 3284
rect 147640 3272 147646 3324
rect 150434 3272 150440 3324
rect 150492 3312 150498 3324
rect 151722 3312 151728 3324
rect 150492 3284 151728 3312
rect 150492 3272 150498 3284
rect 151722 3272 151728 3284
rect 151780 3272 151786 3324
rect 151832 3312 151860 3352
rect 152844 3352 191748 3380
rect 152844 3312 152872 3352
rect 191742 3340 191748 3352
rect 191800 3340 191806 3392
rect 192018 3340 192024 3392
rect 192076 3380 192082 3392
rect 193122 3380 193128 3392
rect 192076 3352 193128 3380
rect 192076 3340 192082 3352
rect 193122 3340 193128 3352
rect 193180 3340 193186 3392
rect 217042 3340 217048 3392
rect 217100 3380 217106 3392
rect 217962 3380 217968 3392
rect 217100 3352 217968 3380
rect 217100 3340 217106 3352
rect 217962 3340 217968 3352
rect 218020 3340 218026 3392
rect 224126 3340 224132 3392
rect 224184 3380 224190 3392
rect 224862 3380 224868 3392
rect 224184 3352 224868 3380
rect 224184 3340 224190 3352
rect 224862 3340 224868 3352
rect 224920 3340 224926 3392
rect 225322 3340 225328 3392
rect 225380 3380 225386 3392
rect 226242 3380 226248 3392
rect 225380 3352 226248 3380
rect 225380 3340 225386 3352
rect 226242 3340 226248 3352
rect 226300 3340 226306 3392
rect 227714 3340 227720 3392
rect 227772 3380 227778 3392
rect 229002 3380 229008 3392
rect 227772 3352 229008 3380
rect 227772 3340 227778 3352
rect 229002 3340 229008 3352
rect 229060 3340 229066 3392
rect 231302 3340 231308 3392
rect 231360 3380 231366 3392
rect 231762 3380 231768 3392
rect 231360 3352 231768 3380
rect 231360 3340 231366 3352
rect 231762 3340 231768 3352
rect 231820 3340 231826 3392
rect 233694 3340 233700 3392
rect 233752 3380 233758 3392
rect 234522 3380 234528 3392
rect 233752 3352 234528 3380
rect 233752 3340 233758 3352
rect 234522 3340 234528 3352
rect 234580 3340 234586 3392
rect 234798 3340 234804 3392
rect 234856 3380 234862 3392
rect 235902 3380 235908 3392
rect 234856 3352 235908 3380
rect 234856 3340 234862 3352
rect 235902 3340 235908 3352
rect 235960 3340 235966 3392
rect 239582 3340 239588 3392
rect 239640 3380 239646 3392
rect 240042 3380 240048 3392
rect 239640 3352 240048 3380
rect 239640 3340 239646 3352
rect 240042 3340 240048 3352
rect 240100 3340 240106 3392
rect 241974 3340 241980 3392
rect 242032 3380 242038 3392
rect 242802 3380 242808 3392
rect 242032 3352 242808 3380
rect 242032 3340 242038 3352
rect 242802 3340 242808 3352
rect 242860 3340 242866 3392
rect 243170 3340 243176 3392
rect 243228 3380 243234 3392
rect 244182 3380 244188 3392
rect 243228 3352 244188 3380
rect 243228 3340 243234 3352
rect 244182 3340 244188 3352
rect 244240 3340 244246 3392
rect 249150 3340 249156 3392
rect 249208 3380 249214 3392
rect 249702 3380 249708 3392
rect 249208 3352 249708 3380
rect 249208 3340 249214 3352
rect 249702 3340 249708 3352
rect 249760 3340 249766 3392
rect 264606 3340 264612 3392
rect 264664 3380 264670 3392
rect 378134 3380 378140 3392
rect 264664 3352 378140 3380
rect 264664 3340 264670 3352
rect 378134 3340 378140 3352
rect 378192 3340 378198 3392
rect 384298 3340 384304 3392
rect 384356 3380 384362 3392
rect 393958 3380 393964 3392
rect 384356 3352 393964 3380
rect 384356 3340 384362 3352
rect 393958 3340 393964 3352
rect 394016 3340 394022 3392
rect 402514 3340 402520 3392
rect 402572 3380 402578 3392
rect 418798 3380 418804 3392
rect 402572 3352 418804 3380
rect 402572 3340 402578 3352
rect 418798 3340 418804 3352
rect 418856 3340 418862 3392
rect 425146 3340 425152 3392
rect 425204 3380 425210 3392
rect 444006 3380 444012 3392
rect 425204 3352 444012 3380
rect 425204 3340 425210 3352
rect 444006 3340 444012 3352
rect 444064 3340 444070 3392
rect 151832 3284 152872 3312
rect 257430 3272 257436 3324
rect 257488 3312 257494 3324
rect 364978 3312 364984 3324
rect 257488 3284 364984 3312
rect 257488 3272 257494 3284
rect 364978 3272 364984 3284
rect 365036 3272 365042 3324
rect 371602 3272 371608 3324
rect 371660 3312 371666 3324
rect 439682 3312 439688 3324
rect 371660 3284 439688 3312
rect 371660 3272 371666 3284
rect 439682 3272 439688 3284
rect 439740 3272 439746 3324
rect 444116 3312 444144 3420
rect 444282 3408 444288 3460
rect 444340 3448 444346 3460
rect 483014 3448 483020 3460
rect 444340 3420 483020 3448
rect 444340 3408 444346 3420
rect 483014 3408 483020 3420
rect 483072 3408 483078 3460
rect 483566 3408 483572 3460
rect 483624 3448 483630 3460
rect 483624 3420 494100 3448
rect 483624 3408 483630 3420
rect 444190 3340 444196 3392
rect 444248 3380 444254 3392
rect 493870 3380 493876 3392
rect 444248 3352 493876 3380
rect 444248 3340 444254 3352
rect 493870 3340 493876 3352
rect 493928 3340 493934 3392
rect 494072 3380 494100 3420
rect 494146 3408 494152 3460
rect 494204 3448 494210 3460
rect 495342 3448 495348 3460
rect 494204 3420 495348 3448
rect 494204 3408 494210 3420
rect 495342 3408 495348 3420
rect 495400 3408 495406 3460
rect 495452 3448 495480 3488
rect 507210 3476 507216 3528
rect 507268 3516 507274 3528
rect 507762 3516 507768 3528
rect 507268 3488 507768 3516
rect 507268 3476 507274 3488
rect 507762 3476 507768 3488
rect 507820 3476 507826 3528
rect 510798 3476 510804 3528
rect 510856 3516 510862 3528
rect 511902 3516 511908 3528
rect 510856 3488 511908 3516
rect 510856 3476 510862 3488
rect 511902 3476 511908 3488
rect 511960 3476 511966 3528
rect 512012 3516 512040 3556
rect 514386 3544 514392 3596
rect 514444 3584 514450 3596
rect 519556 3584 519584 3692
rect 527910 3680 527916 3692
rect 527968 3680 527974 3732
rect 560202 3680 560208 3732
rect 560260 3720 560266 3732
rect 578602 3720 578608 3732
rect 560260 3692 578608 3720
rect 560260 3680 560266 3692
rect 578602 3680 578608 3692
rect 578660 3680 578666 3732
rect 521470 3612 521476 3664
rect 521528 3652 521534 3664
rect 530578 3652 530584 3664
rect 521528 3624 530584 3652
rect 521528 3612 521534 3624
rect 530578 3612 530584 3624
rect 530636 3612 530642 3664
rect 561582 3612 561588 3664
rect 561640 3652 561646 3664
rect 580994 3652 581000 3664
rect 561640 3624 581000 3652
rect 561640 3612 561646 3624
rect 580994 3612 581000 3624
rect 581052 3612 581058 3664
rect 514444 3556 519584 3584
rect 514444 3544 514450 3556
rect 523862 3544 523868 3596
rect 523920 3584 523926 3596
rect 526438 3584 526444 3596
rect 523920 3556 526444 3584
rect 523920 3544 523926 3556
rect 526438 3544 526444 3556
rect 526496 3544 526502 3596
rect 536926 3544 536932 3596
rect 536984 3584 536990 3596
rect 544378 3584 544384 3596
rect 536984 3556 544384 3584
rect 536984 3544 536990 3556
rect 544378 3544 544384 3556
rect 544436 3544 544442 3596
rect 554866 3544 554872 3596
rect 554924 3584 554930 3596
rect 555970 3584 555976 3596
rect 554924 3556 555976 3584
rect 554924 3544 554930 3556
rect 555970 3544 555976 3556
rect 556028 3544 556034 3596
rect 556890 3544 556896 3596
rect 556948 3584 556954 3596
rect 561950 3584 561956 3596
rect 556948 3556 561956 3584
rect 556948 3544 556954 3556
rect 561950 3544 561956 3556
rect 562008 3544 562014 3596
rect 563698 3544 563704 3596
rect 563756 3584 563762 3596
rect 583386 3584 583392 3596
rect 563756 3556 583392 3584
rect 563756 3544 563762 3556
rect 583386 3544 583392 3556
rect 583444 3544 583450 3596
rect 514662 3516 514668 3528
rect 512012 3488 514668 3516
rect 514662 3476 514668 3488
rect 514720 3476 514726 3528
rect 534534 3476 534540 3528
rect 534592 3516 534598 3528
rect 535362 3516 535368 3528
rect 534592 3488 535368 3516
rect 534592 3476 534598 3488
rect 535362 3476 535368 3488
rect 535420 3476 535426 3528
rect 544102 3476 544108 3528
rect 544160 3516 544166 3528
rect 545022 3516 545028 3528
rect 544160 3488 545028 3516
rect 544160 3476 544166 3488
rect 545022 3476 545028 3488
rect 545080 3476 545086 3528
rect 545298 3476 545304 3528
rect 545356 3516 545362 3528
rect 546310 3516 546316 3528
rect 545356 3488 546316 3516
rect 545356 3476 545362 3488
rect 546310 3476 546316 3488
rect 546368 3476 546374 3528
rect 550082 3476 550088 3528
rect 550140 3516 550146 3528
rect 550542 3516 550548 3528
rect 550140 3488 550548 3516
rect 550140 3476 550146 3488
rect 550542 3476 550548 3488
rect 550600 3476 550606 3528
rect 551830 3476 551836 3528
rect 551888 3516 551894 3528
rect 552382 3516 552388 3528
rect 551888 3488 552388 3516
rect 551888 3476 551894 3488
rect 552382 3476 552388 3488
rect 552440 3476 552446 3528
rect 555510 3476 555516 3528
rect 555568 3516 555574 3528
rect 557166 3516 557172 3528
rect 555568 3488 557172 3516
rect 555568 3476 555574 3488
rect 557166 3476 557172 3488
rect 557224 3476 557230 3528
rect 560754 3516 560760 3528
rect 557276 3488 560760 3516
rect 495452 3420 499252 3448
rect 499114 3380 499120 3392
rect 494072 3352 499120 3380
rect 499114 3340 499120 3352
rect 499172 3340 499178 3392
rect 499224 3380 499252 3420
rect 500126 3408 500132 3460
rect 500184 3448 500190 3460
rect 524966 3448 524972 3460
rect 500184 3420 524972 3448
rect 500184 3408 500190 3420
rect 524966 3408 524972 3420
rect 525024 3408 525030 3460
rect 526254 3408 526260 3460
rect 526312 3448 526318 3460
rect 535270 3448 535276 3460
rect 526312 3420 535276 3448
rect 526312 3408 526318 3420
rect 535270 3408 535276 3420
rect 535328 3408 535334 3460
rect 539318 3408 539324 3460
rect 539376 3448 539382 3460
rect 545758 3448 545764 3460
rect 539376 3420 545764 3448
rect 539376 3408 539382 3420
rect 545758 3408 545764 3420
rect 545816 3408 545822 3460
rect 556798 3408 556804 3460
rect 556856 3448 556862 3460
rect 557276 3448 557304 3488
rect 560754 3476 560760 3488
rect 560812 3476 560818 3528
rect 563054 3476 563060 3528
rect 563112 3516 563118 3528
rect 564342 3516 564348 3528
rect 563112 3488 564348 3516
rect 563112 3476 563118 3488
rect 564342 3476 564348 3488
rect 564400 3476 564406 3528
rect 582190 3516 582196 3528
rect 564452 3488 582196 3516
rect 556856 3420 557304 3448
rect 556856 3408 556862 3420
rect 561490 3408 561496 3460
rect 561548 3448 561554 3460
rect 564452 3448 564480 3488
rect 582190 3476 582196 3488
rect 582248 3476 582254 3528
rect 561548 3420 564480 3448
rect 561548 3408 561554 3420
rect 564526 3408 564532 3460
rect 564584 3448 564590 3460
rect 579798 3448 579804 3460
rect 564584 3420 579804 3448
rect 564584 3408 564590 3420
rect 579798 3408 579804 3420
rect 579856 3408 579862 3460
rect 500310 3380 500316 3392
rect 499224 3352 500316 3380
rect 500310 3340 500316 3352
rect 500368 3340 500374 3392
rect 546494 3340 546500 3392
rect 546552 3380 546558 3392
rect 547782 3380 547788 3392
rect 546552 3352 547788 3380
rect 546552 3340 546558 3352
rect 547782 3340 547788 3352
rect 547840 3340 547846 3392
rect 556062 3340 556068 3392
rect 556120 3380 556126 3392
rect 566734 3380 566740 3392
rect 556120 3352 566740 3380
rect 556120 3340 556126 3352
rect 566734 3340 566740 3352
rect 566792 3340 566798 3392
rect 454126 3312 454132 3324
rect 444116 3284 454132 3312
rect 454126 3272 454132 3284
rect 454184 3272 454190 3324
rect 467926 3272 467932 3324
rect 467984 3312 467990 3324
rect 523770 3312 523776 3324
rect 467984 3284 523776 3312
rect 467984 3272 467990 3284
rect 523770 3272 523776 3284
rect 523828 3272 523834 3324
rect 532234 3272 532240 3324
rect 532292 3312 532298 3324
rect 536098 3312 536104 3324
rect 532292 3284 536104 3312
rect 532292 3272 532298 3284
rect 536098 3272 536104 3284
rect 536156 3272 536162 3324
rect 557258 3272 557264 3324
rect 557316 3312 557322 3324
rect 567838 3312 567844 3324
rect 557316 3284 567844 3312
rect 557316 3272 557322 3284
rect 567838 3272 567844 3284
rect 567896 3272 567902 3324
rect 7650 3204 7656 3256
rect 7708 3244 7714 3256
rect 11698 3244 11704 3256
rect 7708 3216 11704 3244
rect 7708 3204 7714 3216
rect 11698 3204 11704 3216
rect 11756 3204 11762 3256
rect 144454 3204 144460 3256
rect 144512 3244 144518 3256
rect 150710 3244 150716 3256
rect 144512 3216 150716 3244
rect 144512 3204 144518 3216
rect 150710 3204 150716 3216
rect 150768 3204 150774 3256
rect 205082 3204 205088 3256
rect 205140 3244 205146 3256
rect 282178 3244 282184 3256
rect 205140 3216 282184 3244
rect 205140 3204 205146 3216
rect 282178 3204 282184 3216
rect 282236 3204 282242 3256
rect 289630 3204 289636 3256
rect 289688 3244 289694 3256
rect 298002 3244 298008 3256
rect 289688 3216 298008 3244
rect 289688 3204 289694 3216
rect 298002 3204 298008 3216
rect 298060 3204 298066 3256
rect 310974 3204 310980 3256
rect 311032 3244 311038 3256
rect 316586 3244 316592 3256
rect 311032 3216 316592 3244
rect 311032 3204 311038 3216
rect 316586 3204 316592 3216
rect 316644 3204 316650 3256
rect 328822 3204 328828 3256
rect 328880 3244 328886 3256
rect 329742 3244 329748 3256
rect 328880 3216 329748 3244
rect 328880 3204 328886 3216
rect 329742 3204 329748 3216
rect 329800 3204 329806 3256
rect 330018 3204 330024 3256
rect 330076 3244 330082 3256
rect 333238 3244 333244 3256
rect 330076 3216 333244 3244
rect 330076 3204 330082 3216
rect 333238 3204 333244 3216
rect 333296 3204 333302 3256
rect 335906 3204 335912 3256
rect 335964 3244 335970 3256
rect 340322 3244 340328 3256
rect 335964 3216 340328 3244
rect 335964 3204 335970 3216
rect 340322 3204 340328 3216
rect 340380 3204 340386 3256
rect 364518 3204 364524 3256
rect 364576 3244 364582 3256
rect 364576 3216 432276 3244
rect 364576 3204 364582 3216
rect 19518 3136 19524 3188
rect 19576 3176 19582 3188
rect 22738 3176 22744 3188
rect 19576 3148 22744 3176
rect 19576 3136 19582 3148
rect 22738 3136 22744 3148
rect 22796 3136 22802 3188
rect 27890 3136 27896 3188
rect 27948 3176 27954 3188
rect 28902 3176 28908 3188
rect 27948 3148 28908 3176
rect 27948 3136 27954 3148
rect 28902 3136 28908 3148
rect 28960 3136 28966 3188
rect 157518 3136 157524 3188
rect 157576 3176 157582 3188
rect 158622 3176 158628 3188
rect 157576 3148 158628 3176
rect 157576 3136 157582 3148
rect 158622 3136 158628 3148
rect 158680 3136 158686 3188
rect 240778 3136 240784 3188
rect 240836 3176 240842 3188
rect 311158 3176 311164 3188
rect 240836 3148 311164 3176
rect 240836 3136 240842 3148
rect 311158 3136 311164 3148
rect 311216 3136 311222 3188
rect 360930 3136 360936 3188
rect 360988 3176 360994 3188
rect 421466 3176 421472 3188
rect 360988 3148 421472 3176
rect 360988 3136 360994 3148
rect 421466 3136 421472 3148
rect 421524 3136 421530 3188
rect 422294 3136 422300 3188
rect 422352 3176 422358 3188
rect 431862 3176 431868 3188
rect 422352 3148 431868 3176
rect 422352 3136 422358 3148
rect 431862 3136 431868 3148
rect 431920 3136 431926 3188
rect 432248 3176 432276 3216
rect 432322 3204 432328 3256
rect 432380 3244 432386 3256
rect 433242 3244 433248 3256
rect 432380 3216 433248 3244
rect 432380 3204 432386 3216
rect 433242 3204 433248 3216
rect 433300 3204 433306 3256
rect 439774 3244 439780 3256
rect 433352 3216 439780 3244
rect 433352 3176 433380 3216
rect 439774 3204 439780 3216
rect 439832 3204 439838 3256
rect 444190 3204 444196 3256
rect 444248 3244 444254 3256
rect 504358 3244 504364 3256
rect 444248 3216 504364 3244
rect 444248 3204 444254 3216
rect 504358 3204 504364 3216
rect 504416 3204 504422 3256
rect 540514 3204 540520 3256
rect 540572 3244 540578 3256
rect 546586 3244 546592 3256
rect 540572 3216 546592 3244
rect 540572 3204 540578 3216
rect 546586 3204 546592 3216
rect 546644 3204 546650 3256
rect 432248 3148 433380 3176
rect 435818 3136 435824 3188
rect 435876 3176 435882 3188
rect 500218 3176 500224 3188
rect 435876 3148 500224 3176
rect 435876 3136 435882 3148
rect 500218 3136 500224 3148
rect 500276 3136 500282 3188
rect 528646 3136 528652 3188
rect 528704 3176 528710 3188
rect 531958 3176 531964 3188
rect 528704 3148 531964 3176
rect 528704 3136 528710 3148
rect 531958 3136 531964 3148
rect 532016 3136 532022 3188
rect 559926 3136 559932 3188
rect 559984 3176 559990 3188
rect 564526 3176 564532 3188
rect 559984 3148 564532 3176
rect 559984 3136 559990 3148
rect 564526 3136 564532 3148
rect 564584 3136 564590 3188
rect 364334 3068 364340 3120
rect 364392 3108 364398 3120
rect 378226 3108 378232 3120
rect 364392 3080 378232 3108
rect 364392 3068 364398 3080
rect 378226 3068 378232 3080
rect 378284 3068 378290 3120
rect 388254 3068 388260 3120
rect 388312 3108 388318 3120
rect 389082 3108 389088 3120
rect 388312 3080 389088 3108
rect 388312 3068 388318 3080
rect 389082 3068 389088 3080
rect 389140 3068 389146 3120
rect 403618 3068 403624 3120
rect 403676 3108 403682 3120
rect 413278 3108 413284 3120
rect 403676 3080 413284 3108
rect 403676 3068 403682 3080
rect 413278 3068 413284 3080
rect 413336 3068 413342 3120
rect 421558 3068 421564 3120
rect 421616 3108 421622 3120
rect 474734 3108 474740 3120
rect 421616 3080 474740 3108
rect 421616 3068 421622 3080
rect 474734 3068 474740 3080
rect 474792 3068 474798 3120
rect 2866 3000 2872 3052
rect 2924 3040 2930 3052
rect 8938 3040 8944 3052
rect 2924 3012 8944 3040
rect 2924 3000 2930 3012
rect 8938 3000 8944 3012
rect 8996 3000 9002 3052
rect 26694 3000 26700 3052
rect 26752 3040 26758 3052
rect 27522 3040 27528 3052
rect 26752 3012 27528 3040
rect 26752 3000 26758 3012
rect 27522 3000 27528 3012
rect 27580 3000 27586 3052
rect 190822 3000 190828 3052
rect 190880 3040 190886 3052
rect 263594 3040 263600 3052
rect 190880 3012 263600 3040
rect 190880 3000 190886 3012
rect 263594 3000 263600 3012
rect 263652 3000 263658 3052
rect 337102 3000 337108 3052
rect 337160 3040 337166 3052
rect 338022 3040 338028 3052
rect 337160 3012 338028 3040
rect 337160 3000 337166 3012
rect 338022 3000 338028 3012
rect 338080 3000 338086 3052
rect 382366 3000 382372 3052
rect 382424 3040 382430 3052
rect 426250 3040 426256 3052
rect 382424 3012 426256 3040
rect 382424 3000 382430 3012
rect 426250 3000 426256 3012
rect 426308 3000 426314 3052
rect 431954 3000 431960 3052
rect 432012 3040 432018 3052
rect 439314 3040 439320 3052
rect 432012 3012 439320 3040
rect 432012 3000 432018 3012
rect 439314 3000 439320 3012
rect 439372 3000 439378 3052
rect 439406 3000 439412 3052
rect 439464 3040 439470 3052
rect 448146 3040 448152 3052
rect 439464 3012 448152 3040
rect 439464 3000 439470 3012
rect 448146 3000 448152 3012
rect 448204 3000 448210 3052
rect 450170 3000 450176 3052
rect 450228 3040 450234 3052
rect 468294 3040 468300 3052
rect 450228 3012 468300 3040
rect 450228 3000 450234 3012
rect 468294 3000 468300 3012
rect 468352 3000 468358 3052
rect 158714 2932 158720 2984
rect 158772 2972 158778 2984
rect 160002 2972 160008 2984
rect 158772 2944 160008 2972
rect 158772 2932 158778 2944
rect 160002 2932 160008 2944
rect 160060 2932 160066 2984
rect 251450 2932 251456 2984
rect 251508 2972 251514 2984
rect 300762 2972 300768 2984
rect 251508 2944 300768 2972
rect 251508 2932 251514 2944
rect 300762 2932 300768 2944
rect 300820 2932 300826 2984
rect 319254 2932 319260 2984
rect 319312 2972 319318 2984
rect 320082 2972 320088 2984
rect 319312 2944 320088 2972
rect 319312 2932 319318 2944
rect 320082 2932 320088 2944
rect 320140 2932 320146 2984
rect 383580 2944 383700 2972
rect 115934 2864 115940 2916
rect 115992 2904 115998 2916
rect 117222 2904 117228 2916
rect 115992 2876 117228 2904
rect 115992 2864 115998 2876
rect 117222 2864 117228 2876
rect 117280 2864 117286 2916
rect 183738 2864 183744 2916
rect 183796 2904 183802 2916
rect 256694 2904 256700 2916
rect 183796 2876 256700 2904
rect 183796 2864 183802 2876
rect 256694 2864 256700 2876
rect 256752 2864 256758 2916
rect 343082 2864 343088 2916
rect 343140 2904 343146 2916
rect 356054 2904 356060 2916
rect 343140 2876 356060 2904
rect 343140 2864 343146 2876
rect 356054 2864 356060 2876
rect 356112 2864 356118 2916
rect 369118 2864 369124 2916
rect 369176 2904 369182 2916
rect 374086 2904 374092 2916
rect 369176 2876 374092 2904
rect 369176 2864 369182 2876
rect 374086 2864 374092 2876
rect 374144 2864 374150 2916
rect 262214 2796 262220 2848
rect 262272 2836 262278 2848
rect 318702 2836 318708 2848
rect 262272 2808 318708 2836
rect 262272 2796 262278 2808
rect 318702 2796 318708 2808
rect 318760 2796 318766 2848
rect 378962 2796 378968 2848
rect 379020 2836 379026 2848
rect 383580 2836 383608 2944
rect 383672 2916 383700 2944
rect 398834 2932 398840 2984
rect 398892 2972 398898 2984
rect 412634 2972 412640 2984
rect 398892 2944 412640 2972
rect 398892 2932 398898 2944
rect 412634 2932 412640 2944
rect 412692 2932 412698 2984
rect 439590 2932 439596 2984
rect 439648 2972 439654 2984
rect 450078 2972 450084 2984
rect 439648 2944 450084 2972
rect 439648 2932 439654 2944
rect 450078 2932 450084 2944
rect 450136 2932 450142 2984
rect 453666 2932 453672 2984
rect 453724 2972 453730 2984
rect 461578 2972 461584 2984
rect 453724 2944 461584 2972
rect 453724 2932 453730 2944
rect 461578 2932 461584 2944
rect 461636 2932 461642 2984
rect 383654 2864 383660 2916
rect 383712 2864 383718 2916
rect 383838 2864 383844 2916
rect 383896 2904 383902 2916
rect 398742 2904 398748 2916
rect 383896 2876 398748 2904
rect 383896 2864 383902 2876
rect 398742 2864 398748 2876
rect 398800 2864 398806 2916
rect 541710 2864 541716 2916
rect 541768 2904 541774 2916
rect 548058 2904 548064 2916
rect 541768 2876 548064 2904
rect 541768 2864 541774 2876
rect 548058 2864 548064 2876
rect 548116 2864 548122 2916
rect 555418 2864 555424 2916
rect 555476 2904 555482 2916
rect 558362 2904 558368 2916
rect 555476 2876 558368 2904
rect 555476 2864 555482 2876
rect 558362 2864 558368 2876
rect 558420 2864 558426 2916
rect 379020 2808 383608 2836
rect 379020 2796 379026 2808
rect 414198 2796 414204 2848
rect 414256 2836 414262 2848
rect 414256 2808 426388 2836
rect 414256 2796 414262 2808
rect 426360 2768 426388 2808
rect 442994 2796 443000 2848
rect 443052 2836 443058 2848
rect 444190 2836 444196 2848
rect 443052 2808 444196 2836
rect 443052 2796 443058 2808
rect 444190 2796 444196 2808
rect 444248 2796 444254 2848
rect 431954 2768 431960 2780
rect 426360 2740 431960 2768
rect 431954 2728 431960 2740
rect 432012 2728 432018 2780
rect 441522 2728 441528 2780
rect 441580 2768 441586 2780
rect 441580 2740 456104 2768
rect 441580 2728 441586 2740
rect 300762 2660 300768 2712
rect 300820 2700 300826 2712
rect 454310 2700 454316 2712
rect 300820 2672 454316 2700
rect 300820 2660 300826 2672
rect 454310 2660 454316 2672
rect 454368 2660 454374 2712
rect 456076 2700 456104 2740
rect 483106 2700 483112 2712
rect 456076 2672 483112 2700
rect 483106 2660 483112 2672
rect 483164 2660 483170 2712
rect 333606 2592 333612 2644
rect 333664 2632 333670 2644
rect 480346 2632 480352 2644
rect 333664 2604 480352 2632
rect 333664 2592 333670 2604
rect 480346 2592 480352 2604
rect 480404 2592 480410 2644
rect 308582 2524 308588 2576
rect 308640 2564 308646 2576
rect 472158 2564 472164 2576
rect 308640 2536 472164 2564
rect 308640 2524 308646 2536
rect 472158 2524 472164 2536
rect 472216 2524 472222 2576
rect 274082 2456 274088 2508
rect 274140 2496 274146 2508
rect 461302 2496 461308 2508
rect 274140 2468 461308 2496
rect 274140 2456 274146 2468
rect 461302 2456 461308 2468
rect 461360 2456 461366 2508
rect 244366 2388 244372 2440
rect 244424 2428 244430 2440
rect 451550 2428 451556 2440
rect 244424 2400 451556 2428
rect 244424 2388 244430 2400
rect 451550 2388 451556 2400
rect 451608 2388 451614 2440
rect 237190 2320 237196 2372
rect 237248 2360 237254 2372
rect 448698 2360 448704 2372
rect 237248 2332 448704 2360
rect 237248 2320 237254 2332
rect 448698 2320 448704 2332
rect 448756 2320 448762 2372
rect 201494 2252 201500 2304
rect 201552 2292 201558 2304
rect 437566 2292 437572 2304
rect 201552 2264 437572 2292
rect 201552 2252 201558 2264
rect 437566 2252 437572 2264
rect 437624 2252 437630 2304
rect 194410 2184 194416 2236
rect 194468 2224 194474 2236
rect 434806 2224 434812 2236
rect 194468 2196 434812 2224
rect 194468 2184 194474 2196
rect 434806 2184 434812 2196
rect 434864 2184 434870 2236
rect 162302 2116 162308 2168
rect 162360 2156 162366 2168
rect 425054 2156 425060 2168
rect 162360 2128 425060 2156
rect 162360 2116 162366 2128
rect 425054 2116 425060 2128
rect 425112 2116 425118 2168
rect 431954 2116 431960 2168
rect 432012 2156 432018 2168
rect 441522 2156 441528 2168
rect 432012 2128 441528 2156
rect 432012 2116 432018 2128
rect 441522 2116 441528 2128
rect 441580 2116 441586 2168
rect 133782 2048 133788 2100
rect 133840 2088 133846 2100
rect 415578 2088 415584 2100
rect 133840 2060 415584 2088
rect 133840 2048 133846 2060
rect 415578 2048 415584 2060
rect 415636 2048 415642 2100
rect 417970 2048 417976 2100
rect 418028 2088 418034 2100
rect 508038 2088 508044 2100
rect 418028 2060 508044 2088
rect 418028 2048 418034 2060
rect 508038 2048 508044 2060
rect 508096 2048 508102 2100
rect 345474 1980 345480 2032
rect 345532 2020 345538 2032
rect 484670 2020 484676 2032
rect 345532 1992 484676 2020
rect 345532 1980 345538 1992
rect 484670 1980 484676 1992
rect 484728 1980 484734 2032
rect 318702 1912 318708 1964
rect 318760 1952 318766 1964
rect 456886 1952 456892 1964
rect 318760 1924 456892 1952
rect 318760 1912 318766 1924
rect 456886 1912 456892 1924
rect 456944 1912 456950 1964
rect 379974 1844 379980 1896
rect 380032 1884 380038 1896
rect 495710 1884 495716 1896
rect 380032 1856 495716 1884
rect 380032 1844 380038 1856
rect 495710 1844 495716 1856
rect 495768 1844 495774 1896
rect 390646 1776 390652 1828
rect 390704 1816 390710 1828
rect 493686 1816 493692 1828
rect 390704 1788 493692 1816
rect 390704 1776 390710 1788
rect 493686 1776 493692 1788
rect 493744 1776 493750 1828
rect 401318 1708 401324 1760
rect 401376 1748 401382 1760
rect 502610 1748 502616 1760
rect 401376 1720 502616 1748
rect 401376 1708 401382 1720
rect 502610 1708 502616 1720
rect 502668 1708 502674 1760
rect 263594 1640 263600 1692
rect 263652 1680 263658 1692
rect 434990 1680 434996 1692
rect 263652 1652 434996 1680
rect 263652 1640 263658 1652
rect 434990 1640 434996 1652
rect 435048 1640 435054 1692
rect 366910 892 366916 944
rect 366968 932 366974 944
rect 491478 932 491484 944
rect 366968 904 491484 932
rect 366968 892 366974 904
rect 491478 892 491484 904
rect 491536 892 491542 944
rect 341886 824 341892 876
rect 341944 864 341950 876
rect 483290 864 483296 876
rect 341944 836 483296 864
rect 341944 824 341950 836
rect 483290 824 483296 836
rect 483348 824 483354 876
rect 326430 756 326436 808
rect 326488 796 326494 808
rect 477678 796 477684 808
rect 326488 768 477684 796
rect 326488 756 326494 768
rect 477678 756 477684 768
rect 477736 756 477742 808
rect 322842 688 322848 740
rect 322900 728 322906 740
rect 476206 728 476212 740
rect 322900 700 476212 728
rect 322900 688 322906 700
rect 476206 688 476212 700
rect 476264 688 476270 740
rect 315758 620 315764 672
rect 315816 660 315822 672
rect 474918 660 474924 672
rect 315816 632 474924 660
rect 315816 620 315822 632
rect 474918 620 474924 632
rect 474976 620 474982 672
rect 202506 552 202512 604
rect 202564 592 202570 604
rect 202690 592 202696 604
rect 202564 564 202696 592
rect 202564 552 202570 564
rect 202690 552 202696 564
rect 202748 552 202754 604
rect 220538 552 220544 604
rect 220596 592 220602 604
rect 220722 592 220728 604
rect 220596 564 220728 592
rect 220596 552 220602 564
rect 220722 552 220728 564
rect 220780 552 220786 604
rect 259822 552 259828 604
rect 259880 552 259886 604
rect 265802 552 265808 604
rect 265860 552 265866 604
rect 270494 552 270500 604
rect 270552 552 270558 604
rect 307294 552 307300 604
rect 307352 592 307358 604
rect 307386 592 307392 604
rect 307352 564 307392 592
rect 307352 552 307358 564
rect 307386 552 307392 564
rect 307444 552 307450 604
rect 312170 552 312176 604
rect 312228 592 312234 604
rect 473446 592 473452 604
rect 312228 564 473452 592
rect 312228 552 312234 564
rect 473446 552 473452 564
rect 473504 552 473510 604
rect 496538 552 496544 604
rect 496596 592 496602 604
rect 496722 592 496728 604
rect 496596 564 496728 592
rect 496596 552 496602 564
rect 496722 552 496728 564
rect 496780 552 496786 604
rect 564434 552 564440 604
rect 564492 592 564498 604
rect 565538 592 565544 604
rect 564492 564 565544 592
rect 564492 552 564498 564
rect 565538 552 565544 564
rect 565596 552 565602 604
rect 259840 388 259868 552
rect 265820 456 265848 552
rect 270512 524 270540 552
rect 459830 524 459836 536
rect 270512 496 459836 524
rect 459830 484 459836 496
rect 459888 484 459894 536
rect 458634 456 458640 468
rect 265820 428 458640 456
rect 458634 416 458640 428
rect 458692 416 458698 468
rect 457070 388 457076 400
rect 259840 360 457076 388
rect 457070 348 457076 360
rect 457128 348 457134 400
rect 213638 280 213644 332
rect 213696 320 213702 332
rect 441614 320 441620 332
rect 213696 292 441620 320
rect 213696 280 213702 292
rect 441614 280 441620 292
rect 441672 280 441678 332
rect 199378 212 199384 264
rect 199436 252 199442 264
rect 437658 252 437664 264
rect 199436 224 437664 252
rect 199436 212 199442 224
rect 437658 212 437664 224
rect 437716 212 437722 264
rect 195790 144 195796 196
rect 195848 184 195854 196
rect 436094 184 436100 196
rect 195848 156 436100 184
rect 195848 144 195854 156
rect 436094 144 436100 156
rect 436152 144 436158 196
rect 188614 76 188620 128
rect 188672 116 188678 128
rect 433794 116 433800 128
rect 188672 88 433800 116
rect 188672 76 188678 88
rect 433794 76 433800 88
rect 433852 76 433858 128
rect 170766 8 170772 60
rect 170824 48 170830 60
rect 428090 48 428096 60
rect 170824 20 428096 48
rect 170824 8 170830 20
rect 428090 8 428096 20
rect 428148 8 428154 60
<< via1 >>
rect 287704 700544 287756 700596
rect 332508 700544 332560 700596
rect 305644 700476 305696 700528
rect 397460 700476 397512 700528
rect 313924 700408 313976 700460
rect 413652 700408 413704 700460
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 138664 700340 138716 700392
rect 154120 700340 154172 700392
rect 308404 700340 308456 700392
rect 462320 700340 462372 700392
rect 8116 700272 8168 700324
rect 8944 700272 8996 700324
rect 89168 700272 89220 700324
rect 138756 700272 138808 700324
rect 202788 700272 202840 700324
rect 250904 700272 250956 700324
rect 267648 700272 267700 700324
rect 282276 700272 282328 700324
rect 309784 700272 309836 700324
rect 527180 700272 527232 700324
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 250904 699116 250956 699168
rect 253204 699116 253256 699168
rect 283288 698232 283340 698284
rect 283932 698232 283984 698284
rect 576124 696940 576176 696992
rect 580172 696940 580224 696992
rect 133144 696872 133196 696924
rect 137836 696872 137888 696924
rect 253204 696872 253256 696924
rect 260012 696872 260064 696924
rect 260012 694764 260064 694816
rect 267004 694764 267056 694816
rect 218980 694152 219032 694204
rect 219164 694152 219216 694204
rect 283104 694084 283156 694136
rect 283288 694084 283340 694136
rect 219164 688644 219216 688696
rect 219072 688576 219124 688628
rect 283012 684496 283064 684548
rect 283104 684496 283156 684548
rect 3516 681708 3568 681760
rect 453304 681708 453356 681760
rect 218796 676132 218848 676184
rect 218980 676132 219032 676184
rect 122104 675452 122156 675504
rect 133144 675452 133196 675504
rect 267004 670624 267056 670676
rect 268384 670624 268436 670676
rect 218796 666544 218848 666596
rect 219072 666544 219124 666596
rect 283104 666544 283156 666596
rect 283380 666544 283432 666596
rect 283104 661716 283156 661768
rect 283380 661716 283432 661768
rect 268384 661172 268436 661224
rect 270408 661172 270460 661224
rect 219164 659608 219216 659660
rect 219348 659608 219400 659660
rect 116584 658520 116636 658572
rect 122104 658520 122156 658572
rect 270408 656888 270460 656940
rect 219072 656820 219124 656872
rect 219348 656820 219400 656872
rect 283104 656888 283156 656940
rect 283196 656888 283248 656940
rect 273260 656820 273312 656872
rect 273260 654100 273312 654152
rect 276664 654032 276716 654084
rect 3056 652740 3108 652792
rect 10324 652740 10376 652792
rect 577504 650020 577556 650072
rect 579620 650020 579672 650072
rect 113824 648864 113876 648916
rect 116584 648864 116636 648916
rect 219072 647232 219124 647284
rect 219256 647232 219308 647284
rect 283104 647232 283156 647284
rect 283196 647232 283248 647284
rect 554412 647232 554464 647284
rect 556252 647232 556304 647284
rect 219256 640364 219308 640416
rect 283104 640364 283156 640416
rect 283196 640364 283248 640416
rect 219072 640228 219124 640280
rect 219072 637508 219124 637560
rect 219164 637508 219216 637560
rect 276664 635060 276716 635112
rect 278044 635060 278096 635112
rect 110420 632408 110472 632460
rect 113824 632408 113876 632460
rect 282920 630640 282972 630692
rect 283196 630640 283248 630692
rect 105544 629280 105596 629332
rect 110420 629280 110472 629332
rect 219164 627920 219216 627972
rect 219348 627920 219400 627972
rect 41328 627172 41380 627224
rect 312544 627172 312596 627224
rect 278044 626492 278096 626544
rect 279148 626492 279200 626544
rect 95884 621732 95936 621784
rect 105544 621732 105596 621784
rect 24768 621664 24820 621716
rect 283012 621664 283064 621716
rect 219072 620984 219124 621036
rect 219348 620984 219400 621036
rect 23388 619624 23440 619676
rect 84108 619624 84160 619676
rect 219072 618876 219124 618928
rect 284300 618876 284352 618928
rect 31484 617448 31536 617500
rect 91100 617448 91152 617500
rect 28632 616768 28684 616820
rect 28632 616564 28684 616616
rect 30288 616564 30340 616616
rect 28632 616428 28684 616480
rect 30196 616428 30248 616480
rect 28264 615680 28316 615732
rect 453304 616768 453356 616820
rect 456800 616768 456852 616820
rect 551100 616156 551152 616208
rect 551744 616156 551796 616208
rect 282920 611328 282972 611380
rect 283288 611328 283340 611380
rect 3332 609968 3384 610020
rect 11704 609968 11756 610020
rect 554136 609968 554188 610020
rect 555516 609968 555568 610020
rect 551100 606500 551152 606552
rect 551836 606500 551888 606552
rect 23296 605820 23348 605872
rect 25228 605820 25280 605872
rect 24124 603440 24176 603492
rect 28264 603440 28316 603492
rect 551928 603032 551980 603084
rect 552664 603032 552716 603084
rect 551100 596844 551152 596896
rect 551836 596844 551888 596896
rect 551836 596708 551888 596760
rect 552664 596708 552716 596760
rect 3516 594804 3568 594856
rect 9036 594804 9088 594856
rect 139216 594668 139268 594720
rect 139584 594668 139636 594720
rect 28632 594192 28684 594244
rect 28632 593988 28684 594040
rect 282920 591948 282972 592000
rect 283196 591948 283248 592000
rect 554504 590656 554556 590708
rect 555608 590656 555660 590708
rect 554504 589296 554556 589348
rect 556160 589296 556212 589348
rect 554320 587868 554372 587920
rect 557632 587868 557684 587920
rect 28632 587800 28684 587852
rect 28724 587800 28776 587852
rect 28816 587324 28868 587376
rect 28908 587324 28960 587376
rect 551100 587188 551152 587240
rect 551836 587188 551888 587240
rect 554320 586984 554372 587036
rect 556804 586984 556856 587036
rect 28080 586644 28132 586696
rect 28908 586644 28960 586696
rect 28264 585556 28316 585608
rect 28816 585556 28868 585608
rect 554504 585216 554556 585268
rect 558920 585216 558972 585268
rect 554320 585148 554372 585200
rect 560300 585148 560352 585200
rect 28540 583720 28592 583772
rect 29000 583720 29052 583772
rect 554320 583720 554372 583772
rect 561772 583720 561824 583772
rect 283196 582428 283248 582480
rect 283196 582292 283248 582344
rect 554320 581000 554372 581052
rect 563060 581000 563112 581052
rect 554320 579640 554372 579692
rect 564440 579640 564492 579692
rect 26148 579164 26200 579216
rect 28908 579164 28960 579216
rect 28540 578892 28592 578944
rect 28724 578892 28776 578944
rect 28356 578756 28408 578808
rect 28540 578756 28592 578808
rect 554320 578212 554372 578264
rect 565820 578212 565872 578264
rect 551100 577532 551152 577584
rect 551836 577532 551888 577584
rect 554320 576852 554372 576904
rect 567292 576852 567344 576904
rect 28264 575560 28316 575612
rect 28908 575560 28960 575612
rect 554412 575492 554464 575544
rect 560944 575492 560996 575544
rect 554320 574132 554372 574184
rect 568580 574132 568632 574184
rect 554412 574064 554464 574116
rect 569960 574064 570012 574116
rect 29184 573452 29236 573504
rect 29460 573452 29512 573504
rect 30288 573452 30340 573504
rect 29552 573384 29604 573436
rect 28724 573248 28776 573300
rect 30288 573248 30340 573300
rect 29552 572704 29604 572756
rect 29736 572704 29788 572756
rect 283196 572704 283248 572756
rect 554412 572704 554464 572756
rect 571432 572704 571484 572756
rect 551100 572636 551152 572688
rect 551836 572636 551888 572688
rect 283196 572568 283248 572620
rect 199292 572500 199344 572552
rect 204260 572500 204312 572552
rect 198096 572364 198148 572416
rect 202972 572364 203024 572416
rect 189540 572296 189592 572348
rect 195980 572296 196032 572348
rect 196808 572296 196860 572348
rect 202880 572296 202932 572348
rect 188344 572228 188396 572280
rect 194600 572228 194652 572280
rect 206652 572160 206704 572212
rect 211160 572160 211212 572212
rect 25136 572092 25188 572144
rect 195612 572092 195664 572144
rect 201500 572092 201552 572144
rect 218888 572092 218940 572144
rect 222200 572092 222252 572144
rect 277308 572092 277360 572144
rect 279332 572092 279384 572144
rect 190276 572024 190328 572076
rect 197360 572024 197412 572076
rect 207848 572024 207900 572076
rect 212540 572024 212592 572076
rect 227444 572024 227496 572076
rect 229100 572024 229152 572076
rect 267648 572024 267700 572076
rect 268292 572024 268344 572076
rect 275928 572024 275980 572076
rect 278044 572024 278096 572076
rect 26792 571616 26844 571668
rect 31852 571616 31904 571668
rect 26700 571548 26752 571600
rect 33140 571548 33192 571600
rect 41420 571548 41472 571600
rect 209044 571956 209096 572008
rect 214012 571956 214064 572008
rect 194416 571888 194468 571940
rect 200120 571888 200172 571940
rect 216404 571888 216456 571940
rect 219440 571888 219492 571940
rect 205364 571616 205416 571668
rect 209780 571616 209832 571668
rect 217600 571616 217652 571668
rect 220820 571616 220872 571668
rect 228640 571616 228692 571668
rect 230480 571616 230532 571668
rect 202788 571548 202840 571600
rect 208400 571548 208452 571600
rect 213828 571548 213880 571600
rect 218060 571548 218112 571600
rect 220084 571548 220136 571600
rect 223580 571548 223632 571600
rect 224868 571548 224920 571600
rect 227812 571548 227864 571600
rect 26608 571480 26660 571532
rect 29000 571412 29052 571464
rect 30380 571412 30432 571464
rect 201408 571480 201460 571532
rect 207020 571480 207072 571532
rect 212448 571480 212500 571532
rect 216680 571480 216732 571532
rect 223488 571480 223540 571532
rect 226340 571480 226392 571532
rect 231032 571480 231084 571532
rect 233332 571480 233384 571532
rect 273168 571480 273220 571532
rect 275652 571480 275704 571532
rect 37280 571412 37332 571464
rect 191748 571412 191800 571464
rect 198832 571412 198884 571464
rect 200488 571412 200540 571464
rect 205640 571412 205692 571464
rect 211528 571412 211580 571464
rect 215300 571412 215352 571464
rect 222108 571412 222160 571464
rect 224960 571412 225012 571464
rect 233148 571412 233200 571464
rect 234620 571412 234672 571464
rect 235908 571412 235960 571464
rect 23204 571344 23256 571396
rect 25596 571344 25648 571396
rect 193128 571344 193180 571396
rect 198740 571344 198792 571396
rect 204168 571344 204220 571396
rect 208492 571344 208544 571396
rect 210332 571344 210384 571396
rect 213920 571344 213972 571396
rect 215208 571344 215260 571396
rect 218152 571344 218204 571396
rect 221280 571344 221332 571396
rect 223672 571344 223724 571396
rect 226156 571344 226208 571396
rect 227720 571344 227772 571396
rect 229836 571344 229888 571396
rect 231860 571344 231912 571396
rect 232320 571344 232372 571396
rect 233240 571344 233292 571396
rect 234528 571344 234580 571396
rect 236000 571344 236052 571396
rect 268936 571412 268988 571464
rect 270776 571412 270828 571464
rect 271788 571412 271840 571464
rect 273260 571412 273312 571464
rect 274548 571412 274600 571464
rect 276848 571412 276900 571464
rect 278596 571412 278648 571464
rect 281724 571412 281776 571464
rect 239588 571344 239640 571396
rect 240140 571344 240192 571396
rect 240876 571344 240928 571396
rect 241520 571344 241572 571396
rect 242072 571344 242124 571396
rect 242992 571344 243044 571396
rect 254860 571344 254912 571396
rect 255320 571344 255372 571396
rect 256056 571344 256108 571396
rect 256700 571344 256752 571396
rect 257344 571344 257396 571396
rect 264612 571344 264664 571396
rect 264888 571344 264940 571396
rect 265900 571344 265952 571396
rect 266268 571344 266320 571396
rect 267096 571344 267148 571396
rect 269028 571344 269080 571396
rect 269488 571344 269540 571396
rect 270408 571344 270460 571396
rect 271972 571344 272024 571396
rect 273076 571344 273128 571396
rect 274640 571344 274692 571396
rect 278688 571344 278740 571396
rect 280528 571344 280580 571396
rect 554228 571344 554280 571396
rect 558184 571344 558236 571396
rect 237380 571276 237432 571328
rect 253940 571276 253992 571328
rect 263508 571276 263560 571328
rect 551928 571208 551980 571260
rect 554596 571208 554648 571260
rect 28632 570800 28684 570852
rect 45652 570800 45704 570852
rect 29184 570732 29236 570784
rect 48320 570732 48372 570784
rect 29460 570664 29512 570716
rect 52460 570664 52512 570716
rect 248420 570664 248472 570716
rect 28540 570596 28592 570648
rect 53840 570596 53892 570648
rect 554320 570664 554372 570716
rect 248512 570460 248564 570512
rect 525708 570460 525760 570512
rect 543648 570392 543700 570444
rect 554504 570392 554556 570444
rect 318524 569916 318576 569968
rect 318708 569916 318760 569968
rect 354404 569916 354456 569968
rect 354588 569916 354640 569968
rect 547788 569916 547840 569968
rect 552940 569916 552992 569968
rect 554412 569916 554464 569968
rect 572720 569916 572772 569968
rect 29184 569848 29236 569900
rect 29736 569848 29788 569900
rect 112536 569848 112588 569900
rect 138664 569848 138716 569900
rect 281540 569848 281592 569900
rect 284392 569848 284444 569900
rect 28448 569304 28500 569356
rect 71780 569304 71832 569356
rect 25780 569236 25832 569288
rect 70400 569236 70452 569288
rect 56416 569168 56468 569220
rect 281540 569168 281592 569220
rect 286324 569168 286376 569220
rect 580540 569168 580592 569220
rect 549168 568556 549220 568608
rect 553032 568556 553084 568608
rect 338304 568488 338356 568540
rect 339316 568488 339368 568540
rect 340144 568488 340196 568540
rect 385040 568488 385092 568540
rect 456064 568488 456116 568540
rect 483664 568488 483716 568540
rect 336556 568420 336608 568472
rect 387892 568420 387944 568472
rect 327540 568352 327592 568404
rect 328276 568352 328328 568404
rect 332968 568352 333020 568404
rect 389364 568352 389416 568404
rect 329380 568284 329432 568336
rect 391940 568284 391992 568336
rect 325792 568216 325844 568268
rect 394700 568216 394752 568268
rect 336648 568148 336700 568200
rect 422576 568148 422628 568200
rect 335268 568080 335320 568132
rect 426164 568080 426216 568132
rect 332508 568012 332560 568064
rect 429752 568012 429804 568064
rect 331128 567944 331180 567996
rect 433340 567944 433392 567996
rect 328368 567876 328420 567928
rect 436928 567876 436980 567928
rect 326988 567808 327040 567860
rect 440516 567808 440568 567860
rect 343732 567740 343784 567792
rect 383752 567740 383804 567792
rect 345480 567672 345532 567724
rect 346308 567672 346360 567724
rect 347320 567672 347372 567724
rect 380900 567672 380952 567724
rect 29092 567604 29144 567656
rect 29460 567604 29512 567656
rect 350908 567604 350960 567656
rect 379520 567604 379572 567656
rect 361672 567536 361724 567588
rect 362868 567536 362920 567588
rect 363420 567536 363472 567588
rect 364248 567536 364300 567588
rect 3516 567196 3568 567248
rect 9128 567196 9180 567248
rect 320364 567196 320416 567248
rect 321468 567196 321520 567248
rect 356244 567196 356296 567248
rect 357348 567196 357400 567248
rect 529020 567196 529072 567248
rect 530584 567196 530636 567248
rect 355876 566448 355928 566500
rect 389180 566448 389232 566500
rect 29276 565700 29328 565752
rect 30012 565700 30064 565752
rect 339408 565088 339460 565140
rect 418160 565088 418212 565140
rect 532608 565088 532660 565140
rect 554780 565088 554832 565140
rect 342076 563660 342128 563712
rect 415400 563660 415452 563712
rect 528468 563660 528520 563712
rect 555148 563660 555200 563712
rect 29552 563184 29604 563236
rect 30288 563184 30340 563236
rect 551100 563048 551152 563100
rect 551836 563048 551888 563100
rect 346216 562300 346268 562352
rect 407120 562300 407172 562352
rect 538128 562300 538180 562352
rect 555516 562300 555568 562352
rect 347688 560940 347740 560992
rect 404360 560940 404412 560992
rect 533988 560940 534040 560992
rect 555332 560940 555384 560992
rect 29184 560260 29236 560312
rect 29736 560260 29788 560312
rect 350448 559512 350500 559564
rect 400220 559512 400272 559564
rect 529848 559512 529900 559564
rect 555056 559512 555108 559564
rect 283196 558900 283248 558952
rect 283380 558900 283432 558952
rect 29368 558492 29420 558544
rect 29644 558492 29696 558544
rect 29552 558152 29604 558204
rect 30288 558152 30340 558204
rect 351736 558152 351788 558204
rect 397460 558152 397512 558204
rect 483664 556452 483716 556504
rect 485780 556452 485832 556504
rect 304264 556180 304316 556232
rect 579804 556180 579856 556232
rect 354496 555432 354548 555484
rect 393320 555432 393372 555484
rect 358636 554004 358688 554056
rect 386420 554004 386472 554056
rect 485780 554004 485832 554056
rect 498200 554004 498252 554056
rect 29276 553392 29328 553444
rect 30012 553392 30064 553444
rect 283196 553392 283248 553444
rect 551008 553392 551060 553444
rect 551100 553324 551152 553376
rect 283288 553256 283340 553308
rect 324136 552644 324188 552696
rect 443000 552644 443052 552696
rect 540888 552644 540940 552696
rect 555240 552644 555292 552696
rect 3148 552032 3200 552084
rect 312544 552032 312596 552084
rect 329748 551284 329800 551336
rect 434720 551284 434772 551336
rect 498200 551284 498252 551336
rect 504364 551284 504416 551336
rect 536748 551284 536800 551336
rect 554964 551284 555016 551336
rect 29460 550536 29512 550588
rect 29736 550536 29788 550588
rect 332416 549856 332468 549908
rect 430580 549856 430632 549908
rect 551008 549244 551060 549296
rect 551100 549244 551152 549296
rect 333888 548496 333940 548548
rect 427820 548496 427872 548548
rect 549076 547680 549128 547732
rect 552756 547680 552808 547732
rect 26148 547476 26200 547528
rect 35900 547476 35952 547528
rect 26884 547408 26936 547460
rect 46940 547408 46992 547460
rect 26976 547340 27028 547392
rect 55312 547340 55364 547392
rect 28172 547272 28224 547324
rect 62120 547272 62172 547324
rect 27068 547204 27120 547256
rect 64880 547204 64932 547256
rect 531228 547204 531280 547256
rect 551652 547204 551704 547256
rect 27988 547136 28040 547188
rect 80060 547136 80112 547188
rect 336556 547136 336608 547188
rect 423680 547136 423732 547188
rect 527088 547136 527140 547188
rect 551560 547136 551612 547188
rect 550548 547068 550600 547120
rect 552848 547068 552900 547120
rect 366916 545776 366968 545828
rect 374000 545776 374052 545828
rect 322848 545708 322900 545760
rect 396080 545708 396132 545760
rect 326896 544348 326948 544400
rect 437480 544348 437532 544400
rect 283288 543804 283340 543856
rect 368388 543736 368440 543788
rect 369860 543736 369912 543788
rect 29368 543668 29420 543720
rect 30012 543668 30064 543720
rect 283104 543668 283156 543720
rect 367008 543260 367060 543312
rect 369860 543260 369912 543312
rect 324228 542988 324280 543040
rect 394884 542988 394936 543040
rect 364248 541696 364300 541748
rect 371332 541696 371384 541748
rect 325608 541628 325660 541680
rect 441620 541628 441672 541680
rect 29460 540948 29512 541000
rect 29736 540948 29788 541000
rect 360108 540268 360160 540320
rect 374000 540268 374052 540320
rect 343548 540200 343600 540252
rect 411260 540200 411312 540252
rect 29276 538840 29328 538892
rect 29552 538840 29604 538892
rect 357348 538840 357400 538892
rect 375472 538840 375524 538892
rect 524328 538840 524380 538892
rect 554872 538840 554924 538892
rect 3516 538228 3568 538280
rect 10416 538228 10468 538280
rect 353208 537480 353260 537532
rect 378232 537480 378284 537532
rect 165436 537344 165488 537396
rect 431040 537344 431092 537396
rect 163228 537276 163280 537328
rect 433340 537276 433392 537328
rect 158904 537208 158956 537260
rect 437572 537208 437624 537260
rect 156788 537140 156840 537192
rect 439688 537140 439740 537192
rect 152464 537072 152516 537124
rect 444380 537072 444432 537124
rect 150348 537004 150400 537056
rect 446128 537004 446180 537056
rect 148140 536936 148192 536988
rect 448704 536936 448756 536988
rect 146024 536868 146076 536920
rect 450452 536868 450504 536920
rect 112628 536800 112680 536852
rect 483848 536800 483900 536852
rect 363788 536256 363840 536308
rect 376760 536256 376812 536308
rect 317328 536188 317380 536240
rect 400220 536188 400272 536240
rect 194508 536120 194560 536172
rect 401968 536120 402020 536172
rect 193404 536052 193456 536104
rect 403164 536052 403216 536104
rect 154672 535984 154724 536036
rect 441804 535984 441856 536036
rect 139492 535916 139544 535968
rect 456984 535916 457036 535968
rect 137376 535848 137428 535900
rect 459100 535848 459152 535900
rect 127716 535780 127768 535832
rect 468760 535780 468812 535832
rect 125508 535712 125560 535764
rect 470968 535712 471020 535764
rect 123392 535644 123444 535696
rect 473452 535644 473504 535696
rect 121184 535576 121236 535628
rect 475292 535576 475344 535628
rect 117964 535508 118016 535560
rect 478880 535508 478932 535560
rect 109316 535440 109368 535492
rect 483664 535440 483716 535492
rect 364892 535100 364944 535152
rect 28356 534964 28408 535016
rect 37188 534964 37240 535016
rect 25412 534896 25464 534948
rect 34980 534896 35032 534948
rect 362868 534896 362920 534948
rect 372896 535032 372948 535084
rect 365628 534964 365680 535016
rect 370688 534964 370740 535016
rect 375380 534964 375432 535016
rect 367008 534896 367060 534948
rect 371240 534896 371292 534948
rect 25688 534828 25740 534880
rect 39304 534828 39356 534880
rect 358728 534828 358780 534880
rect 375380 534828 375432 534880
rect 28080 534760 28132 534812
rect 41420 534760 41472 534812
rect 362776 534760 362828 534812
rect 379612 534760 379664 534812
rect 25872 534692 25924 534744
rect 43628 534692 43680 534744
rect 360568 534692 360620 534744
rect 382280 534692 382332 534744
rect 192392 534624 192444 534676
rect 404452 534624 404504 534676
rect 189080 534556 189132 534608
rect 407396 534556 407448 534608
rect 185860 534488 185912 534540
rect 410616 534488 410668 534540
rect 179420 534420 179472 534472
rect 417056 534420 417108 534472
rect 177304 534352 177356 534404
rect 419632 534352 419684 534404
rect 172980 534284 173032 534336
rect 423680 534284 423732 534336
rect 170772 534216 170824 534268
rect 425704 534216 425756 534268
rect 166448 534148 166500 534200
rect 430028 534148 430080 534200
rect 29368 534080 29420 534132
rect 30012 534080 30064 534132
rect 164332 534080 164384 534132
rect 432144 534080 432196 534132
rect 342168 534012 342220 534064
rect 385132 534012 385184 534064
rect 339316 533944 339368 533996
rect 386880 533944 386932 533996
rect 335176 533876 335228 533928
rect 389180 533876 389232 533928
rect 30196 533808 30248 533860
rect 52276 533808 52328 533860
rect 331036 533808 331088 533860
rect 391204 533808 391256 533860
rect 518716 533808 518768 533860
rect 553860 533808 553912 533860
rect 25964 533740 26016 533792
rect 50068 533740 50120 533792
rect 328276 533740 328328 533792
rect 393320 533740 393372 533792
rect 516876 533740 516928 533792
rect 553768 533740 553820 533792
rect 30012 533672 30064 533724
rect 60832 533672 60884 533724
rect 318708 533672 318760 533724
rect 398932 533672 398984 533724
rect 514668 533672 514720 533724
rect 551192 533672 551244 533724
rect 26056 533604 26108 533656
rect 58716 533604 58768 533656
rect 322848 533604 322900 533656
rect 445760 533604 445812 533656
rect 512552 533604 512604 533656
rect 553676 533604 553728 533656
rect 27160 533536 27212 533588
rect 69480 533536 69532 533588
rect 321284 533536 321336 533588
rect 447140 533536 447192 533588
rect 510436 533536 510488 533588
rect 553584 533536 553636 533588
rect 27252 533468 27304 533520
rect 73804 533468 73856 533520
rect 320732 533468 320784 533520
rect 448520 533468 448572 533520
rect 530584 533468 530636 533520
rect 574376 533468 574428 533520
rect 27344 533400 27396 533452
rect 78128 533400 78180 533452
rect 319628 533400 319680 533452
rect 451280 533400 451332 533452
rect 508228 533400 508280 533452
rect 553492 533400 553544 533452
rect 27620 533332 27672 533384
rect 80244 533332 80296 533384
rect 318524 533332 318576 533384
rect 452660 533332 452712 533384
rect 503628 533332 503680 533384
rect 553400 533332 553452 533384
rect 346308 533264 346360 533316
rect 382556 533264 382608 533316
rect 349068 533196 349120 533248
rect 380440 533196 380492 533248
rect 354588 533128 354640 533180
rect 377220 533128 377272 533180
rect 188068 532788 188120 532840
rect 408592 532788 408644 532840
rect 168656 532720 168708 532772
rect 427912 532720 427964 532772
rect 357256 532652 357308 532704
rect 387800 532652 387852 532704
rect 504364 532652 504416 532704
rect 508504 532652 508556 532704
rect 355232 532584 355284 532636
rect 392032 532584 392084 532636
rect 353024 532516 353076 532568
rect 394792 532516 394844 532568
rect 261300 532448 261352 532500
rect 262128 532448 262180 532500
rect 262404 532448 262456 532500
rect 263416 532448 263468 532500
rect 350908 532448 350960 532500
rect 398840 532448 398892 532500
rect 348700 532380 348752 532432
rect 401600 532380 401652 532432
rect 346308 532312 346360 532364
rect 405740 532312 405792 532364
rect 344376 532244 344428 532296
rect 409880 532244 409932 532296
rect 342168 532176 342220 532228
rect 412640 532176 412692 532228
rect 30288 532108 30340 532160
rect 40408 532108 40460 532160
rect 340052 532108 340104 532160
rect 416780 532108 416832 532160
rect 521200 532108 521252 532160
rect 553952 532108 554004 532160
rect 27436 532040 27488 532092
rect 87788 532040 87840 532092
rect 321468 532040 321520 532092
rect 397644 532040 397696 532092
rect 401508 532040 401560 532092
rect 455420 532040 455472 532092
rect 517980 532040 518032 532092
rect 551284 532040 551336 532092
rect 27528 531972 27580 532024
rect 89996 531972 90048 532024
rect 337936 531972 337988 532024
rect 419540 531972 419592 532024
rect 513656 531972 513708 532024
rect 550732 531972 550784 532024
rect 359464 531904 359516 531956
rect 383660 531904 383712 531956
rect 361488 531836 361540 531888
rect 380992 531836 381044 531888
rect 178316 531768 178368 531820
rect 340144 531768 340196 531820
rect 176200 531700 176252 531752
rect 343640 531700 343692 531752
rect 173992 531632 174044 531684
rect 349068 531632 349120 531684
rect 171876 531564 171928 531616
rect 351920 531564 351972 531616
rect 169760 531496 169812 531548
rect 357348 531496 357400 531548
rect 183744 531428 183796 531480
rect 412732 531428 412784 531480
rect 147036 531360 147088 531412
rect 449440 531360 449492 531412
rect 142804 531292 142856 531344
rect 454040 531292 454092 531344
rect 544844 531292 544896 531344
rect 551744 531292 551796 531344
rect 30104 531224 30156 531276
rect 51172 531224 51224 531276
rect 331496 531224 331548 531276
rect 332416 531224 332468 531276
rect 334716 531224 334768 531276
rect 335268 531224 335320 531276
rect 335820 531224 335872 531276
rect 336556 531224 336608 531276
rect 341156 531224 341208 531276
rect 342076 531224 342128 531276
rect 345480 531224 345532 531276
rect 346216 531224 346268 531276
rect 349804 531224 349856 531276
rect 350448 531224 350500 531276
rect 354036 531224 354088 531276
rect 354496 531224 354548 531276
rect 365996 531224 366048 531276
rect 366916 531224 366968 531276
rect 483664 531224 483716 531276
rect 487160 531224 487212 531276
rect 526536 531224 526588 531276
rect 527088 531224 527140 531276
rect 527640 531224 527692 531276
rect 528468 531224 528520 531276
rect 530860 531224 530912 531276
rect 531228 531224 531280 531276
rect 531964 531224 532016 531276
rect 532608 531224 532660 531276
rect 536288 531224 536340 531276
rect 536748 531224 536800 531276
rect 545580 531224 545632 531276
rect 552020 531224 552072 531276
rect 553216 531224 553268 531276
rect 554044 531224 554096 531276
rect 29920 531156 29972 531208
rect 55496 531156 55548 531208
rect 24584 531088 24636 531140
rect 25320 531088 25372 531140
rect 25504 531088 25556 531140
rect 27436 531088 27488 531140
rect 27896 531088 27948 531140
rect 57612 531088 57664 531140
rect 119068 531088 119120 531140
rect 477500 531088 477552 531140
rect 543556 531088 543608 531140
rect 552480 531156 552532 531208
rect 551376 531088 551428 531140
rect 551928 531088 551980 531140
rect 29828 531020 29880 531072
rect 59820 531020 59872 531072
rect 198740 531020 198792 531072
rect 199660 531020 199712 531072
rect 213920 531020 213972 531072
rect 214748 531020 214800 531072
rect 227720 531020 227772 531072
rect 228732 531020 228784 531072
rect 233240 531020 233292 531072
rect 234068 531020 234120 531072
rect 242900 531020 242952 531072
rect 243820 531020 243872 531072
rect 248420 531020 248472 531072
rect 249156 531020 249208 531072
rect 266728 531020 266780 531072
rect 267648 531020 267700 531072
rect 267832 531020 267884 531072
rect 269028 531020 269080 531072
rect 272064 531020 272116 531072
rect 273076 531020 273128 531072
rect 276388 531020 276440 531072
rect 277308 531020 277360 531072
rect 277492 531020 277544 531072
rect 278688 531020 278740 531072
rect 325056 531020 325108 531072
rect 325608 531020 325660 531072
rect 329288 531020 329340 531072
rect 329748 531020 329800 531072
rect 330392 531020 330444 531072
rect 331128 531020 331180 531072
rect 357348 531020 357400 531072
rect 426716 531020 426768 531072
rect 541624 531020 541676 531072
rect 27804 530952 27856 531004
rect 61936 530952 61988 531004
rect 271052 530952 271104 531004
rect 271788 530952 271840 531004
rect 351920 530952 351972 531004
rect 424600 530952 424652 531004
rect 539508 530952 539560 531004
rect 545764 530952 545816 531004
rect 545948 531020 546000 531072
rect 552572 531020 552624 531072
rect 552388 530952 552440 531004
rect 29736 530884 29788 530936
rect 64052 530884 64104 530936
rect 326068 530884 326120 530936
rect 326988 530884 327040 530936
rect 349068 530884 349120 530936
rect 422484 530884 422536 530936
rect 537300 530884 537352 530936
rect 552204 530884 552256 530936
rect 29552 530816 29604 530868
rect 66260 530816 66312 530868
rect 343640 530816 343692 530868
rect 420276 530816 420328 530868
rect 523316 530816 523368 530868
rect 524328 530816 524380 530868
rect 535184 530816 535236 530868
rect 545672 530816 545724 530868
rect 545764 530816 545816 530868
rect 552296 530816 552348 530868
rect 27712 530748 27764 530800
rect 68376 530748 68428 530800
rect 340144 530748 340196 530800
rect 418252 530748 418304 530800
rect 533068 530748 533120 530800
rect 551468 530748 551520 530800
rect 25228 530680 25280 530732
rect 67364 530680 67416 530732
rect 186964 530680 187016 530732
rect 409880 530680 409932 530732
rect 528468 530680 528520 530732
rect 545580 530680 545632 530732
rect 545672 530680 545724 530732
rect 552112 530680 552164 530732
rect 555424 530680 555476 530732
rect 562600 530680 562652 530732
rect 23296 530612 23348 530664
rect 22100 530544 22152 530596
rect 23388 530544 23440 530596
rect 24768 530612 24820 530664
rect 77024 530612 77076 530664
rect 184848 530612 184900 530664
rect 411628 530612 411680 530664
rect 522212 530612 522264 530664
rect 551284 530612 551336 530664
rect 85672 530544 85724 530596
rect 182640 530544 182692 530596
rect 414020 530544 414072 530596
rect 505008 530544 505060 530596
rect 556252 530544 556304 530596
rect 558184 530544 558236 530596
rect 572260 530544 572312 530596
rect 24676 530476 24728 530528
rect 44732 530476 44784 530528
rect 115848 530476 115900 530528
rect 348884 530476 348936 530528
rect 29276 530408 29328 530460
rect 46848 530408 46900 530460
rect 180524 530408 180576 530460
rect 415952 530408 416004 530460
rect 25044 530340 25096 530392
rect 32864 530340 32916 530392
rect 133052 530340 133104 530392
rect 463792 530340 463844 530392
rect 130936 530272 130988 530324
rect 465540 530272 465592 530324
rect 128728 530204 128780 530256
rect 467840 530204 467892 530256
rect 24952 530136 25004 530188
rect 29644 530136 29696 530188
rect 126612 530136 126664 530188
rect 469864 530136 469916 530188
rect 542728 530136 542780 530188
rect 543648 530136 543700 530188
rect 547052 530136 547104 530188
rect 547788 530136 547840 530188
rect 548156 530136 548208 530188
rect 549076 530136 549128 530188
rect 124404 530068 124456 530120
rect 472072 530068 472124 530120
rect 122288 530000 122340 530052
rect 474188 530000 474240 530052
rect 419448 529932 419500 529984
rect 429292 529932 429344 529984
rect 556804 529932 556856 529984
rect 558276 529932 558328 529984
rect 560944 529932 560996 529984
rect 567936 529932 567988 529984
rect 348884 529592 348936 529644
rect 480628 529592 480680 529644
rect 191288 529524 191340 529576
rect 405188 529524 405240 529576
rect 175096 529456 175148 529508
rect 421380 529456 421432 529508
rect 167552 529388 167604 529440
rect 419448 529388 419500 529440
rect 155684 529320 155736 529372
rect 440792 529320 440844 529372
rect 149244 529252 149296 529304
rect 447232 529252 447284 529304
rect 144920 529184 144972 529236
rect 451556 529184 451608 529236
rect 140596 529116 140648 529168
rect 455880 529116 455932 529168
rect 136272 529048 136324 529100
rect 460526 529048 460578 529100
rect 134156 528980 134208 529032
rect 462642 528980 462694 529032
rect 120448 528912 120500 528964
rect 476304 528912 476356 528964
rect 117136 528844 117188 528896
rect 479616 528844 479668 528896
rect 114008 528776 114060 528828
rect 483020 528776 483072 528828
rect 110696 528708 110748 528760
rect 398840 528708 398892 528760
rect 399208 528708 399260 528760
rect 486056 528708 486108 528760
rect 108672 528640 108724 528692
rect 398932 528640 398984 528692
rect 403624 528640 403676 528692
rect 488356 528640 488408 528692
rect 107568 528572 107620 528624
rect 251916 528504 251968 528556
rect 254216 528504 254268 528556
rect 315396 528504 315448 528556
rect 319628 528504 319680 528556
rect 153936 528368 153988 528420
rect 159364 528368 159416 528420
rect 175188 528368 175240 528420
rect 144184 528164 144236 528216
rect 151728 528164 151780 528216
rect 162768 528232 162820 528284
rect 175188 528232 175240 528284
rect 159364 528164 159416 528216
rect 160376 528164 160428 528216
rect 175924 528164 175976 528216
rect 182180 528232 182232 528284
rect 177948 528164 178000 528216
rect 184204 528436 184256 528488
rect 195428 528436 195480 528488
rect 198004 528436 198056 528488
rect 234160 528436 234212 528488
rect 235080 528436 235132 528488
rect 262220 528436 262272 528488
rect 263048 528436 263100 528488
rect 318064 528436 318116 528488
rect 322020 528436 322072 528488
rect 190368 528368 190420 528420
rect 251824 528368 251876 528420
rect 253848 528368 253900 528420
rect 324136 528368 324188 528420
rect 324228 528368 324280 528420
rect 385684 528368 385736 528420
rect 184112 528300 184164 528352
rect 185952 528300 186004 528352
rect 385776 528300 385828 528352
rect 183928 528232 183980 528284
rect 315212 528232 315264 528284
rect 319628 528232 319680 528284
rect 323952 528232 324004 528284
rect 324228 528232 324280 528284
rect 385960 528232 386012 528284
rect 184112 528164 184164 528216
rect 184204 528164 184256 528216
rect 195428 528164 195480 528216
rect 198004 528164 198056 528216
rect 207020 528164 207072 528216
rect 207572 528164 207624 528216
rect 234160 528164 234212 528216
rect 235080 528164 235132 528216
rect 251824 528164 251876 528216
rect 251916 528164 251968 528216
rect 254216 528164 254268 528216
rect 254308 528164 254360 528216
rect 262220 528164 262272 528216
rect 263048 528164 263100 528216
rect 315396 528164 315448 528216
rect 320088 528164 320140 528216
rect 322020 528164 322072 528216
rect 324136 528164 324188 528216
rect 385408 528164 385460 528216
rect 385868 528164 385920 528216
rect 318064 528096 318116 528148
rect 302148 528028 302200 528080
rect 398840 528504 398892 528556
rect 411260 528572 411312 528624
rect 411444 528572 411496 528624
rect 489276 528572 489328 528624
rect 398932 528436 398984 528488
rect 403624 528436 403676 528488
rect 403716 528436 403768 528488
rect 408224 528436 408276 528488
rect 386236 528368 386288 528420
rect 406292 528368 406344 528420
rect 422300 528368 422352 528420
rect 431868 528368 431920 528420
rect 434720 528368 434772 528420
rect 434812 528368 434864 528420
rect 443368 528436 443420 528488
rect 386328 528300 386380 528352
rect 414940 528300 414992 528352
rect 422208 528300 422260 528352
rect 386512 528232 386564 528284
rect 434260 528232 434312 528284
rect 386420 528164 386472 528216
rect 387340 528164 387392 528216
rect 436468 528164 436520 528216
rect 442816 528164 442868 528216
rect 443368 528164 443420 528216
rect 444932 528164 444984 528216
rect 452752 528164 452804 528216
rect 282828 527960 282880 528012
rect 302240 527960 302292 528012
rect 278688 527892 278740 527944
rect 288532 527892 288584 527944
rect 288532 527756 288584 527808
rect 302148 527824 302200 527876
rect 302424 527960 302476 528012
rect 315304 527824 315356 527876
rect 282828 527484 282880 527536
rect 278688 527348 278740 527400
rect 282828 527076 282880 527128
rect 283104 527076 283156 527128
rect 283012 511980 283064 512032
rect 283104 511980 283156 512032
rect 2872 509260 2924 509312
rect 15844 509260 15896 509312
rect 416596 503004 416648 503056
rect 418160 503004 418212 503056
rect 418804 503004 418856 503056
rect 420276 503004 420328 503056
rect 574008 503004 574060 503056
rect 580448 503004 580500 503056
rect 412088 502936 412140 502988
rect 580356 502936 580408 502988
rect 481272 502868 481324 502920
rect 484308 502868 484360 502920
rect 487160 502868 487212 502920
rect 459468 502664 459520 502716
rect 461216 502664 461268 502716
rect 282920 502324 282972 502376
rect 283196 502324 283248 502376
rect 573364 502324 573416 502376
rect 574008 502324 574060 502376
rect 417424 501576 417476 501628
rect 580540 501576 580592 501628
rect 173900 501168 173952 501220
rect 174820 501168 174872 501220
rect 183652 501168 183704 501220
rect 184572 501168 184624 501220
rect 561680 501168 561732 501220
rect 562600 501168 562652 501220
rect 27528 500896 27580 500948
rect 29644 500896 29696 500948
rect 31668 500896 31720 500948
rect 31760 500896 31812 500948
rect 51172 500896 51224 500948
rect 52368 500896 52420 500948
rect 55496 500896 55548 500948
rect 56508 500896 56560 500948
rect 95424 500896 95476 500948
rect 96436 500896 96488 500948
rect 99656 500896 99708 500948
rect 100668 500896 100720 500948
rect 100760 500896 100812 500948
rect 102048 500896 102100 500948
rect 103980 500896 104032 500948
rect 104808 500896 104860 500948
rect 105084 500896 105136 500948
rect 106924 500896 106976 500948
rect 136272 500896 136324 500948
rect 153660 500896 153712 500948
rect 194600 500896 194652 500948
rect 195612 500896 195664 500948
rect 201500 500896 201552 500948
rect 203156 500896 203208 500948
rect 204904 500896 204956 500948
rect 208492 500896 208544 500948
rect 213828 500896 213880 500948
rect 216036 500896 216088 500948
rect 223488 500896 223540 500948
rect 224684 500896 224736 500948
rect 229100 500896 229152 500948
rect 230112 500896 230164 500948
rect 233056 500896 233108 500948
rect 234344 500896 234396 500948
rect 235908 500896 235960 500948
rect 236552 500896 236604 500948
rect 251180 500896 251232 500948
rect 253756 500896 253808 500948
rect 253940 500896 253992 500948
rect 255964 500896 256016 500948
rect 262220 500896 262272 500948
rect 263508 500896 263560 500948
rect 263600 500896 263652 500948
rect 264520 500896 264572 500948
rect 269120 500896 269172 500948
rect 269948 500896 270000 500948
rect 271972 500896 272024 500948
rect 273168 500896 273220 500948
rect 277584 500896 277636 500948
rect 278596 500896 278648 500948
rect 317328 500896 317380 500948
rect 317880 500896 317932 500948
rect 340144 500896 340196 500948
rect 340788 500896 340840 500948
rect 341156 500896 341208 500948
rect 342076 500896 342128 500948
rect 343180 500896 343232 500948
rect 343732 500896 343784 500948
rect 345480 500896 345532 500948
rect 346216 500896 346268 500948
rect 349804 500896 349856 500948
rect 350448 500896 350500 500948
rect 350908 500896 350960 500948
rect 351828 500896 351880 500948
rect 354128 500896 354180 500948
rect 354588 500896 354640 500948
rect 359464 500896 359516 500948
rect 360108 500896 360160 500948
rect 364892 500896 364944 500948
rect 365628 500896 365680 500948
rect 365996 500896 366048 500948
rect 367008 500896 367060 500948
rect 375656 500896 375708 500948
rect 376576 500896 376628 500948
rect 379980 500896 380032 500948
rect 380716 500896 380768 500948
rect 384304 500896 384356 500948
rect 384948 500896 385000 500948
rect 385408 500896 385460 500948
rect 386328 500896 386380 500948
rect 400496 500896 400548 500948
rect 401508 500896 401560 500948
rect 404728 500896 404780 500948
rect 411628 500896 411680 500948
rect 420828 500896 420880 500948
rect 423128 500896 423180 500948
rect 424968 500896 425020 500948
rect 427084 500896 427136 500948
rect 429292 500896 429344 500948
rect 431408 500896 431460 500948
rect 433432 500896 433484 500948
rect 435548 500896 435600 500948
rect 437572 500896 437624 500948
rect 439688 500896 439740 500948
rect 441988 500896 442040 500948
rect 444380 500896 444432 500948
rect 446312 500896 446364 500948
rect 448520 500896 448572 500948
rect 450452 500896 450504 500948
rect 453304 500896 453356 500948
rect 455328 500896 455380 500948
rect 457352 500896 457404 500948
rect 461860 500896 461912 500948
rect 464068 500896 464120 500948
rect 465908 500896 465960 500948
rect 468116 500896 468168 500948
rect 470232 500896 470284 500948
rect 472716 500896 472768 500948
rect 474648 500896 474700 500948
rect 477776 500896 477828 500948
rect 480812 500896 480864 500948
rect 502892 500896 502944 500948
rect 503628 500896 503680 500948
rect 511448 500896 511500 500948
rect 511908 500896 511960 500948
rect 516876 500896 516928 500948
rect 517428 500896 517480 500948
rect 523316 500896 523368 500948
rect 524328 500896 524380 500948
rect 545948 500896 546000 500948
rect 552112 500896 552164 500948
rect 552388 500896 552440 500948
rect 553492 500896 553544 500948
rect 45744 500828 45796 500880
rect 53932 500828 53984 500880
rect 95332 500828 95384 500880
rect 96528 500828 96580 500880
rect 137376 500828 137428 500880
rect 155132 500828 155184 500880
rect 195060 500828 195112 500880
rect 197728 500828 197780 500880
rect 205640 500828 205692 500880
rect 209596 500828 209648 500880
rect 214656 500828 214708 500880
rect 217140 500828 217192 500880
rect 403716 500828 403768 500880
rect 409880 500828 409932 500880
rect 543648 500828 543700 500880
rect 553768 500828 553820 500880
rect 80060 500760 80112 500812
rect 81348 500760 81400 500812
rect 134156 500760 134208 500812
rect 153844 500760 153896 500812
rect 191840 500760 191892 500812
rect 199936 500760 199988 500812
rect 267740 500760 267792 500812
rect 268844 500760 268896 500812
rect 355232 500760 355284 500812
rect 355968 500760 356020 500812
rect 541624 500760 541676 500812
rect 553860 500760 553912 500812
rect 41420 500692 41472 500744
rect 47032 500692 47084 500744
rect 135260 500692 135312 500744
rect 155316 500692 155368 500744
rect 224868 500692 224920 500744
rect 225788 500692 225840 500744
rect 230480 500692 230532 500744
rect 232228 500692 232280 500744
rect 320272 500692 320324 500744
rect 321100 500692 321152 500744
rect 539508 500692 539560 500744
rect 552020 500692 552072 500744
rect 552112 500692 552164 500744
rect 553676 500692 553728 500744
rect 131948 500624 132000 500676
rect 155500 500624 155552 500676
rect 191932 500624 191984 500676
rect 196624 500624 196676 500676
rect 197176 500624 197228 500676
rect 202052 500624 202104 500676
rect 258264 500624 258316 500676
rect 260288 500624 260340 500676
rect 260840 500624 260892 500676
rect 262404 500624 262456 500676
rect 360568 500624 360620 500676
rect 361396 500624 361448 500676
rect 370320 500624 370372 500676
rect 371056 500624 371108 500676
rect 512552 500624 512604 500676
rect 513288 500624 513340 500676
rect 513656 500624 513708 500676
rect 514668 500624 514720 500676
rect 537300 500624 537352 500676
rect 553952 500624 554004 500676
rect 129832 500556 129884 500608
rect 154764 500556 154816 500608
rect 201592 500556 201644 500608
rect 206376 500556 206428 500608
rect 207112 500556 207164 500608
rect 211712 500556 211764 500608
rect 215392 500556 215444 500608
rect 219256 500556 219308 500608
rect 219532 500556 219584 500608
rect 222568 500556 222620 500608
rect 535184 500556 535236 500608
rect 554044 500556 554096 500608
rect 20628 500488 20680 500540
rect 25320 500488 25372 500540
rect 97540 500488 97592 500540
rect 115204 500488 115256 500540
rect 127716 500488 127768 500540
rect 154856 500488 154908 500540
rect 196440 500488 196492 500540
rect 200948 500488 201000 500540
rect 257528 500488 257580 500540
rect 259184 500488 259236 500540
rect 363788 500488 363840 500540
rect 364248 500488 364300 500540
rect 369216 500488 369268 500540
rect 369768 500488 369820 500540
rect 531964 500488 532016 500540
rect 532608 500488 532660 500540
rect 533068 500488 533120 500540
rect 551192 500488 551244 500540
rect 551376 500488 551428 500540
rect 551928 500488 551980 500540
rect 22100 500420 22152 500472
rect 23388 500420 23440 500472
rect 42524 500420 42576 500472
rect 47584 500420 47636 500472
rect 93216 500420 93268 500472
rect 113824 500420 113876 500472
rect 125508 500420 125560 500472
rect 155224 500420 155276 500472
rect 187424 500420 187476 500472
rect 192392 500420 192444 500472
rect 203892 500420 203944 500472
rect 207480 500420 207532 500472
rect 211160 500420 211212 500472
rect 215024 500420 215076 500472
rect 218152 500420 218204 500472
rect 221464 500420 221516 500472
rect 224224 500420 224276 500472
rect 226800 500420 226852 500472
rect 528468 500420 528520 500472
rect 43628 500352 43680 500404
rect 48964 500352 49016 500404
rect 88892 500352 88944 500404
rect 112444 500352 112496 500404
rect 123392 500352 123444 500404
rect 154948 500352 155000 500404
rect 187608 500352 187660 500404
rect 193404 500352 193456 500404
rect 209136 500352 209188 500404
rect 212816 500352 212868 500404
rect 215208 500352 215260 500404
rect 218244 500352 218296 500404
rect 322848 500352 322900 500404
rect 323308 500352 323360 500404
rect 398288 500352 398340 500404
rect 398748 500352 398800 500404
rect 497464 500352 497516 500404
rect 498108 500352 498160 500404
rect 507124 500352 507176 500404
rect 507768 500352 507820 500404
rect 526536 500352 526588 500404
rect 551284 500352 551336 500404
rect 551376 500352 551428 500404
rect 44732 500284 44784 500336
rect 52552 500284 52604 500336
rect 84568 500284 84620 500336
rect 109684 500284 109736 500336
rect 121184 500284 121236 500336
rect 153292 500284 153344 500336
rect 195888 500284 195940 500336
rect 198832 500284 198884 500336
rect 199476 500284 199528 500336
rect 204168 500284 204220 500336
rect 209872 500284 209924 500336
rect 213920 500284 213972 500336
rect 255320 500284 255372 500336
rect 256976 500284 257028 500336
rect 524236 500284 524288 500336
rect 547972 500284 548024 500336
rect 555056 500352 555108 500404
rect 80244 500216 80296 500268
rect 108304 500216 108356 500268
rect 120172 500216 120224 500268
rect 153384 500216 153436 500268
rect 187516 500216 187568 500268
rect 194508 500216 194560 500268
rect 259460 500216 259512 500268
rect 261300 500216 261352 500268
rect 289728 500216 289780 500268
rect 416136 500216 416188 500268
rect 498568 500216 498620 500268
rect 499488 500216 499540 500268
rect 522212 500216 522264 500268
rect 553308 500284 553360 500336
rect 554228 500284 554280 500336
rect 548156 500216 548208 500268
rect 553584 500216 553636 500268
rect 556804 500216 556856 500268
rect 571340 500216 571392 500268
rect 61936 500148 61988 500200
rect 138480 500148 138532 500200
rect 146852 500148 146904 500200
rect 527640 500148 527692 500200
rect 528468 500148 528520 500200
rect 536288 500148 536340 500200
rect 536748 500148 536800 500200
rect 547052 500148 547104 500200
rect 552664 500148 552716 500200
rect 80244 500080 80296 500132
rect 139492 500080 139544 500132
rect 155040 500080 155092 500132
rect 220820 500080 220872 500132
rect 223580 500080 223632 500132
rect 547972 500080 548024 500132
rect 554964 500080 555016 500132
rect 140596 500012 140648 500064
rect 153752 500012 153804 500064
rect 551192 500012 551244 500064
rect 555424 500012 555476 500064
rect 142804 499944 142856 499996
rect 154028 499944 154080 499996
rect 223580 499944 223632 499996
rect 229008 499944 229060 499996
rect 374552 499944 374604 499996
rect 375288 499944 375340 499996
rect 378876 499944 378928 499996
rect 379428 499944 379480 499996
rect 389640 499944 389692 499996
rect 390468 499944 390520 499996
rect 393964 499944 394016 499996
rect 394608 499944 394660 499996
rect 395068 499944 395120 499996
rect 395896 499944 395948 499996
rect 399392 499944 399444 499996
rect 400128 499944 400180 499996
rect 501788 499944 501840 499996
rect 502248 499944 502300 499996
rect 388628 499876 388680 499928
rect 389088 499876 389140 499928
rect 92112 499808 92164 499860
rect 93768 499808 93820 499860
rect 344376 499808 344428 499860
rect 344928 499808 344980 499860
rect 50068 499740 50120 499792
rect 50988 499740 51040 499792
rect 144920 499740 144972 499792
rect 153936 499740 153988 499792
rect 200120 499740 200172 499792
rect 205272 499740 205324 499792
rect 234528 499740 234580 499792
rect 235448 499740 235500 499792
rect 206376 499672 206428 499724
rect 210700 499672 210752 499724
rect 216680 499604 216732 499656
rect 220360 499604 220412 499656
rect 252652 499604 252704 499656
rect 254860 499604 254912 499656
rect 24768 499536 24820 499588
rect 27436 499536 27488 499588
rect 32036 499536 32088 499588
rect 32864 499536 32916 499588
rect 34980 499536 35032 499588
rect 35808 499536 35860 499588
rect 36084 499536 36136 499588
rect 37188 499536 37240 499588
rect 40408 499536 40460 499588
rect 41328 499536 41380 499588
rect 60832 499536 60884 499588
rect 62028 499536 62080 499588
rect 65156 499536 65208 499588
rect 66168 499536 66220 499588
rect 69480 499536 69532 499588
rect 70308 499536 70360 499588
rect 71780 499536 71832 499588
rect 72700 499536 72752 499588
rect 75920 499536 75972 499588
rect 77208 499536 77260 499588
rect 247040 499536 247092 499588
rect 249432 499536 249484 499588
rect 256792 499536 256844 499588
rect 258080 499536 258132 499588
rect 266544 499536 266596 499588
rect 267832 499536 267884 499588
rect 560944 499536 560996 499588
rect 567200 499536 567252 499588
rect 164240 499128 164292 499180
rect 165068 499128 165120 499180
rect 80060 498856 80112 498908
rect 113180 498856 113232 498908
rect 66260 498788 66312 498840
rect 88340 498788 88392 498840
rect 89812 498788 89864 498840
rect 126980 498788 127032 498840
rect 194600 498788 194652 498840
rect 280160 498788 280212 498840
rect 501604 498788 501656 498840
rect 574100 498788 574152 498840
rect 104900 498108 104952 498160
rect 153200 498108 153252 498160
rect 132500 497632 132552 497684
rect 157432 497632 157484 497684
rect 70584 497564 70636 497616
rect 95240 497564 95292 497616
rect 121460 497564 121512 497616
rect 155592 497564 155644 497616
rect 82820 497496 82872 497548
rect 115940 497496 115992 497548
rect 118700 497496 118752 497548
rect 153476 497496 153528 497548
rect 93860 497428 93912 497480
rect 133880 497428 133932 497480
rect 299388 496068 299440 496120
rect 414020 496068 414072 496120
rect 3516 495456 3568 495508
rect 298100 495456 298152 495508
rect 299388 495456 299440 495508
rect 571340 495456 571392 495508
rect 573456 495456 573508 495508
rect 74540 494844 74592 494896
rect 102140 494844 102192 494896
rect 85672 494776 85724 494828
rect 120080 494776 120132 494828
rect 63500 494708 63552 494760
rect 84200 494708 84252 494760
rect 95424 494708 95476 494760
rect 138664 494708 138716 494760
rect 194508 493960 194560 494012
rect 197176 493960 197228 494012
rect 202880 493960 202932 494012
rect 205640 493960 205692 494012
rect 208860 493960 208912 494012
rect 211160 493960 211212 494012
rect 213644 493960 213696 494012
rect 215392 493960 215444 494012
rect 218428 493960 218480 494012
rect 220820 493960 220872 494012
rect 235172 493960 235224 494012
rect 237564 493960 237616 494012
rect 241152 493960 241204 494012
rect 243084 493960 243136 494012
rect 245936 493960 245988 494012
rect 248420 493960 248472 494012
rect 258264 493960 258316 494012
rect 259092 493960 259144 494012
rect 259460 493960 259512 494012
rect 260288 493960 260340 494012
rect 232780 493892 232832 493944
rect 235908 493892 235960 493944
rect 198096 493824 198148 493876
rect 200120 493824 200172 493876
rect 220820 493824 220872 493876
rect 224868 493824 224920 493876
rect 227996 493824 228048 493876
rect 230480 493824 230532 493876
rect 237564 493824 237616 493876
rect 240140 493824 240192 493876
rect 193312 493756 193364 493808
rect 196440 493756 196492 493808
rect 199292 493756 199344 493808
rect 201592 493756 201644 493808
rect 201684 493756 201736 493808
rect 204904 493756 204956 493808
rect 211252 493756 211304 493808
rect 214656 493756 214708 493808
rect 236368 493756 236420 493808
rect 238760 493756 238812 493808
rect 248328 493756 248380 493808
rect 249800 493892 249852 493944
rect 249524 493756 249576 493808
rect 251272 493756 251324 493808
rect 188620 493688 188672 493740
rect 191932 493688 191984 493740
rect 200488 493688 200540 493740
rect 203892 493688 203944 493740
rect 210056 493688 210108 493740
rect 213828 493688 213880 493740
rect 195704 493620 195756 493672
rect 201500 493620 201552 493672
rect 204076 493620 204128 493672
rect 206376 493620 206428 493672
rect 206468 493620 206520 493672
rect 209136 493620 209188 493672
rect 222016 493620 222068 493672
rect 224224 493620 224276 493672
rect 231584 493620 231636 493672
rect 234528 493620 234580 493672
rect 196900 493552 196952 493604
rect 199476 493552 199528 493604
rect 217232 493552 217284 493604
rect 219532 493552 219584 493604
rect 219624 493552 219676 493604
rect 223488 493552 223540 493604
rect 225604 493552 225656 493604
rect 229008 493552 229060 493604
rect 233976 493552 234028 493604
rect 237288 493552 237340 493604
rect 205272 493484 205324 493536
rect 207112 493484 207164 493536
rect 212448 493484 212500 493536
rect 215208 493484 215260 493536
rect 216036 493484 216088 493536
rect 218152 493484 218204 493536
rect 239956 493484 240008 493536
rect 242808 493484 242860 493536
rect 71780 493416 71832 493468
rect 98000 493416 98052 493468
rect 229192 493416 229244 493468
rect 233148 493416 233200 493468
rect 238760 493416 238812 493468
rect 241520 493416 241572 493468
rect 243544 493416 243596 493468
rect 245660 493416 245712 493468
rect 78680 493348 78732 493400
rect 109040 493348 109092 493400
rect 189724 493348 189776 493400
rect 195060 493348 195112 493400
rect 59360 493280 59412 493332
rect 77300 493280 77352 493332
rect 93768 493280 93820 493332
rect 131120 493280 131172 493332
rect 207664 493280 207716 493332
rect 209872 493280 209924 493332
rect 244740 493280 244792 493332
rect 247224 493280 247276 493332
rect 563704 493280 563756 493332
rect 571340 493280 571392 493332
rect 214840 493212 214892 493264
rect 216680 493212 216732 493264
rect 226800 493212 226852 493264
rect 230388 493212 230440 493264
rect 242348 493212 242400 493264
rect 244280 493212 244332 493264
rect 277584 493144 277636 493196
rect 279424 493144 279476 493196
rect 230388 493076 230440 493128
rect 233056 493076 233108 493128
rect 266452 493076 266504 493128
rect 267464 493076 267516 493128
rect 250720 492940 250772 492992
rect 252744 492940 252796 492992
rect 223212 492872 223264 492924
rect 227904 492872 227956 492924
rect 190920 492804 190972 492856
rect 195888 492804 195940 492856
rect 271972 492804 272024 492856
rect 273444 492804 273496 492856
rect 223580 492736 223632 492788
rect 224408 492736 224460 492788
rect 146024 492668 146076 492720
rect 154120 492668 154172 492720
rect 154304 492668 154356 492720
rect 154396 492668 154448 492720
rect 155684 492600 155736 492652
rect 156144 492600 156196 492652
rect 158904 492600 158956 492652
rect 158996 492600 159048 492652
rect 68928 492056 68980 492108
rect 92112 492056 92164 492108
rect 77116 491988 77168 492040
rect 106464 491988 106516 492040
rect 57888 491920 57940 491972
rect 74172 491920 74224 491972
rect 88248 491920 88300 491972
rect 124312 491920 124364 491972
rect 154304 491240 154356 491292
rect 154488 491240 154540 491292
rect 11704 490560 11756 490612
rect 443644 490560 443696 490612
rect 35808 489812 35860 489864
rect 36544 489812 36596 489864
rect 82728 489812 82780 489864
rect 115020 489812 115072 489864
rect 115204 489812 115256 489864
rect 140504 489812 140556 489864
rect 52368 489744 52420 489796
rect 63132 489744 63184 489796
rect 86868 489744 86920 489796
rect 122564 489744 122616 489796
rect 55128 489676 55180 489728
rect 68744 489676 68796 489728
rect 90916 489676 90968 489728
rect 129740 489676 129792 489728
rect 62028 489608 62080 489660
rect 79508 489608 79560 489660
rect 96528 489608 96580 489660
rect 136916 489608 136968 489660
rect 49608 489540 49660 489592
rect 59820 489540 59872 489592
rect 63408 489540 63460 489592
rect 83096 489540 83148 489592
rect 100668 489540 100720 489592
rect 144092 489540 144144 489592
rect 22192 489472 22244 489524
rect 26332 489472 26384 489524
rect 50988 489472 51040 489524
rect 61660 489472 61712 489524
rect 66168 489472 66220 489524
rect 86684 489472 86736 489524
rect 99288 489472 99340 489524
rect 142252 489472 142304 489524
rect 53748 489404 53800 489456
rect 66996 489404 67048 489456
rect 67456 489404 67508 489456
rect 90272 489404 90324 489456
rect 102048 489404 102100 489456
rect 145840 489404 145892 489456
rect 25780 489336 25832 489388
rect 27620 489336 27672 489388
rect 52276 489336 52328 489388
rect 65156 489336 65208 489388
rect 70308 489336 70360 489388
rect 93860 489336 93912 489388
rect 106924 489336 106976 489388
rect 153016 489336 153068 489388
rect 48228 489268 48280 489320
rect 58072 489268 58124 489320
rect 59268 489268 59320 489320
rect 75920 489268 75972 489320
rect 77208 489268 77260 489320
rect 104624 489268 104676 489320
rect 104808 489268 104860 489320
rect 151268 489268 151320 489320
rect 37096 489200 37148 489252
rect 40132 489200 40184 489252
rect 56508 489200 56560 489252
rect 70584 489200 70636 489252
rect 71688 489200 71740 489252
rect 97448 489200 97500 489252
rect 103428 489200 103480 489252
rect 149428 489200 149480 489252
rect 37188 489132 37240 489184
rect 38292 489132 38344 489184
rect 46848 489132 46900 489184
rect 56232 489132 56284 489184
rect 56416 489132 56468 489184
rect 72332 489132 72384 489184
rect 74448 489132 74500 489184
rect 101036 489132 101088 489184
rect 101956 489132 102008 489184
rect 147680 489132 147732 489184
rect 78588 489064 78640 489116
rect 108212 489064 108264 489116
rect 113824 489064 113876 489116
rect 133328 489064 133380 489116
rect 112444 488996 112496 489048
rect 126152 488996 126204 489048
rect 109684 488928 109736 488980
rect 118976 488928 119028 488980
rect 39948 488656 40000 488708
rect 43720 488656 43772 488708
rect 18604 488588 18656 488640
rect 23572 488588 23624 488640
rect 38568 488588 38620 488640
rect 41880 488588 41932 488640
rect 48964 488588 49016 488640
rect 50896 488588 50948 488640
rect 16856 488520 16908 488572
rect 22284 488520 22336 488572
rect 23940 488520 23992 488572
rect 24768 488520 24820 488572
rect 29368 488520 29420 488572
rect 30288 488520 30340 488572
rect 41328 488520 41380 488572
rect 45468 488520 45520 488572
rect 47584 488520 47636 488572
rect 49056 488520 49108 488572
rect 108304 488520 108356 488572
rect 111800 488520 111852 488572
rect 23388 486412 23440 486464
rect 156052 486412 156104 486464
rect 283012 485800 283064 485852
rect 158904 485732 158956 485784
rect 158996 485732 159048 485784
rect 283104 485732 283156 485784
rect 3424 485052 3476 485104
rect 185584 485052 185636 485104
rect 283104 482944 283156 482996
rect 283288 482944 283340 482996
rect 560392 482808 560444 482860
rect 563704 482808 563756 482860
rect 154304 481652 154356 481704
rect 154488 481652 154540 481704
rect 3148 480224 3200 480276
rect 11704 480224 11756 480276
rect 183652 480224 183704 480276
rect 183836 480224 183888 480276
rect 559564 479476 559616 479528
rect 560392 479476 560444 479528
rect 344928 477436 344980 477488
rect 346032 477436 346084 477488
rect 353208 477436 353260 477488
rect 355784 477436 355836 477488
rect 362868 477436 362920 477488
rect 366732 477436 366784 477488
rect 369768 477436 369820 477488
rect 374092 477436 374144 477488
rect 354588 477368 354640 477420
rect 356980 477368 357032 477420
rect 390468 477300 390520 477352
rect 397276 477300 397328 477352
rect 382188 477164 382240 477216
rect 388720 477164 388772 477216
rect 391848 477164 391900 477216
rect 399760 477164 399812 477216
rect 400128 477164 400180 477216
rect 408316 477164 408368 477216
rect 393228 477096 393280 477148
rect 400956 477096 401008 477148
rect 401508 477096 401560 477148
rect 409512 477096 409564 477148
rect 531228 477096 531280 477148
rect 552756 477096 552808 477148
rect 364248 477028 364300 477080
rect 368020 477028 368072 477080
rect 375288 477028 375340 477080
rect 380164 477028 380216 477080
rect 386236 477028 386288 477080
rect 392492 477028 392544 477080
rect 395896 477028 395948 477080
rect 403440 477028 403492 477080
rect 521568 477028 521620 477080
rect 553216 477028 553268 477080
rect 361488 476960 361540 477012
rect 365536 476960 365588 477012
rect 372528 476960 372580 477012
rect 377772 476960 377824 477012
rect 395988 476960 396040 477012
rect 404636 476960 404688 477012
rect 518808 476960 518860 477012
rect 351828 476892 351880 476944
rect 353300 476892 353352 476944
rect 355876 476892 355928 476944
rect 359464 476892 359516 476944
rect 368388 476892 368440 476944
rect 372896 476892 372948 476944
rect 373908 476892 373960 476944
rect 378968 476892 379020 476944
rect 380808 476892 380860 476944
rect 387524 476892 387576 476944
rect 389088 476892 389140 476944
rect 396080 476892 396132 476944
rect 397368 476892 397420 476944
rect 405832 476892 405884 476944
rect 517428 476892 517480 476944
rect 547328 476892 547380 476944
rect 551928 476960 551980 477012
rect 554136 476960 554188 477012
rect 552112 476892 552164 476944
rect 316684 476824 316736 476876
rect 317328 476824 317380 476876
rect 317880 476824 317932 476876
rect 318708 476824 318760 476876
rect 319076 476824 319128 476876
rect 320088 476824 320140 476876
rect 332600 476824 332652 476876
rect 333796 476824 333848 476876
rect 335360 476824 335412 476876
rect 336188 476824 336240 476876
rect 336648 476824 336700 476876
rect 337476 476824 337528 476876
rect 342168 476824 342220 476876
rect 343548 476824 343600 476876
rect 346216 476824 346268 476876
rect 347228 476824 347280 476876
rect 350448 476824 350500 476876
rect 352104 476824 352156 476876
rect 355968 476824 356020 476876
rect 358176 476824 358228 476876
rect 358728 476824 358780 476876
rect 361856 476824 361908 476876
rect 371056 476824 371108 476876
rect 375288 476824 375340 476876
rect 376576 476824 376628 476876
rect 381452 476824 381504 476876
rect 386328 476824 386380 476876
rect 392400 476824 392452 476876
rect 392492 476824 392544 476876
rect 393688 476824 393740 476876
rect 398748 476824 398800 476876
rect 407120 476824 407172 476876
rect 514576 476824 514628 476876
rect 551928 476824 551980 476876
rect 351736 476756 351788 476808
rect 354588 476756 354640 476808
rect 383568 476756 383620 476808
rect 390008 476756 390060 476808
rect 390376 476756 390428 476808
rect 398564 476756 398616 476808
rect 401416 476756 401468 476808
rect 410708 476756 410760 476808
rect 510528 476756 510580 476808
rect 553124 476756 553176 476808
rect 361396 476688 361448 476740
rect 364340 476688 364392 476740
rect 371148 476688 371200 476740
rect 376576 476688 376628 476740
rect 394608 476688 394660 476740
rect 402244 476688 402296 476740
rect 365628 476620 365680 476672
rect 369216 476620 369268 476672
rect 333980 476552 334032 476604
rect 334992 476552 335044 476604
rect 349068 476552 349120 476604
rect 350908 476552 350960 476604
rect 357348 476552 357400 476604
rect 360660 476552 360712 476604
rect 366916 476552 366968 476604
rect 371608 476552 371660 476604
rect 547328 476552 547380 476604
rect 553308 476552 553360 476604
rect 360108 476484 360160 476536
rect 363052 476484 363104 476536
rect 331404 476416 331456 476468
rect 332508 476416 332560 476468
rect 378048 476416 378100 476468
rect 383844 476416 383896 476468
rect 387708 476416 387760 476468
rect 394884 476416 394936 476468
rect 347688 476348 347740 476400
rect 349620 476348 349672 476400
rect 367008 476348 367060 476400
rect 370412 476348 370464 476400
rect 379428 476348 379480 476400
rect 385132 476348 385184 476400
rect 346308 476280 346360 476332
rect 348424 476280 348476 476332
rect 552664 476280 552716 476332
rect 555240 476280 555292 476332
rect 380716 476212 380768 476264
rect 386328 476212 386380 476264
rect 376668 476144 376720 476196
rect 382648 476144 382700 476196
rect 384948 476144 385000 476196
rect 391204 476144 391256 476196
rect 158812 476076 158864 476128
rect 158996 476076 159048 476128
rect 538128 475736 538180 475788
rect 551744 475736 551796 475788
rect 536748 475668 536800 475720
rect 554320 475668 554372 475720
rect 532608 475600 532660 475652
rect 551652 475600 551704 475652
rect 528468 475532 528520 475584
rect 525708 475464 525760 475516
rect 549168 475532 549220 475584
rect 551560 475532 551612 475584
rect 524328 475396 524380 475448
rect 547420 475396 547472 475448
rect 552848 475464 552900 475516
rect 552940 475396 552992 475448
rect 499488 475328 499540 475380
rect 552572 475328 552624 475380
rect 499304 474716 499356 474768
rect 501604 474716 501656 474768
rect 547420 474512 547472 474564
rect 555332 474512 555384 474564
rect 545028 474444 545080 474496
rect 553400 474444 553452 474496
rect 540888 474376 540940 474428
rect 555608 474376 555660 474428
rect 533988 474308 534040 474360
rect 551836 474308 551888 474360
rect 529848 474240 529900 474292
rect 555792 474240 555844 474292
rect 516048 474172 516100 474224
rect 552664 474172 552716 474224
rect 514668 474104 514720 474156
rect 555884 474104 555936 474156
rect 511908 474036 511960 474088
rect 498108 473968 498160 474020
rect 552388 473968 552440 474020
rect 554688 474036 554740 474088
rect 555148 474036 555200 474088
rect 556068 473968 556120 474020
rect 481640 473696 481692 473748
rect 490656 473696 490708 473748
rect 520556 473628 520608 473680
rect 522672 473628 522724 473680
rect 505008 473560 505060 473612
rect 512644 473560 512696 473612
rect 520464 473560 520516 473612
rect 522856 473560 522908 473612
rect 154304 473492 154356 473544
rect 491852 473424 491904 473476
rect 493140 473424 493192 473476
rect 508504 473424 508556 473476
rect 154304 473356 154356 473408
rect 283012 473356 283064 473408
rect 283288 473356 283340 473408
rect 314660 473356 314712 473408
rect 315948 473356 316000 473408
rect 447784 473356 447836 473408
rect 155776 473288 155828 473340
rect 156144 473288 156196 473340
rect 158904 473288 158956 473340
rect 158996 473288 159048 473340
rect 283012 473220 283064 473272
rect 283196 473220 283248 473272
rect 520464 473424 520516 473476
rect 520556 473424 520608 473476
rect 520740 473424 520792 473476
rect 522672 473424 522724 473476
rect 522856 473424 522908 473476
rect 542912 473424 542964 473476
rect 551468 473288 551520 473340
rect 553032 472880 553084 472932
rect 552204 472812 552256 472864
rect 552112 472608 552164 472660
rect 553032 472540 553084 472592
rect 552112 472404 552164 472456
rect 551560 472268 551612 472320
rect 552112 472268 552164 472320
rect 551468 472200 551520 472252
rect 552204 472200 552256 472252
rect 551560 472132 551612 472184
rect 551744 472132 551796 472184
rect 154304 471928 154356 471980
rect 154488 471928 154540 471980
rect 551744 471996 551796 472048
rect 552756 471996 552808 472048
rect 555700 471928 555752 471980
rect 552756 471860 552808 471912
rect 553216 471860 553268 471912
rect 551652 471792 551704 471844
rect 552480 471724 552532 471776
rect 552940 471724 552992 471776
rect 552940 471520 552992 471572
rect 553032 471520 553084 471572
rect 551744 471180 551796 471232
rect 551836 470636 551888 470688
rect 552296 470636 552348 470688
rect 552388 469956 552440 470008
rect 552848 469956 552900 470008
rect 554872 469140 554924 469192
rect 555332 469140 555384 469192
rect 555332 469004 555384 469056
rect 555608 469004 555660 469056
rect 555608 468868 555660 468920
rect 555792 468868 555844 468920
rect 552940 468392 552992 468444
rect 553216 468392 553268 468444
rect 558552 467780 558604 467832
rect 559564 467780 559616 467832
rect 158996 466420 159048 466472
rect 552664 466420 552716 466472
rect 552756 466420 552808 466472
rect 158904 466352 158956 466404
rect 551744 466352 551796 466404
rect 552480 466352 552532 466404
rect 553124 466352 553176 466404
rect 551744 466148 551796 466200
rect 552664 463700 552716 463752
rect 552756 463700 552808 463752
rect 154304 462340 154356 462392
rect 154488 462340 154540 462392
rect 556896 462340 556948 462392
rect 558552 462340 558604 462392
rect 563704 462340 563756 462392
rect 580172 462340 580224 462392
rect 552388 461592 552440 461644
rect 552572 461592 552624 461644
rect 183652 460912 183704 460964
rect 183836 460912 183888 460964
rect 551836 460844 551888 460896
rect 553032 460844 553084 460896
rect 551744 460708 551796 460760
rect 552388 460708 552440 460760
rect 552388 460572 552440 460624
rect 553124 460572 553176 460624
rect 551744 459824 551796 459876
rect 551928 459824 551980 459876
rect 551744 459280 551796 459332
rect 552480 459280 552532 459332
rect 158812 456764 158864 456816
rect 158996 456764 159048 456816
rect 551744 456764 551796 456816
rect 552664 456764 552716 456816
rect 551744 456288 551796 456340
rect 552756 456288 552808 456340
rect 551744 454860 551796 454912
rect 552480 454860 552532 454912
rect 551744 454724 551796 454776
rect 553032 454724 553084 454776
rect 552020 454112 552072 454164
rect 552480 454112 552532 454164
rect 155776 453976 155828 454028
rect 155868 453976 155920 454028
rect 158904 453976 158956 454028
rect 158996 453976 159048 454028
rect 154304 452548 154356 452600
rect 154488 452548 154540 452600
rect 552204 452004 552256 452056
rect 552572 452004 552624 452056
rect 552204 451868 552256 451920
rect 552480 451868 552532 451920
rect 3424 451256 3476 451308
rect 11796 451256 11848 451308
rect 155868 447108 155920 447160
rect 155776 447040 155828 447092
rect 158996 447108 159048 447160
rect 282920 447108 282972 447160
rect 158904 447040 158956 447092
rect 283012 447040 283064 447092
rect 9128 444320 9180 444372
rect 12624 444320 12676 444372
rect 282736 444320 282788 444372
rect 283012 444320 283064 444372
rect 154304 442960 154356 443012
rect 154488 442960 154540 443012
rect 183652 441600 183704 441652
rect 183836 441600 183888 441652
rect 289636 438880 289688 438932
rect 313280 438880 313332 438932
rect 554872 438880 554924 438932
rect 556896 438880 556948 438932
rect 3516 437452 3568 437504
rect 13084 437452 13136 437504
rect 158812 437452 158864 437504
rect 158996 437452 159048 437504
rect 554780 437248 554832 437300
rect 557632 437248 557684 437300
rect 551744 436908 551796 436960
rect 554872 436908 554924 436960
rect 554780 436500 554832 436552
rect 557724 436500 557776 436552
rect 554872 436024 554924 436076
rect 560300 436024 560352 436076
rect 554780 435956 554832 436008
rect 558920 435956 558972 436008
rect 158904 434664 158956 434716
rect 158996 434664 159048 434716
rect 554872 434664 554924 434716
rect 561680 434664 561732 434716
rect 554780 434596 554832 434648
rect 561772 434596 561824 434648
rect 154304 433236 154356 433288
rect 154488 433236 154540 433288
rect 554872 433236 554924 433288
rect 564440 433236 564492 433288
rect 554780 433168 554832 433220
rect 563060 433168 563112 433220
rect 554964 431876 555016 431928
rect 567292 431876 567344 431928
rect 554780 431808 554832 431860
rect 565820 431808 565872 431860
rect 554872 431740 554924 431792
rect 560944 431740 560996 431792
rect 554872 430516 554924 430568
rect 569960 430516 570012 430568
rect 554780 430448 554832 430500
rect 568580 430448 568632 430500
rect 155776 429836 155828 429888
rect 156052 429836 156104 429888
rect 554780 429088 554832 429140
rect 571616 429088 571668 429140
rect 554872 428884 554924 428936
rect 556804 428884 556856 428936
rect 158996 427796 159048 427848
rect 282920 427796 282972 427848
rect 158904 427728 158956 427780
rect 283012 427728 283064 427780
rect 554780 427728 554832 427780
rect 572720 427728 572772 427780
rect 447784 426368 447836 426420
rect 499304 426368 499356 426420
rect 551468 426368 551520 426420
rect 155776 425144 155828 425196
rect 156052 425144 156104 425196
rect 155776 425008 155828 425060
rect 155868 425008 155920 425060
rect 3424 423648 3476 423700
rect 14464 423648 14516 423700
rect 154304 423648 154356 423700
rect 154488 423648 154540 423700
rect 183652 422288 183704 422340
rect 183836 422288 183888 422340
rect 281632 421540 281684 421592
rect 282184 421540 282236 421592
rect 292580 421540 292632 421592
rect 155868 418140 155920 418192
rect 158812 418140 158864 418192
rect 158996 418140 159048 418192
rect 155776 418072 155828 418124
rect 304356 415420 304408 415472
rect 580172 415420 580224 415472
rect 155868 415352 155920 415404
rect 156144 415352 156196 415404
rect 158904 415352 158956 415404
rect 159180 415352 159232 415404
rect 282920 415352 282972 415404
rect 283104 415352 283156 415404
rect 154304 413924 154356 413976
rect 154488 413924 154540 413976
rect 158996 405696 159048 405748
rect 159180 405696 159232 405748
rect 282920 405696 282972 405748
rect 283196 405696 283248 405748
rect 154304 404336 154356 404388
rect 154488 404336 154540 404388
rect 183652 402976 183704 403028
rect 183836 402976 183888 403028
rect 140688 401548 140740 401600
rect 153752 401548 153804 401600
rect 140596 401480 140648 401532
rect 155040 401480 155092 401532
rect 139308 401412 139360 401464
rect 154212 401412 154264 401464
rect 136548 401344 136600 401396
rect 153660 401344 153712 401396
rect 137928 401276 137980 401328
rect 155132 401276 155184 401328
rect 135168 401208 135220 401260
rect 153844 401208 153896 401260
rect 136456 401140 136508 401192
rect 155316 401140 155368 401192
rect 132408 401072 132460 401124
rect 155500 401072 155552 401124
rect 133788 401004 133840 401056
rect 157432 401004 157484 401056
rect 125416 400936 125468 400988
rect 155224 400936 155276 400988
rect 122748 400868 122800 400920
rect 155592 400868 155644 400920
rect 142068 400800 142120 400852
rect 153568 400800 153620 400852
rect 143448 400732 143500 400784
rect 154028 400732 154080 400784
rect 144828 400664 144880 400716
rect 155408 400664 155460 400716
rect 146208 400596 146260 400648
rect 154120 400596 154172 400648
rect 146116 400256 146168 400308
rect 153936 400256 153988 400308
rect 154120 394612 154172 394664
rect 154304 394612 154356 394664
rect 155776 394612 155828 394664
rect 155868 394612 155920 394664
rect 158812 386316 158864 386368
rect 158996 386316 159048 386368
rect 154120 385024 154172 385076
rect 154304 385024 154356 385076
rect 183652 383664 183704 383716
rect 183836 383664 183888 383716
rect 155868 379516 155920 379568
rect 155684 379448 155736 379500
rect 282184 377204 282236 377256
rect 284392 377204 284444 377256
rect 78588 376728 78640 376780
rect 186964 376728 187016 376780
rect 154120 375300 154172 375352
rect 154304 375300 154356 375352
rect 304448 368500 304500 368552
rect 580172 368500 580224 368552
rect 153844 365712 153896 365764
rect 154120 365712 154172 365764
rect 183652 364352 183704 364404
rect 183836 364352 183888 364404
rect 155500 362244 155552 362296
rect 155776 362244 155828 362296
rect 186964 360136 187016 360188
rect 282184 360136 282236 360188
rect 187424 357484 187476 357536
rect 191932 357484 191984 357536
rect 153844 357416 153896 357468
rect 153936 357416 153988 357468
rect 155500 357416 155552 357468
rect 155592 357416 155644 357468
rect 274640 356396 274692 356448
rect 275652 356396 275704 356448
rect 194416 355988 194468 356040
rect 198924 355988 198976 356040
rect 201408 355988 201460 356040
rect 206928 355988 206980 356040
rect 210332 355988 210384 356040
rect 214748 355988 214800 356040
rect 215208 355988 215260 356040
rect 218980 355988 219032 356040
rect 221280 355988 221332 356040
rect 222844 355988 222896 356040
rect 226156 355988 226208 356040
rect 226984 355988 227036 356040
rect 227444 355988 227496 356040
rect 228180 355988 228232 356040
rect 229836 355988 229888 356040
rect 230480 355988 230532 356040
rect 233148 355988 233200 356040
rect 233700 355988 233752 356040
rect 234528 355988 234580 356040
rect 235908 355988 235960 356040
rect 237196 355988 237248 356040
rect 238300 355988 238352 356040
rect 239588 355988 239640 356040
rect 240508 355988 240560 356040
rect 258080 355988 258132 356040
rect 258540 355988 258592 356040
rect 261576 355988 261628 356040
rect 262220 355988 262272 356040
rect 262680 355988 262732 356040
rect 263600 355988 263652 356040
rect 193128 355920 193180 355972
rect 199660 355920 199712 355972
rect 213828 355920 213880 355972
rect 218060 355920 218112 355972
rect 232320 355920 232372 355972
rect 234068 355920 234120 355972
rect 235816 355920 235868 355972
rect 237288 355920 237340 355972
rect 211528 355852 211580 355904
rect 215668 355852 215720 355904
rect 224868 355852 224920 355904
rect 227720 355852 227772 355904
rect 204168 355784 204220 355836
rect 209228 355784 209280 355836
rect 222108 355784 222160 355836
rect 225420 355784 225472 355836
rect 242072 355784 242124 355836
rect 242808 355784 242860 355836
rect 281448 355784 281500 355836
rect 281724 355784 281776 355836
rect 199292 355716 199344 355768
rect 204996 355716 205048 355768
rect 198096 355648 198148 355700
rect 203892 355648 203944 355700
rect 240876 355648 240928 355700
rect 241704 355648 241756 355700
rect 255320 355648 255372 355700
rect 256056 355648 256108 355700
rect 217600 355580 217652 355632
rect 221188 355580 221240 355632
rect 200488 355512 200540 355564
rect 206100 355512 206152 355564
rect 263416 355512 263468 355564
rect 264612 355512 264664 355564
rect 189540 355444 189592 355496
rect 196348 355444 196400 355496
rect 207848 355376 207900 355428
rect 212632 355376 212684 355428
rect 218888 355376 218940 355428
rect 222384 355376 222436 355428
rect 231032 355376 231084 355428
rect 233148 355376 233200 355428
rect 256700 355376 256752 355428
rect 257344 355376 257396 355428
rect 266084 355376 266136 355428
rect 267096 355376 267148 355428
rect 190368 355308 190420 355360
rect 197268 355308 197320 355360
rect 209044 355308 209096 355360
rect 214012 355308 214064 355360
rect 243268 355308 243320 355360
rect 243820 355308 243872 355360
rect 244096 355308 244148 355360
rect 244924 355308 244976 355360
rect 220084 355240 220136 355292
rect 223672 355240 223724 355292
rect 264888 355240 264940 355292
rect 265900 355240 265952 355292
rect 202788 355172 202840 355224
rect 208308 355172 208360 355224
rect 254124 355104 254176 355156
rect 254860 355104 254912 355156
rect 268200 355104 268252 355156
rect 269488 355104 269540 355156
rect 212356 354968 212408 355020
rect 216772 354968 216824 355020
rect 191748 354832 191800 354884
rect 194968 354832 195020 354884
rect 196808 354832 196860 354884
rect 201500 354832 201552 354884
rect 223396 354832 223448 354884
rect 226524 354832 226576 354884
rect 206652 354764 206704 354816
rect 211436 354764 211488 354816
rect 238392 354764 238444 354816
rect 239404 354764 239456 354816
rect 248052 354764 248104 354816
rect 248512 354764 248564 354816
rect 188344 354696 188396 354748
rect 193220 354696 193272 354748
rect 195612 354696 195664 354748
rect 201408 354696 201460 354748
rect 205364 354696 205416 354748
rect 210332 354696 210384 354748
rect 216404 354696 216456 354748
rect 220084 354696 220136 354748
rect 228640 354696 228692 354748
rect 230388 354696 230440 354748
rect 260564 354696 260616 354748
rect 261024 354696 261076 354748
rect 267096 354696 267148 354748
rect 268292 354696 268344 354748
rect 39948 354628 40000 354680
rect 50988 354628 51040 354680
rect 51448 354628 51500 354680
rect 63592 354628 63644 354680
rect 48320 354560 48372 354612
rect 59636 354560 59688 354612
rect 61568 354560 61620 354612
rect 70400 354560 70452 354612
rect 33508 354492 33560 354544
rect 38660 354492 38712 354544
rect 45008 354492 45060 354544
rect 56968 354492 57020 354544
rect 58624 354492 58676 354544
rect 68928 354492 68980 354544
rect 70860 354492 70912 354544
rect 80060 354492 80112 354544
rect 35624 354424 35676 354476
rect 40316 354424 40368 354476
rect 46480 354424 46532 354476
rect 58072 354424 58124 354476
rect 68008 354424 68060 354476
rect 80152 354424 80204 354476
rect 39304 354356 39356 354408
rect 49700 354356 49752 354408
rect 50712 354356 50764 354408
rect 62212 354356 62264 354408
rect 64788 354356 64840 354408
rect 79324 354356 79376 354408
rect 46848 354288 46900 354340
rect 58624 354288 58676 354340
rect 62028 354288 62080 354340
rect 78588 354288 78640 354340
rect 25596 354220 25648 354272
rect 29276 354220 29328 354272
rect 45468 354220 45520 354272
rect 57152 354220 57204 354272
rect 59268 354220 59320 354272
rect 77208 354220 77260 354272
rect 34244 354152 34296 354204
rect 39212 354152 39264 354204
rect 42708 354152 42760 354204
rect 55128 354152 55180 354204
rect 56508 354152 56560 354204
rect 76012 354152 76064 354204
rect 37832 354084 37884 354136
rect 42800 354084 42852 354136
rect 47860 354084 47912 354136
rect 59360 354084 59412 354136
rect 64420 354084 64472 354136
rect 87420 354084 87472 354136
rect 34980 354016 35032 354068
rect 40040 354016 40092 354068
rect 44088 354016 44140 354068
rect 57244 354016 57296 354068
rect 67272 354016 67324 354068
rect 91836 354016 91888 354068
rect 26148 353948 26200 354000
rect 30380 353948 30432 354000
rect 31668 353948 31720 354000
rect 36728 353948 36780 354000
rect 38384 353948 38436 354000
rect 48596 353948 48648 354000
rect 49332 353948 49384 354000
rect 64972 353948 65024 354000
rect 70124 353948 70176 354000
rect 96068 353948 96120 354000
rect 50068 353880 50120 353932
rect 62120 353880 62172 353932
rect 32772 353812 32824 353864
rect 37832 353812 37884 353864
rect 55772 353812 55824 353864
rect 67548 353812 67600 353864
rect 29920 353744 29972 353796
rect 35808 353744 35860 353796
rect 41328 353744 41380 353796
rect 53012 353744 53064 353796
rect 54300 353744 54352 353796
rect 63500 353744 63552 353796
rect 30288 353676 30340 353728
rect 34520 353676 34572 353728
rect 42156 353676 42208 353728
rect 54116 353676 54168 353728
rect 40684 353608 40736 353660
rect 51908 353608 51960 353660
rect 27068 353540 27120 353592
rect 31852 353540 31904 353592
rect 37096 353540 37148 353592
rect 42248 353540 42300 353592
rect 43536 353540 43588 353592
rect 56140 353540 56192 353592
rect 24768 353472 24820 353524
rect 28172 353472 28224 353524
rect 28908 353472 28960 353524
rect 34428 353472 34480 353524
rect 22008 353404 22060 353456
rect 23940 353404 23992 353456
rect 24216 353404 24268 353456
rect 27068 353404 27120 353456
rect 31392 353404 31444 353456
rect 37096 353404 37148 353456
rect 21272 353336 21324 353388
rect 22836 353336 22888 353388
rect 23388 353336 23440 353388
rect 26240 353336 26292 353388
rect 28448 353336 28500 353388
rect 33508 353336 33560 353388
rect 20628 353268 20680 353320
rect 22192 353268 22244 353320
rect 22744 353268 22796 353320
rect 25044 353268 25096 353320
rect 27528 353268 27580 353320
rect 32588 353268 32640 353320
rect 36360 353268 36412 353320
rect 41420 353268 41472 353320
rect 63500 353132 63552 353184
rect 72332 353132 72384 353184
rect 67548 353064 67600 353116
rect 74724 353064 74776 353116
rect 68928 352996 68980 353048
rect 78772 352996 78824 353048
rect 70400 352928 70452 352980
rect 83188 352928 83240 352980
rect 57060 352860 57112 352912
rect 76748 352860 76800 352912
rect 60096 352792 60148 352844
rect 80980 352792 81032 352844
rect 62948 352724 63000 352776
rect 85580 352724 85632 352776
rect 65800 352656 65852 352708
rect 89720 352656 89772 352708
rect 68744 352588 68796 352640
rect 94044 352588 94096 352640
rect 52920 352520 52972 352572
rect 70400 352520 70452 352572
rect 71596 352520 71648 352572
rect 98276 352520 98328 352572
rect 58072 351840 58124 351892
rect 60740 351840 60792 351892
rect 36728 351772 36780 351824
rect 39028 351772 39080 351824
rect 57796 351704 57848 351756
rect 77852 351840 77904 351892
rect 80060 351840 80112 351892
rect 97172 351840 97224 351892
rect 138848 351840 138900 351892
rect 139308 351840 139360 351892
rect 139768 351840 139820 351892
rect 140596 351840 140648 351892
rect 142988 351840 143040 351892
rect 143448 351840 143500 351892
rect 144184 351840 144236 351892
rect 144828 351840 144880 351892
rect 145288 351840 145340 351892
rect 146116 351840 146168 351892
rect 155960 351840 156012 351892
rect 156420 351840 156472 351892
rect 158812 351840 158864 351892
rect 159732 351840 159784 351892
rect 160100 351840 160152 351892
rect 160836 351840 160888 351892
rect 161480 351840 161532 351892
rect 161940 351840 161992 351892
rect 164240 351840 164292 351892
rect 165068 351840 165120 351892
rect 165620 351840 165672 351892
rect 166172 351840 166224 351892
rect 187516 351840 187568 351892
rect 194140 351840 194192 351892
rect 198924 351840 198976 351892
rect 200580 351840 200632 351892
rect 275744 351840 275796 351892
rect 277400 351840 277452 351892
rect 60648 351636 60700 351688
rect 82084 351772 82136 351824
rect 63408 351704 63460 351756
rect 86316 351704 86368 351756
rect 66168 351636 66220 351688
rect 90732 351636 90784 351688
rect 38660 351568 38712 351620
rect 41512 351568 41564 351620
rect 59636 351568 59688 351620
rect 63684 351568 63736 351620
rect 63776 351568 63828 351620
rect 66996 351568 67048 351620
rect 69388 351568 69440 351620
rect 95240 351568 95292 351620
rect 127992 351568 128044 351620
rect 34520 351500 34572 351552
rect 36820 351500 36872 351552
rect 37832 351500 37884 351552
rect 40132 351500 40184 351552
rect 73712 351500 73764 351552
rect 101404 351500 101456 351552
rect 123760 351500 123812 351552
rect 40316 351432 40368 351484
rect 44364 351432 44416 351484
rect 56968 351432 57020 351484
rect 58348 351432 58400 351484
rect 59360 351432 59412 351484
rect 62764 351432 62816 351484
rect 63592 351432 63644 351484
rect 68100 351432 68152 351484
rect 72240 351432 72292 351484
rect 99380 351432 99432 351484
rect 129096 351432 129148 351484
rect 129648 351432 129700 351484
rect 41420 351364 41472 351416
rect 43444 351364 43496 351416
rect 58624 351364 58676 351416
rect 61660 351364 61712 351416
rect 62212 351364 62264 351416
rect 63776 351364 63828 351416
rect 75184 351364 75236 351416
rect 103704 351364 103756 351416
rect 133328 351568 133380 351620
rect 133788 351568 133840 351620
rect 135536 351568 135588 351620
rect 136456 351568 136508 351620
rect 130200 351500 130252 351552
rect 154764 351500 154816 351552
rect 271328 351500 271380 351552
rect 273260 351500 273312 351552
rect 154856 351432 154908 351484
rect 169944 351432 169996 351484
rect 170404 351432 170456 351484
rect 171140 351432 171192 351484
rect 171600 351432 171652 351484
rect 175280 351432 175332 351484
rect 175924 351432 175976 351484
rect 176660 351432 176712 351484
rect 177120 351432 177172 351484
rect 179512 351432 179564 351484
rect 180156 351432 180208 351484
rect 180800 351432 180852 351484
rect 181260 351432 181312 351484
rect 184940 351432 184992 351484
rect 185492 351432 185544 351484
rect 194968 351432 195020 351484
rect 198740 351432 198792 351484
rect 269028 351432 269080 351484
rect 270500 351432 270552 351484
rect 273076 351432 273128 351484
rect 274640 351432 274692 351484
rect 278688 351432 278740 351484
rect 281448 351432 281500 351484
rect 154948 351364 155000 351416
rect 270224 351364 270276 351416
rect 271880 351364 271932 351416
rect 274548 351364 274600 351416
rect 276204 351364 276256 351416
rect 277768 351364 277820 351416
rect 280160 351364 280212 351416
rect 42800 351296 42852 351348
rect 47676 351296 47728 351348
rect 52184 351296 52236 351348
rect 69204 351296 69256 351348
rect 72976 351296 73028 351348
rect 100852 351296 100904 351348
rect 121368 351296 121420 351348
rect 153292 351296 153344 351348
rect 276664 351296 276716 351348
rect 278780 351296 278832 351348
rect 40040 351228 40092 351280
rect 43260 351228 43312 351280
rect 39212 351160 39264 351212
rect 42156 351160 42208 351212
rect 42248 351160 42300 351212
rect 46572 351228 46624 351280
rect 53656 351228 53708 351280
rect 71228 351228 71280 351280
rect 74448 351228 74500 351280
rect 102508 351228 102560 351280
rect 120448 351228 120500 351280
rect 153384 351228 153436 351280
rect 43444 351160 43496 351212
rect 45652 351160 45704 351212
rect 55036 351160 55088 351212
rect 73436 351160 73488 351212
rect 75828 351160 75880 351212
rect 104900 351160 104952 351212
rect 119344 351160 119396 351212
rect 153476 351160 153528 351212
rect 193220 351160 193272 351212
rect 195244 351160 195296 351212
rect 228180 351160 228232 351212
rect 229836 351160 229888 351212
rect 57152 351092 57204 351144
rect 59452 351092 59504 351144
rect 77208 351092 77260 351144
rect 80060 351092 80112 351144
rect 80152 351092 80204 351144
rect 92940 351092 92992 351144
rect 62120 351024 62172 351076
rect 66352 351024 66404 351076
rect 78588 351024 78640 351076
rect 84384 351024 84436 351076
rect 187608 351024 187660 351076
rect 193220 351024 193272 351076
rect 79324 350956 79376 351008
rect 88524 350956 88576 351008
rect 173900 350956 173952 351008
rect 174820 350956 174872 351008
rect 124680 350888 124732 350940
rect 125508 350888 125560 350940
rect 134432 350888 134484 350940
rect 135168 350888 135220 350940
rect 183652 350888 183704 350940
rect 184572 350888 184624 350940
rect 201500 350888 201552 350940
rect 202880 350888 202932 350940
rect 226984 350888 227036 350940
rect 228732 350888 228784 350940
rect 230480 350888 230532 350940
rect 231860 350888 231912 350940
rect 233700 350888 233752 350940
rect 235172 350888 235224 350940
rect 272432 350888 272484 350940
rect 274732 350888 274784 350940
rect 37096 350752 37148 350804
rect 37924 350752 37976 350804
rect 222844 350752 222896 350804
rect 224316 350752 224368 350804
rect 115756 350684 115808 350736
rect 149060 350684 149112 350736
rect 112904 350616 112956 350668
rect 146300 350616 146352 350668
rect 106188 350548 106240 350600
rect 153200 350548 153252 350600
rect 3148 336744 3200 336796
rect 6184 336744 6236 336796
rect 303620 327020 303672 327072
rect 417424 327020 417476 327072
rect 303620 325592 303672 325644
rect 563704 325592 563756 325644
rect 21364 323484 21416 323536
rect 22192 323484 22244 323536
rect 22192 321580 22244 321632
rect 303620 321580 303672 321632
rect 580172 321580 580224 321632
rect 26884 321512 26936 321564
rect 100760 321172 100812 321224
rect 106280 321172 106332 321224
rect 111524 321104 111576 321156
rect 117964 321104 118016 321156
rect 231768 321104 231820 321156
rect 235448 321104 235500 321156
rect 92112 321036 92164 321088
rect 96620 321036 96672 321088
rect 108304 321036 108356 321088
rect 115204 321036 115256 321088
rect 228272 321036 228324 321088
rect 232228 321036 232280 321088
rect 101772 320968 101824 321020
rect 106372 320968 106424 321020
rect 109316 320968 109368 321020
rect 119344 320968 119396 321020
rect 75920 320900 75972 320952
rect 78680 320900 78732 320952
rect 93216 320900 93268 320952
rect 98000 320900 98052 320952
rect 102876 320900 102928 320952
rect 108948 320900 109000 320952
rect 115848 320900 115900 320952
rect 126244 320900 126296 320952
rect 24768 320832 24820 320884
rect 26332 320832 26384 320884
rect 34888 320832 34940 320884
rect 35808 320832 35860 320884
rect 54392 320832 54444 320884
rect 55312 320832 55364 320884
rect 64052 320832 64104 320884
rect 64880 320832 64932 320884
rect 72700 320832 72752 320884
rect 74540 320832 74592 320884
rect 82452 320832 82504 320884
rect 85120 320832 85172 320884
rect 85672 320832 85724 320884
rect 89628 320832 89680 320884
rect 106096 320832 106148 320884
rect 121552 320832 121604 320884
rect 198740 320832 198792 320884
rect 202052 320832 202104 320884
rect 247408 320832 247460 320884
rect 249432 320832 249484 320884
rect 73804 320764 73856 320816
rect 75920 320764 75972 320816
rect 110420 320764 110472 320816
rect 113824 320764 113876 320816
rect 146024 320764 146076 320816
rect 152464 320764 152516 320816
rect 227076 320764 227128 320816
rect 231124 320764 231176 320816
rect 246120 320764 246172 320816
rect 248420 320764 248472 320816
rect 256516 320764 256568 320816
rect 258080 320764 258132 320816
rect 83464 320696 83516 320748
rect 85672 320696 85724 320748
rect 248328 320696 248380 320748
rect 250536 320696 250588 320748
rect 226248 320628 226300 320680
rect 230112 320628 230164 320680
rect 98552 320560 98604 320612
rect 103520 320560 103572 320612
rect 204260 320560 204312 320612
rect 206376 320560 206428 320612
rect 208400 320560 208452 320612
rect 210700 320560 210752 320612
rect 202880 320492 202932 320544
rect 205272 320492 205324 320544
rect 23296 320424 23348 320476
rect 25320 320424 25372 320476
rect 91008 320424 91060 320476
rect 95240 320424 95292 320476
rect 99656 320424 99708 320476
rect 104900 320424 104952 320476
rect 195980 320424 196032 320476
rect 198832 320424 198884 320476
rect 235448 320424 235500 320476
rect 238668 320424 238720 320476
rect 78128 320356 78180 320408
rect 81256 320356 81308 320408
rect 88892 320356 88944 320408
rect 92388 320356 92440 320408
rect 94228 320356 94280 320408
rect 99564 320356 99616 320408
rect 236644 320356 236696 320408
rect 239772 320356 239824 320408
rect 25320 320288 25372 320340
rect 27436 320288 27488 320340
rect 66260 320288 66312 320340
rect 67640 320288 67692 320340
rect 71596 320288 71648 320340
rect 73896 320288 73948 320340
rect 80244 320288 80296 320340
rect 83004 320288 83056 320340
rect 86684 320288 86736 320340
rect 91100 320288 91152 320340
rect 97540 320288 97592 320340
rect 102140 320288 102192 320340
rect 103980 320288 104032 320340
rect 109776 320288 109828 320340
rect 184848 320288 184900 320340
rect 186964 320288 187016 320340
rect 198832 320288 198884 320340
rect 200948 320288 201000 320340
rect 229284 320288 229336 320340
rect 233332 320288 233384 320340
rect 238668 320288 238720 320340
rect 241888 320288 241940 320340
rect 242624 320288 242676 320340
rect 245200 320288 245252 320340
rect 253388 320288 253440 320340
rect 254860 320288 254912 320340
rect 27712 320220 27764 320272
rect 29644 320220 29696 320272
rect 30288 320220 30340 320272
rect 31760 320220 31812 320272
rect 33692 320220 33744 320272
rect 34980 320220 35032 320272
rect 61936 320220 61988 320272
rect 63500 320220 63552 320272
rect 68376 320220 68428 320272
rect 70400 320220 70452 320272
rect 70584 320220 70636 320272
rect 73252 320220 73304 320272
rect 77024 320220 77076 320272
rect 79968 320220 80020 320272
rect 81348 320220 81400 320272
rect 82820 320220 82872 320272
rect 89996 320220 90048 320272
rect 92756 320220 92808 320272
rect 96436 320220 96488 320272
rect 100760 320220 100812 320272
rect 105084 320220 105136 320272
rect 110420 320220 110472 320272
rect 163228 320220 163280 320272
rect 167644 320220 167696 320272
rect 181536 320220 181588 320272
rect 184204 320220 184256 320272
rect 192484 320220 192536 320272
rect 196624 320220 196676 320272
rect 202144 320220 202196 320272
rect 204168 320220 204220 320272
rect 233148 320220 233200 320272
rect 236552 320220 236604 320272
rect 237840 320220 237892 320272
rect 240876 320220 240928 320272
rect 241428 320220 241480 320272
rect 244096 320220 244148 320272
rect 245016 320220 245068 320272
rect 247316 320220 247368 320272
rect 251088 320220 251140 320272
rect 252744 320220 252796 320272
rect 254584 320220 254636 320272
rect 255964 320220 256016 320272
rect 257988 320220 258040 320272
rect 259184 320220 259236 320272
rect 22008 320152 22060 320204
rect 24216 320152 24268 320204
rect 26516 320152 26568 320204
rect 28540 320152 28592 320204
rect 28908 320152 28960 320204
rect 30656 320152 30708 320204
rect 31668 320152 31720 320204
rect 32864 320152 32916 320204
rect 33048 320152 33100 320204
rect 33876 320152 33928 320204
rect 35900 320152 35952 320204
rect 37188 320152 37240 320204
rect 37280 320152 37332 320204
rect 38200 320152 38252 320204
rect 38568 320152 38620 320204
rect 39304 320152 39356 320204
rect 42524 320152 42576 320204
rect 42800 320152 42852 320204
rect 43628 320152 43680 320204
rect 46940 320152 46992 320204
rect 47952 320152 48004 320204
rect 59820 320152 59872 320204
rect 60740 320152 60792 320204
rect 60832 320152 60884 320204
rect 62120 320152 62172 320204
rect 63040 320152 63092 320204
rect 64328 320152 64380 320204
rect 65156 320152 65208 320204
rect 66260 320152 66312 320204
rect 67364 320152 67416 320204
rect 69020 320152 69072 320204
rect 69480 320152 69532 320204
rect 71780 320152 71832 320204
rect 74908 320152 74960 320204
rect 77300 320152 77352 320204
rect 79140 320152 79192 320204
rect 81624 320152 81676 320204
rect 84568 320152 84620 320204
rect 87696 320152 87748 320204
rect 87788 320152 87840 320204
rect 90180 320152 90232 320204
rect 95332 320152 95384 320204
rect 98736 320152 98788 320204
rect 107200 320152 107252 320204
rect 112444 320152 112496 320204
rect 114744 320152 114796 320204
rect 115848 320152 115900 320204
rect 119068 320152 119120 320204
rect 119988 320152 120040 320204
rect 120172 320152 120224 320204
rect 121276 320152 121328 320204
rect 124404 320152 124456 320204
rect 125508 320152 125560 320204
rect 128728 320152 128780 320204
rect 129648 320152 129700 320204
rect 129832 320152 129884 320204
rect 130936 320152 130988 320204
rect 133052 320152 133104 320204
rect 133788 320152 133840 320204
rect 134156 320152 134208 320204
rect 135168 320152 135220 320204
rect 135260 320152 135312 320204
rect 136456 320152 136508 320204
rect 138480 320152 138532 320204
rect 139308 320152 139360 320204
rect 139492 320152 139544 320204
rect 141424 320152 141476 320204
rect 143816 320152 143868 320204
rect 144828 320152 144880 320204
rect 144920 320152 144972 320204
rect 146208 320152 146260 320204
rect 148140 320152 148192 320204
rect 148968 320152 149020 320204
rect 149244 320152 149296 320204
rect 150256 320152 150308 320204
rect 153568 320152 153620 320204
rect 154488 320152 154540 320204
rect 154672 320152 154724 320204
rect 155868 320152 155920 320204
rect 157892 320152 157944 320204
rect 158628 320152 158680 320204
rect 158904 320152 158956 320204
rect 160008 320152 160060 320204
rect 164332 320152 164384 320204
rect 165436 320152 165488 320204
rect 168656 320152 168708 320204
rect 169668 320152 169720 320204
rect 169760 320152 169812 320204
rect 170956 320152 171008 320204
rect 172980 320152 173032 320204
rect 173808 320152 173860 320204
rect 173992 320152 174044 320204
rect 175188 320152 175240 320204
rect 178316 320152 178368 320204
rect 179328 320152 179380 320204
rect 179420 320152 179472 320204
rect 180616 320152 180668 320204
rect 182640 320152 182692 320204
rect 183468 320152 183520 320204
rect 183744 320152 183796 320204
rect 184848 320152 184900 320204
rect 197452 320152 197504 320204
rect 199936 320152 199988 320204
rect 201132 320152 201184 320204
rect 203156 320152 203208 320204
rect 207112 320152 207164 320204
rect 209596 320152 209648 320204
rect 219900 320152 219952 320204
rect 224684 320152 224736 320204
rect 224868 320152 224920 320204
rect 229008 320152 229060 320204
rect 230296 320152 230348 320204
rect 234344 320152 234396 320204
rect 234528 320152 234580 320204
rect 237656 320152 237708 320204
rect 240048 320152 240100 320204
rect 242992 320152 243044 320204
rect 243820 320152 243872 320204
rect 246212 320152 246264 320204
rect 249708 320152 249760 320204
rect 251640 320152 251692 320204
rect 252468 320152 252520 320204
rect 253756 320152 253808 320204
rect 255780 320152 255832 320204
rect 256976 320152 257028 320204
rect 259368 320152 259420 320204
rect 260288 320152 260340 320204
rect 41420 320084 41472 320136
rect 263508 320152 263560 320204
rect 263600 320152 263652 320204
rect 264520 320152 264572 320204
rect 267740 320152 267792 320204
rect 268844 320152 268896 320204
rect 269120 320152 269172 320204
rect 269948 320152 270000 320204
rect 262220 320016 262272 320068
rect 22100 319404 22152 319456
rect 113180 319404 113232 319456
rect 113640 319404 113692 319456
rect 128452 319404 128504 319456
rect 195612 319404 195664 319456
rect 280160 319404 280212 319456
rect 20628 318724 20680 318776
rect 23112 318724 23164 318776
rect 90180 318724 90232 318776
rect 92296 318724 92348 318776
rect 192392 318724 192444 318776
rect 197452 318724 197504 318776
rect 201960 318724 202012 318776
rect 208308 318724 208360 318776
rect 211528 318724 211580 318776
rect 217140 318724 217192 318776
rect 223488 318724 223540 318776
rect 227904 318724 227956 318776
rect 200764 318656 200816 318708
rect 206928 318656 206980 318708
rect 220636 318656 220688 318708
rect 225788 318656 225840 318708
rect 202788 318588 202840 318640
rect 207112 318588 207164 318640
rect 92388 318520 92440 318572
rect 93492 318520 93544 318572
rect 98736 318520 98788 318572
rect 100668 318520 100720 318572
rect 106372 318520 106424 318572
rect 107844 318520 107896 318572
rect 194508 318452 194560 318504
rect 198740 318452 198792 318504
rect 209136 318452 209188 318504
rect 215024 318452 215076 318504
rect 85120 318384 85172 318436
rect 86316 318384 86368 318436
rect 85672 318316 85724 318368
rect 87512 318316 87564 318368
rect 195888 318316 195940 318368
rect 201132 318316 201184 318368
rect 204168 318316 204220 318368
rect 208400 318316 208452 318368
rect 191196 318248 191248 318300
rect 195980 318248 196032 318300
rect 199568 318248 199620 318300
rect 204260 318248 204312 318300
rect 217508 318248 217560 318300
rect 222568 318248 222620 318300
rect 87696 318180 87748 318232
rect 88708 318180 88760 318232
rect 207940 318180 207992 318232
rect 213828 318180 213880 318232
rect 198372 318112 198424 318164
rect 202880 318112 202932 318164
rect 190000 318044 190052 318096
rect 197268 318044 197320 318096
rect 218704 318044 218756 318096
rect 223580 318044 223632 318096
rect 213828 317908 213880 317960
rect 219256 317908 219308 317960
rect 222016 317908 222068 317960
rect 226800 317908 226852 317960
rect 193588 317840 193640 317892
rect 198832 317840 198884 317892
rect 210332 317704 210384 317756
rect 216036 317704 216088 317756
rect 206744 317568 206796 317620
rect 212448 317568 212500 317620
rect 216312 317568 216364 317620
rect 221464 317568 221516 317620
rect 82820 317500 82872 317552
rect 85120 317500 85172 317552
rect 197176 317500 197228 317552
rect 202144 317500 202196 317552
rect 205548 317500 205600 317552
rect 211068 317500 211120 317552
rect 217968 317500 218020 317552
rect 92756 317432 92808 317484
rect 94688 317432 94740 317484
rect 188620 317432 188672 317484
rect 192484 317432 192536 317484
rect 212448 317432 212500 317484
rect 215116 317432 215168 317484
rect 220360 317432 220412 317484
rect 2780 316684 2832 316736
rect 3424 316684 3476 316736
rect 288900 316684 288952 316736
rect 26884 315324 26936 315376
rect 111800 315324 111852 315376
rect 15844 315256 15896 315308
rect 185584 315256 185636 315308
rect 111800 313624 111852 313676
rect 113548 313624 113600 313676
rect 303620 311856 303672 311908
rect 336004 311856 336056 311908
rect 113548 311584 113600 311636
rect 116584 311584 116636 311636
rect 303620 310496 303672 310548
rect 341524 310496 341576 310548
rect 303620 309136 303672 309188
rect 340144 309136 340196 309188
rect 303620 306348 303672 306400
rect 560944 306348 560996 306400
rect 282184 305600 282236 305652
rect 300860 305600 300912 305652
rect 296168 303560 296220 303612
rect 580356 303560 580408 303612
rect 3424 293972 3476 294024
rect 15844 293972 15896 294024
rect 11796 275952 11848 276004
rect 17132 275952 17184 276004
rect 304356 275952 304408 276004
rect 580172 275952 580224 276004
rect 117228 236648 117280 236700
rect 132500 236648 132552 236700
rect 113916 235900 113968 235952
rect 281540 235900 281592 235952
rect 180616 235220 180668 235272
rect 194600 235220 194652 235272
rect 10508 233860 10560 233912
rect 299480 233860 299532 233912
rect 146208 232500 146260 232552
rect 160100 232500 160152 232552
rect 227628 232500 227680 232552
rect 313924 232500 313976 232552
rect 143448 231072 143500 231124
rect 157524 231072 157576 231124
rect 166908 231072 166960 231124
rect 180892 231072 180944 231124
rect 214748 231072 214800 231124
rect 305644 231072 305696 231124
rect 140688 229712 140740 229764
rect 155960 229712 156012 229764
rect 159916 229712 159968 229764
rect 175280 229712 175332 229764
rect 214564 229712 214616 229764
rect 308404 229712 308456 229764
rect 304264 229032 304316 229084
rect 579988 229032 580040 229084
rect 139308 228352 139360 228404
rect 154304 228352 154356 228404
rect 155776 228352 155828 228404
rect 171416 228352 171468 228404
rect 175096 228352 175148 228404
rect 190644 228352 190696 228404
rect 214932 228352 214984 228404
rect 287704 228352 287756 228404
rect 135168 227060 135220 227112
rect 149980 227060 150032 227112
rect 162768 227060 162820 227112
rect 177764 227060 177816 227112
rect 15844 226992 15896 227044
rect 120080 226992 120132 227044
rect 121276 226992 121328 227044
rect 136088 226992 136140 227044
rect 147588 226992 147640 227044
rect 162860 226992 162912 227044
rect 214656 226992 214708 227044
rect 309784 226992 309836 227044
rect 14464 225564 14516 225616
rect 411996 225564 412048 225616
rect 119344 224884 119396 224936
rect 125416 224884 125468 224936
rect 125508 224884 125560 224936
rect 133696 224884 133748 224936
rect 133788 224884 133840 224936
rect 139400 224884 139452 224936
rect 144828 224884 144880 224936
rect 159640 224884 159692 224936
rect 160008 224884 160060 224936
rect 174636 224884 174688 224936
rect 176568 224884 176620 224936
rect 191748 224884 191800 224936
rect 115204 224816 115256 224868
rect 124312 224816 124364 224868
rect 130936 224816 130988 224868
rect 145748 224816 145800 224868
rect 152464 224816 152516 224868
rect 161756 224816 161808 224868
rect 169668 224816 169720 224868
rect 183836 224816 183888 224868
rect 184204 224816 184256 224868
rect 197084 224816 197136 224868
rect 119988 224748 120040 224800
rect 126152 224748 126204 224800
rect 126244 224748 126296 224800
rect 131764 224748 131816 224800
rect 136456 224748 136508 224800
rect 151084 224748 151136 224800
rect 154488 224748 154540 224800
rect 169208 224748 169260 224800
rect 172428 224748 172480 224800
rect 117964 224680 118016 224732
rect 127532 224680 127584 224732
rect 128268 224680 128320 224732
rect 143540 224680 143592 224732
rect 153108 224680 153160 224732
rect 168196 224680 168248 224732
rect 175188 224680 175240 224732
rect 184020 224680 184072 224732
rect 186964 224748 187016 224800
rect 200304 224748 200356 224800
rect 187424 224680 187476 224732
rect 115848 224612 115900 224664
rect 130752 224612 130804 224664
rect 132408 224612 132460 224664
rect 147864 224612 147916 224664
rect 148968 224612 149020 224664
rect 163872 224612 163924 224664
rect 177948 224612 178000 224664
rect 192760 224612 192812 224664
rect 113824 224544 113876 224596
rect 126428 224544 126480 224596
rect 126888 224544 126940 224596
rect 142528 224544 142580 224596
rect 150256 224544 150308 224596
rect 164976 224544 165028 224596
rect 165436 224544 165488 224596
rect 179972 224544 180024 224596
rect 184848 224544 184900 224596
rect 199200 224544 199252 224596
rect 113088 224476 113140 224528
rect 128636 224476 128688 224528
rect 131028 224476 131080 224528
rect 146760 224476 146812 224528
rect 151728 224476 151780 224528
rect 167092 224476 167144 224528
rect 168288 224476 168340 224528
rect 183192 224476 183244 224528
rect 183468 224476 183520 224528
rect 198096 224476 198148 224528
rect 118608 224408 118660 224460
rect 133972 224408 134024 224460
rect 136548 224408 136600 224460
rect 152096 224408 152148 224460
rect 155868 224408 155920 224460
rect 170312 224408 170364 224460
rect 170956 224408 171008 224460
rect 185308 224408 185360 224460
rect 186228 224408 186280 224460
rect 201316 224408 201368 224460
rect 121368 224340 121420 224392
rect 137192 224340 137244 224392
rect 137928 224340 137980 224392
rect 153200 224340 153252 224392
rect 165528 224340 165580 224392
rect 180984 224340 181036 224392
rect 187608 224340 187660 224392
rect 202420 224340 202472 224392
rect 122748 224272 122800 224324
rect 138204 224272 138256 224324
rect 142068 224272 142120 224324
rect 157432 224272 157484 224324
rect 161388 224272 161440 224324
rect 176752 224272 176804 224324
rect 180708 224272 180760 224324
rect 195980 224272 196032 224324
rect 112444 224204 112496 224256
rect 123208 224204 123260 224256
rect 125232 224204 125284 224256
rect 141424 224204 141476 224256
rect 150348 224204 150400 224256
rect 166080 224204 166132 224256
rect 171048 224204 171100 224256
rect 186320 224204 186372 224256
rect 188436 224204 188488 224256
rect 203432 224204 203484 224256
rect 210976 224204 211028 224256
rect 286324 224204 286376 224256
rect 126152 224068 126204 224120
rect 134984 224068 135036 224120
rect 124128 224000 124180 224052
rect 139308 224136 139360 224188
rect 139400 224136 139452 224188
rect 148876 224136 148928 224188
rect 158628 224136 158680 224188
rect 173532 224136 173584 224188
rect 173808 224136 173860 224188
rect 188528 224136 188580 224188
rect 129648 223932 129700 223984
rect 144644 224068 144696 224120
rect 157248 224068 157300 224120
rect 172428 224068 172480 224120
rect 179328 224068 179380 224120
rect 193864 224068 193916 224120
rect 141332 224000 141384 224052
rect 155316 224000 155368 224052
rect 167644 224000 167696 224052
rect 178868 224000 178920 224052
rect 184020 224000 184072 224052
rect 189540 224000 189592 224052
rect 133696 223864 133748 223916
rect 140320 223864 140372 223916
rect 229744 223592 229796 223644
rect 283380 223592 283432 223644
rect 13084 222844 13136 222896
rect 411904 222844 411956 222896
rect 231124 222436 231176 222488
rect 235264 222436 235316 222488
rect 120724 221484 120776 221536
rect 55220 220872 55272 220924
rect 116400 220872 116452 220924
rect 9128 220804 9180 220856
rect 215116 220804 215168 220856
rect 226340 220804 226392 220856
rect 215116 220124 215168 220176
rect 226432 220124 226484 220176
rect 11704 220056 11756 220108
rect 116676 220056 116728 220108
rect 215208 220056 215260 220108
rect 226340 220056 226392 220108
rect 104808 219376 104860 219428
rect 116124 219444 116176 219496
rect 215116 218764 215168 218816
rect 226340 218764 226392 218816
rect 215208 218696 215260 218748
rect 226432 218696 226484 218748
rect 104808 217948 104860 218000
rect 116400 218016 116452 218068
rect 215116 217268 215168 217320
rect 226340 217268 226392 217320
rect 104808 216588 104860 216640
rect 116400 216656 116452 216708
rect 215116 216588 215168 216640
rect 226432 216588 226484 216640
rect 104808 215908 104860 215960
rect 115940 215908 115992 215960
rect 215116 215908 215168 215960
rect 226340 215908 226392 215960
rect 104808 215228 104860 215280
rect 116400 215296 116452 215348
rect 215116 215228 215168 215280
rect 226432 215228 226484 215280
rect 215208 215160 215260 215212
rect 226340 215160 226392 215212
rect 104808 213868 104860 213920
rect 116400 213936 116452 213988
rect 215116 213868 215168 213920
rect 226432 213868 226484 213920
rect 214380 213800 214432 213852
rect 226340 213800 226392 213852
rect 104440 212440 104492 212492
rect 115940 212508 115992 212560
rect 215116 212440 215168 212492
rect 226432 212440 226484 212492
rect 215208 212372 215260 212424
rect 226340 212372 226392 212424
rect 104808 211080 104860 211132
rect 116308 211148 116360 211200
rect 214196 211080 214248 211132
rect 226524 211080 226576 211132
rect 104808 209720 104860 209772
rect 116308 209788 116360 209840
rect 215116 209720 215168 209772
rect 226156 209720 226208 209772
rect 214196 209652 214248 209704
rect 226248 209652 226300 209704
rect 104808 208292 104860 208344
rect 116032 208360 116084 208412
rect 215116 208292 215168 208344
rect 226064 208292 226116 208344
rect 214288 208224 214340 208276
rect 225972 208224 226024 208276
rect 113088 207068 113140 207120
rect 116032 207068 116084 207120
rect 104808 206864 104860 206916
rect 115940 207000 115992 207052
rect 215116 206932 215168 206984
rect 226064 206932 226116 206984
rect 214380 206864 214432 206916
rect 226248 206864 226300 206916
rect 104716 206796 104768 206848
rect 113088 206796 113140 206848
rect 104808 205572 104860 205624
rect 115940 205640 115992 205692
rect 215116 205572 215168 205624
rect 226156 205572 226208 205624
rect 104808 204212 104860 204264
rect 116400 204280 116452 204332
rect 215208 204212 215260 204264
rect 225972 204212 226024 204264
rect 215116 204144 215168 204196
rect 225880 204144 225932 204196
rect 104808 202784 104860 202836
rect 116308 202852 116360 202904
rect 214288 202784 214340 202836
rect 226064 202784 226116 202836
rect 215116 202716 215168 202768
rect 225788 202716 225840 202768
rect 104808 201424 104860 201476
rect 116124 201492 116176 201544
rect 214380 201424 214432 201476
rect 225604 201424 225656 201476
rect 215116 201356 215168 201408
rect 226064 201356 226116 201408
rect 104808 200064 104860 200116
rect 116124 200200 116176 200252
rect 113272 200132 113324 200184
rect 115940 200132 115992 200184
rect 214104 200064 214156 200116
rect 226248 200064 226300 200116
rect 224040 198772 224092 198824
rect 226432 198772 226484 198824
rect 113180 198704 113232 198756
rect 116400 198704 116452 198756
rect 224132 198704 224184 198756
rect 226340 198704 226392 198756
rect 104808 198636 104860 198688
rect 113272 198636 113324 198688
rect 215116 198636 215168 198688
rect 225972 198636 226024 198688
rect 214104 198568 214156 198620
rect 225696 198568 225748 198620
rect 223948 197412 224000 197464
rect 226432 197412 226484 197464
rect 104808 197276 104860 197328
rect 113088 197276 113140 197328
rect 104532 197208 104584 197260
rect 116400 197344 116452 197396
rect 224316 197344 224368 197396
rect 226340 197344 226392 197396
rect 214380 197276 214432 197328
rect 226156 197276 226208 197328
rect 215116 197208 215168 197260
rect 225880 197208 225932 197260
rect 224224 196052 224276 196104
rect 226616 196052 226668 196104
rect 104808 195916 104860 195968
rect 116400 195984 116452 196036
rect 224592 195984 224644 196036
rect 226708 195984 226760 196036
rect 215208 195916 215260 195968
rect 226064 195916 226116 195968
rect 215116 195848 215168 195900
rect 226248 195848 226300 195900
rect 104808 194488 104860 194540
rect 115940 194556 115992 194608
rect 224408 194556 224460 194608
rect 226340 194556 226392 194608
rect 215116 194488 215168 194540
rect 225788 194488 225840 194540
rect 220268 193264 220320 193316
rect 226432 193264 226484 193316
rect 104440 193128 104492 193180
rect 116124 193196 116176 193248
rect 215944 193196 215996 193248
rect 226340 193196 226392 193248
rect 215116 193128 215168 193180
rect 224040 193128 224092 193180
rect 215208 193060 215260 193112
rect 224132 193060 224184 193112
rect 113180 191972 113232 192024
rect 116400 191972 116452 192024
rect 113272 191904 113324 191956
rect 116032 191904 116084 191956
rect 224868 191904 224920 191956
rect 226432 191904 226484 191956
rect 218152 191836 218204 191888
rect 226340 191836 226392 191888
rect 104808 191768 104860 191820
rect 113180 191768 113232 191820
rect 214288 191768 214340 191820
rect 224316 191768 224368 191820
rect 215116 191700 215168 191752
rect 223948 191700 224000 191752
rect 215300 191088 215352 191140
rect 226616 191088 226668 191140
rect 221464 190884 221516 190936
rect 226340 190884 226392 190936
rect 113364 190612 113416 190664
rect 116492 190612 116544 190664
rect 222844 190476 222896 190528
rect 226340 190476 226392 190528
rect 104716 190408 104768 190460
rect 113272 190408 113324 190460
rect 214380 190408 214432 190460
rect 224592 190408 224644 190460
rect 215116 190340 215168 190392
rect 224224 190340 224276 190392
rect 218060 189728 218112 189780
rect 226984 189728 227036 189780
rect 114192 189048 114244 189100
rect 116400 189048 116452 189100
rect 220084 189048 220136 189100
rect 226340 189048 226392 189100
rect 104808 188980 104860 189032
rect 113364 188980 113416 189032
rect 214012 188980 214064 189032
rect 224408 188980 224460 189032
rect 221648 187756 221700 187808
rect 226432 187756 226484 187808
rect 113180 187688 113232 187740
rect 116216 187688 116268 187740
rect 216036 187688 216088 187740
rect 226340 187688 226392 187740
rect 104808 187620 104860 187672
rect 114192 187620 114244 187672
rect 215116 187552 215168 187604
rect 220268 187552 220320 187604
rect 215208 187144 215260 187196
rect 218060 187144 218112 187196
rect 218796 186464 218848 186516
rect 226340 186464 226392 186516
rect 104808 186260 104860 186312
rect 113088 186260 113140 186312
rect 104532 186192 104584 186244
rect 116308 186328 116360 186380
rect 220176 186328 220228 186380
rect 226340 186328 226392 186380
rect 214472 185648 214524 185700
rect 224868 185648 224920 185700
rect 215300 185580 215352 185632
rect 226524 185580 226576 185632
rect 213920 185512 213972 185564
rect 215944 185512 215996 185564
rect 114468 184968 114520 185020
rect 116400 184968 116452 185020
rect 104808 184832 104860 184884
rect 116032 184900 116084 184952
rect 224224 184900 224276 184952
rect 226340 184900 226392 184952
rect 227168 184832 227220 184884
rect 230848 184832 230900 184884
rect 214196 184764 214248 184816
rect 218152 184764 218204 184816
rect 224316 183608 224368 183660
rect 226524 183608 226576 183660
rect 114376 183540 114428 183592
rect 116400 183540 116452 183592
rect 215024 183540 215076 183592
rect 226340 183540 226392 183592
rect 104808 183472 104860 183524
rect 114468 183472 114520 183524
rect 215116 182520 215168 182572
rect 221464 182520 221516 182572
rect 222936 182248 222988 182300
rect 226524 182248 226576 182300
rect 113180 182180 113232 182232
rect 115940 182180 115992 182232
rect 214840 182180 214892 182232
rect 226340 182180 226392 182232
rect 104808 182112 104860 182164
rect 114376 182112 114428 182164
rect 214196 182112 214248 182164
rect 222844 182112 222896 182164
rect 336004 182112 336056 182164
rect 579988 182112 580040 182164
rect 218888 181432 218940 181484
rect 226432 181432 226484 181484
rect 113272 181092 113324 181144
rect 115940 181092 115992 181144
rect 221556 180888 221608 180940
rect 226340 180888 226392 180940
rect 104808 180752 104860 180804
rect 113180 180752 113232 180804
rect 214012 180752 214064 180804
rect 225788 180752 225840 180804
rect 214104 179732 214156 179784
rect 220084 179732 220136 179784
rect 221464 179460 221516 179512
rect 226432 179460 226484 179512
rect 113916 179392 113968 179444
rect 116400 179392 116452 179444
rect 225696 179392 225748 179444
rect 227628 179392 227680 179444
rect 104808 179324 104860 179376
rect 113272 179324 113324 179376
rect 213920 179188 213972 179240
rect 216036 179188 216088 179240
rect 215944 178644 215996 178696
rect 226340 178644 226392 178696
rect 214104 178576 214156 178628
rect 221648 178576 221700 178628
rect 114192 178032 114244 178084
rect 115940 178032 115992 178084
rect 220084 178032 220136 178084
rect 226432 178032 226484 178084
rect 104164 177964 104216 178016
rect 113916 177964 113968 178016
rect 224960 177964 225012 178016
rect 226984 177964 227036 178016
rect 215024 177488 215076 177540
rect 218796 177488 218848 177540
rect 113916 176740 113968 176792
rect 115940 176740 115992 176792
rect 114468 176672 114520 176724
rect 116400 176672 116452 176724
rect 218704 176672 218756 176724
rect 226340 176672 226392 176724
rect 104164 176604 104216 176656
rect 114192 176604 114244 176656
rect 215116 176604 215168 176656
rect 225604 176604 225656 176656
rect 215116 176128 215168 176180
rect 220176 176128 220228 176180
rect 220268 175584 220320 175636
rect 227168 175584 227220 175636
rect 114284 175244 114336 175296
rect 116400 175244 116452 175296
rect 222844 175244 222896 175296
rect 227444 175244 227496 175296
rect 104440 175176 104492 175228
rect 114468 175176 114520 175228
rect 214104 175176 214156 175228
rect 224960 175176 225012 175228
rect 104808 175108 104860 175160
rect 113916 175108 113968 175160
rect 215116 175108 215168 175160
rect 224224 175108 224276 175160
rect 114376 173884 114428 173936
rect 115940 173884 115992 173936
rect 225604 173884 225656 173936
rect 227352 173884 227404 173936
rect 104808 173816 104860 173868
rect 114284 173816 114336 173868
rect 214288 173816 214340 173868
rect 224316 173816 224368 173868
rect 224316 173272 224368 173324
rect 226708 173272 226760 173324
rect 113180 172524 113232 172576
rect 116400 172524 116452 172576
rect 104440 172456 104492 172508
rect 114376 172456 114428 172508
rect 214288 172456 214340 172508
rect 222936 172456 222988 172508
rect 215024 171980 215076 172032
rect 218888 171980 218940 172032
rect 113272 171572 113324 171624
rect 116124 171572 116176 171624
rect 104808 171028 104860 171080
rect 113180 171028 113232 171080
rect 113916 169804 113968 169856
rect 116308 169804 116360 169856
rect 104256 169736 104308 169788
rect 116400 169736 116452 169788
rect 104808 169668 104860 169720
rect 113272 169668 113324 169720
rect 215116 169668 215168 169720
rect 225696 169668 225748 169720
rect 215116 168580 215168 168632
rect 221556 168580 221608 168632
rect 104808 168376 104860 168428
rect 116400 168376 116452 168428
rect 104164 168308 104216 168360
rect 113916 168308 113968 168360
rect 213920 168036 213972 168088
rect 215944 168036 215996 168088
rect 215300 167628 215352 167680
rect 227076 167628 227128 167680
rect 214288 167560 214340 167612
rect 221464 167560 221516 167612
rect 114468 167016 114520 167068
rect 115940 167016 115992 167068
rect 232228 166948 232280 167000
rect 232596 166948 232648 167000
rect 214380 166812 214432 166864
rect 220084 166812 220136 166864
rect 217232 165792 217284 165844
rect 220268 165792 220320 165844
rect 113824 165588 113876 165640
rect 115940 165588 115992 165640
rect 104624 165520 104676 165572
rect 114468 165520 114520 165572
rect 214104 165520 214156 165572
rect 224316 165520 224368 165572
rect 114468 164228 114520 164280
rect 116124 164228 116176 164280
rect 104808 164160 104860 164212
rect 113824 164160 113876 164212
rect 214380 164160 214432 164212
rect 225604 164160 225656 164212
rect 232320 164160 232372 164212
rect 232596 164160 232648 164212
rect 214932 164092 214984 164144
rect 218704 164092 218756 164144
rect 214932 163344 214984 163396
rect 217232 163344 217284 163396
rect 113180 162868 113232 162920
rect 116400 162868 116452 162920
rect 104808 162800 104860 162852
rect 114468 162800 114520 162852
rect 214288 162800 214340 162852
rect 226984 162800 227036 162852
rect 215116 162732 215168 162784
rect 222844 162732 222896 162784
rect 113272 161984 113324 162036
rect 116216 161984 116268 162036
rect 103704 161440 103756 161492
rect 116400 161440 116452 161492
rect 104808 161372 104860 161424
rect 113180 161372 113232 161424
rect 215116 161372 215168 161424
rect 229744 161372 229796 161424
rect 104256 160080 104308 160132
rect 116400 160080 116452 160132
rect 104808 160012 104860 160064
rect 113272 160012 113324 160064
rect 104808 158720 104860 158772
rect 116400 158720 116452 158772
rect 104348 157360 104400 157412
rect 116400 157360 116452 157412
rect 114284 155932 114336 155984
rect 116032 155932 116084 155984
rect 215116 155932 215168 155984
rect 224684 155932 224736 155984
rect 113456 154640 113508 154692
rect 116032 154640 116084 154692
rect 214380 154640 214432 154692
rect 224592 154640 224644 154692
rect 104164 154572 104216 154624
rect 116400 154572 116452 154624
rect 215116 154572 215168 154624
rect 225604 154572 225656 154624
rect 104624 154504 104676 154556
rect 114284 154504 114336 154556
rect 215208 153280 215260 153332
rect 224868 153280 224920 153332
rect 103796 153212 103848 153264
rect 115940 153212 115992 153264
rect 215116 153212 215168 153264
rect 224776 153212 224828 153264
rect 104808 153144 104860 153196
rect 113456 153144 113508 153196
rect 214012 151852 214064 151904
rect 224500 151852 224552 151904
rect 103704 151784 103756 151836
rect 116400 151784 116452 151836
rect 218704 151784 218756 151836
rect 286140 151784 286192 151836
rect 214380 150492 214432 150544
rect 216680 150492 216732 150544
rect 104348 150424 104400 150476
rect 116400 150424 116452 150476
rect 215116 150424 215168 150476
rect 224040 150424 224092 150476
rect 224684 150356 224736 150408
rect 227444 150356 227496 150408
rect 232136 149676 232188 149728
rect 232504 149676 232556 149728
rect 214380 149200 214432 149252
rect 216864 149200 216916 149252
rect 104440 149064 104492 149116
rect 116400 149064 116452 149116
rect 215116 149064 215168 149116
rect 224224 149064 224276 149116
rect 214748 148996 214800 149048
rect 227444 148996 227496 149048
rect 224592 148928 224644 148980
rect 227536 148928 227588 148980
rect 104808 147636 104860 147688
rect 116400 147636 116452 147688
rect 215116 147636 215168 147688
rect 216772 147636 216824 147688
rect 224868 147568 224920 147620
rect 226708 147568 226760 147620
rect 224776 147500 224828 147552
rect 226524 147500 226576 147552
rect 113640 146344 113692 146396
rect 115940 146344 115992 146396
rect 215208 146344 215260 146396
rect 217692 146344 217744 146396
rect 104164 146276 104216 146328
rect 116400 146276 116452 146328
rect 214840 146276 214892 146328
rect 227628 146276 227680 146328
rect 216680 146208 216732 146260
rect 226708 146208 226760 146260
rect 224500 146140 224552 146192
rect 227444 146140 227496 146192
rect 215208 144984 215260 145036
rect 217416 144984 217468 145036
rect 104532 144916 104584 144968
rect 116032 144916 116084 144968
rect 215024 144916 215076 144968
rect 227260 144916 227312 144968
rect 104624 144848 104676 144900
rect 113640 144848 113692 144900
rect 216864 144848 216916 144900
rect 226524 144848 226576 144900
rect 224040 144780 224092 144832
rect 227444 144780 227496 144832
rect 215208 143624 215260 143676
rect 216680 143624 216732 143676
rect 103520 143556 103572 143608
rect 116400 143556 116452 143608
rect 214472 143556 214524 143608
rect 227536 143556 227588 143608
rect 216772 143488 216824 143540
rect 226892 143488 226944 143540
rect 224224 143420 224276 143472
rect 227444 143420 227496 143472
rect 215208 142196 215260 142248
rect 216772 142196 216824 142248
rect 103704 142128 103756 142180
rect 116400 142128 116452 142180
rect 215116 142128 215168 142180
rect 227352 142128 227404 142180
rect 217692 142060 217744 142112
rect 226708 142060 226760 142112
rect 104348 140768 104400 140820
rect 116400 140768 116452 140820
rect 215116 140768 215168 140820
rect 226708 140768 226760 140820
rect 217416 140700 217468 140752
rect 227076 140700 227128 140752
rect 113548 139476 113600 139528
rect 116308 139476 116360 139528
rect 214380 139476 214432 139528
rect 226616 139476 226668 139528
rect 104808 139408 104860 139460
rect 116400 139408 116452 139460
rect 215116 139408 215168 139460
rect 226524 139408 226576 139460
rect 216680 139340 216732 139392
rect 227444 139340 227496 139392
rect 215116 138048 215168 138100
rect 226800 138048 226852 138100
rect 214472 137980 214524 138032
rect 226432 137980 226484 138032
rect 216772 137912 216824 137964
rect 227444 137912 227496 137964
rect 215116 136688 215168 136740
rect 227260 136688 227312 136740
rect 104716 136620 104768 136672
rect 116400 136620 116452 136672
rect 214288 136620 214340 136672
rect 227444 136620 227496 136672
rect 104348 135260 104400 135312
rect 115940 135260 115992 135312
rect 214196 135260 214248 135312
rect 226524 135260 226576 135312
rect 104808 135192 104860 135244
rect 113548 135192 113600 135244
rect 341524 135192 341576 135244
rect 580172 135192 580224 135244
rect 215116 133968 215168 134020
rect 226708 133968 226760 134020
rect 109868 133900 109920 133952
rect 116400 133900 116452 133952
rect 215208 133900 215260 133952
rect 227536 133900 227588 133952
rect 104808 133832 104860 133884
rect 115848 133832 115900 133884
rect 114560 132880 114612 132932
rect 117136 132880 117188 132932
rect 214012 132540 214064 132592
rect 227352 132540 227404 132592
rect 215116 132472 215168 132524
rect 227444 132472 227496 132524
rect 215116 131180 215168 131232
rect 226524 131180 226576 131232
rect 113732 131112 113784 131164
rect 116124 131112 116176 131164
rect 214380 131112 214432 131164
rect 227076 131112 227128 131164
rect 103980 130704 104032 130756
rect 109868 130704 109920 130756
rect 100760 130364 100812 130416
rect 116400 130364 116452 130416
rect 214196 129752 214248 129804
rect 227536 129752 227588 129804
rect 104808 129684 104860 129736
rect 114560 129684 114612 129736
rect 116400 129276 116452 129328
rect 10416 129208 10468 129260
rect 214196 129004 214248 129056
rect 227444 129004 227496 129056
rect 214012 128324 214064 128376
rect 226340 128324 226392 128376
rect 9036 128256 9088 128308
rect 116400 128256 116452 128308
rect 104808 128188 104860 128240
rect 113732 128188 113784 128240
rect 215116 127576 215168 127628
rect 227444 127576 227496 127628
rect 215116 126964 215168 127016
rect 227444 126964 227496 127016
rect 10324 126896 10376 126948
rect 116400 126896 116452 126948
rect 215116 126216 215168 126268
rect 227444 126216 227496 126268
rect 215116 125604 215168 125656
rect 227444 125604 227496 125656
rect 8944 125536 8996 125588
rect 116400 125536 116452 125588
rect 78220 125468 78272 125520
rect 100760 125468 100812 125520
rect 215116 124856 215168 124908
rect 227260 124856 227312 124908
rect 215116 124108 215168 124160
rect 227260 124108 227312 124160
rect 215116 123428 215168 123480
rect 227260 123428 227312 123480
rect 215116 122748 215168 122800
rect 227444 122748 227496 122800
rect 215116 122068 215168 122120
rect 227444 122068 227496 122120
rect 50988 121456 51040 121508
rect 116400 121456 116452 121508
rect 215116 121388 215168 121440
rect 227444 121388 227496 121440
rect 215116 120708 215168 120760
rect 227444 120708 227496 120760
rect 100024 120096 100076 120148
rect 116400 120096 116452 120148
rect 214196 120028 214248 120080
rect 227444 120028 227496 120080
rect 94780 118668 94832 118720
rect 116400 118668 116452 118720
rect 214288 118600 214340 118652
rect 226340 118600 226392 118652
rect 215116 118532 215168 118584
rect 226432 118532 226484 118584
rect 94688 117308 94740 117360
rect 116400 117308 116452 117360
rect 215208 117240 215260 117292
rect 227444 117240 227496 117292
rect 215116 117172 215168 117224
rect 226248 117172 226300 117224
rect 94872 116016 94924 116068
rect 116308 116016 116360 116068
rect 94596 115948 94648 116000
rect 116400 115948 116452 116000
rect 215208 115880 215260 115932
rect 227444 115880 227496 115932
rect 215116 115812 215168 115864
rect 226156 115812 226208 115864
rect 94504 114520 94556 114572
rect 116400 114520 116452 114572
rect 215116 114452 215168 114504
rect 227076 114452 227128 114504
rect 214012 114384 214064 114436
rect 226248 114384 226300 114436
rect 95884 113160 95936 113212
rect 116400 113160 116452 113212
rect 214380 113092 214432 113144
rect 226156 113092 226208 113144
rect 98644 111800 98696 111852
rect 116400 111800 116452 111852
rect 215208 111732 215260 111784
rect 226248 111732 226300 111784
rect 215116 111664 215168 111716
rect 226064 111664 226116 111716
rect 104164 110440 104216 110492
rect 116400 110440 116452 110492
rect 215116 110372 215168 110424
rect 225972 110372 226024 110424
rect 214472 110304 214524 110356
rect 226156 110304 226208 110356
rect 94964 109012 95016 109064
rect 116400 109012 116452 109064
rect 215208 108944 215260 108996
rect 226248 108944 226300 108996
rect 215116 108876 215168 108928
rect 225788 108876 225840 108928
rect 105544 107720 105596 107772
rect 116308 107720 116360 107772
rect 97264 107652 97316 107704
rect 116400 107652 116452 107704
rect 214196 107584 214248 107636
rect 226064 107584 226116 107636
rect 101404 106292 101456 106344
rect 116400 106292 116452 106344
rect 215116 106224 215168 106276
rect 225696 106224 225748 106276
rect 214380 106156 214432 106208
rect 226156 106156 226208 106208
rect 97356 104864 97408 104916
rect 116400 104864 116452 104916
rect 224776 104864 224828 104916
rect 227444 104864 227496 104916
rect 215116 104796 215168 104848
rect 225604 104796 225656 104848
rect 214380 104728 214432 104780
rect 226248 104728 226300 104780
rect 224868 103640 224920 103692
rect 227444 103640 227496 103692
rect 102784 103504 102836 103556
rect 116400 103504 116452 103556
rect 215116 103436 215168 103488
rect 226064 103436 226116 103488
rect 215208 103368 215260 103420
rect 225788 103368 225840 103420
rect 95976 102144 96028 102196
rect 116308 102144 116360 102196
rect 215116 102076 215168 102128
rect 225880 102076 225932 102128
rect 314200 102076 314252 102128
rect 338396 102076 338448 102128
rect 98736 100716 98788 100768
rect 116400 100716 116452 100768
rect 214472 100648 214524 100700
rect 226156 100648 226208 100700
rect 232136 100648 232188 100700
rect 258080 100648 258132 100700
rect 215116 100580 215168 100632
rect 225972 100580 226024 100632
rect 100116 99356 100168 99408
rect 116400 99356 116452 99408
rect 214656 99288 214708 99340
rect 226248 99288 226300 99340
rect 232136 99288 232188 99340
rect 232504 99288 232556 99340
rect 215116 99220 215168 99272
rect 224776 99220 224828 99272
rect 95148 98948 95200 99000
rect 100024 98948 100076 99000
rect 106924 97996 106976 98048
rect 116400 97996 116452 98048
rect 214104 97928 214156 97980
rect 224868 97928 224920 97980
rect 214564 96976 214616 97028
rect 218704 96976 218756 97028
rect 96068 96636 96120 96688
rect 116400 96636 116452 96688
rect 94688 95208 94740 95260
rect 116308 95208 116360 95260
rect 215116 95140 215168 95192
rect 576124 95140 576176 95192
rect 94596 93848 94648 93900
rect 116400 93848 116452 93900
rect 215208 93780 215260 93832
rect 578884 93780 578936 93832
rect 215116 93712 215168 93764
rect 577504 93712 577556 93764
rect 94872 93644 94924 93696
rect 95884 93644 95936 93696
rect 94412 93304 94464 93356
rect 98644 93304 98696 93356
rect 98828 93100 98880 93152
rect 116676 93100 116728 93152
rect 101496 92488 101548 92540
rect 116400 92488 116452 92540
rect 95148 92420 95200 92472
rect 104164 92420 104216 92472
rect 104256 91060 104308 91112
rect 116400 91060 116452 91112
rect 95056 90992 95108 91044
rect 105544 90992 105596 91044
rect 97448 89700 97500 89752
rect 116400 89700 116452 89752
rect 214472 89700 214524 89752
rect 227352 89700 227404 89752
rect 95148 89292 95200 89344
rect 97264 89292 97316 89344
rect 215116 88408 215168 88460
rect 221464 88408 221516 88460
rect 97540 88340 97592 88392
rect 115940 88340 115992 88392
rect 214104 88340 214156 88392
rect 222844 88340 222896 88392
rect 340144 88272 340196 88324
rect 580172 88272 580224 88324
rect 95148 88204 95200 88256
rect 101404 88204 101456 88256
rect 94412 87864 94464 87916
rect 97356 87864 97408 87916
rect 215024 87048 215076 87100
rect 218704 87048 218756 87100
rect 98644 86980 98696 87032
rect 116400 86980 116452 87032
rect 215116 86980 215168 87032
rect 224224 86980 224276 87032
rect 232320 86912 232372 86964
rect 232504 86912 232556 86964
rect 94504 86708 94556 86760
rect 102784 86708 102836 86760
rect 94044 86164 94096 86216
rect 98736 86164 98788 86216
rect 102876 85552 102928 85604
rect 116124 85552 116176 85604
rect 215116 85552 215168 85604
rect 225604 85552 225656 85604
rect 94872 85484 94924 85536
rect 95976 85484 96028 85536
rect 95148 84804 95200 84856
rect 98828 84804 98880 84856
rect 100024 84804 100076 84856
rect 116400 84804 116452 84856
rect 215208 84192 215260 84244
rect 227076 84192 227128 84244
rect 320824 83512 320876 83564
rect 412088 83512 412140 83564
rect 284484 83444 284536 83496
rect 580264 83444 580316 83496
rect 94228 83376 94280 83428
rect 100116 83376 100168 83428
rect 95884 82832 95936 82884
rect 116400 82832 116452 82884
rect 215944 82832 215996 82884
rect 248144 82832 248196 82884
rect 95148 82764 95200 82816
rect 106924 82764 106976 82816
rect 94964 81404 95016 81456
rect 97540 81404 97592 81456
rect 98736 81404 98788 81456
rect 115940 81404 115992 81456
rect 214196 81404 214248 81456
rect 227168 81404 227220 81456
rect 94412 81336 94464 81388
rect 96068 81336 96120 81388
rect 214564 81336 214616 81388
rect 227444 81336 227496 81388
rect 214748 81268 214800 81320
rect 227536 81268 227588 81320
rect 95240 80656 95292 80708
rect 116584 80656 116636 80708
rect 97264 80044 97316 80096
rect 116400 80044 116452 80096
rect 214012 80044 214064 80096
rect 216128 80044 216180 80096
rect 232320 80044 232372 80096
rect 221464 79976 221516 80028
rect 227444 79976 227496 80028
rect 232320 79908 232372 79960
rect 96068 79296 96120 79348
rect 117044 79296 117096 79348
rect 215116 78752 215168 78804
rect 221556 78752 221608 78804
rect 102784 78684 102836 78736
rect 116400 78684 116452 78736
rect 94412 78616 94464 78668
rect 101496 78616 101548 78668
rect 218704 78616 218756 78668
rect 227536 78616 227588 78668
rect 222844 78548 222896 78600
rect 227444 78548 227496 78600
rect 94228 77936 94280 77988
rect 104256 77936 104308 77988
rect 101404 77256 101456 77308
rect 116400 77256 116452 77308
rect 214748 77256 214800 77308
rect 218796 77256 218848 77308
rect 215208 77188 215260 77240
rect 227536 77188 227588 77240
rect 224224 77120 224276 77172
rect 227444 77120 227496 77172
rect 94044 76848 94096 76900
rect 102876 76848 102928 76900
rect 95976 75896 96028 75948
rect 116400 75896 116452 75948
rect 215208 75896 215260 75948
rect 218060 75896 218112 75948
rect 214656 75828 214708 75880
rect 227444 75828 227496 75880
rect 94596 75692 94648 75744
rect 97448 75692 97500 75744
rect 215208 74604 215260 74656
rect 216036 74604 216088 74656
rect 94596 74536 94648 74588
rect 116400 74536 116452 74588
rect 214840 74468 214892 74520
rect 227444 74468 227496 74520
rect 95148 74196 95200 74248
rect 98644 74196 98696 74248
rect 96620 73788 96672 73840
rect 116584 73788 116636 73840
rect 214840 73448 214892 73500
rect 215116 73448 215168 73500
rect 215116 73312 215168 73364
rect 220728 73312 220780 73364
rect 98828 73176 98880 73228
rect 116400 73176 116452 73228
rect 214932 73108 214984 73160
rect 227444 73108 227496 73160
rect 216128 73040 216180 73092
rect 227536 73040 227588 73092
rect 94412 72632 94464 72684
rect 100024 72632 100076 72684
rect 94780 71748 94832 71800
rect 116400 71748 116452 71800
rect 94228 71680 94280 71732
rect 96068 71680 96120 71732
rect 215024 71680 215076 71732
rect 227444 71680 227496 71732
rect 221556 71612 221608 71664
rect 227536 71612 227588 71664
rect 95056 70456 95108 70508
rect 98736 70456 98788 70508
rect 100024 70456 100076 70508
rect 116308 70456 116360 70508
rect 215116 70456 215168 70508
rect 224132 70456 224184 70508
rect 94504 70388 94556 70440
rect 116400 70388 116452 70440
rect 214104 70388 214156 70440
rect 224868 70388 224920 70440
rect 214564 70320 214616 70372
rect 227444 70320 227496 70372
rect 94872 70252 94924 70304
rect 95884 70252 95936 70304
rect 218796 70252 218848 70304
rect 226524 70252 226576 70304
rect 95148 69844 95200 69896
rect 102784 69844 102836 69896
rect 214932 69096 214984 69148
rect 224408 69096 224460 69148
rect 96068 69028 96120 69080
rect 116400 69028 116452 69080
rect 215116 69028 215168 69080
rect 224592 69028 224644 69080
rect 214472 68960 214524 69012
rect 227444 68960 227496 69012
rect 218060 68892 218112 68944
rect 227536 68892 227588 68944
rect 94044 68552 94096 68604
rect 97264 68552 97316 68604
rect 215208 67668 215260 67720
rect 224224 67668 224276 67720
rect 94688 67600 94740 67652
rect 116400 67600 116452 67652
rect 215116 67600 215168 67652
rect 224776 67600 224828 67652
rect 214840 67532 214892 67584
rect 227444 67532 227496 67584
rect 95148 67464 95200 67516
rect 96620 67464 96672 67516
rect 216036 67464 216088 67516
rect 227536 67464 227588 67516
rect 97264 66240 97316 66292
rect 116400 66240 116452 66292
rect 215116 66240 215168 66292
rect 224684 66240 224736 66292
rect 214288 66172 214340 66224
rect 227444 66172 227496 66224
rect 220728 66104 220780 66156
rect 227536 66104 227588 66156
rect 94412 65968 94464 66020
rect 95976 65968 96028 66020
rect 94136 65900 94188 65952
rect 101404 65900 101456 65952
rect 213920 65152 213972 65204
rect 216864 65152 216916 65204
rect 94872 64880 94924 64932
rect 116400 64880 116452 64932
rect 214012 64880 214064 64932
rect 224500 64880 224552 64932
rect 214656 64676 214708 64728
rect 227260 64676 227312 64728
rect 224868 64472 224920 64524
rect 227444 64472 227496 64524
rect 224132 64200 224184 64252
rect 227536 64200 227588 64252
rect 214104 63588 214156 63640
rect 216956 63588 217008 63640
rect 95240 63520 95292 63572
rect 115940 63520 115992 63572
rect 215116 63520 215168 63572
rect 224316 63520 224368 63572
rect 224592 63452 224644 63504
rect 227076 63452 227128 63504
rect 224408 63384 224460 63436
rect 227444 63384 227496 63436
rect 95148 63180 95200 63232
rect 98828 63180 98880 63232
rect 487620 62772 487672 62824
rect 573364 62772 573416 62824
rect 214380 62160 214432 62212
rect 216680 62160 216732 62212
rect 94596 62092 94648 62144
rect 116400 62092 116452 62144
rect 215116 62092 215168 62144
rect 224132 62092 224184 62144
rect 224776 62024 224828 62076
rect 226708 62024 226760 62076
rect 224224 61956 224276 62008
rect 227444 61956 227496 62008
rect 94320 61752 94372 61804
rect 100024 61752 100076 61804
rect 214748 60800 214800 60852
rect 216772 60800 216824 60852
rect 94780 60732 94832 60784
rect 116400 60732 116452 60784
rect 215116 60732 215168 60784
rect 224408 60732 224460 60784
rect 216864 60664 216916 60716
rect 227536 60664 227588 60716
rect 224684 60596 224736 60648
rect 227444 60596 227496 60648
rect 96160 59984 96212 60036
rect 116492 59984 116544 60036
rect 94320 59848 94372 59900
rect 96068 59848 96120 59900
rect 97356 59372 97408 59424
rect 116400 59372 116452 59424
rect 214380 59372 214432 59424
rect 217324 59372 217376 59424
rect 216956 59304 217008 59356
rect 227536 59304 227588 59356
rect 224500 59236 224552 59288
rect 227444 59236 227496 59288
rect 214288 58012 214340 58064
rect 217692 58012 217744 58064
rect 94964 57944 95016 57996
rect 116400 57944 116452 57996
rect 214380 57944 214432 57996
rect 217784 57944 217836 57996
rect 94412 57876 94464 57928
rect 97264 57876 97316 57928
rect 216680 57876 216732 57928
rect 227444 57876 227496 57928
rect 224316 57808 224368 57860
rect 227260 57808 227312 57860
rect 213920 56652 213972 56704
rect 216864 56652 216916 56704
rect 95240 56584 95292 56636
rect 116308 56584 116360 56636
rect 214012 56584 214064 56636
rect 216680 56584 216732 56636
rect 216772 56516 216824 56568
rect 227444 56516 227496 56568
rect 224132 56448 224184 56500
rect 227260 56448 227312 56500
rect 94044 55292 94096 55344
rect 116308 55292 116360 55344
rect 94136 55224 94188 55276
rect 116400 55224 116452 55276
rect 215116 55224 215168 55276
rect 227536 55224 227588 55276
rect 217324 55156 217376 55208
rect 224408 55156 224460 55208
rect 227444 55156 227496 55208
rect 226524 55020 226576 55072
rect 94596 54680 94648 54732
rect 96160 54680 96212 54732
rect 214748 53864 214800 53916
rect 226524 53864 226576 53916
rect 94872 53796 94924 53848
rect 116400 53796 116452 53848
rect 215116 53796 215168 53848
rect 226984 53796 227036 53848
rect 217784 53728 217836 53780
rect 227444 53728 227496 53780
rect 217692 53660 217744 53712
rect 227260 53660 227312 53712
rect 215116 52504 215168 52556
rect 226800 52504 226852 52556
rect 94780 52436 94832 52488
rect 116400 52436 116452 52488
rect 214748 52436 214800 52488
rect 226708 52436 226760 52488
rect 95148 52368 95200 52420
rect 97356 52368 97408 52420
rect 216680 52368 216732 52420
rect 227444 52368 227496 52420
rect 216864 52300 216916 52352
rect 227260 52300 227312 52352
rect 215116 51144 215168 51196
rect 226616 51144 226668 51196
rect 95056 51076 95108 51128
rect 115940 51076 115992 51128
rect 214564 51076 214616 51128
rect 226340 51076 226392 51128
rect 214380 49784 214432 49836
rect 227352 49784 227404 49836
rect 95148 49716 95200 49768
rect 116400 49716 116452 49768
rect 215116 49716 215168 49768
rect 227076 49716 227128 49768
rect 94964 48356 95016 48408
rect 116124 48356 116176 48408
rect 94412 48288 94464 48340
rect 116400 48288 116452 48340
rect 215116 48288 215168 48340
rect 227536 48288 227588 48340
rect 214748 46996 214800 47048
rect 227444 46996 227496 47048
rect 94136 46928 94188 46980
rect 116400 46928 116452 46980
rect 214012 46928 214064 46980
rect 227628 46928 227680 46980
rect 215116 45636 215168 45688
rect 226708 45636 226760 45688
rect 93952 45568 94004 45620
rect 116400 45568 116452 45620
rect 215208 45568 215260 45620
rect 227076 45568 227128 45620
rect 215116 44208 215168 44260
rect 227352 44208 227404 44260
rect 95056 44140 95108 44192
rect 116400 44140 116452 44192
rect 214472 44140 214524 44192
rect 227444 44140 227496 44192
rect 94596 42780 94648 42832
rect 115940 42780 115992 42832
rect 214380 42780 214432 42832
rect 226432 42780 226484 42832
rect 215116 41488 215168 41540
rect 226616 41488 226668 41540
rect 95148 41420 95200 41472
rect 116400 41420 116452 41472
rect 214104 41420 214156 41472
rect 226340 41420 226392 41472
rect 560944 41352 560996 41404
rect 580172 41352 580224 41404
rect 94504 40128 94556 40180
rect 116308 40128 116360 40180
rect 215116 40128 215168 40180
rect 226892 40128 226944 40180
rect 95056 40060 95108 40112
rect 116400 40060 116452 40112
rect 214656 40060 214708 40112
rect 227076 40060 227128 40112
rect 214472 38700 214524 38752
rect 227444 38700 227496 38752
rect 94596 38632 94648 38684
rect 116400 38632 116452 38684
rect 215116 38632 215168 38684
rect 227536 38632 227588 38684
rect 93860 37272 93912 37324
rect 116400 37272 116452 37324
rect 215116 37272 215168 37324
rect 227444 37272 227496 37324
rect 214564 35980 214616 36032
rect 227536 35980 227588 36032
rect 93952 35912 94004 35964
rect 116400 35912 116452 35964
rect 215116 35912 215168 35964
rect 227444 35912 227496 35964
rect 3424 35844 3476 35896
rect 9128 35844 9180 35896
rect 215116 34552 215168 34604
rect 227352 34552 227404 34604
rect 95148 34484 95200 34536
rect 116400 34484 116452 34536
rect 214656 34484 214708 34536
rect 227444 34484 227496 34536
rect 215116 33192 215168 33244
rect 227536 33192 227588 33244
rect 95148 33124 95200 33176
rect 116308 33124 116360 33176
rect 214564 33124 214616 33176
rect 227444 33124 227496 33176
rect 213920 32512 213972 32564
rect 215944 32512 215996 32564
rect 95148 32376 95200 32428
rect 116400 32376 116452 32428
rect 215116 32376 215168 32428
rect 227444 32376 227496 32428
rect 71688 31764 71740 31816
rect 116400 31764 116452 31816
rect 29920 30268 29972 30320
rect 32312 30268 32364 30320
rect 119988 30268 120040 30320
rect 231952 30268 232004 30320
rect 284576 30268 284628 30320
rect 115848 30200 115900 30252
rect 203248 30200 203300 30252
rect 107568 30132 107620 30184
rect 198096 30132 198148 30184
rect 51724 30064 51776 30116
rect 143356 30064 143408 30116
rect 57244 29996 57296 30048
rect 148600 29996 148652 30048
rect 32404 29928 32456 29980
rect 134708 29928 134760 29980
rect 28264 29860 28316 29912
rect 131212 29860 131264 29912
rect 164884 29860 164936 29912
rect 185032 29860 185084 29912
rect 24124 29792 24176 29844
rect 127716 29792 127768 29844
rect 159364 29792 159416 29844
rect 179788 29792 179840 29844
rect 31024 29724 31076 29776
rect 140780 29724 140832 29776
rect 166264 29724 166316 29776
rect 190276 29724 190328 29776
rect 22744 29656 22796 29708
rect 133788 29656 133840 29708
rect 169024 29656 169076 29708
rect 195428 29656 195480 29708
rect 25504 29588 25556 29640
rect 137284 29588 137336 29640
rect 171784 29588 171836 29640
rect 200672 29588 200724 29640
rect 118608 29520 118660 29572
rect 205824 29520 205876 29572
rect 61384 29452 61436 29504
rect 123392 29452 123444 29504
rect 123484 29452 123536 29504
rect 208492 29452 208544 29504
rect 69664 29384 69716 29436
rect 124312 29384 124364 29436
rect 126244 29384 126296 29436
rect 211068 29384 211120 29436
rect 142804 28976 142856 29028
rect 146024 28976 146076 29028
rect 199016 28908 199068 28960
rect 199108 28908 199160 28960
rect 135260 28840 135312 28892
rect 136180 28840 136232 28892
rect 138112 28840 138164 28892
rect 138756 28840 138808 28892
rect 113088 28364 113140 28416
rect 201500 28364 201552 28416
rect 50988 28296 51040 28348
rect 156420 28296 156472 28348
rect 8944 28228 8996 28280
rect 121644 28228 121696 28280
rect 125508 28228 125560 28280
rect 210240 28228 210292 28280
rect 117228 27072 117280 27124
rect 204168 27072 204220 27124
rect 107476 27004 107528 27056
rect 197176 27004 197228 27056
rect 62028 26936 62080 26988
rect 164240 26936 164292 26988
rect 11704 26868 11756 26920
rect 125140 26868 125192 26920
rect 125876 26732 125928 26784
rect 126612 26732 126664 26784
rect 154580 26732 154632 26784
rect 155132 26732 155184 26784
rect 186504 26256 186556 26308
rect 187332 26256 187384 26308
rect 85488 25644 85540 25696
rect 181536 25644 181588 25696
rect 68928 25576 68980 25628
rect 169392 25576 169444 25628
rect 59268 25508 59320 25560
rect 161572 25508 161624 25560
rect 96528 24216 96580 24268
rect 189172 24216 189224 24268
rect 63408 24148 63460 24200
rect 164240 24148 164292 24200
rect 57888 24080 57940 24132
rect 161480 24080 161532 24132
rect 182180 23740 182232 23792
rect 182916 23740 182968 23792
rect 89628 22856 89680 22908
rect 184204 22856 184256 22908
rect 64788 22788 64840 22840
rect 165896 22788 165948 22840
rect 56508 22720 56560 22772
rect 158812 22720 158864 22772
rect 175464 22040 175516 22092
rect 175556 21972 175608 22024
rect 100668 21564 100720 21616
rect 192116 21564 192168 21616
rect 82728 21496 82780 21548
rect 178132 21496 178184 21548
rect 72976 21428 73028 21480
rect 171232 21428 171284 21480
rect 52368 21360 52420 21412
rect 156052 21360 156104 21412
rect 119988 20136 120040 20188
rect 205824 20136 205876 20188
rect 75828 20068 75880 20120
rect 173900 20068 173952 20120
rect 48228 20000 48280 20052
rect 154672 20000 154724 20052
rect 10968 19932 11020 19984
rect 125876 19932 125928 19984
rect 199108 19320 199160 19372
rect 199200 19320 199252 19372
rect 148048 19252 148100 19304
rect 152004 19252 152056 19304
rect 208492 19252 208544 19304
rect 208676 19252 208728 19304
rect 79968 18640 80020 18692
rect 176660 18640 176712 18692
rect 30288 18572 30340 18624
rect 140872 18572 140924 18624
rect 129648 17960 129700 18012
rect 406476 17960 406528 18012
rect 414388 17620 414440 17672
rect 414296 17416 414348 17468
rect 287060 17348 287112 17400
rect 296536 17348 296588 17400
rect 393964 17348 394016 17400
rect 410524 17348 410576 17400
rect 410616 17348 410668 17400
rect 38568 17280 38620 17332
rect 147772 17280 147824 17332
rect 246948 17280 247000 17332
rect 270500 17280 270552 17332
rect 300768 17280 300820 17332
rect 414388 17280 414440 17332
rect 17868 17212 17920 17264
rect 131304 17212 131356 17264
rect 278688 17212 278740 17264
rect 414296 17212 414348 17264
rect 267648 17144 267700 17196
rect 393964 17144 394016 17196
rect 270592 17076 270644 17128
rect 287060 17076 287112 17128
rect 296536 17076 296588 17128
rect 217968 17008 218020 17060
rect 424600 17008 424652 17060
rect 439412 17008 439464 17060
rect 459100 17008 459152 17060
rect 462596 17008 462648 17060
rect 470048 17008 470100 17060
rect 202788 16940 202840 16992
rect 418712 16940 418764 16992
rect 425612 16940 425664 16992
rect 193128 16872 193180 16924
rect 430028 16872 430080 16924
rect 184848 16804 184900 16856
rect 429936 16804 429988 16856
rect 164148 16736 164200 16788
rect 425796 16736 425848 16788
rect 160008 16668 160060 16720
rect 424232 16668 424284 16720
rect 435364 16736 435416 16788
rect 443000 16736 443052 16788
rect 438400 16668 438452 16720
rect 132408 16600 132460 16652
rect 415400 16600 415452 16652
rect 418712 16600 418764 16652
rect 425612 16600 425664 16652
rect 429936 16600 429988 16652
rect 432696 16600 432748 16652
rect 430028 16532 430080 16584
rect 434996 16532 435048 16584
rect 479064 16396 479116 16448
rect 479800 16396 479852 16448
rect 534356 16396 534408 16448
rect 535000 16396 535052 16448
rect 187608 16192 187660 16244
rect 433708 16192 433760 16244
rect 180708 16124 180760 16176
rect 431408 16124 431460 16176
rect 387708 16056 387760 16108
rect 498108 16056 498160 16108
rect 376208 15988 376260 16040
rect 494704 15988 494756 16040
rect 55128 15920 55180 15972
rect 158720 15920 158772 15972
rect 311164 15920 311216 15972
rect 451004 15920 451056 15972
rect 34428 15852 34480 15904
rect 143540 15852 143592 15904
rect 339408 15852 339460 15904
rect 482376 15852 482428 15904
rect 326344 15784 326396 15836
rect 471704 15784 471756 15836
rect 333244 15716 333296 15768
rect 479708 15716 479760 15768
rect 282184 15648 282236 15700
rect 439504 15648 439556 15700
rect 275284 15580 275336 15632
rect 437204 15580 437256 15632
rect 280068 15512 280120 15564
rect 463240 15512 463292 15564
rect 259368 15444 259420 15496
rect 456708 15444 456760 15496
rect 248328 15376 248380 15428
rect 453304 15376 453356 15428
rect 234528 15308 234580 15360
rect 448704 15308 448756 15360
rect 405648 15240 405700 15292
rect 503904 15240 503956 15292
rect 398748 15172 398800 15224
rect 501604 15172 501656 15224
rect 368664 15104 368716 15156
rect 476304 15104 476356 15156
rect 525064 15104 525116 15156
rect 534540 15104 534592 15156
rect 535368 15104 535420 15156
rect 545672 15104 545724 15156
rect 390468 15036 390520 15088
rect 498844 15036 498896 15088
rect 527916 15036 527968 15088
rect 539140 15036 539192 15088
rect 368388 14968 368440 15020
rect 491944 14968 491996 15020
rect 530584 14968 530636 15020
rect 541440 14968 541492 15020
rect 357348 14900 357400 14952
rect 488540 14900 488592 14952
rect 511908 14900 511960 14952
rect 537944 14900 537996 14952
rect 350172 14832 350224 14884
rect 486240 14832 486292 14884
rect 491944 14832 491996 14884
rect 520740 14832 520792 14884
rect 527824 14832 527876 14884
rect 540244 14832 540296 14884
rect 329748 14764 329800 14816
rect 479340 14764 479392 14816
rect 482928 14764 482980 14816
rect 528744 14764 528796 14816
rect 531964 14764 532016 14816
rect 543740 14764 543792 14816
rect 93768 14696 93820 14748
rect 186504 14696 186556 14748
rect 314568 14696 314620 14748
rect 474740 14696 474792 14748
rect 478788 14696 478840 14748
rect 527640 14696 527692 14748
rect 531228 14696 531280 14748
rect 544476 14696 544528 14748
rect 66168 14628 66220 14680
rect 167000 14628 167052 14680
rect 250536 14628 250588 14680
rect 419448 14628 419500 14680
rect 147588 14560 147640 14612
rect 420644 14628 420696 14680
rect 426992 14628 427044 14680
rect 435640 14628 435692 14680
rect 440424 14628 440476 14680
rect 444472 14628 444524 14680
rect 464988 14628 465040 14680
rect 523040 14628 523092 14680
rect 528468 14628 528520 14680
rect 543372 14628 543424 14680
rect 555608 14628 555660 14680
rect 561680 14628 561732 14680
rect 419632 14560 419684 14612
rect 483204 14560 483256 14612
rect 503628 14560 503680 14612
rect 535644 14560 535696 14612
rect 536748 14560 536800 14612
rect 546040 14560 546092 14612
rect 554872 14560 554924 14612
rect 563152 14560 563204 14612
rect 154488 14492 154540 14544
rect 28908 14424 28960 14476
rect 139400 14424 139452 14476
rect 143448 14424 143500 14476
rect 419540 14424 419592 14476
rect 420920 14492 420972 14544
rect 422944 14424 422996 14476
rect 423128 14424 423180 14476
rect 426440 14424 426492 14476
rect 428464 14492 428516 14544
rect 431040 14492 431092 14544
rect 433248 14492 433300 14544
rect 512644 14492 512696 14544
rect 525708 14492 525760 14544
rect 542544 14492 542596 14544
rect 555240 14492 555292 14544
rect 563060 14492 563112 14544
rect 506204 14424 506256 14476
rect 507768 14424 507820 14476
rect 536840 14424 536892 14476
rect 538128 14424 538180 14476
rect 546776 14424 546828 14476
rect 557908 14424 557960 14476
rect 570604 14424 570656 14476
rect 397368 14356 397420 14408
rect 501144 14356 501196 14408
rect 523960 14356 524012 14408
rect 408408 14288 408460 14340
rect 504640 14288 504692 14340
rect 528652 14356 528704 14408
rect 529296 14356 529348 14408
rect 536104 14356 536156 14408
rect 544844 14356 544896 14408
rect 532240 14288 532292 14340
rect 553676 14288 553728 14340
rect 556988 14288 557040 14340
rect 378048 14220 378100 14272
rect 467840 14220 467892 14272
rect 471980 14220 472032 14272
rect 525340 14220 525392 14272
rect 554044 14220 554096 14272
rect 556620 14220 556672 14272
rect 384120 14152 384172 14204
rect 418344 14152 418396 14204
rect 418528 14152 418580 14204
rect 506940 14152 506992 14204
rect 543648 14152 543700 14204
rect 548340 14152 548392 14204
rect 554504 14152 554556 14204
rect 556896 14152 556948 14204
rect 419540 14084 419592 14136
rect 482008 14084 482060 14136
rect 545028 14084 545080 14136
rect 548708 14084 548760 14136
rect 552204 14084 552256 14136
rect 555240 14084 555292 14136
rect 411260 14016 411312 14068
rect 419448 14016 419500 14068
rect 425244 14016 425296 14068
rect 546316 14016 546368 14068
rect 549076 14016 549128 14068
rect 552940 14016 552992 14068
rect 555516 14016 555568 14068
rect 422208 13948 422260 14000
rect 547696 13948 547748 14000
rect 549904 13948 549956 14000
rect 553308 13948 553360 14000
rect 555424 13948 555476 14000
rect 559840 13948 559892 14000
rect 560208 13948 560260 14000
rect 425060 13880 425112 13932
rect 428740 13880 428792 13932
rect 544384 13880 544436 13932
rect 546408 13880 546460 13932
rect 547788 13880 547840 13932
rect 549444 13880 549496 13932
rect 551376 13880 551428 13932
rect 551836 13880 551888 13932
rect 552572 13880 552624 13932
rect 554872 13880 554924 13932
rect 557540 13880 557592 13932
rect 558736 13880 558788 13932
rect 559104 13880 559156 13932
rect 560024 13880 560076 13932
rect 375196 13744 375248 13796
rect 545764 13812 545816 13864
rect 547144 13812 547196 13864
rect 549168 13812 549220 13864
rect 550272 13812 550324 13864
rect 551744 13812 551796 13864
rect 553400 13812 553452 13864
rect 556344 13812 556396 13864
rect 557264 13812 557316 13864
rect 558276 13812 558328 13864
rect 558828 13812 558880 13864
rect 559472 13812 559524 13864
rect 560116 13812 560168 13864
rect 560576 13812 560628 13864
rect 561588 13812 561640 13864
rect 493876 13744 493928 13796
rect 293868 13676 293920 13728
rect 378048 13676 378100 13728
rect 378140 13676 378192 13728
rect 495072 13676 495124 13728
rect 320088 13608 320140 13660
rect 368664 13608 368716 13660
rect 371148 13608 371200 13660
rect 492772 13608 492824 13660
rect 364248 13540 364300 13592
rect 490472 13540 490524 13592
rect 360108 13472 360160 13524
rect 489276 13472 489328 13524
rect 504364 13472 504416 13524
rect 516140 13472 516192 13524
rect 269028 13404 269080 13456
rect 459744 13404 459796 13456
rect 499120 13404 499172 13456
rect 511540 13404 511592 13456
rect 226248 13336 226300 13388
rect 445944 13336 445996 13388
rect 500224 13336 500276 13388
rect 513840 13336 513892 13388
rect 190368 13268 190420 13320
rect 434444 13268 434496 13320
rect 456984 13268 457036 13320
rect 457444 13268 457496 13320
rect 496728 13268 496780 13320
rect 533344 13268 533396 13320
rect 140688 13200 140740 13252
rect 384120 13200 384172 13252
rect 384488 13200 384540 13252
rect 497372 13200 497424 13252
rect 498108 13200 498160 13252
rect 533804 13200 533856 13252
rect 42708 13132 42760 13184
rect 149336 13132 149388 13184
rect 153108 13132 153160 13184
rect 409144 13132 409196 13184
rect 436744 13132 436796 13184
rect 466644 13132 466696 13184
rect 495348 13132 495400 13184
rect 532608 13132 532660 13184
rect 533988 13132 534040 13184
rect 545304 13132 545356 13184
rect 22008 13064 22060 13116
rect 135352 13064 135404 13116
rect 150348 13064 150400 13116
rect 421472 13064 421524 13116
rect 424968 13064 425020 13116
rect 509976 13064 510028 13116
rect 517428 13064 517480 13116
rect 539876 13064 539928 13116
rect 382188 12996 382240 13048
rect 496176 12996 496228 13048
rect 389088 12928 389140 12980
rect 498476 12928 498528 12980
rect 391848 12860 391900 12912
rect 407028 12792 407080 12844
rect 490564 12792 490616 12844
rect 415308 12724 415360 12776
rect 422576 12724 422628 12776
rect 422760 12724 422812 12776
rect 447048 12724 447100 12776
rect 476028 12724 476080 12776
rect 490748 12792 490800 12844
rect 504272 12792 504324 12844
rect 561680 12792 561732 12844
rect 564440 12792 564492 12844
rect 395988 12656 396040 12708
rect 409144 12588 409196 12640
rect 415308 12588 415360 12640
rect 421564 12656 421616 12708
rect 427084 12656 427136 12708
rect 428004 12656 428056 12708
rect 444380 12656 444432 12708
rect 422300 12520 422352 12572
rect 444380 12520 444432 12572
rect 489644 12656 489696 12708
rect 499672 12724 499724 12776
rect 500776 12656 500828 12708
rect 427084 12452 427136 12504
rect 428004 12452 428056 12504
rect 447048 12452 447100 12504
rect 466184 12588 466236 12640
rect 471888 12588 471940 12640
rect 476028 12588 476080 12640
rect 320456 12384 320508 12436
rect 476672 12384 476724 12436
rect 313372 12316 313424 12368
rect 299112 12112 299164 12164
rect 316684 12248 316736 12300
rect 316960 12316 317012 12368
rect 475476 12316 475528 12368
rect 474372 12248 474424 12300
rect 484492 12248 484544 12300
rect 485044 12248 485096 12300
rect 306196 12180 306248 12232
rect 472072 12180 472124 12232
rect 473452 12180 473504 12232
rect 474004 12180 474056 12232
rect 501236 12180 501288 12232
rect 534908 12180 534960 12232
rect 302608 12112 302660 12164
rect 470876 12112 470928 12164
rect 484308 12112 484360 12164
rect 529204 12112 529256 12164
rect 325608 12044 325660 12096
rect 335360 12044 335412 12096
rect 342996 12044 343048 12096
rect 355324 12044 355376 12096
rect 364156 12044 364208 12096
rect 374644 12044 374696 12096
rect 384304 12044 384356 12096
rect 393964 12044 394016 12096
rect 403624 12044 403676 12096
rect 413284 12044 413336 12096
rect 422208 12044 422260 12096
rect 431960 12044 432012 12096
rect 442264 12044 442316 12096
rect 461492 12044 461544 12096
rect 295524 11976 295576 12028
rect 468576 12044 468628 12096
rect 478696 12044 478748 12096
rect 527272 12044 527324 12096
rect 291936 11908 291988 11960
rect 467472 11976 467524 12028
rect 473912 11976 473964 12028
rect 526076 11976 526128 12028
rect 472716 11908 472768 11960
rect 525432 11908 525484 11960
rect 46848 11840 46900 11892
rect 148048 11840 148100 11892
rect 288348 11840 288400 11892
rect 466276 11840 466328 11892
rect 470508 11840 470560 11892
rect 524972 11840 525024 11892
rect 27528 11772 27580 11824
rect 138112 11772 138164 11824
rect 284760 11772 284812 11824
rect 465172 11772 465224 11824
rect 466828 11772 466880 11824
rect 523776 11772 523828 11824
rect 529848 11772 529900 11824
rect 544108 11772 544160 11824
rect 133788 11704 133840 11756
rect 416044 11704 416096 11756
rect 416688 11704 416740 11756
rect 507308 11704 507360 11756
rect 526444 11704 526496 11756
rect 542176 11704 542228 11756
rect 556804 11704 556856 11756
rect 568580 11704 568632 11756
rect 324228 11636 324280 11688
rect 477500 11636 477552 11688
rect 483112 11636 483164 11688
rect 483664 11636 483716 11688
rect 512092 11636 512144 11688
rect 512920 11636 512972 11688
rect 316684 11568 316736 11620
rect 325608 11568 325660 11620
rect 335360 11568 335412 11620
rect 342996 11568 343048 11620
rect 349068 11568 349120 11620
rect 485872 11568 485924 11620
rect 336004 11500 336056 11552
rect 473176 11500 473228 11552
rect 355324 11432 355376 11484
rect 364156 11432 364208 11484
rect 374644 11432 374696 11484
rect 384304 11432 384356 11484
rect 400220 11432 400272 11484
rect 502340 11432 502392 11484
rect 393964 11364 394016 11416
rect 403624 11364 403676 11416
rect 409696 11364 409748 11416
rect 505376 11364 505428 11416
rect 413284 11296 413336 11348
rect 422208 11296 422260 11348
rect 425060 11296 425112 11348
rect 425520 11296 425572 11348
rect 434812 11296 434864 11348
rect 435732 11296 435784 11348
rect 468300 11296 468352 11348
rect 518440 11296 518492 11348
rect 431960 11228 432012 11280
rect 442264 11228 442316 11280
rect 461492 11228 461544 11280
rect 469772 11228 469824 11280
rect 441712 11024 441764 11076
rect 441988 11024 442040 11076
rect 281264 10956 281316 11008
rect 463976 10956 464028 11008
rect 489920 10956 489972 11008
rect 509148 10956 509200 11008
rect 263508 10888 263560 10940
rect 458272 10888 458324 10940
rect 506388 10888 506440 10940
rect 536472 10888 536524 10940
rect 253848 10820 253900 10872
rect 454776 10820 454828 10872
rect 474740 10820 474792 10872
rect 509240 10820 509292 10872
rect 249708 10752 249760 10804
rect 453672 10752 453724 10804
rect 487068 10752 487120 10804
rect 489920 10752 489972 10804
rect 509148 10752 509200 10804
rect 530308 10820 530360 10872
rect 245568 10684 245620 10736
rect 452476 10684 452528 10736
rect 452660 10684 452712 10736
rect 480444 10684 480496 10736
rect 481548 10684 481600 10736
rect 528376 10684 528428 10736
rect 240048 10616 240100 10668
rect 450544 10616 450596 10668
rect 456064 10616 456116 10668
rect 520280 10616 520332 10668
rect 235908 10548 235960 10600
rect 448796 10548 448848 10600
rect 452476 10548 452528 10600
rect 518900 10548 518952 10600
rect 231768 10480 231820 10532
rect 447600 10480 447652 10532
rect 448152 10480 448204 10532
rect 514944 10480 514996 10532
rect 86132 10412 86184 10464
rect 182272 10412 182324 10464
rect 229008 10412 229060 10464
rect 446772 10412 446824 10464
rect 448980 10412 449032 10464
rect 518072 10412 518124 10464
rect 31668 10344 31720 10396
rect 142252 10344 142304 10396
rect 220728 10344 220780 10396
rect 440424 10344 440476 10396
rect 440608 10344 440660 10396
rect 515404 10344 515456 10396
rect 9036 10276 9088 10328
rect 120080 10276 120132 10328
rect 135168 10276 135220 10328
rect 416872 10276 416924 10328
rect 417056 10276 417108 10328
rect 507676 10276 507728 10328
rect 522672 10276 522724 10328
rect 541808 10276 541860 10328
rect 322848 10208 322900 10260
rect 477040 10208 477092 10260
rect 352564 10140 352616 10192
rect 486976 10140 487028 10192
rect 364984 10072 365036 10124
rect 456340 10072 456392 10124
rect 418804 10004 418856 10056
rect 503076 10004 503128 10056
rect 338028 9936 338080 9988
rect 419540 9936 419592 9988
rect 442356 9936 442408 9988
rect 515772 9936 515824 9988
rect 445760 9868 445812 9920
rect 473544 9868 473596 9920
rect 450084 9800 450136 9852
rect 475844 9800 475896 9852
rect 208492 9664 208544 9716
rect 208768 9664 208820 9716
rect 376208 9664 376260 9716
rect 376392 9664 376444 9716
rect 451832 9664 451884 9716
rect 452108 9664 452160 9716
rect 458640 9664 458692 9716
rect 459008 9664 459060 9716
rect 459928 9664 459980 9716
rect 460572 9664 460624 9716
rect 470600 9664 470652 9716
rect 471244 9664 471296 9716
rect 471520 9664 471572 9716
rect 471980 9664 472032 9716
rect 472164 9664 472216 9716
rect 472808 9664 472860 9716
rect 497096 9664 497148 9716
rect 497740 9664 497792 9716
rect 530124 9664 530176 9716
rect 530676 9664 530728 9716
rect 202788 9596 202840 9648
rect 253756 9596 253808 9648
rect 455144 9596 455196 9648
rect 509240 9596 509292 9648
rect 517244 9596 517296 9648
rect 202512 9528 202564 9580
rect 228916 9528 228968 9580
rect 447140 9528 447192 9580
rect 218152 9460 218204 9512
rect 443644 9460 443696 9512
rect 454132 9460 454184 9512
rect 493140 9460 493192 9512
rect 204352 9392 204404 9444
rect 436468 9392 436520 9444
rect 439780 9392 439832 9444
rect 490840 9392 490892 9444
rect 510620 9392 510672 9444
rect 521844 9392 521896 9444
rect 203892 9324 203944 9376
rect 439044 9324 439096 9376
rect 445392 9324 445444 9376
rect 516876 9324 516928 9376
rect 186044 9256 186096 9308
rect 433340 9256 433392 9308
rect 438216 9256 438268 9308
rect 514576 9256 514628 9308
rect 514668 9256 514720 9308
rect 519544 9256 519596 9308
rect 531320 9256 531372 9308
rect 540888 9256 540940 9308
rect 541072 9256 541124 9308
rect 181352 9188 181404 9240
rect 431040 9188 431092 9240
rect 431132 9188 431184 9240
rect 512276 9188 512328 9240
rect 69480 9120 69532 9172
rect 169760 9120 169812 9172
rect 182548 9120 182600 9172
rect 432144 9120 432196 9172
rect 434628 9120 434680 9172
rect 513472 9120 513524 9172
rect 520280 9120 520332 9172
rect 531320 9120 531372 9172
rect 168196 9052 168248 9104
rect 427268 9052 427320 9104
rect 427544 9052 427596 9104
rect 511172 9052 511224 9104
rect 540888 9052 540940 9104
rect 151544 8984 151596 9036
rect 411260 8984 411312 9036
rect 414480 8984 414532 9036
rect 418528 8984 418580 9036
rect 419172 8984 419224 9036
rect 508504 8984 508556 9036
rect 519084 8984 519136 9036
rect 540704 8984 540756 9036
rect 23112 8916 23164 8968
rect 135260 8916 135312 8968
rect 156328 8916 156380 8968
rect 423772 8916 423824 8968
rect 426348 8916 426400 8968
rect 510804 8916 510856 8968
rect 513196 8916 513248 8968
rect 538772 8916 538824 8968
rect 334716 8848 334768 8900
rect 481272 8848 481324 8900
rect 345664 8780 345716 8832
rect 481640 8780 481692 8832
rect 510804 8780 510856 8832
rect 511816 8780 511868 8832
rect 399024 8712 399076 8764
rect 501972 8712 502024 8764
rect 412088 8644 412140 8696
rect 420920 8644 420972 8696
rect 422760 8644 422812 8696
rect 509608 8644 509660 8696
rect 371424 8576 371476 8628
rect 454040 8576 454092 8628
rect 433340 8508 433392 8560
rect 464344 8508 464396 8560
rect 307208 8304 307260 8356
rect 307392 8304 307444 8356
rect 384488 8304 384540 8356
rect 384672 8304 384724 8356
rect 372804 8236 372856 8288
rect 493508 8236 493560 8288
rect 369216 8168 369268 8220
rect 492404 8168 492456 8220
rect 113548 8100 113600 8152
rect 201592 8100 201644 8152
rect 365720 8100 365772 8152
rect 491208 8100 491260 8152
rect 117136 8032 117188 8084
rect 204260 8032 204312 8084
rect 362132 8032 362184 8084
rect 490104 8032 490156 8084
rect 109960 7964 110012 8016
rect 199200 7964 199252 8016
rect 358544 7964 358596 8016
rect 488908 7964 488960 8016
rect 102784 7896 102836 7948
rect 194692 7896 194744 7948
rect 354956 7896 355008 7948
rect 487804 7896 487856 7948
rect 99288 7828 99340 7880
rect 191840 7828 191892 7880
rect 351368 7828 351420 7880
rect 486608 7828 486660 7880
rect 493876 7828 493928 7880
rect 510344 7964 510396 8016
rect 509608 7828 509660 7880
rect 537576 7828 537628 7880
rect 92112 7760 92164 7812
rect 186320 7760 186372 7812
rect 347872 7760 347924 7812
rect 485504 7760 485556 7812
rect 490564 7760 490616 7812
rect 531504 7760 531556 7812
rect 34980 7692 35032 7744
rect 145012 7692 145064 7744
rect 344284 7692 344336 7744
rect 484032 7692 484084 7744
rect 489368 7692 489420 7744
rect 531044 7692 531096 7744
rect 18328 7624 18380 7676
rect 132592 7624 132644 7676
rect 285956 7624 286008 7676
rect 456800 7624 456852 7676
rect 456892 7624 456944 7676
rect 457628 7624 457680 7676
rect 485780 7624 485832 7676
rect 529940 7624 529992 7676
rect 13636 7556 13688 7608
rect 128544 7556 128596 7608
rect 159916 7556 159968 7608
rect 424876 7556 424928 7608
rect 426256 7556 426308 7608
rect 496544 7556 496596 7608
rect 504824 7556 504876 7608
rect 535828 7556 535880 7608
rect 383568 7488 383620 7540
rect 497004 7488 497056 7540
rect 408500 7420 408552 7472
rect 504732 7420 504784 7472
rect 413192 7352 413244 7404
rect 506572 7352 506624 7404
rect 340696 7284 340748 7336
rect 419632 7284 419684 7336
rect 420368 7284 420420 7336
rect 508872 7284 508924 7336
rect 385040 7216 385092 7268
rect 461216 7216 461268 7268
rect 437572 7148 437624 7200
rect 438032 7148 438084 7200
rect 448704 7148 448756 7200
rect 449624 7148 449676 7200
rect 456800 7148 456852 7200
rect 465540 7148 465592 7200
rect 429476 6876 429528 6928
rect 430120 6876 430172 6928
rect 476212 6876 476264 6928
rect 477224 6876 477276 6928
rect 67180 6808 67232 6860
rect 168380 6808 168432 6860
rect 297916 6808 297968 6860
rect 469404 6808 469456 6860
rect 493692 6808 493744 6860
rect 498936 6808 498988 6860
rect 63592 6740 63644 6792
rect 165620 6740 165672 6792
rect 294328 6740 294380 6792
rect 467932 6740 467984 6792
rect 502432 6740 502484 6792
rect 534356 6740 534408 6792
rect 60004 6672 60056 6724
rect 162860 6672 162912 6724
rect 290740 6672 290792 6724
rect 466920 6672 466972 6724
rect 498936 6672 498988 6724
rect 534172 6672 534224 6724
rect 52828 6604 52880 6656
rect 157340 6604 157392 6656
rect 287152 6604 287204 6656
rect 465632 6604 465684 6656
rect 495256 6604 495308 6656
rect 532884 6604 532936 6656
rect 56416 6536 56468 6588
rect 160100 6536 160152 6588
rect 283656 6536 283708 6588
rect 464436 6536 464488 6588
rect 491760 6536 491812 6588
rect 531688 6536 531740 6588
rect 49332 6468 49384 6520
rect 154580 6468 154632 6520
rect 279976 6468 280028 6520
rect 463332 6468 463384 6520
rect 488172 6468 488224 6520
rect 530124 6468 530176 6520
rect 44548 6400 44600 6452
rect 151820 6400 151872 6452
rect 276480 6400 276532 6452
rect 40960 6332 41012 6384
rect 149060 6332 149112 6384
rect 269304 6332 269356 6384
rect 459836 6332 459888 6384
rect 462320 6400 462372 6452
rect 484492 6400 484544 6452
rect 484584 6400 484636 6452
rect 528652 6400 528704 6452
rect 462412 6332 462464 6384
rect 479892 6332 479944 6384
rect 527732 6332 527784 6384
rect 37372 6264 37424 6316
rect 146300 6264 146352 6316
rect 161112 6264 161164 6316
rect 250536 6264 250588 6316
rect 261024 6264 261076 6316
rect 456984 6264 457036 6316
rect 476304 6264 476356 6316
rect 526628 6264 526680 6316
rect 8852 6196 8904 6248
rect 125600 6196 125652 6248
rect 221740 6196 221792 6248
rect 444656 6196 444708 6248
rect 463240 6196 463292 6248
rect 522396 6196 522448 6248
rect 4068 6128 4120 6180
rect 121644 6128 121696 6180
rect 206284 6128 206336 6180
rect 439596 6128 439648 6180
rect 459652 6128 459704 6180
rect 521200 6128 521252 6180
rect 70676 6060 70728 6112
rect 171140 6060 171192 6112
rect 301412 6060 301464 6112
rect 470232 6060 470284 6112
rect 74264 5992 74316 6044
rect 172612 5992 172664 6044
rect 327632 5992 327684 6044
rect 478972 5992 479024 6044
rect 77852 5924 77904 5976
rect 175556 5924 175608 5976
rect 353760 5924 353812 5976
rect 487160 5924 487212 5976
rect 356152 5856 356204 5908
rect 487252 5856 487304 5908
rect 394240 5788 394292 5840
rect 500132 5788 500184 5840
rect 439044 5720 439096 5772
rect 477592 5720 477644 5772
rect 457260 5652 457312 5704
rect 491944 5652 491996 5704
rect 455972 5584 456024 5636
rect 481732 5584 481784 5636
rect 535276 5584 535328 5636
rect 542728 5584 542780 5636
rect 570604 5516 570656 5568
rect 572628 5516 572680 5568
rect 108764 5448 108816 5500
rect 198740 5448 198792 5500
rect 263600 5448 263652 5500
rect 421104 5448 421156 5500
rect 437020 5448 437072 5500
rect 513564 5448 513616 5500
rect 101588 5380 101640 5432
rect 193220 5380 193272 5432
rect 303804 5380 303856 5432
rect 470600 5380 470652 5432
rect 508412 5380 508464 5432
rect 537024 5380 537076 5432
rect 98092 5312 98144 5364
rect 190460 5312 190512 5364
rect 256240 5312 256292 5364
rect 455788 5312 455840 5364
rect 465632 5312 465684 5364
rect 523132 5312 523184 5364
rect 94504 5244 94556 5296
rect 187700 5244 187752 5296
rect 255044 5244 255096 5296
rect 455512 5244 455564 5296
rect 462044 5244 462096 5296
rect 522028 5244 522080 5296
rect 87328 5176 87380 5228
rect 182180 5176 182232 5228
rect 236000 5176 236052 5228
rect 449164 5176 449216 5228
rect 458456 5176 458508 5228
rect 520924 5176 520976 5228
rect 90916 5108 90968 5160
rect 185124 5108 185176 5160
rect 230112 5108 230164 5160
rect 447416 5108 447468 5160
rect 454868 5108 454920 5160
rect 519636 5108 519688 5160
rect 83832 5040 83884 5092
rect 179512 5040 179564 5092
rect 226524 5040 226576 5092
rect 446128 5040 446180 5092
rect 451280 5040 451332 5092
rect 518624 5040 518676 5092
rect 80244 4972 80296 5024
rect 178040 4972 178092 5024
rect 219348 4972 219400 5024
rect 443828 4972 443880 5024
rect 447784 4972 447836 5024
rect 517612 4972 517664 5024
rect 76656 4904 76708 4956
rect 175280 4904 175332 4956
rect 215852 4904 215904 4956
rect 442724 4904 442776 4956
rect 443920 4904 443972 4956
rect 516324 4904 516376 4956
rect 73068 4836 73120 4888
rect 172520 4836 172572 4888
rect 178960 4836 179012 4888
rect 428464 4836 428516 4888
rect 433524 4836 433576 4888
rect 512092 4836 512144 4888
rect 515588 4836 515640 4888
rect 539232 4836 539284 4888
rect 12440 4768 12492 4820
rect 128360 4768 128412 4820
rect 167092 4768 167144 4820
rect 426532 4768 426584 4820
rect 429936 4768 429988 4820
rect 510804 4768 510856 4820
rect 512000 4768 512052 4820
rect 538404 4768 538456 4820
rect 105176 4700 105228 4752
rect 195980 4700 196032 4752
rect 331220 4700 331272 4752
rect 479064 4700 479116 4752
rect 482284 4700 482336 4752
rect 482928 4700 482980 4752
rect 120632 4632 120684 4684
rect 207020 4632 207072 4684
rect 375288 4632 375340 4684
rect 494152 4632 494204 4684
rect 123024 4564 123076 4616
rect 208768 4564 208820 4616
rect 403716 4564 403768 4616
rect 503168 4564 503220 4616
rect 378140 4496 378192 4548
rect 458364 4496 458416 4548
rect 469128 4496 469180 4548
rect 524604 4496 524656 4548
rect 411168 4428 411220 4480
rect 422300 4428 422352 4480
rect 427084 4428 427136 4480
rect 461768 4428 461820 4480
rect 384856 4360 384908 4412
rect 393228 4360 393280 4412
rect 443000 4360 443052 4412
rect 468668 4360 468720 4412
rect 1676 4088 1728 4140
rect 9036 4088 9088 4140
rect 81440 4088 81492 4140
rect 82728 4088 82780 4140
rect 84936 4088 84988 4140
rect 85488 4088 85540 4140
rect 88524 4088 88576 4140
rect 89628 4088 89680 4140
rect 93308 4088 93360 4140
rect 93768 4088 93820 4140
rect 95700 4088 95752 4140
rect 96528 4088 96580 4140
rect 103520 4088 103572 4140
rect 112996 4088 113048 4140
rect 121828 4088 121880 4140
rect 123484 4088 123536 4140
rect 137284 4088 137336 4140
rect 198188 4088 198240 4140
rect 200396 4088 200448 4140
rect 201408 4088 201460 4140
rect 214656 4088 214708 4140
rect 215208 4088 215260 4140
rect 271696 4088 271748 4140
rect 381176 4088 381228 4140
rect 382188 4088 382240 4140
rect 385040 4088 385092 4140
rect 111156 4020 111208 4072
rect 171600 4020 171652 4072
rect 171784 4020 171836 4072
rect 172428 4020 172480 4072
rect 198004 4020 198056 4072
rect 275284 4020 275336 4072
rect 277676 4020 277728 4072
rect 278688 4020 278740 4072
rect 278872 4020 278924 4072
rect 280068 4020 280120 4072
rect 293132 4020 293184 4072
rect 293868 4020 293920 4072
rect 300308 4020 300360 4072
rect 300768 4020 300820 4072
rect 313924 4020 313976 4072
rect 323032 4020 323084 4072
rect 325240 4020 325292 4072
rect 389272 4224 389324 4276
rect 387064 4088 387116 4140
rect 387708 4088 387760 4140
rect 389456 4088 389508 4140
rect 390468 4088 390520 4140
rect 395436 4088 395488 4140
rect 395988 4088 396040 4140
rect 396632 4088 396684 4140
rect 397368 4088 397420 4140
rect 397460 4088 397512 4140
rect 499764 4088 499816 4140
rect 516784 4088 516836 4140
rect 517428 4088 517480 4140
rect 525064 4088 525116 4140
rect 525708 4088 525760 4140
rect 527456 4088 527508 4140
rect 528468 4088 528520 4140
rect 533436 4088 533488 4140
rect 533988 4088 534040 4140
rect 542912 4088 542964 4140
rect 543648 4088 543700 4140
rect 558736 4088 558788 4140
rect 571432 4088 571484 4140
rect 389272 4020 389324 4072
rect 439044 4020 439096 4072
rect 441804 4020 441856 4072
rect 442356 4020 442408 4072
rect 446588 4020 446640 4072
rect 509240 4020 509292 4072
rect 557356 4020 557408 4072
rect 570236 4020 570288 4072
rect 39764 3952 39816 4004
rect 57244 3952 57296 4004
rect 103980 3952 104032 4004
rect 169024 3952 169076 4004
rect 172980 3952 173032 4004
rect 250444 3952 250496 4004
rect 250536 3952 250588 4004
rect 258448 3952 258500 4004
rect 258540 3952 258592 4004
rect 263600 3952 263652 4004
rect 267740 3952 267792 4004
rect 282736 3952 282788 4004
rect 305000 3952 305052 4004
rect 326344 3952 326396 4004
rect 17132 3884 17184 3936
rect 24124 3884 24176 3936
rect 32680 3884 32732 3936
rect 51724 3884 51776 3936
rect 96896 3884 96948 3936
rect 166264 3884 166316 3936
rect 196808 3884 196860 3936
rect 204352 3884 204404 3936
rect 208676 3884 208728 3936
rect 282828 3884 282880 3936
rect 282920 3884 282972 3936
rect 289820 3884 289872 3936
rect 309784 3884 309836 3936
rect 336004 3952 336056 4004
rect 339500 3952 339552 4004
rect 5264 3816 5316 3868
rect 61384 3816 61436 3868
rect 82636 3816 82688 3868
rect 6460 3748 6512 3800
rect 69664 3748 69716 3800
rect 89812 3816 89864 3868
rect 164884 3816 164936 3868
rect 209872 3816 209924 3868
rect 307760 3816 307812 3868
rect 318064 3816 318116 3868
rect 103520 3748 103572 3800
rect 112996 3748 113048 3800
rect 113180 3748 113232 3800
rect 122748 3748 122800 3800
rect 132500 3748 132552 3800
rect 145840 3748 145892 3800
rect 159364 3748 159416 3800
rect 165896 3748 165948 3800
rect 246304 3748 246356 3800
rect 252652 3748 252704 3800
rect 253848 3748 253900 3800
rect 258448 3748 258500 3800
rect 267740 3748 267792 3800
rect 307668 3748 307720 3800
rect 313924 3748 313976 3800
rect 46940 3680 46992 3732
rect 145932 3680 145984 3732
rect 149244 3680 149296 3732
rect 150348 3680 150400 3732
rect 153936 3680 153988 3732
rect 154488 3680 154540 3732
rect 174176 3680 174228 3732
rect 273168 3680 273220 3732
rect 321652 3680 321704 3732
rect 322848 3680 322900 3732
rect 323032 3816 323084 3868
rect 335268 3884 335320 3936
rect 337752 3884 337804 3936
rect 340144 3884 340196 3936
rect 340328 3952 340380 4004
rect 345664 3952 345716 4004
rect 346676 3952 346728 4004
rect 364340 3952 364392 4004
rect 370412 3952 370464 4004
rect 371148 3952 371200 4004
rect 374000 3952 374052 4004
rect 375196 3952 375248 4004
rect 377588 3952 377640 4004
rect 378048 3952 378100 4004
rect 378232 3952 378284 4004
rect 384304 3952 384356 4004
rect 393964 3952 394016 4004
rect 403624 3952 403676 4004
rect 404912 3952 404964 4004
rect 405648 3952 405700 4004
rect 406108 3952 406160 4004
rect 407028 3952 407080 4004
rect 407304 3952 407356 4004
rect 408408 3952 408460 4004
rect 413284 3952 413336 4004
rect 422300 3952 422352 4004
rect 431868 3952 431920 4004
rect 431960 3952 432012 4004
rect 439320 3952 439372 4004
rect 462320 3952 462372 4004
rect 464436 3952 464488 4004
rect 464988 3952 465040 4004
rect 492956 3952 493008 4004
rect 523960 3952 524012 4004
rect 535736 3952 535788 4004
rect 536748 3952 536800 4004
rect 558828 3952 558880 4004
rect 573824 3952 573876 4004
rect 455972 3884 456024 3936
rect 475108 3884 475160 3936
rect 526260 3884 526312 3936
rect 558644 3884 558696 3936
rect 575020 3884 575072 3936
rect 332416 3816 332468 3868
rect 452660 3816 452712 3868
rect 460848 3816 460900 3868
rect 510620 3816 510672 3868
rect 517888 3816 517940 3868
rect 527824 3816 527876 3868
rect 556988 3816 557040 3868
rect 559564 3816 559616 3868
rect 560024 3816 560076 3868
rect 576216 3816 576268 3868
rect 335268 3748 335320 3800
rect 371424 3748 371476 3800
rect 385868 3748 385920 3800
rect 497096 3748 497148 3800
rect 560116 3748 560168 3800
rect 577412 3748 577464 3800
rect 439596 3680 439648 3732
rect 469036 3680 469088 3732
rect 24308 3612 24360 3664
rect 25504 3612 25556 3664
rect 25596 3612 25648 3664
rect 32404 3612 32456 3664
rect 36176 3612 36228 3664
rect 16028 3544 16080 3596
rect 28264 3544 28316 3596
rect 29092 3544 29144 3596
rect 31024 3544 31076 3596
rect 33876 3544 33928 3596
rect 34428 3544 34480 3596
rect 42156 3544 42208 3596
rect 42708 3544 42760 3596
rect 43352 3612 43404 3664
rect 142804 3544 142856 3596
rect 150440 3612 150492 3664
rect 150532 3612 150584 3664
rect 153200 3612 153252 3664
rect 163504 3612 163556 3664
rect 164148 3612 164200 3664
rect 164700 3612 164752 3664
rect 165528 3612 165580 3664
rect 180156 3612 180208 3664
rect 180708 3612 180760 3664
rect 189632 3612 189684 3664
rect 190368 3612 190420 3664
rect 207480 3612 207532 3664
rect 289728 3612 289780 3664
rect 289912 3612 289964 3664
rect 337752 3612 337804 3664
rect 338304 3612 338356 3664
rect 339408 3612 339460 3664
rect 363328 3612 363380 3664
rect 364248 3612 364300 3664
rect 378876 3612 378928 3664
rect 434720 3612 434772 3664
rect 446404 3612 446456 3664
rect 455972 3612 456024 3664
rect 477500 3680 477552 3732
rect 478696 3680 478748 3732
rect 481088 3680 481140 3732
rect 481548 3680 481600 3732
rect 483020 3680 483072 3732
rect 471888 3612 471940 3664
rect 472072 3612 472124 3664
rect 10048 3476 10100 3528
rect 10968 3476 11020 3528
rect 11244 3476 11296 3528
rect 17132 3476 17184 3528
rect 17224 3476 17276 3528
rect 17868 3476 17920 3528
rect 25504 3476 25556 3528
rect 572 3408 624 3460
rect 10508 3408 10560 3460
rect 14832 3408 14884 3460
rect 20720 3340 20772 3392
rect 25596 3340 25648 3392
rect 45744 3340 45796 3392
rect 46848 3340 46900 3392
rect 50528 3340 50580 3392
rect 50988 3340 51040 3392
rect 51632 3340 51684 3392
rect 52368 3340 52420 3392
rect 54024 3340 54076 3392
rect 55128 3340 55180 3392
rect 55220 3340 55272 3392
rect 56508 3340 56560 3392
rect 58808 3340 58860 3392
rect 59268 3340 59320 3392
rect 61200 3340 61252 3392
rect 62028 3340 62080 3392
rect 62396 3340 62448 3392
rect 63408 3340 63460 3392
rect 68284 3340 68336 3392
rect 68928 3340 68980 3392
rect 71872 3340 71924 3392
rect 72976 3340 73028 3392
rect 79048 3340 79100 3392
rect 79968 3340 80020 3392
rect 106372 3340 106424 3392
rect 107476 3340 107528 3392
rect 112352 3340 112404 3392
rect 113088 3340 113140 3392
rect 114744 3340 114796 3392
rect 115848 3340 115900 3392
rect 119436 3340 119488 3392
rect 119988 3340 120040 3392
rect 113180 3272 113232 3324
rect 122748 3272 122800 3324
rect 124220 3408 124272 3460
rect 125508 3408 125560 3460
rect 129004 3408 129056 3460
rect 129648 3408 129700 3460
rect 130200 3408 130252 3460
rect 131028 3408 131080 3460
rect 131396 3408 131448 3460
rect 132408 3408 132460 3460
rect 125416 3340 125468 3392
rect 126244 3340 126296 3392
rect 132592 3476 132644 3528
rect 133788 3476 133840 3528
rect 136088 3476 136140 3528
rect 136548 3476 136600 3528
rect 139676 3476 139728 3528
rect 140688 3476 140740 3528
rect 138204 3340 138256 3392
rect 129832 3272 129884 3324
rect 132500 3272 132552 3324
rect 145840 3408 145892 3460
rect 146116 3408 146168 3460
rect 150532 3476 150584 3528
rect 148048 3408 148100 3460
rect 258540 3544 258592 3596
rect 258632 3544 258684 3596
rect 259368 3544 259420 3596
rect 267004 3544 267056 3596
rect 267648 3544 267700 3596
rect 268108 3544 268160 3596
rect 269028 3544 269080 3596
rect 282736 3544 282788 3596
rect 289636 3544 289688 3596
rect 298100 3544 298152 3596
rect 307668 3544 307720 3596
rect 316592 3544 316644 3596
rect 445760 3544 445812 3596
rect 461584 3544 461636 3596
rect 483480 3680 483532 3732
rect 484308 3680 484360 3732
rect 484400 3680 484452 3732
rect 495532 3612 495584 3664
rect 500316 3544 500368 3596
rect 505284 3544 505336 3596
rect 150716 3476 150768 3528
rect 384856 3476 384908 3528
rect 393044 3476 393096 3528
rect 397460 3476 397512 3528
rect 397828 3476 397880 3528
rect 398748 3476 398800 3528
rect 410892 3476 410944 3528
rect 483204 3476 483256 3528
rect 483388 3476 483440 3528
rect 155132 3408 155184 3460
rect 411168 3408 411220 3460
rect 415676 3408 415728 3460
rect 416688 3408 416740 3460
rect 423956 3408 424008 3460
rect 424968 3408 425020 3460
rect 428740 3408 428792 3460
rect 439504 3408 439556 3460
rect 439688 3408 439740 3460
rect 140872 3340 140924 3392
rect 146852 3272 146904 3324
rect 147588 3272 147640 3324
rect 150440 3272 150492 3324
rect 151728 3272 151780 3324
rect 191748 3340 191800 3392
rect 192024 3340 192076 3392
rect 193128 3340 193180 3392
rect 217048 3340 217100 3392
rect 217968 3340 218020 3392
rect 224132 3340 224184 3392
rect 224868 3340 224920 3392
rect 225328 3340 225380 3392
rect 226248 3340 226300 3392
rect 227720 3340 227772 3392
rect 229008 3340 229060 3392
rect 231308 3340 231360 3392
rect 231768 3340 231820 3392
rect 233700 3340 233752 3392
rect 234528 3340 234580 3392
rect 234804 3340 234856 3392
rect 235908 3340 235960 3392
rect 239588 3340 239640 3392
rect 240048 3340 240100 3392
rect 241980 3340 242032 3392
rect 242808 3340 242860 3392
rect 243176 3340 243228 3392
rect 244188 3340 244240 3392
rect 249156 3340 249208 3392
rect 249708 3340 249760 3392
rect 264612 3340 264664 3392
rect 378140 3340 378192 3392
rect 384304 3340 384356 3392
rect 393964 3340 394016 3392
rect 402520 3340 402572 3392
rect 418804 3340 418856 3392
rect 425152 3340 425204 3392
rect 444012 3340 444064 3392
rect 257436 3272 257488 3324
rect 364984 3272 365036 3324
rect 371608 3272 371660 3324
rect 439688 3272 439740 3324
rect 444288 3408 444340 3460
rect 483020 3408 483072 3460
rect 483572 3408 483624 3460
rect 444196 3340 444248 3392
rect 493876 3340 493928 3392
rect 494152 3408 494204 3460
rect 495348 3408 495400 3460
rect 507216 3476 507268 3528
rect 507768 3476 507820 3528
rect 510804 3476 510856 3528
rect 511908 3476 511960 3528
rect 514392 3544 514444 3596
rect 527916 3680 527968 3732
rect 560208 3680 560260 3732
rect 578608 3680 578660 3732
rect 521476 3612 521528 3664
rect 530584 3612 530636 3664
rect 561588 3612 561640 3664
rect 581000 3612 581052 3664
rect 523868 3544 523920 3596
rect 526444 3544 526496 3596
rect 536932 3544 536984 3596
rect 544384 3544 544436 3596
rect 554872 3544 554924 3596
rect 555976 3544 556028 3596
rect 556896 3544 556948 3596
rect 561956 3544 562008 3596
rect 563704 3544 563756 3596
rect 583392 3544 583444 3596
rect 514668 3476 514720 3528
rect 534540 3476 534592 3528
rect 535368 3476 535420 3528
rect 544108 3476 544160 3528
rect 545028 3476 545080 3528
rect 545304 3476 545356 3528
rect 546316 3476 546368 3528
rect 550088 3476 550140 3528
rect 550548 3476 550600 3528
rect 551836 3476 551888 3528
rect 552388 3476 552440 3528
rect 555516 3476 555568 3528
rect 557172 3476 557224 3528
rect 499120 3340 499172 3392
rect 500132 3408 500184 3460
rect 524972 3408 525024 3460
rect 526260 3408 526312 3460
rect 535276 3408 535328 3460
rect 539324 3408 539376 3460
rect 545764 3408 545816 3460
rect 556804 3408 556856 3460
rect 560760 3476 560812 3528
rect 563060 3476 563112 3528
rect 564348 3476 564400 3528
rect 561496 3408 561548 3460
rect 582196 3476 582248 3528
rect 564532 3408 564584 3460
rect 579804 3408 579856 3460
rect 500316 3340 500368 3392
rect 546500 3340 546552 3392
rect 547788 3340 547840 3392
rect 556068 3340 556120 3392
rect 566740 3340 566792 3392
rect 454132 3272 454184 3324
rect 467932 3272 467984 3324
rect 523776 3272 523828 3324
rect 532240 3272 532292 3324
rect 536104 3272 536156 3324
rect 557264 3272 557316 3324
rect 567844 3272 567896 3324
rect 7656 3204 7708 3256
rect 11704 3204 11756 3256
rect 144460 3204 144512 3256
rect 150716 3204 150768 3256
rect 205088 3204 205140 3256
rect 282184 3204 282236 3256
rect 289636 3204 289688 3256
rect 298008 3204 298060 3256
rect 310980 3204 311032 3256
rect 316592 3204 316644 3256
rect 328828 3204 328880 3256
rect 329748 3204 329800 3256
rect 330024 3204 330076 3256
rect 333244 3204 333296 3256
rect 335912 3204 335964 3256
rect 340328 3204 340380 3256
rect 364524 3204 364576 3256
rect 19524 3136 19576 3188
rect 22744 3136 22796 3188
rect 27896 3136 27948 3188
rect 28908 3136 28960 3188
rect 157524 3136 157576 3188
rect 158628 3136 158680 3188
rect 240784 3136 240836 3188
rect 311164 3136 311216 3188
rect 360936 3136 360988 3188
rect 421472 3136 421524 3188
rect 422300 3136 422352 3188
rect 431868 3136 431920 3188
rect 432328 3204 432380 3256
rect 433248 3204 433300 3256
rect 439780 3204 439832 3256
rect 444196 3204 444248 3256
rect 504364 3204 504416 3256
rect 540520 3204 540572 3256
rect 546592 3204 546644 3256
rect 435824 3136 435876 3188
rect 500224 3136 500276 3188
rect 528652 3136 528704 3188
rect 531964 3136 532016 3188
rect 559932 3136 559984 3188
rect 564532 3136 564584 3188
rect 364340 3068 364392 3120
rect 378232 3068 378284 3120
rect 388260 3068 388312 3120
rect 389088 3068 389140 3120
rect 403624 3068 403676 3120
rect 413284 3068 413336 3120
rect 421564 3068 421616 3120
rect 474740 3068 474792 3120
rect 2872 3000 2924 3052
rect 8944 3000 8996 3052
rect 26700 3000 26752 3052
rect 27528 3000 27580 3052
rect 190828 3000 190880 3052
rect 263600 3000 263652 3052
rect 337108 3000 337160 3052
rect 338028 3000 338080 3052
rect 382372 3000 382424 3052
rect 426256 3000 426308 3052
rect 431960 3000 432012 3052
rect 439320 3000 439372 3052
rect 439412 3000 439464 3052
rect 448152 3000 448204 3052
rect 450176 3000 450228 3052
rect 468300 3000 468352 3052
rect 158720 2932 158772 2984
rect 160008 2932 160060 2984
rect 251456 2932 251508 2984
rect 300768 2932 300820 2984
rect 319260 2932 319312 2984
rect 320088 2932 320140 2984
rect 115940 2864 115992 2916
rect 117228 2864 117280 2916
rect 183744 2864 183796 2916
rect 256700 2864 256752 2916
rect 343088 2864 343140 2916
rect 356060 2864 356112 2916
rect 369124 2864 369176 2916
rect 374092 2864 374144 2916
rect 262220 2796 262272 2848
rect 318708 2796 318760 2848
rect 378968 2796 379020 2848
rect 398840 2932 398892 2984
rect 412640 2932 412692 2984
rect 439596 2932 439648 2984
rect 450084 2932 450136 2984
rect 453672 2932 453724 2984
rect 461584 2932 461636 2984
rect 383660 2864 383712 2916
rect 383844 2864 383896 2916
rect 398748 2864 398800 2916
rect 541716 2864 541768 2916
rect 548064 2864 548116 2916
rect 555424 2864 555476 2916
rect 558368 2864 558420 2916
rect 414204 2796 414256 2848
rect 443000 2796 443052 2848
rect 444196 2796 444248 2848
rect 431960 2728 432012 2780
rect 441528 2728 441580 2780
rect 300768 2660 300820 2712
rect 454316 2660 454368 2712
rect 483112 2660 483164 2712
rect 333612 2592 333664 2644
rect 480352 2592 480404 2644
rect 308588 2524 308640 2576
rect 472164 2524 472216 2576
rect 274088 2456 274140 2508
rect 461308 2456 461360 2508
rect 244372 2388 244424 2440
rect 451556 2388 451608 2440
rect 237196 2320 237248 2372
rect 448704 2320 448756 2372
rect 201500 2252 201552 2304
rect 437572 2252 437624 2304
rect 194416 2184 194468 2236
rect 434812 2184 434864 2236
rect 162308 2116 162360 2168
rect 425060 2116 425112 2168
rect 431960 2116 432012 2168
rect 441528 2116 441580 2168
rect 133788 2048 133840 2100
rect 415584 2048 415636 2100
rect 417976 2048 418028 2100
rect 508044 2048 508096 2100
rect 345480 1980 345532 2032
rect 484676 1980 484728 2032
rect 318708 1912 318760 1964
rect 456892 1912 456944 1964
rect 379980 1844 380032 1896
rect 495716 1844 495768 1896
rect 390652 1776 390704 1828
rect 493692 1776 493744 1828
rect 401324 1708 401376 1760
rect 502616 1708 502668 1760
rect 263600 1640 263652 1692
rect 434996 1640 435048 1692
rect 366916 892 366968 944
rect 491484 892 491536 944
rect 341892 824 341944 876
rect 483296 824 483348 876
rect 326436 756 326488 808
rect 477684 756 477736 808
rect 322848 688 322900 740
rect 476212 688 476264 740
rect 315764 620 315816 672
rect 474924 620 474976 672
rect 202512 552 202564 604
rect 202696 552 202748 604
rect 220544 552 220596 604
rect 220728 552 220780 604
rect 259828 552 259880 604
rect 265808 552 265860 604
rect 270500 552 270552 604
rect 307300 552 307352 604
rect 307392 552 307444 604
rect 312176 552 312228 604
rect 473452 552 473504 604
rect 496544 552 496596 604
rect 496728 552 496780 604
rect 564440 552 564492 604
rect 565544 552 565596 604
rect 459836 484 459888 536
rect 458640 416 458692 468
rect 457076 348 457128 400
rect 213644 280 213696 332
rect 441620 280 441672 332
rect 199384 212 199436 264
rect 437664 212 437716 264
rect 195796 144 195848 196
rect 436100 144 436152 196
rect 188620 76 188672 128
rect 433800 76 433852 128
rect 170772 8 170824 60
rect 428096 8 428148 60
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700330 8156 703520
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 8944 700324 8996 700330
rect 8944 700266 8996 700272
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3528 681766 3556 682207
rect 3516 681760 3568 681766
rect 3516 681702 3568 681708
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 3422 624880 3478 624889
rect 3422 624815 3478 624824
rect 3330 610464 3386 610473
rect 3330 610399 3386 610408
rect 3344 610026 3372 610399
rect 3332 610020 3384 610026
rect 3332 609962 3384 609968
rect 3146 553072 3202 553081
rect 3146 553007 3202 553016
rect 3160 552090 3188 553007
rect 3148 552084 3200 552090
rect 3148 552026 3200 552032
rect 2870 509960 2926 509969
rect 2870 509895 2926 509904
rect 2884 509318 2912 509895
rect 2872 509312 2924 509318
rect 2872 509254 2924 509260
rect 3436 485110 3464 624815
rect 3514 596048 3570 596057
rect 3514 595983 3570 595992
rect 3528 594862 3556 595983
rect 3516 594856 3568 594862
rect 3516 594798 3568 594804
rect 3514 567352 3570 567361
rect 3514 567287 3570 567296
rect 3528 567254 3556 567287
rect 3516 567248 3568 567254
rect 3516 567190 3568 567196
rect 3514 538656 3570 538665
rect 3514 538591 3570 538600
rect 3528 538286 3556 538591
rect 3516 538280 3568 538286
rect 3516 538222 3568 538228
rect 3514 495544 3570 495553
rect 3514 495479 3516 495488
rect 3568 495479 3570 495488
rect 3516 495450 3568 495456
rect 3424 485104 3476 485110
rect 3424 485046 3476 485052
rect 3146 481128 3202 481137
rect 3146 481063 3202 481072
rect 3160 480282 3188 481063
rect 3148 480276 3200 480282
rect 3148 480218 3200 480224
rect 3422 452432 3478 452441
rect 3422 452367 3478 452376
rect 3436 451314 3464 452367
rect 3424 451308 3476 451314
rect 3424 451250 3476 451256
rect 3514 438016 3570 438025
rect 3514 437951 3570 437960
rect 3528 437510 3556 437951
rect 3516 437504 3568 437510
rect 3516 437446 3568 437452
rect 3422 423736 3478 423745
rect 3422 423671 3424 423680
rect 3476 423671 3478 423680
rect 3424 423642 3476 423648
rect 4802 395040 4858 395049
rect 4802 394975 4858 394984
rect 2778 380624 2834 380633
rect 2778 380559 2834 380568
rect 2792 366217 2820 380559
rect 2778 366208 2834 366217
rect 2778 366143 2834 366152
rect 2792 323105 2820 366143
rect 3146 337512 3202 337521
rect 3146 337447 3202 337456
rect 3160 336802 3188 337447
rect 3148 336796 3200 336802
rect 3148 336738 3200 336744
rect 2778 323096 2834 323105
rect 2778 323031 2834 323040
rect 2792 316742 2820 323031
rect 2780 316736 2832 316742
rect 2780 316678 2832 316684
rect 3424 316736 3476 316742
rect 3424 316678 3476 316684
rect 3436 309097 3464 316678
rect 2778 309088 2834 309097
rect 2778 309023 2834 309032
rect 3422 309088 3478 309097
rect 3422 309023 3478 309032
rect 2792 308825 2820 309023
rect 2778 308816 2834 308825
rect 2778 308751 2834 308760
rect 2792 280129 2820 308751
rect 3422 294400 3478 294409
rect 3422 294335 3478 294344
rect 3436 294030 3464 294335
rect 3424 294024 3476 294030
rect 3424 293966 3476 293972
rect 2778 280120 2834 280129
rect 2778 280055 2834 280064
rect 2792 265713 2820 280055
rect 2778 265704 2834 265713
rect 2778 265639 2834 265648
rect 2792 237017 2820 265639
rect 2778 237008 2834 237017
rect 2778 236943 2834 236952
rect 2792 222601 2820 236943
rect 2778 222592 2834 222601
rect 2778 222527 2834 222536
rect 2792 193905 2820 222527
rect 2778 193896 2834 193905
rect 2778 193831 2834 193840
rect 2792 179489 2820 193831
rect 2778 179480 2834 179489
rect 2778 179415 2834 179424
rect 2792 150793 2820 179415
rect 4816 173777 4844 394975
rect 6184 336796 6236 336802
rect 6184 336738 6236 336744
rect 4802 173768 4858 173777
rect 4802 173703 4858 173712
rect 2778 150784 2834 150793
rect 2778 150719 2834 150728
rect 2792 136377 2820 150719
rect 2778 136368 2834 136377
rect 2778 136303 2834 136312
rect 2792 107681 2820 136303
rect 2778 107672 2834 107681
rect 2778 107607 2834 107616
rect 2792 93265 2820 107607
rect 2778 93256 2834 93265
rect 2778 93191 2834 93200
rect 2792 64569 2820 93191
rect 6196 65521 6224 336738
rect 8956 125594 8984 700266
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 72988 700369 73016 703520
rect 41328 700334 41380 700340
rect 72974 700360 73030 700369
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 10324 652792 10376 652798
rect 10324 652734 10376 652740
rect 9036 594856 9088 594862
rect 9036 594798 9088 594804
rect 9048 128314 9076 594798
rect 9128 567248 9180 567254
rect 9128 567190 9180 567196
rect 9140 444378 9168 567190
rect 9128 444372 9180 444378
rect 9128 444314 9180 444320
rect 9128 220856 9180 220862
rect 9128 220798 9180 220804
rect 9036 128308 9088 128314
rect 9036 128250 9088 128256
rect 8944 125588 8996 125594
rect 8944 125530 8996 125536
rect 6182 65512 6238 65521
rect 6182 65447 6238 65456
rect 2778 64560 2834 64569
rect 2778 64495 2834 64504
rect 2792 50153 2820 64495
rect 2778 50144 2834 50153
rect 2778 50079 2834 50088
rect 2792 21457 2820 50079
rect 9140 35902 9168 220798
rect 10336 126954 10364 652734
rect 24780 621722 24808 699654
rect 41340 627230 41368 700334
rect 89180 700330 89208 703520
rect 72974 700295 73030 700304
rect 89168 700324 89220 700330
rect 89168 700266 89220 700272
rect 137848 696930 137876 703520
rect 154132 700398 154160 703520
rect 138664 700392 138716 700398
rect 138664 700334 138716 700340
rect 154120 700392 154172 700398
rect 154120 700334 154172 700340
rect 133144 696924 133196 696930
rect 133144 696866 133196 696872
rect 137836 696924 137888 696930
rect 137836 696866 137888 696872
rect 133156 675510 133184 696866
rect 122104 675504 122156 675510
rect 122104 675446 122156 675452
rect 133144 675504 133196 675510
rect 133144 675446 133196 675452
rect 122116 658578 122144 675446
rect 116584 658572 116636 658578
rect 116584 658514 116636 658520
rect 122104 658572 122156 658578
rect 122104 658514 122156 658520
rect 116596 648922 116624 658514
rect 113824 648916 113876 648922
rect 113824 648858 113876 648864
rect 116584 648916 116636 648922
rect 116584 648858 116636 648864
rect 113836 632466 113864 648858
rect 110420 632460 110472 632466
rect 110420 632402 110472 632408
rect 113824 632460 113876 632466
rect 113824 632402 113876 632408
rect 110432 629338 110460 632402
rect 105544 629332 105596 629338
rect 105544 629274 105596 629280
rect 110420 629332 110472 629338
rect 110420 629274 110472 629280
rect 41328 627224 41380 627230
rect 41328 627166 41380 627172
rect 105556 621790 105584 629274
rect 95884 621784 95936 621790
rect 95884 621726 95936 621732
rect 105544 621784 105596 621790
rect 105544 621726 105596 621732
rect 24768 621716 24820 621722
rect 24768 621658 24820 621664
rect 23388 619676 23440 619682
rect 23388 619618 23440 619624
rect 84108 619676 84160 619682
rect 84108 619618 84160 619624
rect 11704 610020 11756 610026
rect 11704 609962 11756 609968
rect 10416 538280 10468 538286
rect 10416 538222 10468 538228
rect 10428 129266 10456 538222
rect 11716 490618 11744 609962
rect 23296 605872 23348 605878
rect 23296 605814 23348 605820
rect 23204 571396 23256 571402
rect 23204 571338 23256 571344
rect 22100 530596 22152 530602
rect 22100 530538 22152 530544
rect 22112 528836 22140 530538
rect 23216 528850 23244 571338
rect 23308 530670 23336 605814
rect 23296 530664 23348 530670
rect 23296 530606 23348 530612
rect 23400 530602 23428 619618
rect 30194 617808 30250 617817
rect 30194 617743 30250 617752
rect 28630 616992 28686 617001
rect 28630 616927 28686 616936
rect 28644 616826 28672 616927
rect 28632 616820 28684 616826
rect 28632 616762 28684 616768
rect 28632 616616 28684 616622
rect 28630 616584 28632 616593
rect 28684 616584 28686 616593
rect 28630 616519 28686 616528
rect 30208 616486 30236 617743
rect 30286 617672 30342 617681
rect 84120 617658 84148 619618
rect 95896 619585 95924 621726
rect 91098 619576 91154 619585
rect 91098 619511 91154 619520
rect 95882 619576 95938 619585
rect 95882 619511 95938 619520
rect 84120 617630 84180 617658
rect 30286 617607 30342 617616
rect 30300 616622 30328 617607
rect 31482 617536 31538 617545
rect 91112 617506 91140 619511
rect 31482 617471 31484 617480
rect 31536 617471 31538 617480
rect 91100 617500 91152 617506
rect 31484 617442 31536 617448
rect 91100 617442 91152 617448
rect 30288 616616 30340 616622
rect 30288 616558 30340 616564
rect 28632 616480 28684 616486
rect 28632 616422 28684 616428
rect 30196 616480 30248 616486
rect 30196 616422 30248 616428
rect 28644 615913 28672 616422
rect 28630 615904 28686 615913
rect 28630 615839 28686 615848
rect 28264 615732 28316 615738
rect 28264 615674 28316 615680
rect 27526 608968 27582 608977
rect 27526 608903 27582 608912
rect 27434 607744 27490 607753
rect 27434 607679 27490 607688
rect 25226 606656 25282 606665
rect 25226 606591 25282 606600
rect 25240 605878 25268 606591
rect 25228 605872 25280 605878
rect 25228 605814 25280 605820
rect 24124 603492 24176 603498
rect 24124 603434 24176 603440
rect 24136 571985 24164 603434
rect 27342 602440 27398 602449
rect 27342 602375 27398 602384
rect 24766 601760 24822 601769
rect 24766 601695 24822 601704
rect 24674 583808 24730 583817
rect 24674 583743 24730 583752
rect 24582 572928 24638 572937
rect 24582 572863 24638 572872
rect 24490 572384 24546 572393
rect 24490 572319 24546 572328
rect 24122 571976 24178 571985
rect 24122 571911 24178 571920
rect 23388 530596 23440 530602
rect 23388 530538 23440 530544
rect 24504 528850 24532 572319
rect 24596 531146 24624 572863
rect 24584 531140 24636 531146
rect 24584 531082 24636 531088
rect 24688 530534 24716 583743
rect 24780 530670 24808 601695
rect 27250 599992 27306 600001
rect 27250 599927 27306 599936
rect 25778 598768 25834 598777
rect 25778 598703 25834 598712
rect 25226 596456 25282 596465
rect 25226 596391 25282 596400
rect 25134 582584 25190 582593
rect 25134 582519 25190 582528
rect 25042 577144 25098 577153
rect 25042 577079 25098 577088
rect 24950 575376 25006 575385
rect 24950 575311 25006 575320
rect 24768 530664 24820 530670
rect 24768 530606 24820 530612
rect 24676 530528 24728 530534
rect 24676 530470 24728 530476
rect 24964 530194 24992 575311
rect 25056 530398 25084 577079
rect 25148 572150 25176 582519
rect 25136 572144 25188 572150
rect 25136 572086 25188 572092
rect 25240 530738 25268 596391
rect 25318 587752 25374 587761
rect 25318 587687 25374 587696
rect 25332 570625 25360 587687
rect 25686 580816 25742 580825
rect 25686 580751 25742 580760
rect 25410 578368 25466 578377
rect 25410 578303 25466 578312
rect 25318 570616 25374 570625
rect 25318 570551 25374 570560
rect 25424 534954 25452 578303
rect 25502 574152 25558 574161
rect 25502 574087 25558 574096
rect 25412 534948 25464 534954
rect 25412 534890 25464 534896
rect 25516 531146 25544 574087
rect 25594 571840 25650 571849
rect 25594 571775 25650 571784
rect 25608 571402 25636 571775
rect 25596 571396 25648 571402
rect 25596 571338 25648 571344
rect 25700 534886 25728 580751
rect 25792 569294 25820 598703
rect 27158 597544 27214 597553
rect 27158 597479 27214 597488
rect 27066 595232 27122 595241
rect 27066 595167 27122 595176
rect 26054 591560 26110 591569
rect 26054 591495 26110 591504
rect 25962 586800 26018 586809
rect 25962 586735 26018 586744
rect 25870 583128 25926 583137
rect 25870 583063 25926 583072
rect 25780 569288 25832 569294
rect 25780 569230 25832 569236
rect 25688 534880 25740 534886
rect 25688 534822 25740 534828
rect 25884 534750 25912 583063
rect 25872 534744 25924 534750
rect 25872 534686 25924 534692
rect 25976 533798 26004 586735
rect 25964 533792 26016 533798
rect 25964 533734 26016 533740
rect 26068 533662 26096 591495
rect 26974 590336 27030 590345
rect 26974 590271 27030 590280
rect 26882 585576 26938 585585
rect 26882 585511 26938 585520
rect 26146 585032 26202 585041
rect 26146 584967 26202 584976
rect 26160 579222 26188 584967
rect 26606 580136 26662 580145
rect 26606 580071 26662 580080
rect 26148 579216 26200 579222
rect 26148 579158 26200 579164
rect 26146 578912 26202 578921
rect 26146 578847 26202 578856
rect 26160 547534 26188 578847
rect 26330 573608 26386 573617
rect 26330 573543 26386 573552
rect 26148 547528 26200 547534
rect 26148 547470 26200 547476
rect 26056 533656 26108 533662
rect 26056 533598 26108 533604
rect 25320 531140 25372 531146
rect 25320 531082 25372 531088
rect 25504 531140 25556 531146
rect 25504 531082 25556 531088
rect 25228 530732 25280 530738
rect 25228 530674 25280 530680
rect 25044 530392 25096 530398
rect 25044 530334 25096 530340
rect 24952 530188 25004 530194
rect 24952 530130 25004 530136
rect 23138 528822 23244 528850
rect 24242 528822 24532 528850
rect 25332 528836 25360 531082
rect 26344 528836 26372 573543
rect 26620 571538 26648 580071
rect 26698 577824 26754 577833
rect 26698 577759 26754 577768
rect 26712 571606 26740 577759
rect 26790 576600 26846 576609
rect 26790 576535 26846 576544
rect 26804 571674 26832 576535
rect 26792 571668 26844 571674
rect 26792 571610 26844 571616
rect 26700 571600 26752 571606
rect 26700 571542 26752 571548
rect 26608 571532 26660 571538
rect 26608 571474 26660 571480
rect 26896 547466 26924 585511
rect 26884 547460 26936 547466
rect 26884 547402 26936 547408
rect 26988 547398 27016 590271
rect 26976 547392 27028 547398
rect 26976 547334 27028 547340
rect 27080 547262 27108 595167
rect 27068 547256 27120 547262
rect 27068 547198 27120 547204
rect 27172 533594 27200 597479
rect 27160 533588 27212 533594
rect 27160 533530 27212 533536
rect 27264 533526 27292 599927
rect 27252 533520 27304 533526
rect 27252 533462 27304 533468
rect 27356 533458 27384 602375
rect 27344 533452 27396 533458
rect 27344 533394 27396 533400
rect 27448 532098 27476 607679
rect 27436 532092 27488 532098
rect 27436 532034 27488 532040
rect 27540 532030 27568 608903
rect 27986 603800 28042 603809
rect 27986 603735 28042 603744
rect 27618 603664 27674 603673
rect 27618 603599 27674 603608
rect 27632 533390 27660 603599
rect 27710 597000 27766 597009
rect 27710 596935 27766 596944
rect 27620 533384 27672 533390
rect 27620 533326 27672 533332
rect 27528 532024 27580 532030
rect 27528 531966 27580 531972
rect 27436 531140 27488 531146
rect 27436 531082 27488 531088
rect 27448 528836 27476 531082
rect 27724 530806 27752 596935
rect 27802 593328 27858 593337
rect 27802 593263 27858 593272
rect 27816 531010 27844 593263
rect 27894 590744 27950 590753
rect 27894 590679 27950 590688
rect 27908 531146 27936 590679
rect 28000 547194 28028 603735
rect 28276 603498 28304 615674
rect 28354 604888 28410 604897
rect 28354 604823 28410 604832
rect 28264 603492 28316 603498
rect 28264 603434 28316 603440
rect 28368 596737 28396 604823
rect 28538 600128 28594 600137
rect 28538 600063 28594 600072
rect 28446 599040 28502 599049
rect 28446 598975 28502 598984
rect 28354 596728 28410 596737
rect 28354 596663 28410 596672
rect 28262 595368 28318 595377
rect 28262 595303 28318 595312
rect 28170 593464 28226 593473
rect 28170 593399 28226 593408
rect 28078 591696 28134 591705
rect 28078 591631 28134 591640
rect 28092 586702 28120 591631
rect 28080 586696 28132 586702
rect 28080 586638 28132 586644
rect 28078 581496 28134 581505
rect 28078 581431 28134 581440
rect 27988 547188 28040 547194
rect 27988 547130 28040 547136
rect 28092 534818 28120 581431
rect 28184 547330 28212 593399
rect 28276 585614 28304 595303
rect 28354 594688 28410 594697
rect 28354 594623 28410 594632
rect 28368 591977 28396 594623
rect 28354 591968 28410 591977
rect 28354 591903 28410 591912
rect 28354 588704 28410 588713
rect 28354 588639 28410 588648
rect 28264 585608 28316 585614
rect 28264 585550 28316 585556
rect 28262 579048 28318 579057
rect 28262 578983 28318 578992
rect 28276 576178 28304 578983
rect 28368 578814 28396 588639
rect 28356 578808 28408 578814
rect 28356 578750 28408 578756
rect 28276 576150 28396 576178
rect 28262 575648 28318 575657
rect 28262 575583 28264 575592
rect 28316 575583 28318 575592
rect 28264 575554 28316 575560
rect 28262 574288 28318 574297
rect 28262 574223 28318 574232
rect 28172 547324 28224 547330
rect 28172 547266 28224 547272
rect 28080 534812 28132 534818
rect 28080 534754 28132 534760
rect 27896 531140 27948 531146
rect 27896 531082 27948 531088
rect 27804 531004 27856 531010
rect 27804 530946 27856 530952
rect 27712 530800 27764 530806
rect 27712 530742 27764 530748
rect 28276 528850 28304 574223
rect 28368 535022 28396 576150
rect 28460 569362 28488 598975
rect 28552 593473 28580 600063
rect 28630 598360 28686 598369
rect 28630 598295 28686 598304
rect 28644 594250 28672 598295
rect 28632 594244 28684 594250
rect 28632 594186 28684 594192
rect 28630 594144 28686 594153
rect 28686 594102 30328 594130
rect 28630 594079 28686 594088
rect 28632 594040 28684 594046
rect 28632 593982 28684 593988
rect 28538 593464 28594 593473
rect 28538 593399 28594 593408
rect 28644 592498 28672 593982
rect 28552 592470 28672 592498
rect 28552 591297 28580 592470
rect 28630 592376 28686 592385
rect 28686 592334 28764 592362
rect 28630 592311 28686 592320
rect 28538 591288 28594 591297
rect 28538 591223 28594 591232
rect 28630 589384 28686 589393
rect 28630 589319 28686 589328
rect 28538 588160 28594 588169
rect 28538 588095 28594 588104
rect 28552 583778 28580 588095
rect 28644 587858 28672 589319
rect 28736 587858 28764 592334
rect 28632 587852 28684 587858
rect 28632 587794 28684 587800
rect 28724 587852 28776 587858
rect 28724 587794 28776 587800
rect 28630 587752 28686 587761
rect 28686 587710 30236 587738
rect 28630 587687 28686 587696
rect 28630 587480 28686 587489
rect 28686 587438 29776 587466
rect 28630 587415 28686 587424
rect 28816 587376 28868 587382
rect 28816 587318 28868 587324
rect 28908 587376 28960 587382
rect 28960 587336 29592 587364
rect 28908 587318 28960 587324
rect 28828 586922 28856 587318
rect 29564 587058 29592 587336
rect 29748 587194 29776 587438
rect 29748 587166 30144 587194
rect 29564 587030 30052 587058
rect 28828 586894 29776 586922
rect 28908 586696 28960 586702
rect 28908 586638 28960 586644
rect 28920 585970 28948 586638
rect 28920 585942 29592 585970
rect 28630 585712 28686 585721
rect 28686 585670 28764 585698
rect 28630 585647 28686 585656
rect 28736 585018 28764 585670
rect 28816 585608 28868 585614
rect 28868 585556 29224 585562
rect 28816 585550 29224 585556
rect 28828 585534 29224 585550
rect 28736 584990 29132 585018
rect 28630 583944 28686 583953
rect 28630 583879 28686 583888
rect 28540 583772 28592 583778
rect 28540 583714 28592 583720
rect 28538 580952 28594 580961
rect 28538 580887 28594 580896
rect 28552 578950 28580 580887
rect 28540 578944 28592 578950
rect 28540 578886 28592 578892
rect 28540 578808 28592 578814
rect 28540 578750 28592 578756
rect 28552 570654 28580 578750
rect 28644 570858 28672 583879
rect 29000 583772 29052 583778
rect 29000 583714 29052 583720
rect 29012 579306 29040 583714
rect 29104 582434 29132 584990
rect 29196 584066 29224 585534
rect 29564 584610 29592 585942
rect 29748 584746 29776 586894
rect 29748 584718 29960 584746
rect 29564 584582 29868 584610
rect 29196 584038 29684 584066
rect 29104 582406 29224 582434
rect 29196 579442 29224 582406
rect 29196 579414 29316 579442
rect 29012 579278 29224 579306
rect 28908 579216 28960 579222
rect 28960 579164 29132 579170
rect 28908 579158 29132 579164
rect 28920 579142 29132 579158
rect 28724 578944 28776 578950
rect 28724 578886 28776 578892
rect 28736 573306 28764 578886
rect 28908 575612 28960 575618
rect 28908 575554 28960 575560
rect 28920 575498 28948 575554
rect 28920 575470 29040 575498
rect 28724 573300 28776 573306
rect 28724 573242 28776 573248
rect 29012 571470 29040 575470
rect 29000 571464 29052 571470
rect 29000 571406 29052 571412
rect 28632 570852 28684 570858
rect 28632 570794 28684 570800
rect 28540 570648 28592 570654
rect 28540 570590 28592 570596
rect 28448 569356 28500 569362
rect 28448 569298 28500 569304
rect 29104 567662 29132 579142
rect 29196 573510 29224 579278
rect 29184 573504 29236 573510
rect 29184 573446 29236 573452
rect 29288 573322 29316 579414
rect 29460 573504 29512 573510
rect 29460 573446 29512 573452
rect 29196 573294 29316 573322
rect 29196 570790 29224 573294
rect 29184 570784 29236 570790
rect 29184 570726 29236 570732
rect 29472 570722 29500 573446
rect 29552 573436 29604 573442
rect 29552 573378 29604 573384
rect 29564 572762 29592 573378
rect 29552 572756 29604 572762
rect 29552 572698 29604 572704
rect 29460 570716 29512 570722
rect 29460 570658 29512 570664
rect 29184 569900 29236 569906
rect 29184 569842 29236 569848
rect 29092 567656 29144 567662
rect 29092 567598 29144 567604
rect 29090 567488 29146 567497
rect 29090 567423 29146 567432
rect 29104 558385 29132 567423
rect 29196 560318 29224 569842
rect 29656 567882 29684 584038
rect 29736 572756 29788 572762
rect 29736 572698 29788 572704
rect 29748 569906 29776 572698
rect 29736 569900 29788 569906
rect 29736 569842 29788 569848
rect 29380 567854 29684 567882
rect 29276 565752 29328 565758
rect 29276 565694 29328 565700
rect 29184 560312 29236 560318
rect 29184 560254 29236 560260
rect 29090 558376 29146 558385
rect 29090 558311 29146 558320
rect 29288 553450 29316 565694
rect 29380 558550 29408 567854
rect 29460 567656 29512 567662
rect 29460 567598 29512 567604
rect 29368 558544 29420 558550
rect 29368 558486 29420 558492
rect 29472 558090 29500 567598
rect 29552 563236 29604 563242
rect 29552 563178 29604 563184
rect 29564 558210 29592 563178
rect 29736 560312 29788 560318
rect 29736 560254 29788 560260
rect 29644 558544 29696 558550
rect 29644 558486 29696 558492
rect 29552 558204 29604 558210
rect 29552 558146 29604 558152
rect 29472 558062 29592 558090
rect 29276 553444 29328 553450
rect 29276 553386 29328 553392
rect 29460 550588 29512 550594
rect 29460 550530 29512 550536
rect 29182 547632 29238 547641
rect 29182 547567 29238 547576
rect 28356 535016 28408 535022
rect 28356 534958 28408 534964
rect 29196 531593 29224 547567
rect 29368 543720 29420 543726
rect 29368 543662 29420 543668
rect 29276 538892 29328 538898
rect 29276 538834 29328 538840
rect 29182 531584 29238 531593
rect 29182 531519 29238 531528
rect 29288 530466 29316 538834
rect 29380 534138 29408 543662
rect 29472 541006 29500 550530
rect 29460 541000 29512 541006
rect 29460 540942 29512 540948
rect 29564 538898 29592 558062
rect 29552 538892 29604 538898
rect 29552 538834 29604 538840
rect 29656 536602 29684 558486
rect 29748 550594 29776 560254
rect 29736 550588 29788 550594
rect 29736 550530 29788 550536
rect 29736 541000 29788 541006
rect 29736 540942 29788 540948
rect 29564 536574 29684 536602
rect 29368 534132 29420 534138
rect 29368 534074 29420 534080
rect 29564 530874 29592 536574
rect 29748 530942 29776 540942
rect 29840 531078 29868 584582
rect 29932 531214 29960 584718
rect 30024 565758 30052 587030
rect 30012 565752 30064 565758
rect 30012 565694 30064 565700
rect 30010 557424 30066 557433
rect 30010 557359 30066 557368
rect 30024 557161 30052 557359
rect 30010 557152 30066 557161
rect 30010 557087 30066 557096
rect 30012 553444 30064 553450
rect 30012 553386 30064 553392
rect 30024 543726 30052 553386
rect 30012 543720 30064 543726
rect 30012 543662 30064 543668
rect 30012 534132 30064 534138
rect 30012 534074 30064 534080
rect 30024 533730 30052 534074
rect 30012 533724 30064 533730
rect 30012 533666 30064 533672
rect 30116 531282 30144 587166
rect 30208 533866 30236 587710
rect 30300 573510 30328 594102
rect 30288 573504 30340 573510
rect 30288 573446 30340 573452
rect 30288 573300 30340 573306
rect 30288 573242 30340 573248
rect 30300 563242 30328 573242
rect 31852 571668 31904 571674
rect 31852 571610 31904 571616
rect 30380 571464 30432 571470
rect 30380 571406 30432 571412
rect 30288 563236 30340 563242
rect 30288 563178 30340 563184
rect 30288 558204 30340 558210
rect 30288 558146 30340 558152
rect 30196 533860 30248 533866
rect 30196 533802 30248 533808
rect 30300 532166 30328 558146
rect 30288 532160 30340 532166
rect 30288 532102 30340 532108
rect 30104 531276 30156 531282
rect 30104 531218 30156 531224
rect 29920 531208 29972 531214
rect 29920 531150 29972 531156
rect 29828 531072 29880 531078
rect 29828 531014 29880 531020
rect 29736 530936 29788 530942
rect 29736 530878 29788 530884
rect 29552 530868 29604 530874
rect 29552 530810 29604 530816
rect 29276 530460 29328 530466
rect 29276 530402 29328 530408
rect 29644 530188 29696 530194
rect 29644 530130 29696 530136
rect 28276 528822 28566 528850
rect 29656 528836 29684 530130
rect 30392 528850 30420 571406
rect 30470 540968 30526 540977
rect 30470 540903 30526 540912
rect 30484 533633 30512 540903
rect 30470 533624 30526 533633
rect 30470 533559 30526 533568
rect 31864 528850 31892 571610
rect 33140 571600 33192 571606
rect 33140 571542 33192 571548
rect 41420 571600 41472 571606
rect 41420 571542 41472 571548
rect 32864 530392 32916 530398
rect 32864 530334 32916 530340
rect 30392 528822 30682 528850
rect 31786 528822 31892 528850
rect 32876 528836 32904 530334
rect 33152 528714 33180 571542
rect 37280 571464 37332 571470
rect 37280 571406 37332 571412
rect 35900 547528 35952 547534
rect 35900 547470 35952 547476
rect 34980 534948 35032 534954
rect 34980 534890 35032 534896
rect 34992 528836 35020 534890
rect 35912 528850 35940 547470
rect 37188 535016 37240 535022
rect 37188 534958 37240 534964
rect 35912 528822 36110 528850
rect 37200 528836 37228 534958
rect 37292 528986 37320 571406
rect 41432 534970 41460 571542
rect 56120 571526 56456 571554
rect 112240 571526 112576 571554
rect 45652 570852 45704 570858
rect 45652 570794 45704 570800
rect 41432 534942 42196 534970
rect 39304 534880 39356 534886
rect 39304 534822 39356 534828
rect 37292 528958 37964 528986
rect 37936 528850 37964 528958
rect 37936 528822 38226 528850
rect 39316 528836 39344 534822
rect 41420 534812 41472 534818
rect 41420 534754 41472 534760
rect 40408 532160 40460 532166
rect 40408 532102 40460 532108
rect 40420 528836 40448 532102
rect 41432 528836 41460 534754
rect 42168 528850 42196 534942
rect 43628 534744 43680 534750
rect 43628 534686 43680 534692
rect 42168 528822 42550 528850
rect 43640 528836 43668 534686
rect 44732 530528 44784 530534
rect 44732 530470 44784 530476
rect 44744 528836 44772 530470
rect 45664 528850 45692 570794
rect 48320 570784 48372 570790
rect 48320 570726 48372 570732
rect 46940 547460 46992 547466
rect 46940 547402 46992 547408
rect 46848 530460 46900 530466
rect 46848 530402 46900 530408
rect 45664 528822 45770 528850
rect 46860 528836 46888 530402
rect 46952 528986 46980 547402
rect 48332 528986 48360 570726
rect 52460 570716 52512 570722
rect 52460 570658 52512 570664
rect 52276 533860 52328 533866
rect 52276 533802 52328 533808
rect 50068 533792 50120 533798
rect 50068 533734 50120 533740
rect 46952 528958 47716 528986
rect 48332 528958 48636 528986
rect 47688 528850 47716 528958
rect 48608 528850 48636 528958
rect 47688 528822 47978 528850
rect 48608 528822 48990 528850
rect 50080 528836 50108 533734
rect 51172 531276 51224 531282
rect 51172 531218 51224 531224
rect 51184 528836 51212 531218
rect 52288 528836 52316 533802
rect 52472 528986 52500 570658
rect 53840 570648 53892 570654
rect 53840 570590 53892 570596
rect 53852 528986 53880 570590
rect 56428 569226 56456 571526
rect 76010 570616 76066 570625
rect 76010 570551 76066 570560
rect 71780 569356 71832 569362
rect 71780 569298 71832 569304
rect 70400 569288 70452 569294
rect 70400 569230 70452 569236
rect 56416 569220 56468 569226
rect 56416 569162 56468 569168
rect 55312 547392 55364 547398
rect 55312 547334 55364 547340
rect 55324 531298 55352 547334
rect 62120 547324 62172 547330
rect 62120 547266 62172 547272
rect 60832 533724 60884 533730
rect 60832 533666 60884 533672
rect 58716 533656 58768 533662
rect 58716 533598 58768 533604
rect 55324 531270 56180 531298
rect 55496 531208 55548 531214
rect 55496 531150 55548 531156
rect 52472 528958 53052 528986
rect 53852 528958 54156 528986
rect 53024 528850 53052 528958
rect 54128 528850 54156 528958
rect 53024 528822 53314 528850
rect 54128 528822 54418 528850
rect 55508 528836 55536 531150
rect 56152 528850 56180 531270
rect 57612 531140 57664 531146
rect 57612 531082 57664 531088
rect 56152 528822 56534 528850
rect 57624 528836 57652 531082
rect 58728 528836 58756 533598
rect 59820 531072 59872 531078
rect 59820 531014 59872 531020
rect 59832 528836 59860 531014
rect 60844 528836 60872 533666
rect 61936 531004 61988 531010
rect 61936 530946 61988 530952
rect 61948 528836 61976 530946
rect 62132 528986 62160 547266
rect 64880 547256 64932 547262
rect 64880 547198 64932 547204
rect 64052 530936 64104 530942
rect 64052 530878 64104 530884
rect 62132 528958 62804 528986
rect 62776 528850 62804 528958
rect 62776 528822 63066 528850
rect 64064 528836 64092 530878
rect 64892 528850 64920 547198
rect 69480 533588 69532 533594
rect 69480 533530 69532 533536
rect 66260 530868 66312 530874
rect 66260 530810 66312 530816
rect 64892 528822 65182 528850
rect 66272 528836 66300 530810
rect 68376 530800 68428 530806
rect 68376 530742 68428 530748
rect 67364 530732 67416 530738
rect 67364 530674 67416 530680
rect 67376 528836 67404 530674
rect 68388 528836 68416 530742
rect 69492 528836 69520 533530
rect 70412 531026 70440 569230
rect 70412 530998 71268 531026
rect 70582 530904 70638 530913
rect 70582 530839 70638 530848
rect 70596 528836 70624 530839
rect 71240 528850 71268 530998
rect 71792 529938 71820 569298
rect 73804 533520 73856 533526
rect 73804 533462 73856 533468
rect 71792 529910 72372 529938
rect 72344 528850 72372 529910
rect 71240 528822 71622 528850
rect 72344 528822 72726 528850
rect 73816 528836 73844 533462
rect 74906 531720 74962 531729
rect 74906 531655 74962 531664
rect 74920 528836 74948 531655
rect 76024 528850 76052 570551
rect 112548 569906 112576 571526
rect 138676 569906 138704 700334
rect 202800 700330 202828 703520
rect 138756 700324 138808 700330
rect 138756 700266 138808 700272
rect 202788 700324 202840 700330
rect 202788 700266 202840 700272
rect 138768 605826 138796 700266
rect 218992 694210 219020 703520
rect 267660 700330 267688 703520
rect 283852 703474 283880 703520
rect 283852 703446 283972 703474
rect 250904 700324 250956 700330
rect 250904 700266 250956 700272
rect 267648 700324 267700 700330
rect 267648 700266 267700 700272
rect 282276 700324 282328 700330
rect 282276 700266 282328 700272
rect 250916 699174 250944 700266
rect 250904 699168 250956 699174
rect 250904 699110 250956 699116
rect 253204 699168 253256 699174
rect 253204 699110 253256 699116
rect 253216 696930 253244 699110
rect 253204 696924 253256 696930
rect 253204 696866 253256 696872
rect 260012 696924 260064 696930
rect 260012 696866 260064 696872
rect 260024 694822 260052 696866
rect 260012 694816 260064 694822
rect 260012 694758 260064 694764
rect 267004 694816 267056 694822
rect 267004 694758 267056 694764
rect 218980 694204 219032 694210
rect 218980 694146 219032 694152
rect 219164 694204 219216 694210
rect 219164 694146 219216 694152
rect 219176 688702 219204 694146
rect 219164 688696 219216 688702
rect 219164 688638 219216 688644
rect 219072 688628 219124 688634
rect 219072 688570 219124 688576
rect 219084 679153 219112 688570
rect 219070 679144 219126 679153
rect 219070 679079 219126 679088
rect 218978 676288 219034 676297
rect 218978 676223 219034 676232
rect 218992 676190 219020 676223
rect 218796 676184 218848 676190
rect 218796 676126 218848 676132
rect 218980 676184 219032 676190
rect 218980 676126 219032 676132
rect 218808 666602 218836 676126
rect 267016 670682 267044 694758
rect 267004 670676 267056 670682
rect 267004 670618 267056 670624
rect 268384 670676 268436 670682
rect 268384 670618 268436 670624
rect 218796 666596 218848 666602
rect 218796 666538 218848 666544
rect 219072 666596 219124 666602
rect 219072 666538 219124 666544
rect 219084 659682 219112 666538
rect 268396 661230 268424 670618
rect 268384 661224 268436 661230
rect 268384 661166 268436 661172
rect 270408 661224 270460 661230
rect 270408 661166 270460 661172
rect 219084 659666 219204 659682
rect 219084 659660 219216 659666
rect 219084 659654 219164 659660
rect 219164 659602 219216 659608
rect 219348 659660 219400 659666
rect 219348 659602 219400 659608
rect 219360 656878 219388 659602
rect 270420 656946 270448 661166
rect 270408 656940 270460 656946
rect 270408 656882 270460 656888
rect 219072 656872 219124 656878
rect 219072 656814 219124 656820
rect 219348 656872 219400 656878
rect 219348 656814 219400 656820
rect 273260 656872 273312 656878
rect 273260 656814 273312 656820
rect 219084 647290 219112 656814
rect 273272 654158 273300 656814
rect 273260 654152 273312 654158
rect 273260 654094 273312 654100
rect 276664 654084 276716 654090
rect 276664 654026 276716 654032
rect 219072 647284 219124 647290
rect 219072 647226 219124 647232
rect 219256 647284 219308 647290
rect 219256 647226 219308 647232
rect 219268 640422 219296 647226
rect 219256 640416 219308 640422
rect 219256 640358 219308 640364
rect 219072 640280 219124 640286
rect 219072 640222 219124 640228
rect 219084 637566 219112 640222
rect 219072 637560 219124 637566
rect 219072 637502 219124 637508
rect 219164 637560 219216 637566
rect 219164 637502 219216 637508
rect 219176 627978 219204 637502
rect 276676 635118 276704 654026
rect 276664 635112 276716 635118
rect 276664 635054 276716 635060
rect 278044 635112 278096 635118
rect 278044 635054 278096 635060
rect 219164 627972 219216 627978
rect 219164 627914 219216 627920
rect 219348 627972 219400 627978
rect 219348 627914 219400 627920
rect 219360 621042 219388 627914
rect 278056 626550 278084 635054
rect 278044 626544 278096 626550
rect 278044 626486 278096 626492
rect 279148 626544 279200 626550
rect 279148 626486 279200 626492
rect 219072 621036 219124 621042
rect 219072 620978 219124 620984
rect 219348 621036 219400 621042
rect 219348 620978 219400 620984
rect 219084 618934 219112 620978
rect 279160 619585 279188 626486
rect 279146 619576 279202 619585
rect 279146 619511 279202 619520
rect 219072 618928 219124 618934
rect 219072 618870 219124 618876
rect 138768 605798 138888 605826
rect 138860 605418 138888 605798
rect 138860 605390 139164 605418
rect 139136 594674 139164 605390
rect 139582 594824 139638 594833
rect 139582 594759 139638 594768
rect 139596 594726 139624 594759
rect 139216 594720 139268 594726
rect 139136 594668 139216 594674
rect 139136 594662 139268 594668
rect 139584 594720 139636 594726
rect 139584 594662 139636 594668
rect 139136 594646 139256 594662
rect 188048 574110 188384 574138
rect 189244 574110 189580 574138
rect 188356 572286 188384 574110
rect 189552 572354 189580 574110
rect 190288 574110 190440 574138
rect 191636 574110 191788 574138
rect 192924 574110 193168 574138
rect 194120 574110 194456 574138
rect 195316 574110 195652 574138
rect 196512 574110 196848 574138
rect 197800 574110 198136 574138
rect 198996 574110 199332 574138
rect 200192 574110 200528 574138
rect 189540 572348 189592 572354
rect 189540 572290 189592 572296
rect 188344 572280 188396 572286
rect 188344 572222 188396 572228
rect 190288 572082 190316 574110
rect 190276 572076 190328 572082
rect 190276 572018 190328 572024
rect 191760 571470 191788 574110
rect 191748 571464 191800 571470
rect 191748 571406 191800 571412
rect 193140 571402 193168 574110
rect 194428 571946 194456 574110
rect 194600 572280 194652 572286
rect 194600 572222 194652 572228
rect 194416 571940 194468 571946
rect 194416 571882 194468 571888
rect 193128 571396 193180 571402
rect 193128 571338 193180 571344
rect 112536 569900 112588 569906
rect 112536 569842 112588 569848
rect 138664 569900 138716 569906
rect 138664 569842 138716 569848
rect 80060 547188 80112 547194
rect 80060 547130 80112 547136
rect 78678 547088 78734 547097
rect 78678 547023 78734 547032
rect 78128 533452 78180 533458
rect 78128 533394 78180 533400
rect 77024 530664 77076 530670
rect 77024 530606 77076 530612
rect 75946 528822 76052 528850
rect 77036 528836 77064 530606
rect 78140 528836 78168 533394
rect 78692 528850 78720 547023
rect 80072 533474 80100 547130
rect 165436 537396 165488 537402
rect 165436 537338 165488 537344
rect 163228 537328 163280 537334
rect 163228 537270 163280 537276
rect 158904 537260 158956 537266
rect 158904 537202 158956 537208
rect 156788 537192 156840 537198
rect 156788 537134 156840 537140
rect 152464 537124 152516 537130
rect 152464 537066 152516 537072
rect 150348 537056 150400 537062
rect 150348 536998 150400 537004
rect 148140 536988 148192 536994
rect 148140 536930 148192 536936
rect 146024 536920 146076 536926
rect 146024 536862 146076 536868
rect 112628 536852 112680 536858
rect 112628 536794 112680 536800
rect 109316 535492 109368 535498
rect 109316 535434 109368 535440
rect 91006 534984 91062 534993
rect 91006 534919 91062 534928
rect 88890 534848 88946 534857
rect 88890 534783 88946 534792
rect 84566 533896 84622 533905
rect 84566 533831 84622 533840
rect 80072 533446 80836 533474
rect 80244 533384 80296 533390
rect 80244 533326 80296 533332
rect 78692 528822 79166 528850
rect 80256 528836 80284 533326
rect 80808 528714 80836 533446
rect 83462 531856 83518 531865
rect 83462 531791 83518 531800
rect 82450 530768 82506 530777
rect 82450 530703 82506 530712
rect 82464 528836 82492 530703
rect 83476 528836 83504 531791
rect 84580 528836 84608 533831
rect 86682 533760 86738 533769
rect 86682 533695 86738 533704
rect 85672 530596 85724 530602
rect 85672 530538 85724 530544
rect 85684 528836 85712 530538
rect 86696 528836 86724 533695
rect 87788 532092 87840 532098
rect 87788 532034 87840 532040
rect 87800 528836 87828 532034
rect 88904 528836 88932 534783
rect 89996 532024 90048 532030
rect 89996 531966 90048 531972
rect 90008 528836 90036 531966
rect 91020 528836 91048 534919
rect 93214 534712 93270 534721
rect 93214 534647 93270 534656
rect 92110 532672 92166 532681
rect 92110 532607 92166 532616
rect 92124 528836 92152 532607
rect 93228 528836 93256 534647
rect 101770 533624 101826 533633
rect 101770 533559 101826 533568
rect 94226 532536 94282 532545
rect 94226 532471 94282 532480
rect 94240 528836 94268 532471
rect 96434 532400 96490 532409
rect 96434 532335 96490 532344
rect 95330 531312 95386 531321
rect 95330 531247 95386 531256
rect 95344 528836 95372 531247
rect 96448 528836 96476 532335
rect 98550 532264 98606 532273
rect 98550 532199 98606 532208
rect 97538 530632 97594 530641
rect 97538 530567 97594 530576
rect 97552 528836 97580 530567
rect 98564 528836 98592 532199
rect 99654 532128 99710 532137
rect 99654 532063 99710 532072
rect 99668 528836 99696 532063
rect 100758 531992 100814 532001
rect 100758 531927 100814 531936
rect 100772 528836 100800 531927
rect 101784 528836 101812 533559
rect 102874 533488 102930 533497
rect 102874 533423 102930 533432
rect 102888 528836 102916 533423
rect 103978 533352 104034 533361
rect 103978 533287 104034 533296
rect 103992 528836 104020 533287
rect 105082 531312 105138 531321
rect 105082 531247 105138 531256
rect 105096 528836 105124 531247
rect 106094 529952 106150 529961
rect 106094 529887 106150 529896
rect 106108 528836 106136 529887
rect 109328 528836 109356 535434
rect 111522 531448 111578 531457
rect 111522 531383 111578 531392
rect 111536 528836 111564 531383
rect 112640 528836 112668 536794
rect 139492 535968 139544 535974
rect 139492 535910 139544 535916
rect 137376 535900 137428 535906
rect 137376 535842 137428 535848
rect 127716 535832 127768 535838
rect 127716 535774 127768 535780
rect 125508 535764 125560 535770
rect 125508 535706 125560 535712
rect 123392 535696 123444 535702
rect 123392 535638 123444 535644
rect 121184 535628 121236 535634
rect 121184 535570 121236 535576
rect 117964 535560 118016 535566
rect 117964 535502 118016 535508
rect 114742 534168 114798 534177
rect 114742 534103 114798 534112
rect 113666 528834 114048 528850
rect 114756 528836 114784 534103
rect 115848 530528 115900 530534
rect 115848 530470 115900 530476
rect 115860 528836 115888 530470
rect 117136 528896 117188 528902
rect 116886 528844 117136 528850
rect 116886 528838 117188 528844
rect 113666 528828 114060 528834
rect 113666 528822 114008 528828
rect 116886 528822 117176 528838
rect 117976 528836 118004 535502
rect 119068 531140 119120 531146
rect 119068 531082 119120 531088
rect 119080 528836 119108 531082
rect 120448 528964 120500 528970
rect 120448 528906 120500 528912
rect 120460 528850 120488 528906
rect 120198 528822 120488 528850
rect 121196 528836 121224 535570
rect 122288 530052 122340 530058
rect 122288 529994 122340 530000
rect 122300 528836 122328 529994
rect 123404 528836 123432 535638
rect 124404 530120 124456 530126
rect 124404 530062 124456 530068
rect 124416 528836 124444 530062
rect 125520 528836 125548 535706
rect 126612 530188 126664 530194
rect 126612 530130 126664 530136
rect 126624 528836 126652 530130
rect 127728 528836 127756 535774
rect 131946 534304 132002 534313
rect 131946 534239 132002 534248
rect 129830 532808 129886 532817
rect 129830 532743 129886 532752
rect 128728 530256 128780 530262
rect 128728 530198 128780 530204
rect 128740 528836 128768 530198
rect 129844 528836 129872 532743
rect 130936 530324 130988 530330
rect 130936 530266 130988 530272
rect 130948 528836 130976 530266
rect 131960 528836 131988 534239
rect 135258 531584 135314 531593
rect 135258 531519 135314 531528
rect 133052 530392 133104 530398
rect 133052 530334 133104 530340
rect 133064 528836 133092 530334
rect 134156 529032 134208 529038
rect 134156 528974 134208 528980
rect 134168 528836 134196 528974
rect 135272 528836 135300 531519
rect 136272 529100 136324 529106
rect 136272 529042 136324 529048
rect 136284 528836 136312 529042
rect 137388 528836 137416 535842
rect 138478 531720 138534 531729
rect 138478 531655 138534 531664
rect 138492 528836 138520 531655
rect 139504 528836 139532 535910
rect 141698 534440 141754 534449
rect 141698 534375 141754 534384
rect 140596 529168 140648 529174
rect 140596 529110 140648 529116
rect 140608 528836 140636 529110
rect 141712 528836 141740 534375
rect 142804 531344 142856 531350
rect 142804 531286 142856 531292
rect 142816 528836 142844 531286
rect 144920 529236 144972 529242
rect 144920 529178 144972 529184
rect 144932 528836 144960 529178
rect 146036 528836 146064 536862
rect 147036 531412 147088 531418
rect 147036 531354 147088 531360
rect 147048 528836 147076 531354
rect 148152 528836 148180 536930
rect 149244 529304 149296 529310
rect 149244 529246 149296 529252
rect 149256 528836 149284 529246
rect 150360 528836 150388 536998
rect 152476 528836 152504 537066
rect 154672 536036 154724 536042
rect 154672 535978 154724 535984
rect 154684 528836 154712 535978
rect 155684 529372 155736 529378
rect 155684 529314 155736 529320
rect 155696 528836 155724 529314
rect 156800 528836 156828 537134
rect 157890 532944 157946 532953
rect 157890 532879 157946 532888
rect 157904 528836 157932 532879
rect 158916 528836 158944 537202
rect 161110 533080 161166 533089
rect 161110 533015 161166 533024
rect 161124 528836 161152 533015
rect 163240 528836 163268 537270
rect 164332 534132 164384 534138
rect 164332 534074 164384 534080
rect 164344 528836 164372 534074
rect 165448 528836 165476 537338
rect 194508 536172 194560 536178
rect 194508 536114 194560 536120
rect 193404 536104 193456 536110
rect 193404 536046 193456 536052
rect 192392 534676 192444 534682
rect 192392 534618 192444 534624
rect 189080 534608 189132 534614
rect 189080 534550 189132 534556
rect 185860 534540 185912 534546
rect 185860 534482 185912 534488
rect 179420 534472 179472 534478
rect 179420 534414 179472 534420
rect 177304 534404 177356 534410
rect 177304 534346 177356 534352
rect 172980 534336 173032 534342
rect 172980 534278 173032 534284
rect 170772 534268 170824 534274
rect 170772 534210 170824 534216
rect 166448 534200 166500 534206
rect 166448 534142 166500 534148
rect 166460 528836 166488 534142
rect 168656 532772 168708 532778
rect 168656 532714 168708 532720
rect 167552 529440 167604 529446
rect 167552 529382 167604 529388
rect 167564 528836 167592 529382
rect 168668 528836 168696 532714
rect 169760 531548 169812 531554
rect 169760 531490 169812 531496
rect 169772 528836 169800 531490
rect 170784 528836 170812 534210
rect 171876 531616 171928 531622
rect 171876 531558 171928 531564
rect 171888 528836 171916 531558
rect 172992 528836 173020 534278
rect 176200 531752 176252 531758
rect 176200 531694 176252 531700
rect 173992 531684 174044 531690
rect 173992 531626 174044 531632
rect 174004 528836 174032 531626
rect 175096 529508 175148 529514
rect 175096 529450 175148 529456
rect 175108 528836 175136 529450
rect 176212 528836 176240 531694
rect 177316 528836 177344 534346
rect 178316 531820 178368 531826
rect 178316 531762 178368 531768
rect 178328 528836 178356 531762
rect 179432 528836 179460 534414
rect 183744 531480 183796 531486
rect 183744 531422 183796 531428
rect 182640 530596 182692 530602
rect 182640 530538 182692 530544
rect 180524 530460 180576 530466
rect 180524 530402 180576 530408
rect 180536 528836 180564 530402
rect 182652 528836 182680 530538
rect 183756 528836 183784 531422
rect 184848 530664 184900 530670
rect 184848 530606 184900 530612
rect 184860 528836 184888 530606
rect 185872 528836 185900 534482
rect 188068 532840 188120 532846
rect 188068 532782 188120 532788
rect 186964 530732 187016 530738
rect 186964 530674 187016 530680
rect 186976 528836 187004 530674
rect 188080 528836 188108 532782
rect 189092 528836 189120 534550
rect 191288 529576 191340 529582
rect 191288 529518 191340 529524
rect 191300 528836 191328 529518
rect 192404 528836 192432 534618
rect 193416 528836 193444 536046
rect 194520 528836 194548 536114
rect 114008 528770 114060 528776
rect 110696 528760 110748 528766
rect 33152 528686 33902 528714
rect 80808 528686 81374 528714
rect 108330 528698 108712 528714
rect 110446 528708 110696 528714
rect 110446 528702 110748 528708
rect 194612 528714 194640 572222
rect 195624 572150 195652 574110
rect 196820 572354 196848 574110
rect 198108 572422 198136 574110
rect 199304 572558 199332 574110
rect 199292 572552 199344 572558
rect 199292 572494 199344 572500
rect 198096 572416 198148 572422
rect 198096 572358 198148 572364
rect 195980 572348 196032 572354
rect 195980 572290 196032 572296
rect 196808 572348 196860 572354
rect 196808 572290 196860 572296
rect 195612 572144 195664 572150
rect 195612 572086 195664 572092
rect 195992 528714 196020 572290
rect 197360 572076 197412 572082
rect 197360 572018 197412 572024
rect 197372 528850 197400 572018
rect 200120 571940 200172 571946
rect 200120 571882 200172 571888
rect 198832 571464 198884 571470
rect 198832 571406 198884 571412
rect 198740 571396 198792 571402
rect 198740 571338 198792 571344
rect 198752 531078 198780 571338
rect 198740 531072 198792 531078
rect 198740 531014 198792 531020
rect 197372 528822 197754 528850
rect 198844 528836 198872 571406
rect 199660 531072 199712 531078
rect 199660 531014 199712 531020
rect 199672 528850 199700 531014
rect 199672 528822 199962 528850
rect 200132 528714 200160 571882
rect 200500 571470 200528 574110
rect 201420 574110 201480 574138
rect 202676 574110 202828 574138
rect 203872 574110 204208 574138
rect 205068 574110 205404 574138
rect 206356 574110 206692 574138
rect 207552 574110 207888 574138
rect 208748 574110 209084 574138
rect 210036 574110 210372 574138
rect 211232 574110 211568 574138
rect 212428 574110 212488 574138
rect 213624 574110 213868 574138
rect 214912 574110 215248 574138
rect 216108 574110 216444 574138
rect 217304 574110 217640 574138
rect 218592 574110 218928 574138
rect 219788 574110 220124 574138
rect 220984 574110 221320 574138
rect 201420 571538 201448 574110
rect 201500 572144 201552 572150
rect 201500 572086 201552 572092
rect 201408 571532 201460 571538
rect 201408 571474 201460 571480
rect 200488 571464 200540 571470
rect 200488 571406 200540 571412
rect 201512 528714 201540 572086
rect 202800 571606 202828 574110
rect 202972 572416 203024 572422
rect 202972 572358 203024 572364
rect 202880 572348 202932 572354
rect 202880 572290 202932 572296
rect 202788 571600 202840 571606
rect 202788 571542 202840 571548
rect 202892 528850 202920 572290
rect 202984 528986 203012 572358
rect 204180 571402 204208 574110
rect 204260 572552 204312 572558
rect 204260 572494 204312 572500
rect 204168 571396 204220 571402
rect 204168 571338 204220 571344
rect 204272 528986 204300 572494
rect 205376 571674 205404 574110
rect 206664 572218 206692 574110
rect 206652 572212 206704 572218
rect 206652 572154 206704 572160
rect 207860 572082 207888 574110
rect 207848 572076 207900 572082
rect 207848 572018 207900 572024
rect 209056 572014 209084 574110
rect 209044 572008 209096 572014
rect 209044 571950 209096 571956
rect 205364 571668 205416 571674
rect 205364 571610 205416 571616
rect 209780 571668 209832 571674
rect 209780 571610 209832 571616
rect 208400 571600 208452 571606
rect 208400 571542 208452 571548
rect 207020 571532 207072 571538
rect 207020 571474 207072 571480
rect 205640 571464 205692 571470
rect 205640 571406 205692 571412
rect 205652 528986 205680 571406
rect 202984 528958 203748 528986
rect 204272 528958 204852 528986
rect 205652 528958 205956 528986
rect 202892 528822 203182 528850
rect 203720 528714 203748 528958
rect 204824 528714 204852 528958
rect 205928 528714 205956 528958
rect 207032 528714 207060 571474
rect 208412 528850 208440 571542
rect 208492 571396 208544 571402
rect 208492 571338 208544 571344
rect 208504 529258 208532 571338
rect 208504 529230 209084 529258
rect 208412 528822 208518 528850
rect 209056 528714 209084 529230
rect 209792 528714 209820 571610
rect 210344 571402 210372 574110
rect 211160 572212 211212 572218
rect 211160 572154 211212 572160
rect 210332 571396 210384 571402
rect 210332 571338 210384 571344
rect 211172 528714 211200 572154
rect 211540 571470 211568 574110
rect 212460 571538 212488 574110
rect 212540 572076 212592 572082
rect 212540 572018 212592 572024
rect 212448 571532 212500 571538
rect 212448 571474 212500 571480
rect 211528 571464 211580 571470
rect 211528 571406 211580 571412
rect 212552 528850 212580 572018
rect 213840 571606 213868 574110
rect 214012 572008 214064 572014
rect 214012 571950 214064 571956
rect 213828 571600 213880 571606
rect 213828 571542 213880 571548
rect 213920 571396 213972 571402
rect 213920 571338 213972 571344
rect 213932 531078 213960 571338
rect 213920 531072 213972 531078
rect 213920 531014 213972 531020
rect 214024 528850 214052 571950
rect 215220 571402 215248 574110
rect 216416 571946 216444 574110
rect 216404 571940 216456 571946
rect 216404 571882 216456 571888
rect 217612 571674 217640 574110
rect 218900 572150 218928 574110
rect 218888 572144 218940 572150
rect 218888 572086 218940 572092
rect 219440 571940 219492 571946
rect 219440 571882 219492 571888
rect 217600 571668 217652 571674
rect 217600 571610 217652 571616
rect 218060 571600 218112 571606
rect 218060 571542 218112 571548
rect 216680 571532 216732 571538
rect 216680 571474 216732 571480
rect 215300 571464 215352 571470
rect 215300 571406 215352 571412
rect 215208 571396 215260 571402
rect 215208 571338 215260 571344
rect 214748 531072 214800 531078
rect 214748 531014 214800 531020
rect 212552 528822 212842 528850
rect 213946 528822 214052 528850
rect 214760 528850 214788 531014
rect 214760 528822 215050 528850
rect 215312 528714 215340 571406
rect 216692 528850 216720 571474
rect 218072 528850 218100 571542
rect 218152 571396 218204 571402
rect 218152 571338 218204 571344
rect 218164 528986 218192 571338
rect 218164 528958 218836 528986
rect 216692 528822 217166 528850
rect 218072 528822 218270 528850
rect 218808 528714 218836 528958
rect 219452 528714 219480 571882
rect 220096 571606 220124 574110
rect 220820 571668 220872 571674
rect 220820 571610 220872 571616
rect 220084 571600 220136 571606
rect 220084 571542 220136 571548
rect 220832 528714 220860 571610
rect 221292 571402 221320 574110
rect 222120 574110 222180 574138
rect 223468 574110 223528 574138
rect 224664 574110 224908 574138
rect 225860 574110 226196 574138
rect 227148 574110 227484 574138
rect 228344 574110 228680 574138
rect 229540 574110 229876 574138
rect 230736 574110 231072 574138
rect 232024 574110 232360 574138
rect 222120 571470 222148 574110
rect 222200 572144 222252 572150
rect 222200 572086 222252 572092
rect 222108 571464 222160 571470
rect 222108 571406 222160 571412
rect 221280 571396 221332 571402
rect 221280 571338 221332 571344
rect 222212 528850 222240 572086
rect 223500 571538 223528 574110
rect 224880 571606 224908 574110
rect 223580 571600 223632 571606
rect 223580 571542 223632 571548
rect 224868 571600 224920 571606
rect 224868 571542 224920 571548
rect 223488 571532 223540 571538
rect 223488 571474 223540 571480
rect 222212 528822 222594 528850
rect 223592 528836 223620 571542
rect 224960 571464 225012 571470
rect 224960 571406 225012 571412
rect 223672 571396 223724 571402
rect 223672 571338 223724 571344
rect 223684 528714 223712 571338
rect 224972 528986 225000 571406
rect 226168 571402 226196 574110
rect 227456 572082 227484 574110
rect 227444 572076 227496 572082
rect 227444 572018 227496 572024
rect 228652 571674 228680 574110
rect 229100 572076 229152 572082
rect 229100 572018 229152 572024
rect 228640 571668 228692 571674
rect 228640 571610 228692 571616
rect 227812 571600 227864 571606
rect 227812 571542 227864 571548
rect 226340 571532 226392 571538
rect 226340 571474 226392 571480
rect 226156 571396 226208 571402
rect 226156 571338 226208 571344
rect 224972 528958 225276 528986
rect 225248 528714 225276 528958
rect 226352 528714 226380 571474
rect 227720 571396 227772 571402
rect 227720 571338 227772 571344
rect 227732 531078 227760 571338
rect 227720 531072 227772 531078
rect 227720 531014 227772 531020
rect 227824 528850 227852 571542
rect 228732 531072 228784 531078
rect 228732 531014 228784 531020
rect 228744 528850 228772 531014
rect 229112 528986 229140 572018
rect 229848 571402 229876 574110
rect 230480 571668 230532 571674
rect 230480 571610 230532 571616
rect 229836 571396 229888 571402
rect 229836 571338 229888 571344
rect 229112 528958 229692 528986
rect 227824 528822 227930 528850
rect 228744 528822 229034 528850
rect 229664 528714 229692 528958
rect 230492 528714 230520 571610
rect 231044 571538 231072 574110
rect 231032 571532 231084 571538
rect 231032 571474 231084 571480
rect 232332 571402 232360 574110
rect 233160 574110 233220 574138
rect 234416 574110 234568 574138
rect 235704 574110 235948 574138
rect 236900 574110 237328 574138
rect 238096 574110 238616 574138
rect 239292 574110 239628 574138
rect 240580 574110 240916 574138
rect 241776 574110 242112 574138
rect 233160 571470 233188 574110
rect 233332 571532 233384 571538
rect 233332 571474 233384 571480
rect 233148 571464 233200 571470
rect 233148 571406 233200 571412
rect 231860 571396 231912 571402
rect 231860 571338 231912 571344
rect 232320 571396 232372 571402
rect 232320 571338 232372 571344
rect 233240 571396 233292 571402
rect 233240 571338 233292 571344
rect 231872 528850 231900 571338
rect 233252 531078 233280 571338
rect 233240 531072 233292 531078
rect 233240 531014 233292 531020
rect 231872 528822 232254 528850
rect 233344 528836 233372 571474
rect 234540 571402 234568 574110
rect 235920 571470 235948 574110
rect 234620 571464 234672 571470
rect 234620 571406 234672 571412
rect 235908 571464 235960 571470
rect 235908 571406 235960 571412
rect 237300 571418 237328 574110
rect 238588 572098 238616 574110
rect 238588 572070 238800 572098
rect 234528 571396 234580 571402
rect 234528 571338 234580 571344
rect 234068 531072 234120 531078
rect 234068 531014 234120 531020
rect 234080 528850 234108 531014
rect 234080 528822 234370 528850
rect 234632 528714 234660 571406
rect 236000 571396 236052 571402
rect 237300 571390 237512 571418
rect 236000 571338 236052 571344
rect 236012 528714 236040 571338
rect 237380 571328 237432 571334
rect 237380 571270 237432 571276
rect 237392 528850 237420 571270
rect 237484 528986 237512 571390
rect 237484 528958 238156 528986
rect 237392 528822 237682 528850
rect 238128 528714 238156 528958
rect 238772 528714 238800 572070
rect 239600 571402 239628 574110
rect 240888 571402 240916 574110
rect 242084 571402 242112 574110
rect 242912 574110 242972 574138
rect 244168 574110 244228 574138
rect 245456 574110 245608 574138
rect 246652 574110 246988 574138
rect 247848 574110 248368 574138
rect 239588 571396 239640 571402
rect 239588 571338 239640 571344
rect 240140 571396 240192 571402
rect 240140 571338 240192 571344
rect 240876 571396 240928 571402
rect 240876 571338 240928 571344
rect 241520 571396 241572 571402
rect 241520 571338 241572 571344
rect 242072 571396 242124 571402
rect 242072 571338 242124 571344
rect 240152 528714 240180 571338
rect 241532 528850 241560 571338
rect 242912 531078 242940 574110
rect 244200 571418 244228 574110
rect 245580 571418 245608 574110
rect 246960 571418 246988 574110
rect 248340 572098 248368 574110
rect 248524 574110 249136 574138
rect 249812 574110 250332 574138
rect 251192 574110 251528 574138
rect 252664 574110 252724 574138
rect 253952 574110 254012 574138
rect 254872 574110 255208 574138
rect 256068 574110 256404 574138
rect 257356 574110 257692 574138
rect 258184 574110 258888 574138
rect 259472 574110 260084 574138
rect 260852 574110 261280 574138
rect 262232 574110 262568 574138
rect 263612 574110 263764 574138
rect 264624 574110 264960 574138
rect 265912 574110 266248 574138
rect 267108 574110 267444 574138
rect 268304 574110 268640 574138
rect 269500 574110 269836 574138
rect 270788 574110 271124 574138
rect 271984 574110 272320 574138
rect 273272 574110 273516 574138
rect 274652 574110 274804 574138
rect 275664 574110 276000 574138
rect 276860 574110 277196 574138
rect 278056 574110 278392 574138
rect 279344 574110 279680 574138
rect 280540 574110 280876 574138
rect 281736 574110 282072 574138
rect 248340 572070 248460 572098
rect 242992 571396 243044 571402
rect 244200 571390 244320 571418
rect 245580 571390 245700 571418
rect 246960 571390 247080 571418
rect 242992 571338 243044 571344
rect 242900 531072 242952 531078
rect 242900 531014 242952 531020
rect 241532 528822 241914 528850
rect 243004 528836 243032 571338
rect 243820 531072 243872 531078
rect 243820 531014 243872 531020
rect 243832 528850 243860 531014
rect 243832 528822 244122 528850
rect 244292 528714 244320 571390
rect 245672 528714 245700 571390
rect 247052 528850 247080 571390
rect 248432 570722 248460 572070
rect 248420 570716 248472 570722
rect 248420 570658 248472 570664
rect 248524 570602 248552 574110
rect 248432 570574 248552 570602
rect 248432 531078 248460 570574
rect 248512 570512 248564 570518
rect 248512 570454 248564 570460
rect 248420 531072 248472 531078
rect 248420 531014 248472 531020
rect 248524 528850 248552 570454
rect 249156 531072 249208 531078
rect 249156 531014 249208 531020
rect 247052 528822 247342 528850
rect 248446 528822 248552 528850
rect 249168 528850 249196 531014
rect 249168 528822 249458 528850
rect 249812 528714 249840 574110
rect 251192 528714 251220 574110
rect 252664 528850 252692 574110
rect 253952 571418 253980 574110
rect 253860 571390 253980 571418
rect 254872 571402 254900 574110
rect 256068 571402 256096 574110
rect 257356 571402 257384 574110
rect 254860 571396 254912 571402
rect 253860 528850 253888 571390
rect 254860 571338 254912 571344
rect 255320 571396 255372 571402
rect 255320 571338 255372 571344
rect 256056 571396 256108 571402
rect 256056 571338 256108 571344
rect 256700 571396 256752 571402
rect 256700 571338 256752 571344
rect 257344 571396 257396 571402
rect 257344 571338 257396 571344
rect 253940 571328 253992 571334
rect 253940 571270 253992 571276
rect 252664 528822 252770 528850
rect 253782 528822 253888 528850
rect 253952 528714 253980 571270
rect 255332 528714 255360 571338
rect 256712 528850 256740 571338
rect 258184 528850 258212 574110
rect 259472 571418 259500 574110
rect 260852 571418 260880 574110
rect 262232 571418 262260 574110
rect 263612 571418 263640 574110
rect 259380 571390 259500 571418
rect 260760 571390 260880 571418
rect 262140 571390 262260 571418
rect 263428 571390 263640 571418
rect 264624 571402 264652 574110
rect 265912 571402 265940 574110
rect 267108 571402 267136 574110
rect 268304 572082 268332 574110
rect 267648 572076 267700 572082
rect 267648 572018 267700 572024
rect 268292 572076 268344 572082
rect 268292 572018 268344 572024
rect 264612 571396 264664 571402
rect 259380 528850 259408 571390
rect 260760 528850 260788 571390
rect 262140 532506 262168 571390
rect 263428 532506 263456 571390
rect 264612 571338 264664 571344
rect 264888 571396 264940 571402
rect 264888 571338 264940 571344
rect 265900 571396 265952 571402
rect 265900 571338 265952 571344
rect 266268 571396 266320 571402
rect 266268 571338 266320 571344
rect 267096 571396 267148 571402
rect 267096 571338 267148 571344
rect 263508 571328 263560 571334
rect 263508 571270 263560 571276
rect 261300 532500 261352 532506
rect 261300 532442 261352 532448
rect 262128 532500 262180 532506
rect 262128 532442 262180 532448
rect 262404 532500 262456 532506
rect 262404 532442 262456 532448
rect 263416 532500 263468 532506
rect 263416 532442 263468 532448
rect 256712 528822 257002 528850
rect 258106 528822 258212 528850
rect 259210 528822 259408 528850
rect 260314 528822 260788 528850
rect 261312 528836 261340 532442
rect 262416 528836 262444 532442
rect 263520 528836 263548 571270
rect 264900 528850 264928 571338
rect 264546 528822 264928 528850
rect 266280 528714 266308 571338
rect 267660 531078 267688 572018
rect 268936 571464 268988 571470
rect 268936 571406 268988 571412
rect 266728 531072 266780 531078
rect 266728 531014 266780 531020
rect 267648 531072 267700 531078
rect 267648 531014 267700 531020
rect 267832 531072 267884 531078
rect 267832 531014 267884 531020
rect 266740 528836 266768 531014
rect 267844 528836 267872 531014
rect 268948 528850 268976 571406
rect 269500 571402 269528 574110
rect 270788 571470 270816 574110
rect 270776 571464 270828 571470
rect 270776 571406 270828 571412
rect 271788 571464 271840 571470
rect 271788 571406 271840 571412
rect 269028 571396 269080 571402
rect 269028 571338 269080 571344
rect 269488 571396 269540 571402
rect 269488 571338 269540 571344
rect 270408 571396 270460 571402
rect 270408 571338 270460 571344
rect 269040 531078 269068 571338
rect 269028 531072 269080 531078
rect 269028 531014 269080 531020
rect 268870 528822 268976 528850
rect 270420 528714 270448 571338
rect 271800 531010 271828 571406
rect 271984 571402 272012 574110
rect 273168 571532 273220 571538
rect 273168 571474 273220 571480
rect 271972 571396 272024 571402
rect 271972 571338 272024 571344
rect 273076 571396 273128 571402
rect 273076 571338 273128 571344
rect 273088 531078 273116 571338
rect 272064 531072 272116 531078
rect 272064 531014 272116 531020
rect 273076 531072 273128 531078
rect 273076 531014 273128 531020
rect 271052 531004 271104 531010
rect 271052 530946 271104 530952
rect 271788 531004 271840 531010
rect 271788 530946 271840 530952
rect 271064 528836 271092 530946
rect 272076 528836 272104 531014
rect 273180 528836 273208 571474
rect 273272 571470 273300 574110
rect 273260 571464 273312 571470
rect 273260 571406 273312 571412
rect 274548 571464 274600 571470
rect 274548 571406 274600 571412
rect 274560 528850 274588 571406
rect 274652 571402 274680 574110
rect 275664 571538 275692 574110
rect 275928 572076 275980 572082
rect 275928 572018 275980 572024
rect 275652 571532 275704 571538
rect 275652 571474 275704 571480
rect 274640 571396 274692 571402
rect 274640 571338 274692 571344
rect 274298 528822 274588 528850
rect 275940 528714 275968 572018
rect 276860 571470 276888 574110
rect 277308 572144 277360 572150
rect 277308 572086 277360 572092
rect 276848 571464 276900 571470
rect 276848 571406 276900 571412
rect 277320 531078 277348 572086
rect 278056 572082 278084 574110
rect 279344 572150 279372 574110
rect 279332 572144 279384 572150
rect 279332 572086 279384 572092
rect 278044 572076 278096 572082
rect 278044 572018 278096 572024
rect 278596 571464 278648 571470
rect 278596 571406 278648 571412
rect 276388 531072 276440 531078
rect 276388 531014 276440 531020
rect 277308 531072 277360 531078
rect 277308 531014 277360 531020
rect 277492 531072 277544 531078
rect 277492 531014 277544 531020
rect 276400 528836 276428 531014
rect 277504 528836 277532 531014
rect 278608 528836 278636 571406
rect 280540 571402 280568 574110
rect 281736 571470 281764 574110
rect 281724 571464 281776 571470
rect 281724 571406 281776 571412
rect 278688 571396 278740 571402
rect 278688 571338 278740 571344
rect 280528 571396 280580 571402
rect 280528 571338 280580 571344
rect 278700 531078 278728 571338
rect 281540 569900 281592 569906
rect 281540 569842 281592 569848
rect 281552 569226 281580 569842
rect 281540 569220 281592 569226
rect 281540 569162 281592 569168
rect 278688 531072 278740 531078
rect 278688 531014 278740 531020
rect 108330 528692 108724 528698
rect 108330 528686 108672 528692
rect 110446 528686 110736 528702
rect 194612 528686 195638 528714
rect 195992 528686 196650 528714
rect 200132 528686 200974 528714
rect 201512 528686 202078 528714
rect 203720 528686 204194 528714
rect 204824 528686 205298 528714
rect 205928 528686 206402 528714
rect 207032 528686 207506 528714
rect 209056 528686 209622 528714
rect 209792 528686 210726 528714
rect 211172 528686 211738 528714
rect 215312 528686 216062 528714
rect 218808 528686 219282 528714
rect 219452 528686 220386 528714
rect 220832 528686 221490 528714
rect 223684 528686 224710 528714
rect 225248 528686 225814 528714
rect 226352 528686 226826 528714
rect 229664 528686 230138 528714
rect 230492 528686 231150 528714
rect 234632 528686 235474 528714
rect 236012 528686 236578 528714
rect 238128 528686 238694 528714
rect 238772 528686 239798 528714
rect 240152 528686 240902 528714
rect 244292 528686 245226 528714
rect 245672 528686 246238 528714
rect 249812 528686 250562 528714
rect 251192 528686 251666 528714
rect 253952 528686 254886 528714
rect 255332 528686 255990 528714
rect 265650 528686 266308 528714
rect 269974 528686 270448 528714
rect 275402 528686 275968 528714
rect 108672 528634 108724 528640
rect 107568 528624 107620 528630
rect 107226 528572 107568 528578
rect 107226 528566 107620 528572
rect 107226 528550 107608 528566
rect 251916 528556 251968 528562
rect 251916 528498 251968 528504
rect 254216 528556 254268 528562
rect 254216 528498 254268 528504
rect 184204 528488 184256 528494
rect 182178 528456 182234 528465
rect 153594 528426 153976 528442
rect 153594 528420 153988 528426
rect 153594 528414 153936 528420
rect 153936 528362 153988 528368
rect 159364 528420 159416 528426
rect 159364 528362 159416 528368
rect 175188 528420 175240 528426
rect 182178 528391 182234 528400
rect 183926 528456 183982 528465
rect 195428 528488 195480 528494
rect 184204 528430 184256 528436
rect 183926 528391 183982 528400
rect 175188 528362 175240 528368
rect 159376 528222 159404 528362
rect 175200 528290 175228 528362
rect 175922 528320 175978 528329
rect 162768 528284 162820 528290
rect 162688 528244 162768 528272
rect 144184 528216 144236 528222
rect 143842 528164 144184 528170
rect 151728 528216 151780 528222
rect 143842 528158 144236 528164
rect 151386 528164 151728 528170
rect 151386 528158 151780 528164
rect 159364 528216 159416 528222
rect 160376 528216 160428 528222
rect 159364 528158 159416 528164
rect 160034 528164 160376 528170
rect 162688 528170 162716 528244
rect 162768 528226 162820 528232
rect 175188 528284 175240 528290
rect 175922 528255 175978 528264
rect 177946 528320 178002 528329
rect 181902 528320 181958 528329
rect 181562 528278 181902 528306
rect 177946 528255 178002 528264
rect 182192 528290 182220 528391
rect 183940 528290 183968 528391
rect 184112 528352 184164 528358
rect 184112 528294 184164 528300
rect 181902 528255 181958 528264
rect 182180 528284 182232 528290
rect 175188 528226 175240 528232
rect 175936 528222 175964 528255
rect 177960 528222 177988 528255
rect 182180 528226 182232 528232
rect 183928 528284 183980 528290
rect 183928 528226 183980 528232
rect 184124 528222 184152 528294
rect 184216 528222 184244 528430
rect 190210 528426 190408 528442
rect 195428 528430 195480 528436
rect 198004 528488 198056 528494
rect 198004 528430 198056 528436
rect 234160 528488 234212 528494
rect 234160 528430 234212 528436
rect 235080 528488 235132 528494
rect 235080 528430 235132 528436
rect 251822 528456 251878 528465
rect 190210 528420 190420 528426
rect 190210 528414 190368 528420
rect 190368 528362 190420 528368
rect 185952 528352 186004 528358
rect 185950 528320 185952 528329
rect 186004 528320 186006 528329
rect 185950 528255 186006 528264
rect 195440 528222 195468 528430
rect 198016 528222 198044 528430
rect 207570 528320 207626 528329
rect 207570 528255 207626 528264
rect 160034 528158 160428 528164
rect 143842 528142 144224 528158
rect 151386 528142 151768 528158
rect 160034 528142 160416 528158
rect 162242 528142 162716 528170
rect 175924 528216 175976 528222
rect 175924 528158 175976 528164
rect 177948 528216 178000 528222
rect 177948 528158 178000 528164
rect 184112 528216 184164 528222
rect 184112 528158 184164 528164
rect 184204 528216 184256 528222
rect 184204 528158 184256 528164
rect 195428 528216 195480 528222
rect 195428 528158 195480 528164
rect 198004 528216 198056 528222
rect 198004 528158 198056 528164
rect 207018 528218 207074 528227
rect 207584 528222 207612 528255
rect 234172 528222 234200 528430
rect 235092 528222 235120 528430
rect 251822 528391 251824 528400
rect 251876 528391 251878 528400
rect 251824 528362 251876 528368
rect 251822 528320 251878 528329
rect 251822 528255 251878 528264
rect 251836 528222 251864 528255
rect 251928 528222 251956 528498
rect 253846 528456 253902 528465
rect 253846 528391 253848 528400
rect 253900 528391 253902 528400
rect 253848 528362 253900 528368
rect 254228 528222 254256 528498
rect 262220 528488 262272 528494
rect 262220 528430 262272 528436
rect 263048 528488 263100 528494
rect 263048 528430 263100 528436
rect 254306 528320 254362 528329
rect 254306 528255 254362 528264
rect 254320 528222 254348 528255
rect 262232 528222 262260 528430
rect 263060 528222 263088 528430
rect 207018 528153 207074 528162
rect 207572 528216 207624 528222
rect 207572 528158 207624 528164
rect 234160 528216 234212 528222
rect 234160 528158 234212 528164
rect 235080 528216 235132 528222
rect 235080 528158 235132 528164
rect 251824 528216 251876 528222
rect 251824 528158 251876 528164
rect 251916 528216 251968 528222
rect 251916 528158 251968 528164
rect 254216 528216 254268 528222
rect 254216 528158 254268 528164
rect 254308 528216 254360 528222
rect 254308 528158 254360 528164
rect 262220 528216 262272 528222
rect 262220 528158 262272 528164
rect 263048 528216 263100 528222
rect 263048 528158 263100 528164
rect 278688 527944 278740 527950
rect 278688 527886 278740 527892
rect 278700 527406 278728 527886
rect 278688 527400 278740 527406
rect 278688 527342 278740 527348
rect 281552 515953 281580 569162
rect 281538 515944 281594 515953
rect 281538 515879 281594 515888
rect 15844 509312 15896 509318
rect 15844 509254 15896 509260
rect 11704 490612 11756 490618
rect 11704 490554 11756 490560
rect 11704 480276 11756 480282
rect 11704 480218 11756 480224
rect 10508 233912 10560 233918
rect 10508 233854 10560 233860
rect 10416 129260 10468 129266
rect 10416 129202 10468 129208
rect 10324 126948 10376 126954
rect 10324 126890 10376 126896
rect 3424 35896 3476 35902
rect 3422 35864 3424 35873
rect 9128 35896 9180 35902
rect 3476 35864 3478 35873
rect 9128 35838 9180 35844
rect 3422 35799 3478 35808
rect 8944 28280 8996 28286
rect 8944 28222 8996 28228
rect 2778 21448 2834 21457
rect 2778 21383 2834 21392
rect 2792 7177 2820 21383
rect 2778 7168 2834 7177
rect 2778 7103 2834 7112
rect 8852 6248 8904 6254
rect 8852 6190 8904 6196
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 1676 4140 1728 4146
rect 1676 4082 1728 4088
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 4082
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 2884 480 2912 2994
rect 4080 480 4108 6122
rect 5264 3868 5316 3874
rect 5264 3810 5316 3816
rect 5276 480 5304 3810
rect 6460 3800 6512 3806
rect 6460 3742 6512 3748
rect 6472 480 6500 3742
rect 7656 3256 7708 3262
rect 7656 3198 7708 3204
rect 7668 480 7696 3198
rect 8864 480 8892 6190
rect 8956 3058 8984 28222
rect 9036 10328 9088 10334
rect 9036 10270 9088 10276
rect 9048 4146 9076 10270
rect 9036 4140 9088 4146
rect 9036 4082 9088 4088
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 10060 480 10088 3470
rect 10520 3466 10548 233854
rect 11716 220114 11744 480218
rect 11796 451308 11848 451314
rect 11796 451250 11848 451256
rect 11808 276010 11836 451250
rect 12624 444372 12676 444378
rect 12624 444314 12676 444320
rect 12636 443601 12664 444314
rect 12622 443592 12678 443601
rect 12622 443527 12678 443536
rect 13084 437504 13136 437510
rect 13084 437446 13136 437452
rect 11796 276004 11848 276010
rect 11796 275946 11848 275952
rect 13096 222902 13124 437446
rect 14464 423700 14516 423706
rect 14464 423642 14516 423648
rect 14476 225622 14504 423642
rect 15856 315314 15884 509254
rect 159008 502982 160034 503010
rect 274298 502982 274588 503010
rect 20628 500540 20680 500546
rect 20628 500482 20680 500488
rect 18604 488640 18656 488646
rect 18604 488582 18656 488588
rect 16856 488572 16908 488578
rect 16856 488514 16908 488520
rect 16868 486948 16896 488514
rect 18616 486948 18644 488582
rect 20640 486962 20668 500482
rect 22112 500478 22140 502860
rect 22296 502846 23138 502874
rect 23584 502846 24242 502874
rect 22100 500472 22152 500478
rect 22100 500414 22152 500420
rect 22192 489524 22244 489530
rect 22192 489466 22244 489472
rect 20378 486934 20668 486962
rect 22204 486948 22232 489466
rect 22296 488578 22324 502846
rect 23388 500472 23440 500478
rect 23388 500414 23440 500420
rect 22284 488572 22336 488578
rect 22284 488514 22336 488520
rect 23400 486470 23428 500414
rect 23584 488646 23612 502846
rect 25332 500546 25360 502860
rect 25320 500540 25372 500546
rect 25320 500482 25372 500488
rect 24768 499588 24820 499594
rect 24768 499530 24820 499536
rect 23572 488640 23624 488646
rect 23572 488582 23624 488588
rect 24780 488578 24808 499530
rect 26344 489530 26372 502860
rect 27448 499594 27476 502860
rect 27632 502846 28566 502874
rect 27528 500948 27580 500954
rect 27528 500890 27580 500896
rect 27436 499588 27488 499594
rect 27436 499530 27488 499536
rect 26332 489524 26384 489530
rect 26332 489466 26384 489472
rect 25780 489388 25832 489394
rect 25780 489330 25832 489336
rect 23940 488572 23992 488578
rect 23940 488514 23992 488520
rect 24768 488572 24820 488578
rect 24768 488514 24820 488520
rect 23952 486948 23980 488514
rect 25792 486948 25820 489330
rect 27540 486948 27568 500890
rect 27632 489394 27660 502846
rect 29656 500954 29684 502860
rect 30484 502846 30682 502874
rect 29644 500948 29696 500954
rect 30484 500936 30512 502846
rect 31772 500954 31800 502860
rect 29644 500890 29696 500896
rect 30300 500908 30512 500936
rect 31668 500948 31720 500954
rect 27620 489388 27672 489394
rect 27620 489330 27672 489336
rect 30300 488578 30328 500908
rect 31668 500890 31720 500896
rect 31760 500948 31812 500954
rect 31760 500890 31812 500896
rect 29368 488572 29420 488578
rect 29368 488514 29420 488520
rect 30288 488572 30340 488578
rect 30288 488514 30340 488520
rect 29380 486948 29408 488514
rect 31680 486826 31708 500890
rect 32876 499594 32904 502860
rect 33902 502846 34468 502874
rect 32036 499588 32088 499594
rect 32036 499530 32088 499536
rect 32864 499588 32916 499594
rect 32864 499530 32916 499536
rect 32048 487098 32076 499530
rect 34440 488594 34468 502846
rect 34992 499594 35020 502860
rect 36096 499594 36124 502860
rect 37108 502846 37214 502874
rect 38226 502846 38608 502874
rect 39330 502846 39988 502874
rect 34980 499588 35032 499594
rect 34980 499530 35032 499536
rect 35808 499588 35860 499594
rect 35808 499530 35860 499536
rect 36084 499588 36136 499594
rect 36084 499530 36136 499536
rect 35820 489870 35848 499530
rect 35808 489864 35860 489870
rect 35808 489806 35860 489812
rect 36544 489864 36596 489870
rect 36544 489806 36596 489812
rect 34440 488566 34560 488594
rect 32048 487070 32628 487098
rect 32600 486962 32628 487070
rect 34532 486962 34560 488566
rect 32600 486934 32982 486962
rect 34532 486934 34730 486962
rect 36556 486948 36584 489806
rect 37108 489258 37136 502846
rect 37188 499588 37240 499594
rect 37188 499530 37240 499536
rect 37096 489252 37148 489258
rect 37096 489194 37148 489200
rect 37200 489190 37228 499530
rect 37188 489184 37240 489190
rect 37188 489126 37240 489132
rect 38292 489184 38344 489190
rect 38292 489126 38344 489132
rect 38304 486948 38332 489126
rect 38580 488646 38608 502846
rect 39960 488714 39988 502846
rect 40420 499594 40448 502860
rect 41432 500750 41460 502860
rect 41420 500744 41472 500750
rect 41420 500686 41472 500692
rect 42536 500478 42564 502860
rect 42524 500472 42576 500478
rect 42524 500414 42576 500420
rect 43640 500410 43668 502860
rect 43628 500404 43680 500410
rect 43628 500346 43680 500352
rect 44744 500342 44772 502860
rect 45756 500886 45784 502860
rect 45744 500880 45796 500886
rect 45744 500822 45796 500828
rect 44732 500336 44784 500342
rect 44732 500278 44784 500284
rect 40408 499588 40460 499594
rect 40408 499530 40460 499536
rect 41328 499588 41380 499594
rect 41328 499530 41380 499536
rect 40132 489252 40184 489258
rect 40132 489194 40184 489200
rect 39948 488708 40000 488714
rect 39948 488650 40000 488656
rect 38568 488640 38620 488646
rect 38568 488582 38620 488588
rect 40144 486948 40172 489194
rect 41340 488578 41368 499530
rect 46860 489190 46888 502860
rect 47978 502846 48268 502874
rect 48990 502846 49648 502874
rect 47032 500744 47084 500750
rect 47032 500686 47084 500692
rect 46848 489184 46900 489190
rect 46848 489126 46900 489132
rect 43720 488708 43772 488714
rect 43720 488650 43772 488656
rect 41880 488640 41932 488646
rect 41880 488582 41932 488588
rect 41328 488572 41380 488578
rect 41328 488514 41380 488520
rect 41892 486948 41920 488582
rect 43732 486948 43760 488650
rect 45468 488572 45520 488578
rect 45468 488514 45520 488520
rect 45480 486948 45508 488514
rect 47044 486962 47072 500686
rect 47584 500472 47636 500478
rect 47584 500414 47636 500420
rect 47596 488578 47624 500414
rect 48240 489326 48268 502846
rect 48964 500404 49016 500410
rect 48964 500346 49016 500352
rect 48228 489320 48280 489326
rect 48228 489262 48280 489268
rect 48976 488646 49004 500346
rect 49620 489598 49648 502846
rect 50080 499798 50108 502860
rect 51184 500954 51212 502860
rect 51172 500948 51224 500954
rect 51172 500890 51224 500896
rect 50068 499792 50120 499798
rect 50068 499734 50120 499740
rect 50988 499792 51040 499798
rect 50988 499734 51040 499740
rect 49608 489592 49660 489598
rect 49608 489534 49660 489540
rect 51000 489530 51028 499734
rect 50988 489524 51040 489530
rect 50988 489466 51040 489472
rect 52288 489394 52316 502860
rect 53314 502846 53788 502874
rect 54418 502846 55168 502874
rect 52368 500948 52420 500954
rect 52368 500890 52420 500896
rect 52380 489802 52408 500890
rect 52552 500336 52604 500342
rect 52552 500278 52604 500284
rect 52368 489796 52420 489802
rect 52368 489738 52420 489744
rect 52276 489388 52328 489394
rect 52276 489330 52328 489336
rect 48964 488640 49016 488646
rect 48964 488582 49016 488588
rect 50896 488640 50948 488646
rect 50896 488582 50948 488588
rect 47584 488572 47636 488578
rect 47584 488514 47636 488520
rect 49056 488572 49108 488578
rect 49056 488514 49108 488520
rect 47044 486934 47334 486962
rect 49068 486948 49096 488514
rect 50908 486948 50936 488582
rect 52564 486962 52592 500278
rect 53760 489462 53788 502846
rect 53932 500880 53984 500886
rect 53932 500822 53984 500828
rect 53748 489456 53800 489462
rect 53748 489398 53800 489404
rect 53944 486962 53972 500822
rect 55140 489734 55168 502846
rect 55508 500954 55536 502860
rect 56428 502846 56534 502874
rect 57638 502846 57928 502874
rect 58742 502846 59308 502874
rect 55496 500948 55548 500954
rect 55496 500890 55548 500896
rect 55128 489728 55180 489734
rect 55128 489670 55180 489676
rect 56428 489190 56456 502846
rect 56508 500948 56560 500954
rect 56508 500890 56560 500896
rect 56520 489258 56548 500890
rect 57900 491978 57928 502846
rect 57888 491972 57940 491978
rect 57888 491914 57940 491920
rect 59280 489326 59308 502846
rect 59372 502846 59846 502874
rect 59372 493338 59400 502846
rect 60844 499594 60872 502860
rect 61948 500206 61976 502860
rect 63066 502846 63448 502874
rect 61936 500200 61988 500206
rect 61936 500142 61988 500148
rect 60832 499588 60884 499594
rect 60832 499530 60884 499536
rect 62028 499588 62080 499594
rect 62028 499530 62080 499536
rect 59360 493332 59412 493338
rect 59360 493274 59412 493280
rect 62040 489666 62068 499530
rect 63132 489796 63184 489802
rect 63132 489738 63184 489744
rect 62028 489660 62080 489666
rect 62028 489602 62080 489608
rect 59820 489592 59872 489598
rect 59820 489534 59872 489540
rect 58072 489320 58124 489326
rect 58072 489262 58124 489268
rect 59268 489320 59320 489326
rect 59268 489262 59320 489268
rect 56508 489252 56560 489258
rect 56508 489194 56560 489200
rect 56232 489184 56284 489190
rect 56232 489126 56284 489132
rect 56416 489184 56468 489190
rect 56416 489126 56468 489132
rect 52564 486934 52670 486962
rect 53944 486934 54510 486962
rect 56244 486948 56272 489126
rect 58084 486948 58112 489262
rect 59832 486948 59860 489534
rect 61660 489524 61712 489530
rect 61660 489466 61712 489472
rect 61672 486948 61700 489466
rect 63144 486962 63172 489738
rect 63420 489598 63448 502846
rect 63512 502846 64078 502874
rect 63512 494766 63540 502846
rect 65168 499594 65196 502860
rect 65156 499588 65208 499594
rect 65156 499530 65208 499536
rect 66168 499588 66220 499594
rect 66168 499530 66220 499536
rect 63500 494760 63552 494766
rect 63500 494702 63552 494708
rect 63408 489592 63460 489598
rect 63408 489534 63460 489540
rect 66180 489530 66208 499530
rect 66272 498846 66300 502860
rect 67390 502846 67496 502874
rect 68402 502846 68968 502874
rect 66260 498840 66312 498846
rect 66260 498782 66312 498788
rect 66168 489524 66220 489530
rect 66168 489466 66220 489472
rect 67468 489462 67496 502846
rect 68940 492114 68968 502846
rect 69492 499594 69520 502860
rect 69480 499588 69532 499594
rect 69480 499530 69532 499536
rect 70308 499588 70360 499594
rect 70308 499530 70360 499536
rect 68928 492108 68980 492114
rect 68928 492050 68980 492056
rect 68744 489728 68796 489734
rect 68744 489670 68796 489676
rect 66996 489456 67048 489462
rect 66996 489398 67048 489404
rect 67456 489456 67508 489462
rect 67456 489398 67508 489404
rect 65156 489388 65208 489394
rect 65156 489330 65208 489336
rect 63144 486934 63434 486962
rect 65168 486948 65196 489330
rect 67008 486948 67036 489398
rect 68756 486948 68784 489670
rect 70320 489394 70348 499530
rect 70596 497622 70624 502860
rect 71622 502846 71728 502874
rect 70584 497616 70636 497622
rect 70584 497558 70636 497564
rect 70308 489388 70360 489394
rect 70308 489330 70360 489336
rect 71700 489258 71728 502846
rect 72712 499594 72740 502860
rect 73830 502846 74488 502874
rect 71780 499588 71832 499594
rect 71780 499530 71832 499536
rect 72700 499588 72752 499594
rect 72700 499530 72752 499536
rect 71792 493474 71820 499530
rect 71780 493468 71832 493474
rect 71780 493410 71832 493416
rect 74172 491972 74224 491978
rect 74172 491914 74224 491920
rect 70584 489252 70636 489258
rect 70584 489194 70636 489200
rect 71688 489252 71740 489258
rect 71688 489194 71740 489200
rect 70596 486948 70624 489194
rect 72332 489184 72384 489190
rect 72332 489126 72384 489132
rect 72344 486948 72372 489126
rect 74184 486948 74212 491914
rect 74460 489190 74488 502846
rect 74552 502846 74934 502874
rect 74552 494902 74580 502846
rect 75932 499594 75960 502860
rect 77050 502846 77156 502874
rect 78154 502846 78628 502874
rect 75920 499588 75972 499594
rect 75920 499530 75972 499536
rect 74540 494896 74592 494902
rect 74540 494838 74592 494844
rect 77128 492046 77156 502846
rect 77208 499588 77260 499594
rect 77208 499530 77260 499536
rect 77116 492040 77168 492046
rect 77116 491982 77168 491988
rect 77220 489326 77248 499530
rect 77300 493332 77352 493338
rect 77300 493274 77352 493280
rect 75920 489320 75972 489326
rect 75920 489262 75972 489268
rect 77208 489320 77260 489326
rect 77208 489262 77260 489268
rect 74448 489184 74500 489190
rect 74448 489126 74500 489132
rect 75932 486948 75960 489262
rect 77312 488050 77340 493274
rect 78600 489122 78628 502846
rect 78692 502846 79166 502874
rect 78692 493406 78720 502846
rect 80060 500812 80112 500818
rect 80060 500754 80112 500760
rect 80072 498914 80100 500754
rect 80256 500274 80284 502860
rect 81360 500818 81388 502860
rect 82478 502846 82768 502874
rect 81348 500812 81400 500818
rect 81348 500754 81400 500760
rect 80244 500268 80296 500274
rect 80244 500210 80296 500216
rect 80244 500132 80296 500138
rect 80244 500074 80296 500080
rect 80060 498908 80112 498914
rect 80060 498850 80112 498856
rect 78680 493400 78732 493406
rect 78680 493342 78732 493348
rect 79508 489660 79560 489666
rect 79508 489602 79560 489608
rect 78588 489116 78640 489122
rect 78588 489058 78640 489064
rect 77312 488022 77524 488050
rect 77496 486962 77524 488022
rect 77496 486934 77786 486962
rect 79520 486948 79548 489602
rect 80256 488050 80284 500074
rect 82740 489870 82768 502846
rect 82832 502846 83490 502874
rect 82832 497554 82860 502846
rect 84580 500342 84608 502860
rect 84568 500336 84620 500342
rect 84568 500278 84620 500284
rect 82820 497548 82872 497554
rect 82820 497490 82872 497496
rect 85684 494834 85712 502860
rect 86710 502846 86908 502874
rect 87814 502846 88288 502874
rect 85672 494828 85724 494834
rect 85672 494770 85724 494776
rect 84200 494760 84252 494766
rect 84200 494702 84252 494708
rect 82728 489864 82780 489870
rect 82728 489806 82780 489812
rect 83096 489592 83148 489598
rect 83096 489534 83148 489540
rect 80256 488022 81020 488050
rect 80992 486962 81020 488022
rect 80992 486934 81374 486962
rect 83108 486948 83136 489534
rect 31142 486798 31708 486826
rect 84212 486826 84240 494702
rect 86880 489802 86908 502846
rect 88260 491978 88288 502846
rect 88904 500410 88932 502860
rect 89824 502846 90022 502874
rect 90928 502846 91034 502874
rect 88892 500404 88944 500410
rect 88892 500346 88944 500352
rect 89824 498846 89852 502846
rect 88340 498840 88392 498846
rect 88340 498782 88392 498788
rect 89812 498840 89864 498846
rect 89812 498782 89864 498788
rect 88248 491972 88300 491978
rect 88248 491914 88300 491920
rect 86868 489796 86920 489802
rect 86868 489738 86920 489744
rect 86684 489524 86736 489530
rect 86684 489466 86736 489472
rect 86696 486948 86724 489466
rect 88352 486962 88380 498782
rect 90928 489734 90956 502846
rect 92124 499866 92152 502860
rect 93228 500478 93256 502860
rect 93872 502846 94254 502874
rect 93216 500472 93268 500478
rect 93216 500414 93268 500420
rect 92112 499860 92164 499866
rect 92112 499802 92164 499808
rect 93768 499860 93820 499866
rect 93768 499802 93820 499808
rect 93780 493338 93808 499802
rect 93872 497486 93900 502846
rect 95344 500886 95372 502860
rect 96448 500954 96476 502860
rect 95424 500948 95476 500954
rect 95424 500890 95476 500896
rect 96436 500948 96488 500954
rect 96436 500890 96488 500896
rect 95332 500880 95384 500886
rect 95332 500822 95384 500828
rect 95240 497616 95292 497622
rect 95240 497558 95292 497564
rect 93860 497480 93912 497486
rect 93860 497422 93912 497428
rect 93768 493332 93820 493338
rect 93768 493274 93820 493280
rect 92112 492108 92164 492114
rect 92112 492050 92164 492056
rect 90916 489728 90968 489734
rect 90916 489670 90968 489676
rect 90272 489456 90324 489462
rect 90272 489398 90324 489404
rect 88352 486934 88550 486962
rect 90284 486948 90312 489398
rect 92124 486948 92152 492050
rect 93860 489388 93912 489394
rect 93860 489330 93912 489336
rect 93872 486948 93900 489330
rect 95252 486962 95280 497558
rect 95436 494766 95464 500890
rect 96528 500880 96580 500886
rect 96528 500822 96580 500828
rect 95424 494760 95476 494766
rect 95424 494702 95476 494708
rect 96540 489666 96568 500822
rect 97552 500546 97580 502860
rect 98578 502846 99328 502874
rect 97540 500540 97592 500546
rect 97540 500482 97592 500488
rect 98000 493468 98052 493474
rect 98000 493410 98052 493416
rect 96528 489660 96580 489666
rect 96528 489602 96580 489608
rect 97448 489252 97500 489258
rect 97448 489194 97500 489200
rect 95252 486934 95726 486962
rect 97460 486948 97488 489194
rect 98012 488050 98040 493410
rect 99300 489530 99328 502846
rect 99668 500954 99696 502860
rect 100772 500954 100800 502860
rect 101798 502846 101996 502874
rect 102902 502846 103468 502874
rect 99656 500948 99708 500954
rect 99656 500890 99708 500896
rect 100668 500948 100720 500954
rect 100668 500890 100720 500896
rect 100760 500948 100812 500954
rect 100760 500890 100812 500896
rect 100680 489598 100708 500890
rect 100668 489592 100720 489598
rect 100668 489534 100720 489540
rect 99288 489524 99340 489530
rect 99288 489466 99340 489472
rect 101968 489190 101996 502846
rect 102048 500948 102100 500954
rect 102048 500890 102100 500896
rect 102060 489462 102088 500890
rect 102140 494896 102192 494902
rect 102140 494838 102192 494844
rect 102048 489456 102100 489462
rect 102048 489398 102100 489404
rect 101036 489184 101088 489190
rect 101036 489126 101088 489132
rect 101956 489184 102008 489190
rect 101956 489126 102008 489132
rect 98012 488022 98776 488050
rect 98748 486962 98776 488022
rect 98748 486934 99314 486962
rect 101048 486948 101076 489126
rect 102152 486962 102180 494838
rect 103440 489258 103468 502846
rect 103992 500954 104020 502860
rect 105096 500954 105124 502860
rect 105280 502846 106122 502874
rect 103980 500948 104032 500954
rect 103980 500890 104032 500896
rect 104808 500948 104860 500954
rect 104808 500890 104860 500896
rect 105084 500948 105136 500954
rect 105084 500890 105136 500896
rect 104820 489326 104848 500890
rect 105280 500834 105308 502846
rect 106924 500948 106976 500954
rect 106924 500890 106976 500896
rect 104912 500806 105308 500834
rect 104912 498166 104940 500806
rect 104900 498160 104952 498166
rect 104900 498102 104952 498108
rect 106464 492040 106516 492046
rect 106464 491982 106516 491988
rect 104624 489320 104676 489326
rect 104624 489262 104676 489268
rect 104808 489320 104860 489326
rect 104808 489262 104860 489268
rect 103428 489252 103480 489258
rect 103428 489194 103480 489200
rect 102152 486934 102902 486962
rect 104636 486948 104664 489262
rect 106476 486948 106504 491982
rect 106936 489394 106964 500890
rect 107212 500449 107240 502860
rect 107672 502846 108330 502874
rect 109052 502846 109342 502874
rect 107198 500440 107254 500449
rect 107198 500375 107254 500384
rect 107672 497593 107700 502846
rect 108304 500268 108356 500274
rect 108304 500210 108356 500216
rect 107658 497584 107714 497593
rect 107658 497519 107714 497528
rect 106924 489388 106976 489394
rect 106924 489330 106976 489336
rect 108212 489116 108264 489122
rect 108212 489058 108264 489064
rect 108224 486948 108252 489058
rect 108316 488578 108344 500210
rect 109052 497457 109080 502846
rect 109684 500336 109736 500342
rect 109684 500278 109736 500284
rect 109038 497448 109094 497457
rect 109038 497383 109094 497392
rect 109040 493400 109092 493406
rect 109040 493342 109092 493348
rect 108304 488572 108356 488578
rect 108304 488514 108356 488520
rect 109052 488050 109080 493342
rect 109696 488986 109724 500278
rect 110432 497729 110460 502860
rect 110616 502846 111550 502874
rect 110616 497865 110644 502846
rect 112444 500404 112496 500410
rect 112444 500346 112496 500352
rect 110602 497856 110658 497865
rect 110602 497791 110658 497800
rect 110418 497720 110474 497729
rect 110418 497655 110474 497664
rect 112456 489054 112484 500346
rect 112640 500177 112668 502860
rect 113652 500313 113680 502860
rect 114756 500721 114784 502860
rect 114940 502846 115874 502874
rect 114742 500712 114798 500721
rect 114742 500647 114798 500656
rect 114940 500562 114968 502846
rect 116872 500585 116900 502860
rect 114572 500534 114968 500562
rect 116858 500576 116914 500585
rect 115204 500540 115256 500546
rect 113824 500472 113876 500478
rect 113824 500414 113876 500420
rect 113638 500304 113694 500313
rect 113638 500239 113694 500248
rect 112626 500168 112682 500177
rect 112626 500103 112682 500112
rect 113180 498908 113232 498914
rect 113180 498850 113232 498856
rect 112444 489048 112496 489054
rect 112444 488990 112496 488996
rect 109684 488980 109736 488986
rect 109684 488922 109736 488928
rect 111800 488572 111852 488578
rect 111800 488514 111852 488520
rect 109052 488022 109724 488050
rect 109696 486962 109724 488022
rect 109696 486934 109986 486962
rect 111812 486948 111840 488514
rect 113192 486962 113220 498850
rect 113836 489122 113864 500414
rect 114572 498001 114600 500534
rect 116858 500511 116914 500520
rect 115204 500482 115256 500488
rect 114558 497992 114614 498001
rect 114558 497927 114614 497936
rect 115216 489870 115244 500482
rect 117976 500449 118004 502860
rect 118712 502846 119094 502874
rect 117962 500440 118018 500449
rect 117962 500375 118018 500384
rect 118712 497554 118740 502846
rect 120184 500274 120212 502860
rect 121196 500342 121224 502860
rect 121472 502846 122314 502874
rect 121184 500336 121236 500342
rect 121184 500278 121236 500284
rect 120172 500268 120224 500274
rect 120172 500210 120224 500216
rect 121472 497622 121500 502846
rect 123404 500410 123432 502860
rect 124232 502846 124430 502874
rect 123392 500404 123444 500410
rect 123392 500346 123444 500352
rect 124232 498137 124260 502846
rect 125520 500478 125548 502860
rect 125612 502846 126638 502874
rect 125508 500472 125560 500478
rect 125508 500414 125560 500420
rect 124218 498128 124274 498137
rect 124218 498063 124274 498072
rect 121460 497616 121512 497622
rect 121460 497558 121512 497564
rect 115940 497548 115992 497554
rect 115940 497490 115992 497496
rect 118700 497548 118752 497554
rect 118700 497490 118752 497496
rect 115020 489864 115072 489870
rect 115020 489806 115072 489812
rect 115204 489864 115256 489870
rect 115204 489806 115256 489812
rect 113824 489116 113876 489122
rect 113824 489058 113876 489064
rect 115032 486962 115060 489806
rect 115952 488050 115980 497490
rect 125612 497321 125640 502846
rect 127728 500546 127756 502860
rect 128372 502846 128754 502874
rect 127716 500540 127768 500546
rect 127716 500482 127768 500488
rect 126980 498840 127032 498846
rect 126980 498782 127032 498788
rect 125598 497312 125654 497321
rect 125598 497247 125654 497256
rect 120080 494828 120132 494834
rect 120080 494770 120132 494776
rect 118976 488980 119028 488986
rect 118976 488922 119028 488928
rect 115952 488022 116716 488050
rect 113192 486934 113574 486962
rect 115032 486934 115414 486962
rect 116688 486826 116716 488022
rect 118988 486948 119016 488922
rect 120092 486826 120120 494770
rect 124312 491972 124364 491978
rect 124312 491914 124364 491920
rect 122564 489796 122616 489802
rect 122564 489738 122616 489744
rect 122576 486948 122604 489738
rect 124324 486948 124352 491914
rect 126152 489048 126204 489054
rect 126152 488990 126204 488996
rect 126164 486948 126192 488990
rect 126992 486826 127020 498782
rect 128372 497185 128400 502846
rect 129844 500614 129872 502860
rect 130948 500857 130976 502860
rect 130934 500848 130990 500857
rect 130934 500783 130990 500792
rect 131960 500682 131988 502860
rect 132512 502846 133078 502874
rect 131948 500676 132000 500682
rect 131948 500618 132000 500624
rect 129832 500608 129884 500614
rect 129832 500550 129884 500556
rect 132512 497690 132540 502846
rect 134168 500818 134196 502860
rect 134156 500812 134208 500818
rect 134156 500754 134208 500760
rect 135272 500750 135300 502860
rect 136284 500954 136312 502860
rect 136272 500948 136324 500954
rect 136272 500890 136324 500896
rect 137388 500886 137416 502860
rect 137376 500880 137428 500886
rect 137376 500822 137428 500828
rect 135260 500744 135312 500750
rect 135260 500686 135312 500692
rect 138492 500206 138520 502860
rect 138480 500200 138532 500206
rect 138480 500142 138532 500148
rect 139504 500138 139532 502860
rect 139492 500132 139544 500138
rect 139492 500074 139544 500080
rect 140608 500070 140636 502860
rect 141712 500857 141740 502860
rect 141698 500848 141754 500857
rect 141698 500783 141754 500792
rect 142710 500712 142766 500721
rect 142710 500647 142766 500656
rect 140596 500064 140648 500070
rect 140596 500006 140648 500012
rect 142724 499905 142752 500647
rect 142816 500002 142844 502860
rect 142804 499996 142856 500002
rect 142804 499938 142856 499944
rect 142710 499896 142766 499905
rect 142710 499831 142766 499840
rect 143828 499769 143856 502860
rect 144932 499798 144960 502860
rect 144920 499792 144972 499798
rect 143814 499760 143870 499769
rect 144920 499734 144972 499740
rect 143814 499695 143870 499704
rect 132500 497684 132552 497690
rect 132500 497626 132552 497632
rect 133880 497480 133932 497486
rect 133880 497422 133932 497428
rect 128358 497176 128414 497185
rect 128358 497111 128414 497120
rect 131120 493332 131172 493338
rect 131120 493274 131172 493280
rect 129740 489728 129792 489734
rect 129740 489670 129792 489676
rect 129752 486948 129780 489670
rect 131132 486962 131160 493274
rect 133328 489116 133380 489122
rect 133328 489058 133380 489064
rect 131132 486934 131514 486962
rect 133340 486948 133368 489058
rect 133892 488050 133920 497422
rect 138664 494760 138716 494766
rect 138664 494702 138716 494708
rect 136916 489660 136968 489666
rect 136916 489602 136968 489608
rect 133892 488022 134564 488050
rect 134536 486826 134564 488022
rect 136928 486948 136956 489602
rect 138676 486948 138704 494702
rect 146036 492726 146064 502860
rect 146852 500200 146904 500206
rect 146852 500142 146904 500148
rect 146024 492720 146076 492726
rect 146864 492697 146892 500142
rect 147048 499633 147076 502860
rect 148152 499633 148180 502860
rect 149256 499633 149284 502860
rect 150360 499633 150388 502860
rect 151372 499633 151400 502860
rect 152476 499633 152504 502860
rect 153594 502846 154344 502874
rect 154316 502353 154344 502846
rect 154592 502846 154698 502874
rect 154302 502344 154358 502353
rect 154302 502279 154358 502288
rect 154394 502208 154450 502217
rect 154394 502143 154450 502152
rect 153660 500948 153712 500954
rect 153660 500890 153712 500896
rect 153566 500848 153622 500857
rect 153566 500783 153622 500792
rect 153292 500336 153344 500342
rect 153292 500278 153344 500284
rect 147034 499624 147090 499633
rect 147034 499559 147090 499568
rect 148138 499624 148194 499633
rect 148138 499559 148194 499568
rect 149242 499624 149298 499633
rect 149242 499559 149298 499568
rect 150346 499624 150402 499633
rect 150346 499559 150402 499568
rect 151358 499624 151414 499633
rect 151358 499559 151414 499568
rect 152462 499624 152518 499633
rect 152462 499559 152518 499568
rect 153200 498160 153252 498166
rect 153200 498102 153252 498108
rect 153212 497729 153240 498102
rect 153198 497720 153254 497729
rect 153198 497655 153254 497664
rect 146024 492662 146076 492668
rect 146850 492688 146906 492697
rect 146850 492623 146906 492632
rect 140504 489864 140556 489870
rect 140504 489806 140556 489812
rect 140516 486948 140544 489806
rect 144092 489592 144144 489598
rect 144092 489534 144144 489540
rect 142252 489524 142304 489530
rect 142252 489466 142304 489472
rect 142264 486948 142292 489466
rect 144104 486948 144132 489534
rect 145840 489456 145892 489462
rect 145840 489398 145892 489404
rect 145852 486948 145880 489398
rect 153016 489388 153068 489394
rect 153016 489330 153068 489336
rect 151268 489320 151320 489326
rect 151268 489262 151320 489268
rect 149428 489252 149480 489258
rect 149428 489194 149480 489200
rect 147680 489184 147732 489190
rect 147680 489126 147732 489132
rect 147692 486948 147720 489126
rect 149440 486948 149468 489194
rect 151280 486948 151308 489262
rect 153028 486948 153056 489330
rect 84212 486798 84962 486826
rect 116688 486798 117162 486826
rect 120092 486798 120750 486826
rect 126992 486798 127926 486826
rect 134536 486798 135102 486826
rect 23388 486464 23440 486470
rect 23388 486406 23440 486412
rect 140688 401600 140740 401606
rect 140688 401542 140740 401548
rect 140596 401532 140648 401538
rect 140596 401474 140648 401480
rect 139308 401464 139360 401470
rect 131026 401432 131082 401441
rect 139308 401406 139360 401412
rect 131026 401367 131082 401376
rect 136548 401396 136600 401402
rect 129646 401296 129702 401305
rect 129646 401231 129702 401240
rect 126886 401160 126942 401169
rect 126886 401095 126942 401104
rect 125506 401024 125562 401033
rect 125416 400988 125468 400994
rect 125506 400959 125562 400968
rect 125416 400930 125468 400936
rect 122748 400920 122800 400926
rect 118606 400888 118662 400897
rect 122748 400862 122800 400868
rect 118606 400823 118662 400832
rect 78586 377360 78642 377369
rect 78586 377295 78642 377304
rect 78600 376786 78628 377295
rect 78588 376780 78640 376786
rect 78588 376722 78640 376728
rect 21362 357368 21418 357377
rect 21362 357303 21418 357312
rect 20332 357054 20668 357082
rect 20976 357054 21312 357082
rect 20640 353326 20668 357054
rect 21284 353394 21312 357054
rect 21272 353388 21324 353394
rect 21272 353330 21324 353336
rect 20628 353320 20680 353326
rect 20628 353262 20680 353268
rect 21376 323542 21404 357303
rect 21712 357054 22048 357082
rect 22448 357054 22784 357082
rect 23184 357054 23428 357082
rect 23920 357054 24256 357082
rect 24564 357054 24808 357082
rect 25300 357054 25636 357082
rect 26036 357054 26188 357082
rect 26772 357054 27108 357082
rect 22020 353462 22048 357054
rect 22008 353456 22060 353462
rect 22008 353398 22060 353404
rect 22756 353326 22784 357054
rect 23400 353394 23428 357054
rect 24228 353462 24256 357054
rect 24780 353530 24808 357054
rect 25608 354278 25636 357054
rect 25596 354272 25648 354278
rect 25596 354214 25648 354220
rect 26160 354006 26188 357054
rect 26148 354000 26200 354006
rect 26148 353942 26200 353948
rect 27080 353598 27108 357054
rect 27494 356810 27522 357068
rect 28152 357054 28488 357082
rect 27494 356782 27568 356810
rect 27068 353592 27120 353598
rect 27068 353534 27120 353540
rect 24768 353524 24820 353530
rect 24768 353466 24820 353472
rect 23940 353456 23992 353462
rect 23940 353398 23992 353404
rect 24216 353456 24268 353462
rect 24216 353398 24268 353404
rect 27068 353456 27120 353462
rect 27068 353398 27120 353404
rect 22836 353388 22888 353394
rect 22836 353330 22888 353336
rect 23388 353388 23440 353394
rect 23388 353330 23440 353336
rect 22192 353320 22244 353326
rect 22192 353262 22244 353268
rect 22744 353320 22796 353326
rect 22744 353262 22796 353268
rect 22204 348786 22232 353262
rect 22848 348922 22876 353330
rect 23952 348922 23980 353398
rect 26240 353388 26292 353394
rect 26240 353330 26292 353336
rect 25044 353320 25096 353326
rect 25044 353262 25096 353268
rect 25056 348922 25084 353262
rect 26252 348922 26280 353330
rect 27080 348922 27108 353398
rect 27540 353326 27568 356782
rect 28172 353524 28224 353530
rect 28172 353466 28224 353472
rect 27528 353320 27580 353326
rect 27528 353262 27580 353268
rect 28184 348922 28212 353466
rect 28460 353394 28488 357054
rect 28874 356810 28902 357068
rect 29624 357054 29960 357082
rect 28874 356782 28948 356810
rect 28920 353530 28948 356782
rect 29276 354272 29328 354278
rect 29276 354214 29328 354220
rect 28908 353524 28960 353530
rect 28908 353466 28960 353472
rect 28448 353388 28500 353394
rect 28448 353330 28500 353336
rect 29288 348922 29316 354214
rect 29932 353802 29960 357054
rect 30300 357054 30360 357082
rect 31096 357054 31432 357082
rect 29920 353796 29972 353802
rect 29920 353738 29972 353744
rect 30300 353734 30328 357054
rect 30380 354000 30432 354006
rect 30380 353942 30432 353948
rect 30288 353728 30340 353734
rect 30288 353670 30340 353676
rect 30392 348922 30420 353942
rect 31404 353462 31432 357054
rect 31680 357054 31740 357082
rect 32476 357054 32812 357082
rect 33212 357054 33548 357082
rect 33948 357054 34284 357082
rect 34684 357054 35020 357082
rect 35328 357054 35664 357082
rect 36064 357054 36400 357082
rect 36800 357054 37136 357082
rect 37536 357054 37872 357082
rect 38272 357054 38424 357082
rect 39008 357054 39344 357082
rect 39652 357054 39988 357082
rect 40388 357054 40724 357082
rect 41124 357054 41368 357082
rect 41860 357054 42196 357082
rect 42596 357054 42748 357082
rect 43240 357054 43576 357082
rect 43976 357054 44128 357082
rect 44712 357054 45048 357082
rect 31680 354006 31708 357054
rect 31668 354000 31720 354006
rect 31668 353942 31720 353948
rect 32784 353870 32812 357054
rect 33520 354550 33548 357054
rect 33508 354544 33560 354550
rect 33508 354486 33560 354492
rect 34256 354210 34284 357054
rect 34244 354204 34296 354210
rect 34244 354146 34296 354152
rect 34992 354074 35020 357054
rect 35636 354482 35664 357054
rect 35624 354476 35676 354482
rect 35624 354418 35676 354424
rect 34980 354068 35032 354074
rect 34980 354010 35032 354016
rect 32772 353864 32824 353870
rect 32772 353806 32824 353812
rect 35808 353796 35860 353802
rect 35808 353738 35860 353744
rect 34520 353728 34572 353734
rect 34520 353670 34572 353676
rect 31852 353592 31904 353598
rect 31852 353534 31904 353540
rect 31392 353456 31444 353462
rect 31392 353398 31444 353404
rect 22848 348894 23138 348922
rect 23952 348894 24242 348922
rect 25056 348894 25346 348922
rect 26252 348894 26358 348922
rect 27080 348894 27462 348922
rect 28184 348894 28566 348922
rect 29288 348894 29670 348922
rect 30392 348894 30682 348922
rect 31864 348786 31892 353534
rect 34428 353524 34480 353530
rect 34428 353466 34480 353472
rect 33508 353388 33560 353394
rect 33508 353330 33560 353336
rect 32588 353320 32640 353326
rect 32588 353262 32640 353268
rect 32600 348922 32628 353262
rect 33520 348922 33548 353330
rect 34440 350554 34468 353466
rect 34532 351558 34560 353670
rect 34520 351552 34572 351558
rect 34520 351494 34572 351500
rect 35820 350554 35848 353738
rect 36372 353326 36400 357054
rect 36728 354000 36780 354006
rect 36728 353942 36780 353948
rect 36360 353320 36412 353326
rect 36360 353262 36412 353268
rect 36740 351830 36768 353942
rect 37108 353598 37136 357054
rect 37844 354142 37872 357054
rect 37832 354136 37884 354142
rect 37832 354078 37884 354084
rect 38396 354006 38424 357054
rect 38660 354544 38712 354550
rect 38660 354486 38712 354492
rect 38384 354000 38436 354006
rect 38384 353942 38436 353948
rect 37832 353864 37884 353870
rect 37832 353806 37884 353812
rect 37096 353592 37148 353598
rect 37096 353534 37148 353540
rect 37096 353456 37148 353462
rect 37096 353398 37148 353404
rect 36728 351824 36780 351830
rect 36728 351766 36780 351772
rect 36820 351552 36872 351558
rect 36820 351494 36872 351500
rect 34440 350526 34560 350554
rect 35820 350526 35940 350554
rect 34532 348922 34560 350526
rect 35912 348922 35940 350526
rect 36832 348922 36860 351494
rect 37108 350810 37136 353398
rect 37844 351558 37872 353806
rect 38672 351626 38700 354486
rect 39316 354414 39344 357054
rect 39960 354686 39988 357054
rect 39948 354680 40000 354686
rect 39948 354622 40000 354628
rect 40316 354476 40368 354482
rect 40316 354418 40368 354424
rect 39304 354408 39356 354414
rect 39304 354350 39356 354356
rect 39212 354204 39264 354210
rect 39212 354146 39264 354152
rect 39028 351824 39080 351830
rect 39028 351766 39080 351772
rect 38660 351620 38712 351626
rect 38660 351562 38712 351568
rect 37832 351552 37884 351558
rect 37832 351494 37884 351500
rect 37096 350804 37148 350810
rect 37096 350746 37148 350752
rect 37924 350804 37976 350810
rect 37924 350746 37976 350752
rect 37936 348922 37964 350746
rect 39040 348922 39068 351766
rect 39224 351218 39252 354146
rect 40040 354068 40092 354074
rect 40040 354010 40092 354016
rect 40052 351286 40080 354010
rect 40132 351552 40184 351558
rect 40132 351494 40184 351500
rect 40040 351280 40092 351286
rect 40040 351222 40092 351228
rect 39212 351212 39264 351218
rect 39212 351154 39264 351160
rect 40144 348922 40172 351494
rect 40328 351490 40356 354418
rect 40696 353666 40724 357054
rect 41340 353802 41368 357054
rect 41328 353796 41380 353802
rect 41328 353738 41380 353744
rect 42168 353734 42196 357054
rect 42720 354210 42748 357054
rect 42708 354204 42760 354210
rect 42708 354146 42760 354152
rect 42800 354136 42852 354142
rect 42800 354078 42852 354084
rect 42156 353728 42208 353734
rect 42156 353670 42208 353676
rect 40684 353660 40736 353666
rect 40684 353602 40736 353608
rect 42248 353592 42300 353598
rect 42248 353534 42300 353540
rect 41420 353320 41472 353326
rect 41420 353262 41472 353268
rect 40316 351484 40368 351490
rect 40316 351426 40368 351432
rect 41432 351422 41460 353262
rect 41512 351620 41564 351626
rect 41512 351562 41564 351568
rect 41420 351416 41472 351422
rect 41420 351358 41472 351364
rect 32600 348894 32890 348922
rect 33520 348894 33902 348922
rect 34532 348894 35006 348922
rect 35912 348894 36110 348922
rect 36832 348894 37214 348922
rect 37936 348894 38226 348922
rect 39040 348894 39330 348922
rect 40144 348894 40434 348922
rect 41524 348786 41552 351562
rect 42260 351218 42288 353534
rect 42812 351354 42840 354078
rect 43548 353598 43576 357054
rect 44100 354074 44128 357054
rect 45020 354550 45048 357054
rect 45434 356810 45462 357068
rect 46184 357054 46520 357082
rect 45434 356782 45508 356810
rect 45008 354544 45060 354550
rect 45008 354486 45060 354492
rect 45480 354278 45508 356782
rect 46492 354482 46520 357054
rect 46814 356810 46842 357068
rect 47564 357054 47900 357082
rect 46814 356782 46888 356810
rect 46480 354476 46532 354482
rect 46480 354418 46532 354424
rect 46860 354346 46888 356782
rect 46848 354340 46900 354346
rect 46848 354282 46900 354288
rect 45468 354272 45520 354278
rect 45468 354214 45520 354220
rect 47872 354142 47900 357054
rect 48240 357054 48300 357082
rect 49036 357054 49372 357082
rect 49772 357054 50108 357082
rect 50416 357054 50752 357082
rect 51152 357054 51488 357082
rect 51888 357054 52224 357082
rect 52624 357054 52960 357082
rect 53360 357054 53696 357082
rect 54004 357054 54340 357082
rect 54740 357054 55076 357082
rect 55476 357054 55812 357082
rect 56212 357054 56548 357082
rect 56948 357054 57284 357082
rect 57684 357054 57836 357082
rect 58328 357054 58664 357082
rect 59064 357054 59308 357082
rect 59800 357054 60136 357082
rect 60536 357054 60688 357082
rect 61272 357054 61608 357082
rect 61916 357054 62068 357082
rect 62652 357054 62988 357082
rect 48240 354634 48268 357054
rect 48240 354618 48360 354634
rect 48240 354612 48372 354618
rect 48240 354606 48320 354612
rect 48320 354554 48372 354560
rect 47860 354136 47912 354142
rect 47860 354078 47912 354084
rect 44088 354068 44140 354074
rect 44088 354010 44140 354016
rect 49344 354006 49372 357054
rect 49700 354408 49752 354414
rect 49700 354350 49752 354356
rect 48596 354000 48648 354006
rect 48596 353942 48648 353948
rect 49332 354000 49384 354006
rect 49332 353942 49384 353948
rect 43536 353592 43588 353598
rect 43536 353534 43588 353540
rect 44364 351484 44416 351490
rect 44364 351426 44416 351432
rect 43444 351416 43496 351422
rect 43444 351358 43496 351364
rect 42800 351348 42852 351354
rect 42800 351290 42852 351296
rect 43260 351280 43312 351286
rect 43260 351222 43312 351228
rect 42156 351212 42208 351218
rect 42156 351154 42208 351160
rect 42248 351212 42300 351218
rect 42248 351154 42300 351160
rect 42168 348922 42196 351154
rect 43272 348922 43300 351222
rect 43456 351218 43484 351358
rect 43444 351212 43496 351218
rect 43444 351154 43496 351160
rect 44376 348922 44404 351426
rect 47676 351348 47728 351354
rect 47676 351290 47728 351296
rect 46572 351280 46624 351286
rect 46572 351222 46624 351228
rect 45652 351212 45704 351218
rect 45652 351154 45704 351160
rect 45664 348922 45692 351154
rect 46584 348922 46612 351222
rect 47688 348922 47716 351290
rect 48608 348922 48636 353942
rect 49712 348922 49740 354350
rect 50080 353938 50108 357054
rect 50724 354414 50752 357054
rect 51460 354686 51488 357054
rect 50988 354680 51040 354686
rect 50988 354622 51040 354628
rect 51448 354680 51500 354686
rect 51448 354622 51500 354628
rect 50712 354408 50764 354414
rect 50712 354350 50764 354356
rect 50068 353932 50120 353938
rect 50068 353874 50120 353880
rect 51000 351778 51028 354622
rect 51908 353660 51960 353666
rect 51908 353602 51960 353608
rect 51000 351750 51120 351778
rect 51092 348922 51120 351750
rect 51920 348922 51948 353602
rect 52196 351354 52224 357054
rect 52932 352578 52960 357054
rect 53012 353796 53064 353802
rect 53012 353738 53064 353744
rect 52920 352572 52972 352578
rect 52920 352514 52972 352520
rect 52184 351348 52236 351354
rect 52184 351290 52236 351296
rect 53024 348922 53052 353738
rect 53668 351286 53696 357054
rect 54312 353802 54340 357054
rect 54300 353796 54352 353802
rect 54300 353738 54352 353744
rect 54116 353728 54168 353734
rect 54116 353670 54168 353676
rect 53656 351280 53708 351286
rect 53656 351222 53708 351228
rect 54128 348922 54156 353670
rect 55048 351218 55076 357054
rect 55128 354204 55180 354210
rect 55128 354146 55180 354152
rect 55140 351778 55168 354146
rect 55784 353870 55812 357054
rect 56520 354210 56548 357054
rect 56968 354544 57020 354550
rect 56968 354486 57020 354492
rect 56508 354204 56560 354210
rect 56508 354146 56560 354152
rect 55772 353864 55824 353870
rect 55772 353806 55824 353812
rect 56140 353592 56192 353598
rect 56140 353534 56192 353540
rect 55140 351750 55260 351778
rect 55036 351212 55088 351218
rect 55036 351154 55088 351160
rect 55232 348922 55260 351750
rect 56152 348922 56180 353534
rect 56980 351490 57008 354486
rect 57256 354362 57284 357054
rect 57072 354334 57284 354362
rect 57072 352918 57100 354334
rect 57152 354272 57204 354278
rect 57152 354214 57204 354220
rect 57060 352912 57112 352918
rect 57060 352854 57112 352860
rect 56968 351484 57020 351490
rect 56968 351426 57020 351432
rect 57164 351150 57192 354214
rect 57244 354068 57296 354074
rect 57244 354010 57296 354016
rect 57152 351144 57204 351150
rect 57152 351086 57204 351092
rect 57256 348922 57284 354010
rect 57808 351762 57836 357054
rect 58636 354550 58664 357054
rect 58624 354544 58676 354550
rect 58624 354486 58676 354492
rect 58072 354476 58124 354482
rect 58072 354418 58124 354424
rect 58084 351898 58112 354418
rect 58624 354340 58676 354346
rect 58624 354282 58676 354288
rect 58072 351892 58124 351898
rect 58072 351834 58124 351840
rect 57796 351756 57848 351762
rect 57796 351698 57848 351704
rect 58348 351484 58400 351490
rect 58348 351426 58400 351432
rect 58360 348922 58388 351426
rect 58636 351422 58664 354282
rect 59280 354278 59308 357054
rect 59636 354612 59688 354618
rect 59636 354554 59688 354560
rect 59268 354272 59320 354278
rect 59268 354214 59320 354220
rect 59360 354136 59412 354142
rect 59360 354078 59412 354084
rect 59372 351490 59400 354078
rect 59648 351626 59676 354554
rect 60108 352850 60136 357054
rect 60096 352844 60148 352850
rect 60096 352786 60148 352792
rect 60660 351694 60688 357054
rect 61580 354618 61608 357054
rect 61568 354612 61620 354618
rect 61568 354554 61620 354560
rect 62040 354346 62068 357054
rect 62212 354408 62264 354414
rect 62212 354350 62264 354356
rect 62028 354340 62080 354346
rect 62028 354282 62080 354288
rect 62120 353932 62172 353938
rect 62120 353874 62172 353880
rect 60740 351892 60792 351898
rect 60740 351834 60792 351840
rect 60648 351688 60700 351694
rect 60648 351630 60700 351636
rect 59636 351620 59688 351626
rect 59636 351562 59688 351568
rect 59360 351484 59412 351490
rect 59360 351426 59412 351432
rect 58624 351416 58676 351422
rect 58624 351358 58676 351364
rect 59452 351144 59504 351150
rect 59452 351086 59504 351092
rect 59464 348922 59492 351086
rect 60752 348922 60780 351834
rect 61660 351416 61712 351422
rect 61660 351358 61712 351364
rect 61672 348922 61700 351358
rect 62132 351082 62160 353874
rect 62224 351422 62252 354350
rect 62960 352782 62988 357054
rect 63374 356810 63402 357068
rect 64124 357054 64460 357082
rect 63374 356782 63448 356810
rect 62948 352776 63000 352782
rect 62948 352718 63000 352724
rect 63420 351762 63448 356782
rect 63592 354680 63644 354686
rect 63592 354622 63644 354628
rect 63500 353796 63552 353802
rect 63500 353738 63552 353744
rect 63512 353190 63540 353738
rect 63500 353184 63552 353190
rect 63500 353126 63552 353132
rect 63408 351756 63460 351762
rect 63408 351698 63460 351704
rect 63604 351490 63632 354622
rect 64432 354142 64460 357054
rect 64800 357054 64860 357082
rect 65504 357054 65840 357082
rect 64800 354414 64828 357054
rect 64788 354408 64840 354414
rect 64788 354350 64840 354356
rect 64420 354136 64472 354142
rect 64420 354078 64472 354084
rect 64972 354000 65024 354006
rect 64972 353942 65024 353948
rect 63684 351620 63736 351626
rect 63684 351562 63736 351568
rect 63776 351620 63828 351626
rect 63776 351562 63828 351568
rect 62764 351484 62816 351490
rect 62764 351426 62816 351432
rect 63592 351484 63644 351490
rect 63592 351426 63644 351432
rect 62212 351416 62264 351422
rect 62212 351358 62264 351364
rect 62120 351076 62172 351082
rect 62120 351018 62172 351024
rect 62776 348922 62804 351426
rect 63696 348922 63724 351562
rect 63788 351422 63816 351562
rect 63776 351416 63828 351422
rect 63776 351358 63828 351364
rect 64984 348922 65012 353942
rect 65812 352714 65840 357054
rect 66180 357054 66240 357082
rect 66976 357054 67312 357082
rect 67712 357054 68048 357082
rect 68448 357054 68784 357082
rect 69092 357054 69428 357082
rect 69828 357054 70164 357082
rect 70564 357054 70900 357082
rect 71300 357054 71636 357082
rect 72036 357054 72372 357082
rect 72680 357054 73016 357082
rect 73416 357054 73752 357082
rect 74152 357054 74488 357082
rect 74888 357054 75224 357082
rect 75624 357054 75868 357082
rect 65800 352708 65852 352714
rect 65800 352650 65852 352656
rect 66180 351694 66208 357054
rect 67284 354074 67312 357054
rect 68020 354482 68048 357054
rect 68008 354476 68060 354482
rect 68008 354418 68060 354424
rect 67272 354068 67324 354074
rect 67272 354010 67324 354016
rect 67548 353864 67600 353870
rect 67548 353806 67600 353812
rect 67560 353122 67588 353806
rect 67548 353116 67600 353122
rect 67548 353058 67600 353064
rect 68756 352646 68784 357054
rect 68928 354544 68980 354550
rect 68928 354486 68980 354492
rect 68940 353054 68968 354486
rect 68928 353048 68980 353054
rect 68928 352990 68980 352996
rect 68744 352640 68796 352646
rect 68744 352582 68796 352588
rect 66168 351688 66220 351694
rect 66168 351630 66220 351636
rect 69400 351626 69428 357054
rect 70136 354006 70164 357054
rect 70400 354612 70452 354618
rect 70400 354554 70452 354560
rect 70124 354000 70176 354006
rect 70124 353942 70176 353948
rect 70412 352986 70440 354554
rect 70872 354550 70900 357054
rect 70860 354544 70912 354550
rect 70860 354486 70912 354492
rect 70400 352980 70452 352986
rect 70400 352922 70452 352928
rect 71608 352578 71636 357054
rect 72344 353274 72372 357054
rect 72252 353246 72372 353274
rect 70400 352572 70452 352578
rect 70400 352514 70452 352520
rect 71596 352572 71648 352578
rect 71596 352514 71648 352520
rect 66996 351620 67048 351626
rect 66996 351562 67048 351568
rect 69388 351620 69440 351626
rect 69388 351562 69440 351568
rect 66352 351076 66404 351082
rect 66352 351018 66404 351024
rect 42168 348894 42550 348922
rect 43272 348894 43654 348922
rect 44376 348894 44758 348922
rect 45664 348894 45770 348922
rect 46584 348894 46874 348922
rect 47688 348894 47978 348922
rect 48608 348894 48990 348922
rect 49712 348894 50094 348922
rect 51092 348894 51198 348922
rect 51920 348894 52302 348922
rect 53024 348894 53314 348922
rect 54128 348894 54418 348922
rect 55232 348894 55522 348922
rect 56152 348894 56534 348922
rect 57256 348894 57638 348922
rect 58360 348894 58742 348922
rect 59464 348894 59846 348922
rect 60752 348894 60858 348922
rect 61672 348894 61962 348922
rect 62776 348894 63066 348922
rect 63696 348894 64078 348922
rect 64984 348894 65182 348922
rect 66364 348786 66392 351018
rect 67008 348922 67036 351562
rect 68100 351484 68152 351490
rect 68100 351426 68152 351432
rect 68112 348922 68140 351426
rect 69204 351348 69256 351354
rect 69204 351290 69256 351296
rect 69216 348922 69244 351290
rect 70412 348922 70440 352514
rect 72252 351490 72280 353246
rect 72332 353184 72384 353190
rect 72332 353126 72384 353132
rect 72240 351484 72292 351490
rect 72240 351426 72292 351432
rect 71228 351280 71280 351286
rect 71228 351222 71280 351228
rect 71240 348922 71268 351222
rect 72344 348922 72372 353126
rect 72988 351354 73016 357054
rect 73724 351558 73752 357054
rect 73712 351552 73764 351558
rect 73712 351494 73764 351500
rect 72976 351348 73028 351354
rect 72976 351290 73028 351296
rect 74460 351286 74488 357054
rect 74724 353116 74776 353122
rect 74724 353058 74776 353064
rect 74448 351280 74500 351286
rect 74448 351222 74500 351228
rect 73436 351212 73488 351218
rect 73436 351154 73488 351160
rect 73448 348922 73476 351154
rect 74736 348922 74764 353058
rect 75196 351422 75224 357054
rect 75184 351416 75236 351422
rect 75184 351358 75236 351364
rect 75840 351218 75868 357054
rect 80060 354544 80112 354550
rect 80060 354486 80112 354492
rect 79324 354408 79376 354414
rect 79324 354350 79376 354356
rect 78588 354340 78640 354346
rect 78588 354282 78640 354288
rect 77208 354272 77260 354278
rect 77208 354214 77260 354220
rect 76012 354204 76064 354210
rect 76012 354146 76064 354152
rect 75828 351212 75880 351218
rect 75828 351154 75880 351160
rect 67008 348894 67390 348922
rect 68112 348894 68402 348922
rect 69216 348894 69506 348922
rect 70412 348894 70610 348922
rect 71240 348894 71622 348922
rect 72344 348894 72726 348922
rect 73448 348894 73830 348922
rect 74736 348894 74934 348922
rect 76024 348786 76052 354146
rect 76748 352912 76800 352918
rect 76748 352854 76800 352860
rect 76760 348922 76788 352854
rect 77220 351150 77248 354214
rect 77852 351892 77904 351898
rect 77852 351834 77904 351840
rect 77208 351144 77260 351150
rect 77208 351086 77260 351092
rect 77864 348922 77892 351834
rect 78600 351082 78628 354282
rect 78772 353048 78824 353054
rect 78772 352990 78824 352996
rect 78588 351076 78640 351082
rect 78588 351018 78640 351024
rect 78784 348922 78812 352990
rect 79336 351014 79364 354350
rect 80072 351898 80100 354486
rect 80152 354476 80204 354482
rect 80152 354418 80204 354424
rect 80060 351892 80112 351898
rect 80060 351834 80112 351840
rect 80164 351150 80192 354418
rect 87420 354136 87472 354142
rect 87420 354078 87472 354084
rect 83188 352980 83240 352986
rect 83188 352922 83240 352928
rect 80980 352844 81032 352850
rect 80980 352786 81032 352792
rect 80060 351144 80112 351150
rect 80060 351086 80112 351092
rect 80152 351144 80204 351150
rect 80152 351086 80204 351092
rect 79324 351008 79376 351014
rect 79324 350950 79376 350956
rect 80072 348922 80100 351086
rect 80992 348922 81020 352786
rect 82084 351824 82136 351830
rect 82084 351766 82136 351772
rect 82096 348922 82124 351766
rect 83200 348922 83228 352922
rect 85580 352776 85632 352782
rect 85580 352718 85632 352724
rect 84384 351076 84436 351082
rect 84384 351018 84436 351024
rect 84396 348922 84424 351018
rect 85592 348922 85620 352718
rect 86316 351756 86368 351762
rect 86316 351698 86368 351704
rect 86328 348922 86356 351698
rect 87432 348922 87460 354078
rect 91836 354068 91888 354074
rect 91836 354010 91888 354016
rect 89720 352708 89772 352714
rect 89720 352650 89772 352656
rect 88524 351008 88576 351014
rect 88524 350950 88576 350956
rect 88536 348922 88564 350950
rect 89732 348922 89760 352650
rect 90732 351688 90784 351694
rect 90732 351630 90784 351636
rect 90744 348922 90772 351630
rect 91848 348922 91876 354010
rect 96068 354000 96120 354006
rect 96068 353942 96120 353948
rect 94044 352640 94096 352646
rect 94044 352582 94096 352588
rect 92940 351144 92992 351150
rect 92940 351086 92992 351092
rect 92952 348922 92980 351086
rect 94056 348922 94084 352582
rect 95240 351620 95292 351626
rect 95240 351562 95292 351568
rect 95252 348922 95280 351562
rect 96080 348922 96108 353942
rect 98276 352572 98328 352578
rect 98276 352514 98328 352520
rect 97172 351892 97224 351898
rect 97172 351834 97224 351840
rect 97184 348922 97212 351834
rect 98288 348922 98316 352514
rect 114006 351792 114062 351801
rect 114006 351727 114062 351736
rect 111706 351656 111762 351665
rect 111706 351591 111762 351600
rect 101404 351552 101456 351558
rect 101404 351494 101456 351500
rect 110694 351520 110750 351529
rect 99380 351484 99432 351490
rect 99380 351426 99432 351432
rect 99392 348922 99420 351426
rect 100852 351348 100904 351354
rect 100852 351290 100904 351296
rect 76760 348894 77050 348922
rect 77864 348894 78154 348922
rect 78784 348894 79166 348922
rect 80072 348894 80270 348922
rect 80992 348894 81374 348922
rect 82096 348894 82478 348922
rect 83200 348894 83490 348922
rect 84396 348894 84594 348922
rect 85592 348894 85698 348922
rect 86328 348894 86710 348922
rect 87432 348894 87814 348922
rect 88536 348894 88918 348922
rect 89732 348894 90022 348922
rect 90744 348894 91034 348922
rect 91848 348894 92138 348922
rect 92952 348894 93242 348922
rect 94056 348894 94254 348922
rect 95252 348894 95358 348922
rect 96080 348894 96462 348922
rect 97184 348894 97566 348922
rect 98288 348894 98578 348922
rect 99392 348894 99682 348922
rect 100864 348786 100892 351290
rect 101416 348922 101444 351494
rect 110694 351455 110750 351464
rect 103704 351416 103756 351422
rect 103704 351358 103756 351364
rect 108670 351384 108726 351393
rect 102508 351280 102560 351286
rect 102508 351222 102560 351228
rect 102520 348922 102548 351222
rect 103716 348922 103744 351358
rect 108670 351319 108726 351328
rect 104900 351212 104952 351218
rect 104900 351154 104952 351160
rect 104912 348922 104940 351154
rect 107566 351112 107622 351121
rect 107566 351047 107622 351056
rect 106188 350600 106240 350606
rect 106188 350542 106240 350548
rect 101416 348894 101798 348922
rect 102520 348894 102902 348922
rect 103716 348894 104006 348922
rect 104912 348894 105110 348922
rect 106200 348786 106228 350542
rect 107580 348786 107608 351047
rect 108684 348786 108712 351319
rect 109590 351248 109646 351257
rect 109590 351183 109646 351192
rect 109604 348786 109632 351183
rect 110708 348786 110736 351455
rect 111720 348786 111748 351591
rect 112904 350668 112956 350674
rect 112904 350610 112956 350616
rect 112916 348786 112944 350610
rect 114020 348786 114048 351727
rect 117134 350976 117190 350985
rect 117134 350911 117190 350920
rect 115110 350840 115166 350849
rect 115110 350775 115166 350784
rect 115124 348786 115152 350775
rect 115756 350736 115808 350742
rect 115756 350678 115808 350684
rect 115768 348922 115796 350678
rect 115768 348894 115874 348922
rect 117148 348786 117176 350911
rect 118620 349058 118648 400823
rect 122654 351792 122710 351801
rect 122654 351727 122710 351736
rect 121368 351348 121420 351354
rect 121368 351290 121420 351296
rect 120448 351280 120500 351286
rect 120448 351222 120500 351228
rect 119344 351212 119396 351218
rect 119344 351154 119396 351160
rect 118252 349030 118648 349058
rect 118252 348786 118280 349030
rect 119356 348786 119384 351154
rect 120460 348786 120488 351222
rect 121380 348786 121408 351290
rect 122668 350713 122696 351727
rect 122654 350704 122710 350713
rect 122654 350639 122710 350648
rect 122760 348786 122788 400862
rect 123760 351552 123812 351558
rect 123760 351494 123812 351500
rect 123772 348786 123800 351494
rect 124680 350940 124732 350946
rect 124680 350882 124732 350888
rect 124692 348786 124720 350882
rect 125428 348922 125456 400930
rect 125520 350946 125548 400959
rect 125508 350940 125560 350946
rect 125508 350882 125560 350888
rect 125428 348894 125534 348922
rect 126900 348786 126928 401095
rect 127992 351620 128044 351626
rect 127992 351562 128044 351568
rect 128004 348786 128032 351562
rect 129660 351490 129688 401231
rect 130200 351552 130252 351558
rect 130200 351494 130252 351500
rect 129096 351484 129148 351490
rect 129096 351426 129148 351432
rect 129648 351484 129700 351490
rect 129648 351426 129700 351432
rect 129108 348786 129136 351426
rect 130212 348786 130240 351494
rect 131040 348786 131068 401367
rect 136548 401338 136600 401344
rect 135168 401260 135220 401266
rect 135168 401202 135220 401208
rect 132408 401124 132460 401130
rect 132408 401066 132460 401072
rect 132420 349058 132448 401066
rect 133788 401056 133840 401062
rect 133788 400998 133840 401004
rect 133800 351626 133828 400998
rect 133328 351620 133380 351626
rect 133328 351562 133380 351568
rect 133788 351620 133840 351626
rect 133788 351562 133840 351568
rect 132236 349030 132448 349058
rect 132236 348786 132264 349030
rect 133340 348786 133368 351562
rect 135180 350946 135208 401202
rect 136456 401192 136508 401198
rect 136456 401134 136508 401140
rect 136468 351626 136496 401134
rect 135536 351620 135588 351626
rect 135536 351562 135588 351568
rect 136456 351620 136508 351626
rect 136456 351562 136508 351568
rect 134432 350940 134484 350946
rect 134432 350882 134484 350888
rect 135168 350940 135220 350946
rect 135168 350882 135220 350888
rect 134444 348786 134472 350882
rect 135548 348786 135576 351562
rect 136560 348786 136588 401338
rect 137928 401328 137980 401334
rect 137928 401270 137980 401276
rect 137940 348922 137968 401270
rect 139320 351898 139348 401406
rect 140608 351898 140636 401474
rect 138848 351892 138900 351898
rect 138848 351834 138900 351840
rect 139308 351892 139360 351898
rect 139308 351834 139360 351840
rect 139768 351892 139820 351898
rect 139768 351834 139820 351840
rect 140596 351892 140648 351898
rect 140596 351834 140648 351840
rect 137756 348894 137968 348922
rect 137756 348786 137784 348894
rect 138860 348786 138888 351834
rect 139780 348786 139808 351834
rect 140700 348786 140728 401542
rect 142068 400852 142120 400858
rect 142068 400794 142120 400800
rect 142080 348786 142108 400794
rect 143448 400784 143500 400790
rect 143448 400726 143500 400732
rect 143460 351898 143488 400726
rect 144828 400716 144880 400722
rect 144828 400658 144880 400664
rect 144840 351898 144868 400658
rect 146208 400648 146260 400654
rect 146208 400590 146260 400596
rect 146116 400308 146168 400314
rect 146116 400250 146168 400256
rect 146128 351898 146156 400250
rect 142988 351892 143040 351898
rect 142988 351834 143040 351840
rect 143448 351892 143500 351898
rect 143448 351834 143500 351840
rect 144184 351892 144236 351898
rect 144184 351834 144236 351840
rect 144828 351892 144880 351898
rect 144828 351834 144880 351840
rect 145288 351892 145340 351898
rect 145288 351834 145340 351840
rect 146116 351892 146168 351898
rect 146116 351834 146168 351840
rect 142618 351248 142674 351257
rect 142618 351183 142674 351192
rect 142802 351248 142858 351257
rect 142802 351183 142858 351192
rect 142632 350713 142660 351183
rect 142816 350985 142844 351183
rect 142802 350976 142858 350985
rect 142802 350911 142858 350920
rect 142618 350704 142674 350713
rect 142618 350639 142674 350648
rect 143000 348786 143028 351834
rect 144196 348786 144224 351834
rect 145300 348786 145328 351834
rect 146220 348786 146248 400590
rect 147126 389464 147182 389473
rect 147126 389399 147182 389408
rect 147140 386481 147168 389399
rect 147126 386472 147182 386481
rect 147126 386407 147182 386416
rect 147586 351928 147642 351937
rect 147586 351863 147642 351872
rect 146942 351792 146998 351801
rect 146942 351727 146998 351736
rect 147218 351792 147274 351801
rect 147218 351727 147274 351736
rect 146298 350976 146354 350985
rect 146298 350911 146354 350920
rect 146312 350674 146340 350911
rect 146300 350668 146352 350674
rect 146300 350610 146352 350616
rect 146956 348922 146984 351727
rect 147232 351529 147260 351727
rect 147218 351520 147274 351529
rect 147218 351455 147274 351464
rect 147600 350577 147628 351863
rect 147678 351792 147734 351801
rect 147678 351727 147734 351736
rect 148046 351792 148102 351801
rect 148046 351727 148102 351736
rect 149426 351792 149482 351801
rect 149426 351727 149482 351736
rect 150070 351792 150126 351801
rect 150070 351727 150126 351736
rect 151174 351792 151230 351801
rect 151174 351727 151230 351736
rect 152370 351792 152426 351801
rect 152370 351727 152426 351736
rect 147692 351529 147720 351727
rect 147678 351520 147734 351529
rect 147678 351455 147734 351464
rect 147586 350568 147642 350577
rect 147586 350503 147642 350512
rect 148060 348922 148088 351727
rect 149058 350840 149114 350849
rect 149058 350775 149114 350784
rect 149072 350742 149100 350775
rect 149060 350736 149112 350742
rect 149060 350678 149112 350684
rect 146956 348894 147062 348922
rect 148060 348894 148166 348922
rect 149440 348786 149468 351727
rect 150084 348922 150112 351727
rect 151188 348922 151216 351727
rect 152384 348922 152412 351727
rect 153198 351384 153254 351393
rect 153304 351354 153332 500278
rect 153384 500268 153436 500274
rect 153384 500210 153436 500216
rect 153198 351319 153254 351328
rect 153292 351348 153344 351354
rect 153212 350606 153240 351319
rect 153292 351290 153344 351296
rect 153396 351286 153424 500210
rect 153476 497548 153528 497554
rect 153476 497490 153528 497496
rect 153384 351280 153436 351286
rect 153384 351222 153436 351228
rect 153488 351218 153516 497490
rect 153580 400858 153608 500783
rect 153672 401402 153700 500890
rect 153844 500812 153896 500818
rect 153844 500754 153896 500760
rect 153752 500064 153804 500070
rect 153752 500006 153804 500012
rect 153764 401606 153792 500006
rect 153752 401600 153804 401606
rect 153752 401542 153804 401548
rect 153660 401396 153712 401402
rect 153660 401338 153712 401344
rect 153856 401266 153884 500754
rect 154028 499996 154080 500002
rect 154028 499938 154080 499944
rect 153936 499792 153988 499798
rect 153936 499734 153988 499740
rect 153844 401260 153896 401266
rect 153844 401202 153896 401208
rect 153568 400852 153620 400858
rect 153568 400794 153620 400800
rect 153948 400314 153976 499734
rect 154040 400790 154068 499938
rect 154408 492726 154436 502143
rect 154120 492720 154172 492726
rect 154304 492720 154356 492726
rect 154120 492662 154172 492668
rect 154210 492688 154266 492697
rect 154028 400784 154080 400790
rect 154028 400726 154080 400732
rect 154132 400654 154160 492662
rect 154304 492662 154356 492668
rect 154396 492720 154448 492726
rect 154396 492662 154448 492668
rect 154210 492623 154266 492632
rect 154224 401470 154252 492623
rect 154316 491298 154344 492662
rect 154304 491292 154356 491298
rect 154304 491234 154356 491240
rect 154488 491292 154540 491298
rect 154488 491234 154540 491240
rect 154500 481710 154528 491234
rect 154304 481704 154356 481710
rect 154304 481646 154356 481652
rect 154488 481704 154540 481710
rect 154488 481646 154540 481652
rect 154316 473550 154344 481646
rect 154304 473544 154356 473550
rect 154304 473486 154356 473492
rect 154304 473408 154356 473414
rect 154304 473350 154356 473356
rect 154316 471986 154344 473350
rect 154304 471980 154356 471986
rect 154304 471922 154356 471928
rect 154488 471980 154540 471986
rect 154488 471922 154540 471928
rect 154500 462398 154528 471922
rect 154304 462392 154356 462398
rect 154304 462334 154356 462340
rect 154488 462392 154540 462398
rect 154488 462334 154540 462340
rect 154316 452606 154344 462334
rect 154304 452600 154356 452606
rect 154304 452542 154356 452548
rect 154488 452600 154540 452606
rect 154488 452542 154540 452548
rect 154500 443018 154528 452542
rect 154304 443012 154356 443018
rect 154304 442954 154356 442960
rect 154488 443012 154540 443018
rect 154488 442954 154540 442960
rect 154316 433294 154344 442954
rect 154304 433288 154356 433294
rect 154304 433230 154356 433236
rect 154488 433288 154540 433294
rect 154488 433230 154540 433236
rect 154500 423706 154528 433230
rect 154304 423700 154356 423706
rect 154304 423642 154356 423648
rect 154488 423700 154540 423706
rect 154488 423642 154540 423648
rect 154316 413982 154344 423642
rect 154304 413976 154356 413982
rect 154304 413918 154356 413924
rect 154488 413976 154540 413982
rect 154488 413918 154540 413924
rect 154500 404394 154528 413918
rect 154304 404388 154356 404394
rect 154304 404330 154356 404336
rect 154488 404388 154540 404394
rect 154488 404330 154540 404336
rect 154212 401464 154264 401470
rect 154212 401406 154264 401412
rect 154120 400648 154172 400654
rect 154120 400590 154172 400596
rect 153936 400308 153988 400314
rect 153936 400250 153988 400256
rect 154316 394670 154344 404330
rect 154120 394664 154172 394670
rect 154120 394606 154172 394612
rect 154304 394664 154356 394670
rect 154304 394606 154356 394612
rect 154132 385082 154160 394606
rect 154120 385076 154172 385082
rect 154120 385018 154172 385024
rect 154304 385076 154356 385082
rect 154304 385018 154356 385024
rect 154316 375358 154344 385018
rect 154120 375352 154172 375358
rect 154120 375294 154172 375300
rect 154304 375352 154356 375358
rect 154304 375294 154356 375300
rect 154132 365770 154160 375294
rect 153844 365764 153896 365770
rect 153844 365706 153896 365712
rect 154120 365764 154172 365770
rect 154120 365706 154172 365712
rect 153856 357474 153884 365706
rect 153844 357468 153896 357474
rect 153844 357410 153896 357416
rect 153936 357468 153988 357474
rect 153936 357410 153988 357416
rect 153476 351212 153528 351218
rect 153476 351154 153528 351160
rect 153200 350600 153252 350606
rect 153200 350542 153252 350548
rect 150084 348894 150374 348922
rect 151188 348894 151386 348922
rect 152384 348894 152490 348922
rect 153948 348786 153976 357410
rect 154592 348922 154620 502846
rect 155132 500880 155184 500886
rect 155132 500822 155184 500828
rect 154764 500608 154816 500614
rect 154764 500550 154816 500556
rect 154776 351558 154804 500550
rect 154856 500540 154908 500546
rect 154856 500482 154908 500488
rect 154764 351552 154816 351558
rect 154764 351494 154816 351500
rect 154868 351490 154896 500482
rect 154948 500404 155000 500410
rect 154948 500346 155000 500352
rect 154856 351484 154908 351490
rect 154856 351426 154908 351432
rect 154960 351422 154988 500346
rect 155040 500132 155092 500138
rect 155040 500074 155092 500080
rect 155052 401538 155080 500074
rect 155040 401532 155092 401538
rect 155040 401474 155092 401480
rect 155144 401334 155172 500822
rect 155316 500744 155368 500750
rect 155316 500686 155368 500692
rect 155224 500472 155276 500478
rect 155224 500414 155276 500420
rect 155132 401328 155184 401334
rect 155132 401270 155184 401276
rect 155236 400994 155264 500414
rect 155328 401198 155356 500686
rect 155500 500676 155552 500682
rect 155500 500618 155552 500624
rect 155406 499760 155462 499769
rect 155406 499695 155462 499704
rect 155316 401192 155368 401198
rect 155316 401134 155368 401140
rect 155224 400988 155276 400994
rect 155224 400930 155276 400936
rect 155420 400722 155448 499695
rect 155512 401130 155540 500618
rect 155592 497616 155644 497622
rect 155592 497558 155644 497564
rect 155500 401124 155552 401130
rect 155500 401066 155552 401072
rect 155604 400926 155632 497558
rect 155696 492658 155724 502860
rect 155972 502846 156814 502874
rect 157352 502846 157918 502874
rect 158732 502846 158930 502874
rect 155684 492652 155736 492658
rect 155684 492594 155736 492600
rect 155866 483032 155922 483041
rect 155866 482967 155922 482976
rect 155880 476082 155908 482967
rect 155788 476054 155908 476082
rect 155788 473346 155816 476054
rect 155776 473340 155828 473346
rect 155776 473282 155828 473288
rect 155774 463720 155830 463729
rect 155774 463655 155830 463664
rect 155788 454034 155816 463655
rect 155776 454028 155828 454034
rect 155776 453970 155828 453976
rect 155868 454028 155920 454034
rect 155868 453970 155920 453976
rect 155880 447166 155908 453970
rect 155868 447160 155920 447166
rect 155868 447102 155920 447108
rect 155776 447092 155828 447098
rect 155776 447034 155828 447040
rect 155788 444394 155816 447034
rect 155788 444366 155908 444394
rect 155880 437458 155908 444366
rect 155788 437430 155908 437458
rect 155788 429894 155816 437430
rect 155776 429888 155828 429894
rect 155776 429830 155828 429836
rect 155776 425196 155828 425202
rect 155776 425138 155828 425144
rect 155788 425066 155816 425138
rect 155776 425060 155828 425066
rect 155776 425002 155828 425008
rect 155868 425060 155920 425066
rect 155868 425002 155920 425008
rect 155880 418198 155908 425002
rect 155868 418192 155920 418198
rect 155868 418134 155920 418140
rect 155776 418124 155828 418130
rect 155776 418066 155828 418072
rect 155788 415426 155816 418066
rect 155788 415410 155908 415426
rect 155788 415404 155920 415410
rect 155788 415398 155868 415404
rect 155868 415346 155920 415352
rect 155682 405784 155738 405793
rect 155682 405719 155738 405728
rect 155592 400920 155644 400926
rect 155696 400908 155724 405719
rect 155696 400880 155908 400908
rect 155592 400862 155644 400868
rect 155408 400716 155460 400722
rect 155408 400658 155460 400664
rect 155880 396114 155908 400880
rect 155788 396086 155908 396114
rect 155788 394670 155816 396086
rect 155776 394664 155828 394670
rect 155776 394606 155828 394612
rect 155868 394664 155920 394670
rect 155868 394606 155920 394612
rect 155880 379574 155908 394606
rect 155868 379568 155920 379574
rect 155868 379510 155920 379516
rect 155684 379500 155736 379506
rect 155684 379442 155736 379448
rect 155696 376689 155724 379442
rect 155682 376680 155738 376689
rect 155682 376615 155738 376624
rect 155774 369744 155830 369753
rect 155774 369679 155830 369688
rect 155788 362302 155816 369679
rect 155500 362296 155552 362302
rect 155500 362238 155552 362244
rect 155776 362296 155828 362302
rect 155776 362238 155828 362244
rect 155512 357474 155540 362238
rect 155500 357468 155552 357474
rect 155500 357410 155552 357416
rect 155592 357468 155644 357474
rect 155592 357410 155644 357416
rect 154948 351416 155000 351422
rect 154948 351358 155000 351364
rect 155604 348922 155632 357410
rect 155972 351898 156000 502846
rect 156144 492652 156196 492658
rect 156144 492594 156196 492600
rect 156052 486464 156104 486470
rect 156052 486406 156104 486412
rect 156064 465361 156092 486406
rect 156156 483041 156184 492594
rect 156142 483032 156198 483041
rect 156142 482967 156198 482976
rect 156144 473340 156196 473346
rect 156144 473282 156196 473288
rect 156050 465352 156106 465361
rect 156050 465287 156106 465296
rect 156156 463729 156184 473282
rect 156142 463720 156198 463729
rect 156142 463655 156198 463664
rect 156052 429888 156104 429894
rect 156052 429830 156104 429836
rect 156064 425202 156092 429830
rect 156052 425196 156104 425202
rect 156052 425138 156104 425144
rect 156144 415404 156196 415410
rect 156144 415346 156196 415352
rect 156156 405929 156184 415346
rect 156142 405920 156198 405929
rect 156142 405855 156198 405864
rect 155960 351892 156012 351898
rect 155960 351834 156012 351840
rect 156420 351892 156472 351898
rect 156420 351834 156472 351840
rect 156432 348922 156460 351834
rect 154592 348894 154698 348922
rect 155604 348894 155710 348922
rect 156432 348894 156814 348922
rect 22126 348758 22232 348786
rect 31786 348758 31892 348786
rect 41446 348758 41552 348786
rect 66286 348758 66392 348786
rect 75946 348758 76052 348786
rect 100786 348758 100892 348786
rect 106122 348758 106228 348786
rect 107226 348758 107608 348786
rect 108330 348758 108712 348786
rect 109342 348758 109632 348786
rect 110446 348758 110736 348786
rect 111550 348758 111748 348786
rect 112654 348758 112944 348786
rect 113666 348758 114048 348786
rect 114770 348758 115152 348786
rect 116886 348758 117176 348786
rect 117990 348758 118280 348786
rect 119094 348758 119384 348786
rect 120198 348758 120488 348786
rect 121210 348758 121408 348786
rect 122314 348758 122788 348786
rect 123418 348758 123800 348786
rect 124430 348758 124720 348786
rect 126638 348758 126928 348786
rect 127742 348758 128032 348786
rect 128754 348758 129136 348786
rect 129858 348758 130240 348786
rect 130962 348758 131068 348786
rect 131974 348758 132264 348786
rect 133078 348758 133368 348786
rect 134182 348758 134472 348786
rect 135286 348758 135576 348786
rect 136298 348758 136588 348786
rect 137402 348758 137784 348786
rect 138506 348758 138888 348786
rect 139518 348758 139808 348786
rect 140622 348758 140728 348786
rect 141726 348758 142108 348786
rect 142830 348758 143028 348786
rect 143842 348758 144224 348786
rect 144946 348758 145328 348786
rect 146050 348758 146248 348786
rect 149270 348758 149468 348786
rect 153594 348758 153976 348786
rect 157352 348786 157380 502846
rect 157432 497684 157484 497690
rect 157432 497626 157484 497632
rect 157444 401062 157472 497626
rect 157432 401056 157484 401062
rect 157432 400998 157484 401004
rect 158732 348922 158760 502846
rect 159008 499338 159036 502982
rect 158824 499310 159036 499338
rect 160112 502846 161138 502874
rect 161492 502846 162242 502874
rect 162872 502846 163254 502874
rect 158824 495394 158852 499310
rect 158824 495366 158944 495394
rect 158916 492658 158944 495366
rect 158904 492652 158956 492658
rect 158904 492594 158956 492600
rect 158996 492652 159048 492658
rect 158996 492594 159048 492600
rect 159008 485790 159036 492594
rect 158904 485784 158956 485790
rect 158904 485726 158956 485732
rect 158996 485784 159048 485790
rect 158996 485726 159048 485732
rect 158916 483018 158944 485726
rect 158916 482990 159036 483018
rect 159008 476134 159036 482990
rect 158812 476128 158864 476134
rect 158996 476128 159048 476134
rect 158864 476076 158944 476082
rect 158812 476070 158944 476076
rect 158996 476070 159048 476076
rect 158824 476054 158944 476070
rect 158916 473346 158944 476054
rect 158904 473340 158956 473346
rect 158904 473282 158956 473288
rect 158996 473340 159048 473346
rect 158996 473282 159048 473288
rect 159008 466478 159036 473282
rect 158996 466472 159048 466478
rect 158996 466414 159048 466420
rect 158904 466404 158956 466410
rect 158904 466346 158956 466352
rect 158916 463706 158944 466346
rect 158916 463678 159036 463706
rect 159008 456822 159036 463678
rect 158812 456816 158864 456822
rect 158996 456816 159048 456822
rect 158864 456764 158944 456770
rect 158812 456758 158944 456764
rect 158996 456758 159048 456764
rect 158824 456742 158944 456758
rect 158916 454034 158944 456742
rect 158904 454028 158956 454034
rect 158904 453970 158956 453976
rect 158996 454028 159048 454034
rect 158996 453970 159048 453976
rect 159008 447166 159036 453970
rect 158996 447160 159048 447166
rect 158996 447102 159048 447108
rect 158904 447092 158956 447098
rect 158904 447034 158956 447040
rect 158916 444394 158944 447034
rect 158916 444366 159036 444394
rect 159008 437510 159036 444366
rect 158812 437504 158864 437510
rect 158996 437504 159048 437510
rect 158864 437452 158944 437458
rect 158812 437446 158944 437452
rect 158996 437446 159048 437452
rect 158824 437430 158944 437446
rect 158916 434722 158944 437430
rect 158904 434716 158956 434722
rect 158904 434658 158956 434664
rect 158996 434716 159048 434722
rect 158996 434658 159048 434664
rect 159008 427854 159036 434658
rect 158996 427848 159048 427854
rect 158996 427790 159048 427796
rect 158904 427780 158956 427786
rect 158904 427722 158956 427728
rect 158916 425082 158944 427722
rect 158916 425054 159036 425082
rect 159008 418198 159036 425054
rect 158812 418192 158864 418198
rect 158996 418192 159048 418198
rect 158864 418140 158944 418146
rect 158812 418134 158944 418140
rect 158996 418134 159048 418140
rect 158824 418118 158944 418134
rect 158916 415410 158944 418118
rect 158904 415404 158956 415410
rect 158904 415346 158956 415352
rect 159180 415404 159232 415410
rect 159180 415346 159232 415352
rect 159192 405754 159220 415346
rect 158996 405748 159048 405754
rect 158996 405690 159048 405696
rect 159180 405748 159232 405754
rect 159180 405690 159232 405696
rect 159008 398698 159036 405690
rect 158916 398670 159036 398698
rect 158916 389178 158944 398670
rect 158916 389150 159036 389178
rect 159008 386374 159036 389150
rect 158812 386368 158864 386374
rect 158812 386310 158864 386316
rect 158996 386368 159048 386374
rect 158996 386310 159048 386316
rect 158824 379522 158852 386310
rect 158824 379494 158944 379522
rect 158916 369866 158944 379494
rect 158916 369838 159036 369866
rect 159008 360210 159036 369838
rect 158824 360182 159036 360210
rect 158824 351898 158852 360182
rect 160112 351898 160140 502846
rect 161492 351898 161520 502846
rect 158812 351892 158864 351898
rect 158812 351834 158864 351840
rect 159732 351892 159784 351898
rect 159732 351834 159784 351840
rect 160100 351892 160152 351898
rect 160100 351834 160152 351840
rect 160836 351892 160888 351898
rect 160836 351834 160888 351840
rect 161480 351892 161532 351898
rect 161480 351834 161532 351840
rect 161940 351892 161992 351898
rect 161940 351834 161992 351840
rect 159744 348922 159772 351834
rect 160848 348922 160876 351834
rect 161952 348922 161980 351834
rect 162872 348922 162900 502846
rect 164240 499180 164292 499186
rect 164240 499122 164292 499128
rect 164252 351898 164280 499122
rect 164240 351892 164292 351898
rect 164240 351834 164292 351840
rect 164344 349058 164372 502860
rect 165080 502846 165462 502874
rect 165632 502846 166474 502874
rect 167012 502846 167578 502874
rect 168392 502846 168682 502874
rect 169786 502846 169892 502874
rect 165080 499186 165108 502846
rect 165068 499180 165120 499186
rect 165068 499122 165120 499128
rect 165632 351898 165660 502846
rect 165068 351892 165120 351898
rect 165068 351834 165120 351840
rect 165620 351892 165672 351898
rect 165620 351834 165672 351840
rect 166172 351892 166224 351898
rect 166172 351834 166224 351840
rect 164252 349030 164372 349058
rect 164252 348922 164280 349030
rect 165080 348922 165108 351834
rect 166184 348922 166212 351834
rect 158732 348894 158930 348922
rect 159744 348894 160034 348922
rect 160848 348894 161138 348922
rect 161952 348894 162242 348922
rect 162872 348894 163254 348922
rect 164252 348894 164358 348922
rect 165080 348894 165462 348922
rect 166184 348894 166474 348922
rect 167012 348786 167040 502846
rect 168392 348922 168420 502846
rect 168392 348894 168682 348922
rect 169864 348786 169892 502846
rect 169956 502846 170798 502874
rect 171152 502846 171902 502874
rect 172532 502846 173006 502874
rect 169956 351490 169984 502846
rect 171152 351490 171180 502846
rect 169944 351484 169996 351490
rect 169944 351426 169996 351432
rect 170404 351484 170456 351490
rect 170404 351426 170456 351432
rect 171140 351484 171192 351490
rect 171140 351426 171192 351432
rect 171600 351484 171652 351490
rect 171600 351426 171652 351432
rect 170416 348922 170444 351426
rect 171612 348922 171640 351426
rect 172532 348922 172560 502846
rect 173900 501220 173952 501226
rect 173900 501162 173952 501168
rect 173912 351014 173940 501162
rect 173900 351008 173952 351014
rect 173900 350950 173952 350956
rect 174004 349058 174032 502860
rect 174832 502846 175122 502874
rect 175292 502846 176226 502874
rect 176672 502846 177330 502874
rect 178052 502846 178342 502874
rect 174832 501226 174860 502846
rect 174820 501220 174872 501226
rect 174820 501162 174872 501168
rect 175292 351490 175320 502846
rect 176672 351490 176700 502846
rect 175280 351484 175332 351490
rect 175280 351426 175332 351432
rect 175924 351484 175976 351490
rect 175924 351426 175976 351432
rect 176660 351484 176712 351490
rect 176660 351426 176712 351432
rect 177120 351484 177172 351490
rect 177120 351426 177172 351432
rect 174820 351008 174872 351014
rect 174820 350950 174872 350956
rect 173912 349030 174032 349058
rect 173912 348922 173940 349030
rect 174832 348922 174860 350950
rect 175936 348922 175964 351426
rect 177132 348922 177160 351426
rect 178052 348922 178080 502846
rect 179432 349058 179460 502860
rect 179524 502846 180550 502874
rect 180812 502846 181562 502874
rect 182192 502846 182666 502874
rect 183572 502846 183770 502874
rect 184584 502846 184874 502874
rect 184952 502846 185886 502874
rect 186332 502846 186990 502874
rect 187712 502846 188094 502874
rect 179524 351490 179552 502846
rect 180812 351490 180840 502846
rect 179512 351484 179564 351490
rect 179512 351426 179564 351432
rect 180156 351484 180208 351490
rect 180156 351426 180208 351432
rect 180800 351484 180852 351490
rect 180800 351426 180852 351432
rect 181260 351484 181312 351490
rect 181260 351426 181312 351432
rect 179432 349030 179552 349058
rect 170416 348894 170798 348922
rect 171612 348894 171902 348922
rect 172532 348894 173006 348922
rect 173912 348894 174018 348922
rect 174832 348894 175122 348922
rect 175936 348894 176226 348922
rect 177132 348894 177330 348922
rect 178052 348894 178342 348922
rect 179524 348786 179552 349030
rect 180168 348922 180196 351426
rect 181272 348922 181300 351426
rect 182192 348922 182220 502846
rect 183572 348922 183600 502846
rect 184584 501226 184612 502846
rect 183652 501220 183704 501226
rect 183652 501162 183704 501168
rect 184572 501220 184624 501226
rect 184572 501162 184624 501168
rect 183664 499474 183692 501162
rect 183664 499446 183784 499474
rect 183756 489954 183784 499446
rect 183756 489926 183876 489954
rect 183848 480282 183876 489926
rect 183652 480276 183704 480282
rect 183652 480218 183704 480224
rect 183836 480276 183888 480282
rect 183836 480218 183888 480224
rect 183664 480162 183692 480218
rect 183664 480134 183784 480162
rect 183756 470642 183784 480134
rect 183756 470614 183876 470642
rect 183848 460970 183876 470614
rect 183652 460964 183704 460970
rect 183652 460906 183704 460912
rect 183836 460964 183888 460970
rect 183836 460906 183888 460912
rect 183664 460850 183692 460906
rect 183664 460822 183784 460850
rect 183756 451330 183784 460822
rect 183756 451302 183876 451330
rect 183848 441658 183876 451302
rect 183652 441652 183704 441658
rect 183652 441594 183704 441600
rect 183836 441652 183888 441658
rect 183836 441594 183888 441600
rect 183664 441538 183692 441594
rect 183664 441510 183784 441538
rect 183756 432018 183784 441510
rect 183756 431990 183876 432018
rect 183848 422346 183876 431990
rect 183652 422340 183704 422346
rect 183652 422282 183704 422288
rect 183836 422340 183888 422346
rect 183836 422282 183888 422288
rect 183664 422226 183692 422282
rect 183664 422198 183784 422226
rect 183756 412706 183784 422198
rect 183756 412678 183876 412706
rect 183848 403034 183876 412678
rect 183652 403028 183704 403034
rect 183652 402970 183704 402976
rect 183836 403028 183888 403034
rect 183836 402970 183888 402976
rect 183664 402914 183692 402970
rect 183664 402886 183784 402914
rect 183756 393394 183784 402886
rect 183756 393366 183876 393394
rect 183848 383722 183876 393366
rect 183652 383716 183704 383722
rect 183652 383658 183704 383664
rect 183836 383716 183888 383722
rect 183836 383658 183888 383664
rect 183664 383602 183692 383658
rect 183664 383574 183784 383602
rect 183756 374082 183784 383574
rect 183756 374054 183876 374082
rect 183848 364410 183876 374054
rect 183652 364404 183704 364410
rect 183652 364346 183704 364352
rect 183836 364404 183888 364410
rect 183836 364346 183888 364352
rect 183664 350946 183692 364346
rect 184952 351490 184980 502846
rect 185584 485104 185636 485110
rect 185584 485046 185636 485052
rect 185596 450945 185624 485046
rect 185582 450936 185638 450945
rect 185582 450871 185638 450880
rect 184940 351484 184992 351490
rect 184940 351426 184992 351432
rect 185492 351484 185544 351490
rect 185492 351426 185544 351432
rect 183652 350940 183704 350946
rect 183652 350882 183704 350888
rect 184572 350940 184624 350946
rect 184572 350882 184624 350888
rect 184584 348922 184612 350882
rect 185504 348922 185532 351426
rect 180168 348894 180550 348922
rect 181272 348894 181562 348922
rect 182192 348894 182666 348922
rect 183572 348894 183770 348922
rect 184584 348894 184874 348922
rect 185504 348894 185886 348922
rect 157352 348758 157918 348786
rect 167012 348758 167578 348786
rect 169786 348758 169892 348786
rect 179446 348758 179552 348786
rect 186332 348786 186360 502846
rect 187424 500472 187476 500478
rect 187424 500414 187476 500420
rect 186964 376780 187016 376786
rect 186964 376722 187016 376728
rect 186976 360194 187004 376722
rect 186964 360188 187016 360194
rect 186964 360130 187016 360136
rect 187436 357542 187464 500414
rect 187608 500404 187660 500410
rect 187608 500346 187660 500352
rect 187516 500268 187568 500274
rect 187516 500210 187568 500216
rect 187424 357536 187476 357542
rect 187424 357478 187476 357484
rect 187528 351898 187556 500210
rect 187516 351892 187568 351898
rect 187516 351834 187568 351840
rect 187620 351082 187648 500346
rect 187608 351076 187660 351082
rect 187608 351018 187660 351024
rect 187712 348922 187740 502846
rect 189092 500721 189120 502860
rect 190196 500857 190224 502860
rect 191300 500857 191328 502860
rect 190182 500848 190238 500857
rect 190182 500783 190238 500792
rect 191286 500848 191342 500857
rect 191286 500783 191342 500792
rect 191840 500812 191892 500818
rect 191840 500754 191892 500760
rect 189078 500712 189134 500721
rect 189078 500647 189134 500656
rect 188620 493740 188672 493746
rect 188620 493682 188672 493688
rect 188632 491572 188660 493682
rect 189724 493400 189776 493406
rect 189724 493342 189776 493348
rect 189736 491572 189764 493342
rect 190920 492856 190972 492862
rect 190920 492798 190972 492804
rect 190932 491572 190960 492798
rect 191852 491586 191880 500754
rect 191932 500676 191984 500682
rect 191932 500618 191984 500624
rect 191944 493746 191972 500618
rect 192404 500478 192432 502860
rect 192392 500472 192444 500478
rect 192392 500414 192444 500420
rect 193416 500410 193444 502860
rect 193404 500404 193456 500410
rect 193404 500346 193456 500352
rect 194520 500274 194548 502860
rect 195624 500954 195652 502860
rect 194600 500948 194652 500954
rect 194600 500890 194652 500896
rect 195612 500948 195664 500954
rect 195612 500890 195664 500896
rect 194508 500268 194560 500274
rect 194508 500210 194560 500216
rect 194612 498846 194640 500890
rect 195060 500880 195112 500886
rect 195060 500822 195112 500828
rect 194600 498840 194652 498846
rect 194600 498782 194652 498788
rect 194508 494012 194560 494018
rect 194508 493954 194560 493960
rect 193312 493808 193364 493814
rect 193312 493750 193364 493756
rect 191932 493740 191984 493746
rect 191932 493682 191984 493688
rect 191852 491558 192142 491586
rect 193324 491572 193352 493750
rect 194520 491572 194548 493954
rect 195072 493406 195100 500822
rect 196636 500682 196664 502860
rect 197740 500886 197768 502860
rect 197728 500880 197780 500886
rect 197728 500822 197780 500828
rect 196624 500676 196676 500682
rect 196624 500618 196676 500624
rect 197176 500676 197228 500682
rect 197176 500618 197228 500624
rect 196440 500540 196492 500546
rect 196440 500482 196492 500488
rect 195888 500336 195940 500342
rect 195888 500278 195940 500284
rect 195704 493672 195756 493678
rect 195704 493614 195756 493620
rect 195060 493400 195112 493406
rect 195060 493342 195112 493348
rect 195716 491572 195744 493614
rect 195900 492862 195928 500278
rect 196452 493814 196480 500482
rect 197188 494018 197216 500618
rect 198844 500342 198872 502860
rect 199948 500818 199976 502860
rect 199936 500812 199988 500818
rect 199936 500754 199988 500760
rect 200960 500546 200988 502860
rect 201500 500948 201552 500954
rect 201500 500890 201552 500896
rect 200948 500540 201000 500546
rect 200948 500482 201000 500488
rect 198832 500336 198884 500342
rect 198832 500278 198884 500284
rect 199476 500336 199528 500342
rect 199476 500278 199528 500284
rect 197176 494012 197228 494018
rect 197176 493954 197228 493960
rect 198096 493876 198148 493882
rect 198096 493818 198148 493824
rect 196440 493808 196492 493814
rect 196440 493750 196492 493756
rect 196900 493604 196952 493610
rect 196900 493546 196952 493552
rect 195888 492856 195940 492862
rect 195888 492798 195940 492804
rect 196912 491572 196940 493546
rect 198108 491572 198136 493818
rect 199292 493808 199344 493814
rect 199292 493750 199344 493756
rect 199304 491572 199332 493750
rect 199488 493610 199516 500278
rect 200120 499792 200172 499798
rect 200120 499734 200172 499740
rect 200132 493882 200160 499734
rect 200120 493876 200172 493882
rect 200120 493818 200172 493824
rect 200488 493740 200540 493746
rect 200488 493682 200540 493688
rect 199476 493604 199528 493610
rect 199476 493546 199528 493552
rect 200500 491572 200528 493682
rect 201512 493678 201540 500890
rect 202064 500682 202092 502860
rect 203168 500954 203196 502860
rect 203156 500948 203208 500954
rect 203156 500890 203208 500896
rect 202052 500676 202104 500682
rect 202052 500618 202104 500624
rect 201592 500608 201644 500614
rect 201592 500550 201644 500556
rect 201604 493814 201632 500550
rect 203892 500472 203944 500478
rect 203892 500414 203944 500420
rect 202880 494012 202932 494018
rect 202880 493954 202932 493960
rect 201592 493808 201644 493814
rect 201592 493750 201644 493756
rect 201684 493808 201736 493814
rect 201684 493750 201736 493756
rect 201500 493672 201552 493678
rect 201500 493614 201552 493620
rect 201696 491572 201724 493750
rect 202892 491572 202920 493954
rect 203904 493746 203932 500414
rect 204180 500342 204208 502860
rect 204904 500948 204956 500954
rect 204904 500890 204956 500896
rect 204168 500336 204220 500342
rect 204168 500278 204220 500284
rect 204916 493814 204944 500890
rect 205284 499798 205312 502860
rect 205640 500880 205692 500886
rect 205640 500822 205692 500828
rect 205272 499792 205324 499798
rect 205272 499734 205324 499740
rect 205652 494018 205680 500822
rect 206388 500614 206416 502860
rect 206376 500608 206428 500614
rect 206376 500550 206428 500556
rect 207112 500608 207164 500614
rect 207112 500550 207164 500556
rect 206376 499724 206428 499730
rect 206376 499666 206428 499672
rect 205640 494012 205692 494018
rect 205640 493954 205692 493960
rect 204904 493808 204956 493814
rect 204904 493750 204956 493756
rect 203892 493740 203944 493746
rect 203892 493682 203944 493688
rect 206388 493678 206416 499666
rect 204076 493672 204128 493678
rect 204076 493614 204128 493620
rect 206376 493672 206428 493678
rect 206376 493614 206428 493620
rect 206468 493672 206520 493678
rect 206468 493614 206520 493620
rect 204088 491572 204116 493614
rect 205272 493536 205324 493542
rect 205272 493478 205324 493484
rect 205284 491572 205312 493478
rect 206480 491572 206508 493614
rect 207124 493542 207152 500550
rect 207492 500478 207520 502860
rect 208504 500954 208532 502860
rect 208492 500948 208544 500954
rect 208492 500890 208544 500896
rect 209608 500886 209636 502860
rect 209596 500880 209648 500886
rect 209596 500822 209648 500828
rect 207480 500472 207532 500478
rect 207480 500414 207532 500420
rect 209136 500404 209188 500410
rect 209136 500346 209188 500352
rect 208860 494012 208912 494018
rect 208860 493954 208912 493960
rect 207112 493536 207164 493542
rect 207112 493478 207164 493484
rect 207664 493332 207716 493338
rect 207664 493274 207716 493280
rect 207676 491572 207704 493274
rect 208872 491572 208900 493954
rect 209148 493678 209176 500346
rect 209872 500336 209924 500342
rect 209872 500278 209924 500284
rect 209136 493672 209188 493678
rect 209136 493614 209188 493620
rect 209884 493338 209912 500278
rect 210712 499730 210740 502860
rect 211724 500614 211752 502860
rect 211712 500608 211764 500614
rect 211712 500550 211764 500556
rect 211160 500472 211212 500478
rect 211160 500414 211212 500420
rect 210700 499724 210752 499730
rect 210700 499666 210752 499672
rect 211172 494018 211200 500414
rect 212828 500410 212856 502860
rect 213828 500948 213880 500954
rect 213828 500890 213880 500896
rect 212816 500404 212868 500410
rect 212816 500346 212868 500352
rect 211160 494012 211212 494018
rect 211160 493954 211212 493960
rect 213644 494012 213696 494018
rect 213644 493954 213696 493960
rect 211252 493808 211304 493814
rect 211252 493750 211304 493756
rect 210056 493740 210108 493746
rect 210056 493682 210108 493688
rect 209872 493332 209924 493338
rect 209872 493274 209924 493280
rect 210068 491572 210096 493682
rect 211264 491572 211292 493750
rect 212448 493536 212500 493542
rect 212448 493478 212500 493484
rect 212460 491572 212488 493478
rect 213656 491572 213684 493954
rect 213840 493746 213868 500890
rect 213932 500342 213960 502860
rect 214656 500880 214708 500886
rect 214656 500822 214708 500828
rect 213920 500336 213972 500342
rect 213920 500278 213972 500284
rect 214668 493814 214696 500822
rect 215036 500478 215064 502860
rect 216048 500954 216076 502860
rect 216036 500948 216088 500954
rect 216036 500890 216088 500896
rect 217152 500886 217180 502860
rect 217140 500880 217192 500886
rect 217140 500822 217192 500828
rect 215392 500608 215444 500614
rect 215392 500550 215444 500556
rect 215024 500472 215076 500478
rect 215024 500414 215076 500420
rect 215208 500404 215260 500410
rect 215208 500346 215260 500352
rect 214656 493808 214708 493814
rect 214656 493750 214708 493756
rect 213828 493740 213880 493746
rect 213828 493682 213880 493688
rect 215220 493542 215248 500346
rect 215404 494018 215432 500550
rect 218152 500472 218204 500478
rect 218152 500414 218204 500420
rect 216680 499656 216732 499662
rect 216680 499598 216732 499604
rect 215392 494012 215444 494018
rect 215392 493954 215444 493960
rect 215208 493536 215260 493542
rect 215208 493478 215260 493484
rect 216036 493536 216088 493542
rect 216036 493478 216088 493484
rect 214840 493264 214892 493270
rect 214840 493206 214892 493212
rect 214852 491572 214880 493206
rect 216048 491572 216076 493478
rect 216692 493270 216720 499598
rect 217232 493604 217284 493610
rect 217232 493546 217284 493552
rect 216680 493264 216732 493270
rect 216680 493206 216732 493212
rect 217244 491572 217272 493546
rect 218164 493542 218192 500414
rect 218256 500410 218284 502860
rect 219268 500614 219296 502860
rect 219256 500608 219308 500614
rect 219256 500550 219308 500556
rect 219532 500608 219584 500614
rect 219532 500550 219584 500556
rect 218244 500404 218296 500410
rect 218244 500346 218296 500352
rect 218428 494012 218480 494018
rect 218428 493954 218480 493960
rect 218152 493536 218204 493542
rect 218152 493478 218204 493484
rect 218440 491572 218468 493954
rect 219544 493610 219572 500550
rect 220372 499662 220400 502860
rect 221476 500478 221504 502860
rect 222580 500614 222608 502860
rect 223488 500948 223540 500954
rect 223488 500890 223540 500896
rect 222568 500608 222620 500614
rect 222568 500550 222620 500556
rect 221464 500472 221516 500478
rect 221464 500414 221516 500420
rect 220820 500132 220872 500138
rect 220820 500074 220872 500080
rect 220360 499656 220412 499662
rect 220360 499598 220412 499604
rect 220832 494018 220860 500074
rect 220820 494012 220872 494018
rect 220820 493954 220872 493960
rect 220820 493876 220872 493882
rect 220820 493818 220872 493824
rect 219532 493604 219584 493610
rect 219532 493546 219584 493552
rect 219624 493604 219676 493610
rect 219624 493546 219676 493552
rect 219636 491572 219664 493546
rect 220832 491572 220860 493818
rect 222016 493672 222068 493678
rect 222016 493614 222068 493620
rect 222028 491572 222056 493614
rect 223500 493610 223528 500890
rect 223592 500138 223620 502860
rect 224696 500954 224724 502860
rect 224684 500948 224736 500954
rect 224684 500890 224736 500896
rect 225800 500750 225828 502860
rect 224868 500744 224920 500750
rect 224868 500686 224920 500692
rect 225788 500744 225840 500750
rect 225788 500686 225840 500692
rect 224224 500472 224276 500478
rect 224224 500414 224276 500420
rect 223580 500132 223632 500138
rect 223580 500074 223632 500080
rect 223580 499996 223632 500002
rect 223580 499938 223632 499944
rect 223488 493604 223540 493610
rect 223488 493546 223540 493552
rect 223212 492924 223264 492930
rect 223212 492866 223264 492872
rect 223224 491572 223252 492866
rect 223592 492794 223620 499938
rect 224236 493678 224264 500414
rect 224880 493882 224908 500686
rect 226812 500478 226840 502860
rect 226800 500472 226852 500478
rect 226800 500414 226852 500420
rect 224868 493876 224920 493882
rect 224868 493818 224920 493824
rect 224224 493672 224276 493678
rect 224224 493614 224276 493620
rect 225604 493604 225656 493610
rect 225604 493546 225656 493552
rect 223580 492788 223632 492794
rect 223580 492730 223632 492736
rect 224408 492788 224460 492794
rect 224408 492730 224460 492736
rect 224420 491572 224448 492730
rect 225616 491572 225644 493546
rect 226800 493264 226852 493270
rect 226800 493206 226852 493212
rect 226812 491572 226840 493206
rect 227916 492930 227944 502860
rect 229020 500002 229048 502860
rect 230124 500954 230152 502860
rect 230492 502846 231150 502874
rect 229100 500948 229152 500954
rect 229100 500890 229152 500896
rect 230112 500948 230164 500954
rect 230112 500890 230164 500896
rect 229008 499996 229060 500002
rect 229008 499938 229060 499944
rect 229112 499610 229140 500890
rect 230492 500834 230520 502846
rect 229020 499582 229140 499610
rect 230400 500806 230520 500834
rect 227996 493876 228048 493882
rect 227996 493818 228048 493824
rect 227904 492924 227956 492930
rect 227904 492866 227956 492872
rect 228008 491572 228036 493818
rect 229020 493610 229048 499582
rect 229008 493604 229060 493610
rect 229008 493546 229060 493552
rect 229192 493468 229244 493474
rect 229192 493410 229244 493416
rect 229204 491572 229232 493410
rect 230400 493270 230428 500806
rect 232240 500750 232268 502860
rect 233252 502846 233358 502874
rect 233056 500948 233108 500954
rect 233056 500890 233108 500896
rect 230480 500744 230532 500750
rect 230480 500686 230532 500692
rect 232228 500744 232280 500750
rect 232228 500686 232280 500692
rect 230492 493882 230520 500686
rect 232780 493944 232832 493950
rect 232780 493886 232832 493892
rect 230480 493876 230532 493882
rect 230480 493818 230532 493824
rect 231584 493672 231636 493678
rect 231584 493614 231636 493620
rect 230388 493264 230440 493270
rect 230388 493206 230440 493212
rect 230388 493128 230440 493134
rect 230388 493070 230440 493076
rect 230400 491572 230428 493070
rect 231596 491572 231624 493614
rect 232792 491572 232820 493886
rect 233068 493134 233096 500890
rect 233252 500834 233280 502846
rect 234356 500954 234384 502860
rect 234344 500948 234396 500954
rect 234344 500890 234396 500896
rect 233160 500806 233280 500834
rect 233160 493474 233188 500806
rect 235460 499798 235488 502860
rect 236564 500954 236592 502860
rect 237484 502846 237682 502874
rect 237944 502846 238694 502874
rect 238772 502846 239798 502874
rect 240152 502846 240902 502874
rect 241532 502846 241914 502874
rect 235908 500948 235960 500954
rect 235908 500890 235960 500896
rect 236552 500948 236604 500954
rect 236552 500890 236604 500896
rect 234528 499792 234580 499798
rect 234528 499734 234580 499740
rect 235448 499792 235500 499798
rect 235448 499734 235500 499740
rect 234540 493678 234568 499734
rect 235172 494012 235224 494018
rect 235172 493954 235224 493960
rect 234528 493672 234580 493678
rect 234528 493614 234580 493620
rect 233976 493604 234028 493610
rect 233976 493546 234028 493552
rect 233148 493468 233200 493474
rect 233148 493410 233200 493416
rect 233056 493128 233108 493134
rect 233056 493070 233108 493076
rect 233988 491572 234016 493546
rect 235184 491572 235212 493954
rect 235920 493950 235948 500890
rect 237484 500834 237512 502846
rect 237944 501242 237972 502846
rect 237300 500806 237512 500834
rect 237576 501214 237972 501242
rect 235908 493944 235960 493950
rect 235908 493886 235960 493892
rect 236368 493808 236420 493814
rect 236368 493750 236420 493756
rect 236380 491572 236408 493750
rect 237300 493610 237328 500806
rect 237576 494018 237604 501214
rect 237564 494012 237616 494018
rect 237564 493954 237616 493960
rect 237564 493876 237616 493882
rect 237564 493818 237616 493824
rect 237288 493604 237340 493610
rect 237288 493546 237340 493552
rect 237576 491572 237604 493818
rect 238772 493814 238800 502846
rect 240152 493882 240180 502846
rect 241152 494012 241204 494018
rect 241152 493954 241204 493960
rect 240140 493876 240192 493882
rect 240140 493818 240192 493824
rect 238760 493808 238812 493814
rect 238760 493750 238812 493756
rect 239956 493536 240008 493542
rect 239956 493478 240008 493484
rect 238760 493468 238812 493474
rect 238760 493410 238812 493416
rect 238772 491572 238800 493410
rect 239968 491572 239996 493478
rect 241164 491572 241192 493954
rect 241532 493474 241560 502846
rect 243004 500018 243032 502860
rect 242820 499990 243032 500018
rect 243096 502846 244122 502874
rect 244292 502846 245226 502874
rect 245672 502846 246238 502874
rect 247236 502846 247342 502874
rect 242820 493542 242848 499990
rect 243096 494018 243124 502846
rect 243084 494012 243136 494018
rect 243084 493954 243136 493960
rect 242808 493536 242860 493542
rect 242808 493478 242860 493484
rect 241520 493468 241572 493474
rect 241520 493410 241572 493416
rect 243544 493468 243596 493474
rect 243544 493410 243596 493416
rect 242348 493264 242400 493270
rect 242348 493206 242400 493212
rect 242360 491572 242388 493206
rect 243556 491572 243584 493410
rect 244292 493270 244320 502846
rect 245672 493474 245700 502846
rect 247040 499588 247092 499594
rect 247040 499530 247092 499536
rect 245936 494012 245988 494018
rect 245936 493954 245988 493960
rect 245660 493468 245712 493474
rect 245660 493410 245712 493416
rect 244740 493332 244792 493338
rect 244740 493274 244792 493280
rect 244280 493264 244332 493270
rect 244280 493206 244332 493212
rect 244752 491572 244780 493274
rect 245948 491572 245976 493954
rect 247052 491586 247080 499530
rect 247236 493338 247264 502846
rect 248432 494018 248460 502860
rect 249444 499594 249472 502860
rect 249812 502846 250562 502874
rect 251284 502846 251666 502874
rect 249432 499588 249484 499594
rect 249432 499530 249484 499536
rect 248420 494012 248472 494018
rect 248420 493954 248472 493960
rect 249812 493950 249840 502846
rect 251180 500948 251232 500954
rect 251180 500890 251232 500896
rect 249800 493944 249852 493950
rect 249800 493886 249852 493892
rect 248328 493808 248380 493814
rect 248328 493750 248380 493756
rect 249524 493808 249576 493814
rect 249524 493750 249576 493756
rect 247224 493332 247276 493338
rect 247224 493274 247276 493280
rect 247052 491558 247158 491586
rect 248340 491572 248368 493750
rect 249536 491572 249564 493750
rect 250720 492992 250772 492998
rect 250720 492934 250772 492940
rect 250732 491572 250760 492934
rect 251192 492674 251220 500890
rect 251284 493814 251312 502846
rect 252652 499656 252704 499662
rect 252652 499598 252704 499604
rect 251272 493808 251324 493814
rect 251272 493750 251324 493756
rect 251192 492646 251496 492674
rect 251468 491586 251496 492646
rect 252664 491586 252692 499598
rect 252756 492998 252784 502860
rect 253768 500954 253796 502860
rect 253756 500948 253808 500954
rect 253756 500890 253808 500896
rect 253940 500948 253992 500954
rect 253940 500890 253992 500896
rect 252744 492992 252796 492998
rect 252744 492934 252796 492940
rect 253952 491586 253980 500890
rect 254872 499662 254900 502860
rect 255976 500954 256004 502860
rect 255964 500948 256016 500954
rect 255964 500890 256016 500896
rect 256988 500342 257016 502860
rect 257528 500540 257580 500546
rect 257528 500482 257580 500488
rect 255320 500336 255372 500342
rect 255320 500278 255372 500284
rect 256976 500336 257028 500342
rect 256976 500278 257028 500284
rect 254860 499656 254912 499662
rect 254860 499598 254912 499604
rect 255332 491586 255360 500278
rect 256792 499588 256844 499594
rect 256792 499530 256844 499536
rect 256804 491586 256832 499530
rect 251468 491558 251942 491586
rect 252664 491558 253138 491586
rect 253952 491558 254334 491586
rect 255332 491558 255530 491586
rect 256726 491558 256832 491586
rect 257540 491586 257568 500482
rect 258092 499594 258120 502860
rect 258264 500676 258316 500682
rect 258264 500618 258316 500624
rect 258080 499588 258132 499594
rect 258080 499530 258132 499536
rect 258276 494018 258304 500618
rect 259196 500546 259224 502860
rect 260300 500682 260328 502860
rect 260288 500676 260340 500682
rect 260288 500618 260340 500624
rect 260840 500676 260892 500682
rect 260840 500618 260892 500624
rect 259184 500540 259236 500546
rect 259184 500482 259236 500488
rect 259460 500268 259512 500274
rect 259460 500210 259512 500216
rect 259472 494018 259500 500210
rect 258264 494012 258316 494018
rect 258264 493954 258316 493960
rect 259092 494012 259144 494018
rect 259092 493954 259144 493960
rect 259460 494012 259512 494018
rect 259460 493954 259512 493960
rect 260288 494012 260340 494018
rect 260288 493954 260340 493960
rect 257540 491558 257922 491586
rect 259104 491572 259132 493954
rect 260300 491572 260328 493954
rect 260852 493626 260880 500618
rect 261312 500274 261340 502860
rect 262220 500948 262272 500954
rect 262220 500890 262272 500896
rect 261300 500268 261352 500274
rect 261300 500210 261352 500216
rect 262232 493762 262260 500890
rect 262416 500682 262444 502860
rect 263520 500954 263548 502860
rect 264532 500954 264560 502860
rect 264992 502846 265650 502874
rect 266464 502846 266754 502874
rect 263508 500948 263560 500954
rect 263508 500890 263560 500896
rect 263600 500948 263652 500954
rect 263600 500890 263652 500896
rect 264520 500948 264572 500954
rect 264520 500890 264572 500896
rect 262404 500676 262456 500682
rect 262404 500618 262456 500624
rect 262232 493734 262444 493762
rect 260852 493598 261156 493626
rect 261128 491586 261156 493598
rect 262416 491586 262444 493734
rect 263612 491586 263640 500890
rect 264992 491586 265020 502846
rect 266464 500834 266492 502846
rect 266280 500806 266492 500834
rect 267740 500812 267792 500818
rect 261128 491558 261510 491586
rect 262416 491558 262706 491586
rect 263612 491558 263902 491586
rect 264992 491558 265098 491586
rect 266280 491572 266308 500806
rect 267740 500754 267792 500760
rect 266464 499594 266584 499610
rect 266464 499588 266596 499594
rect 266464 499582 266544 499588
rect 266464 493134 266492 499582
rect 266544 499530 266596 499536
rect 266452 493128 266504 493134
rect 266452 493070 266504 493076
rect 267464 493128 267516 493134
rect 267464 493070 267516 493076
rect 267476 491572 267504 493070
rect 267752 492402 267780 500754
rect 267844 499594 267872 502860
rect 268856 500818 268884 502860
rect 269960 500954 269988 502860
rect 270512 502846 271078 502874
rect 271892 502846 272090 502874
rect 269120 500948 269172 500954
rect 269120 500890 269172 500896
rect 269948 500948 270000 500954
rect 269948 500890 270000 500896
rect 268844 500812 268896 500818
rect 268844 500754 268896 500760
rect 267832 499588 267884 499594
rect 267832 499530 267884 499536
rect 269132 494034 269160 500890
rect 270512 494306 270540 502846
rect 270512 494278 270724 494306
rect 269132 494006 269620 494034
rect 267752 492374 268240 492402
rect 268212 491586 268240 492374
rect 269592 491586 269620 494006
rect 270696 491586 270724 494278
rect 271892 491586 271920 502846
rect 273180 500954 273208 502860
rect 271972 500948 272024 500954
rect 271972 500890 272024 500896
rect 273168 500948 273220 500954
rect 273168 500890 273220 500896
rect 271984 492862 272012 500890
rect 274560 493218 274588 502982
rect 274744 502846 275402 502874
rect 276032 502846 276414 502874
rect 277412 502846 277518 502874
rect 274560 493190 274680 493218
rect 271972 492856 272024 492862
rect 271972 492798 272024 492804
rect 273444 492856 273496 492862
rect 273444 492798 273496 492804
rect 268212 491558 268686 491586
rect 269592 491558 269882 491586
rect 270696 491558 271078 491586
rect 271892 491558 272274 491586
rect 273456 491572 273484 492798
rect 274652 491572 274680 493190
rect 274744 491450 274772 502846
rect 276032 491450 276060 502846
rect 277412 491586 277440 502846
rect 278608 500954 278636 502860
rect 277584 500948 277636 500954
rect 277584 500890 277636 500896
rect 278596 500948 278648 500954
rect 278596 500890 278648 500896
rect 277596 493202 277624 500890
rect 280160 498840 280212 498846
rect 280160 498782 280212 498788
rect 277584 493196 277636 493202
rect 277584 493138 277636 493144
rect 279424 493196 279476 493202
rect 279424 493138 279476 493144
rect 277412 491558 278254 491586
rect 279436 491572 279464 493138
rect 274744 491422 275862 491450
rect 276032 491422 277058 491450
rect 280172 471345 280200 498782
rect 280158 471336 280214 471345
rect 280158 471271 280214 471280
rect 281552 430545 281580 515879
rect 281538 430536 281594 430545
rect 281538 430471 281594 430480
rect 282182 430536 282238 430545
rect 282182 430471 282238 430480
rect 282196 421598 282224 430471
rect 281632 421592 281684 421598
rect 281632 421534 281684 421540
rect 282184 421592 282236 421598
rect 282184 421534 282236 421540
rect 281644 421297 281672 421534
rect 281630 421288 281686 421297
rect 281630 421223 281686 421232
rect 282184 377256 282236 377262
rect 282184 377198 282236 377204
rect 282196 360194 282224 377198
rect 282184 360188 282236 360194
rect 282184 360130 282236 360136
rect 245456 358278 245608 358306
rect 188048 358142 188384 358170
rect 189244 358142 189580 358170
rect 188356 354754 188384 358142
rect 189552 355502 189580 358142
rect 190380 358142 190440 358170
rect 191636 358142 191788 358170
rect 192924 358142 193168 358170
rect 194120 358142 194456 358170
rect 195316 358142 195652 358170
rect 196512 358142 196848 358170
rect 197800 358142 198136 358170
rect 198996 358142 199332 358170
rect 200192 358142 200528 358170
rect 189540 355496 189592 355502
rect 189540 355438 189592 355444
rect 190380 355366 190408 358142
rect 190368 355360 190420 355366
rect 190368 355302 190420 355308
rect 191760 354890 191788 358142
rect 191932 357536 191984 357542
rect 191932 357478 191984 357484
rect 191748 354884 191800 354890
rect 191748 354826 191800 354832
rect 188344 354748 188396 354754
rect 188344 354690 188396 354696
rect 189446 351792 189502 351801
rect 189446 351727 189502 351736
rect 191194 351792 191250 351801
rect 191194 351727 191250 351736
rect 187712 348894 188094 348922
rect 189460 348786 189488 351727
rect 189906 351656 189962 351665
rect 189906 351591 189962 351600
rect 189920 348922 189948 351591
rect 191208 348922 191236 351727
rect 191944 349058 191972 357478
rect 193140 355978 193168 358142
rect 194428 356046 194456 358142
rect 194416 356040 194468 356046
rect 194416 355982 194468 355988
rect 193128 355972 193180 355978
rect 193128 355914 193180 355920
rect 194968 354884 195020 354890
rect 194968 354826 195020 354832
rect 193220 354748 193272 354754
rect 193220 354690 193272 354696
rect 193232 351218 193260 354690
rect 194140 351892 194192 351898
rect 194140 351834 194192 351840
rect 193220 351212 193272 351218
rect 193220 351154 193272 351160
rect 193220 351076 193272 351082
rect 193220 351018 193272 351024
rect 191944 349030 192156 349058
rect 192128 348922 192156 349030
rect 193232 348922 193260 351018
rect 194152 348922 194180 351834
rect 194980 351490 195008 354826
rect 195624 354754 195652 358142
rect 196348 355496 196400 355502
rect 196348 355438 196400 355444
rect 195612 354748 195664 354754
rect 195612 354690 195664 354696
rect 194968 351484 195020 351490
rect 194968 351426 195020 351432
rect 195244 351212 195296 351218
rect 195244 351154 195296 351160
rect 195256 348922 195284 351154
rect 196360 348922 196388 355438
rect 196820 354890 196848 358142
rect 198108 355706 198136 358142
rect 198924 356040 198976 356046
rect 198924 355982 198976 355988
rect 198096 355700 198148 355706
rect 198096 355642 198148 355648
rect 197268 355360 197320 355366
rect 197268 355302 197320 355308
rect 196808 354884 196860 354890
rect 196808 354826 196860 354832
rect 197280 350554 197308 355302
rect 198936 351898 198964 355982
rect 199304 355774 199332 358142
rect 199660 355972 199712 355978
rect 199660 355914 199712 355920
rect 199292 355768 199344 355774
rect 199292 355710 199344 355716
rect 198924 351892 198976 351898
rect 198924 351834 198976 351840
rect 198740 351484 198792 351490
rect 198740 351426 198792 351432
rect 197280 350526 197400 350554
rect 197372 348922 197400 350526
rect 198752 348922 198780 351426
rect 199672 348922 199700 355914
rect 200500 355570 200528 358142
rect 201420 358142 201480 358170
rect 202676 358142 202828 358170
rect 203872 358142 204208 358170
rect 205068 358142 205404 358170
rect 206356 358142 206692 358170
rect 207552 358142 207888 358170
rect 208748 358142 209084 358170
rect 210036 358142 210372 358170
rect 211232 358142 211568 358170
rect 201420 356046 201448 358142
rect 201408 356040 201460 356046
rect 201408 355982 201460 355988
rect 200488 355564 200540 355570
rect 200488 355506 200540 355512
rect 202800 355230 202828 358142
rect 204180 355842 204208 358142
rect 204168 355836 204220 355842
rect 204168 355778 204220 355784
rect 204996 355768 205048 355774
rect 204996 355710 205048 355716
rect 203892 355700 203944 355706
rect 203892 355642 203944 355648
rect 202788 355224 202840 355230
rect 202788 355166 202840 355172
rect 201500 354884 201552 354890
rect 201500 354826 201552 354832
rect 201408 354748 201460 354754
rect 201408 354690 201460 354696
rect 200580 351892 200632 351898
rect 200580 351834 200632 351840
rect 200592 348922 200620 351834
rect 201420 350554 201448 354690
rect 201512 350946 201540 354826
rect 201500 350940 201552 350946
rect 201500 350882 201552 350888
rect 202880 350940 202932 350946
rect 202880 350882 202932 350888
rect 201420 350526 201632 350554
rect 201604 348922 201632 350526
rect 202892 348922 202920 350882
rect 203904 348922 203932 355642
rect 205008 348922 205036 355710
rect 205376 354754 205404 358142
rect 206100 355564 206152 355570
rect 206100 355506 206152 355512
rect 205364 354748 205416 354754
rect 205364 354690 205416 354696
rect 206112 348922 206140 355506
rect 206664 354822 206692 358142
rect 206928 356040 206980 356046
rect 206928 355982 206980 355988
rect 206652 354816 206704 354822
rect 206652 354758 206704 354764
rect 206940 350554 206968 355982
rect 207860 355434 207888 358142
rect 207848 355428 207900 355434
rect 207848 355370 207900 355376
rect 209056 355366 209084 358142
rect 210344 356046 210372 358142
rect 210332 356040 210384 356046
rect 210332 355982 210384 355988
rect 211540 355910 211568 358142
rect 212368 358142 212428 358170
rect 213624 358142 213868 358170
rect 214912 358142 215248 358170
rect 216108 358142 216444 358170
rect 217304 358142 217640 358170
rect 218592 358142 218928 358170
rect 219788 358142 220124 358170
rect 220984 358142 221320 358170
rect 211528 355904 211580 355910
rect 211528 355846 211580 355852
rect 209228 355836 209280 355842
rect 209228 355778 209280 355784
rect 209044 355360 209096 355366
rect 209044 355302 209096 355308
rect 208308 355224 208360 355230
rect 208308 355166 208360 355172
rect 208320 350554 208348 355166
rect 206940 350526 207152 350554
rect 208320 350526 208440 350554
rect 207124 348922 207152 350526
rect 208412 348922 208440 350526
rect 209240 348922 209268 355778
rect 212368 355026 212396 358142
rect 213840 355978 213868 358142
rect 215220 356046 215248 358142
rect 214748 356040 214800 356046
rect 214748 355982 214800 355988
rect 215208 356040 215260 356046
rect 215208 355982 215260 355988
rect 213828 355972 213880 355978
rect 213828 355914 213880 355920
rect 212632 355428 212684 355434
rect 212632 355370 212684 355376
rect 212356 355020 212408 355026
rect 212356 354962 212408 354968
rect 211436 354816 211488 354822
rect 211436 354758 211488 354764
rect 210332 354748 210384 354754
rect 210332 354690 210384 354696
rect 210344 348922 210372 354690
rect 211448 348922 211476 354758
rect 212644 348922 212672 355370
rect 214012 355360 214064 355366
rect 214012 355302 214064 355308
rect 189920 348894 190210 348922
rect 191208 348894 191314 348922
rect 192128 348894 192418 348922
rect 193232 348894 193430 348922
rect 194152 348894 194534 348922
rect 195256 348894 195638 348922
rect 196360 348894 196650 348922
rect 197372 348894 197754 348922
rect 198752 348894 198858 348922
rect 199672 348894 199962 348922
rect 200592 348894 200974 348922
rect 201604 348894 202078 348922
rect 202892 348894 203182 348922
rect 203904 348894 204194 348922
rect 205008 348894 205298 348922
rect 206112 348894 206402 348922
rect 207124 348894 207506 348922
rect 208412 348894 208518 348922
rect 209240 348894 209622 348922
rect 210344 348894 210726 348922
rect 211448 348894 211738 348922
rect 212644 348894 212842 348922
rect 214024 348786 214052 355302
rect 214760 348922 214788 355982
rect 215668 355904 215720 355910
rect 215668 355846 215720 355852
rect 215680 348922 215708 355846
rect 216416 354754 216444 358142
rect 217612 355638 217640 358142
rect 218060 355972 218112 355978
rect 218060 355914 218112 355920
rect 217600 355632 217652 355638
rect 217600 355574 217652 355580
rect 216772 355020 216824 355026
rect 216772 354962 216824 354968
rect 216404 354748 216456 354754
rect 216404 354690 216456 354696
rect 216784 348922 216812 354962
rect 218072 348922 218100 355914
rect 218900 355434 218928 358142
rect 218980 356040 219032 356046
rect 218980 355982 219032 355988
rect 218888 355428 218940 355434
rect 218888 355370 218940 355376
rect 218992 348922 219020 355982
rect 220096 355298 220124 358142
rect 221292 356046 221320 358142
rect 222120 358142 222180 358170
rect 223408 358142 223468 358170
rect 224664 358142 224908 358170
rect 225860 358142 226196 358170
rect 227148 358142 227484 358170
rect 228344 358142 228680 358170
rect 229540 358142 229876 358170
rect 230736 358142 231072 358170
rect 232024 358142 232360 358170
rect 221280 356040 221332 356046
rect 221280 355982 221332 355988
rect 222120 355842 222148 358142
rect 222844 356040 222896 356046
rect 222844 355982 222896 355988
rect 222108 355836 222160 355842
rect 222108 355778 222160 355784
rect 221188 355632 221240 355638
rect 221188 355574 221240 355580
rect 220084 355292 220136 355298
rect 220084 355234 220136 355240
rect 220084 354748 220136 354754
rect 220084 354690 220136 354696
rect 220096 348922 220124 354690
rect 221200 348922 221228 355574
rect 222384 355428 222436 355434
rect 222384 355370 222436 355376
rect 222396 348922 222424 355370
rect 222856 350810 222884 355982
rect 223408 354890 223436 358142
rect 224880 355910 224908 358142
rect 226168 356046 226196 358142
rect 227456 356046 227484 358142
rect 226156 356040 226208 356046
rect 226156 355982 226208 355988
rect 226984 356040 227036 356046
rect 226984 355982 227036 355988
rect 227444 356040 227496 356046
rect 227444 355982 227496 355988
rect 228180 356040 228232 356046
rect 228180 355982 228232 355988
rect 224868 355904 224920 355910
rect 224868 355846 224920 355852
rect 225420 355836 225472 355842
rect 225420 355778 225472 355784
rect 223672 355292 223724 355298
rect 223672 355234 223724 355240
rect 223396 354884 223448 354890
rect 223396 354826 223448 354832
rect 222844 350804 222896 350810
rect 222844 350746 222896 350752
rect 214760 348894 215050 348922
rect 215680 348894 216062 348922
rect 216784 348894 217166 348922
rect 218072 348894 218270 348922
rect 218992 348894 219282 348922
rect 220096 348894 220386 348922
rect 221200 348894 221490 348922
rect 222396 348894 222594 348922
rect 223684 348786 223712 355234
rect 224316 350804 224368 350810
rect 224316 350746 224368 350752
rect 224328 348922 224356 350746
rect 225432 348922 225460 355778
rect 226524 354884 226576 354890
rect 226524 354826 226576 354832
rect 226536 348922 226564 354826
rect 226996 350946 227024 355982
rect 227720 355904 227772 355910
rect 227720 355846 227772 355852
rect 226984 350940 227036 350946
rect 226984 350882 227036 350888
rect 227732 348922 227760 355846
rect 228192 351218 228220 355982
rect 228652 354754 228680 358142
rect 229848 356046 229876 358142
rect 229836 356040 229888 356046
rect 229836 355982 229888 355988
rect 230480 356040 230532 356046
rect 230480 355982 230532 355988
rect 228640 354748 228692 354754
rect 228640 354690 228692 354696
rect 230388 354748 230440 354754
rect 230388 354690 230440 354696
rect 228180 351212 228232 351218
rect 228180 351154 228232 351160
rect 229836 351212 229888 351218
rect 229836 351154 229888 351160
rect 228732 350940 228784 350946
rect 228732 350882 228784 350888
rect 228744 348922 228772 350882
rect 229848 348922 229876 351154
rect 230400 350554 230428 354690
rect 230492 350946 230520 355982
rect 231044 355434 231072 358142
rect 232332 355978 232360 358142
rect 233160 358142 233220 358170
rect 234416 358142 234568 358170
rect 235704 358142 235856 358170
rect 236900 358142 237236 358170
rect 238096 358142 238432 358170
rect 239292 358142 239628 358170
rect 240580 358142 240916 358170
rect 241776 358142 242112 358170
rect 242972 358142 243308 358170
rect 233160 356046 233188 358142
rect 234540 356046 234568 358142
rect 233148 356040 233200 356046
rect 233148 355982 233200 355988
rect 233700 356040 233752 356046
rect 233700 355982 233752 355988
rect 234528 356040 234580 356046
rect 234528 355982 234580 355988
rect 232320 355972 232372 355978
rect 232320 355914 232372 355920
rect 231032 355428 231084 355434
rect 231032 355370 231084 355376
rect 233148 355428 233200 355434
rect 233148 355370 233200 355376
rect 230480 350940 230532 350946
rect 230480 350882 230532 350888
rect 231860 350940 231912 350946
rect 231860 350882 231912 350888
rect 230400 350526 230704 350554
rect 230676 348922 230704 350526
rect 231872 348922 231900 350882
rect 233160 350554 233188 355370
rect 233712 350946 233740 355982
rect 235828 355978 235856 358142
rect 237208 356046 237236 358142
rect 235908 356040 235960 356046
rect 235908 355982 235960 355988
rect 237196 356040 237248 356046
rect 237196 355982 237248 355988
rect 238300 356040 238352 356046
rect 238300 355982 238352 355988
rect 234068 355972 234120 355978
rect 234068 355914 234120 355920
rect 235816 355972 235868 355978
rect 235816 355914 235868 355920
rect 233700 350940 233752 350946
rect 233700 350882 233752 350888
rect 233160 350526 233280 350554
rect 233252 348922 233280 350526
rect 234080 348922 234108 355914
rect 235172 350940 235224 350946
rect 235172 350882 235224 350888
rect 235184 348922 235212 350882
rect 235920 350554 235948 355982
rect 237288 355972 237340 355978
rect 237288 355914 237340 355920
rect 237300 350554 237328 355914
rect 235920 350526 236224 350554
rect 237300 350526 237420 350554
rect 236196 348922 236224 350526
rect 237392 348922 237420 350526
rect 238312 348922 238340 355982
rect 238404 354822 238432 358142
rect 239600 356046 239628 358142
rect 239588 356040 239640 356046
rect 239588 355982 239640 355988
rect 240508 356040 240560 356046
rect 240508 355982 240560 355988
rect 238392 354816 238444 354822
rect 238392 354758 238444 354764
rect 239404 354816 239456 354822
rect 239404 354758 239456 354764
rect 239416 348922 239444 354758
rect 240520 348922 240548 355982
rect 240888 355706 240916 358142
rect 242084 355842 242112 358142
rect 242072 355836 242124 355842
rect 242072 355778 242124 355784
rect 242808 355836 242860 355842
rect 242808 355778 242860 355784
rect 240876 355700 240928 355706
rect 240876 355642 240928 355648
rect 241704 355700 241756 355706
rect 241704 355642 241756 355648
rect 241716 348922 241744 355642
rect 242820 354634 242848 355778
rect 243280 355366 243308 358142
rect 244108 358142 244168 358170
rect 244108 355366 244136 358142
rect 245580 356028 245608 358278
rect 246652 358142 246896 358170
rect 247848 358142 248092 358170
rect 246868 356028 246896 358142
rect 245580 356000 245884 356028
rect 246868 356000 247080 356028
rect 243268 355360 243320 355366
rect 243268 355302 243320 355308
rect 243820 355360 243872 355366
rect 243820 355302 243872 355308
rect 244096 355360 244148 355366
rect 244096 355302 244148 355308
rect 244924 355360 244976 355366
rect 244924 355302 244976 355308
rect 242820 354606 242940 354634
rect 242912 348922 242940 354606
rect 243832 348922 243860 355302
rect 244936 348922 244964 355302
rect 245856 348922 245884 356000
rect 247052 348922 247080 356000
rect 248064 354822 248092 358142
rect 249122 357898 249150 358156
rect 250272 358142 250332 358170
rect 251192 358142 251528 358170
rect 252572 358142 252724 358170
rect 249122 357870 249196 357898
rect 248052 354816 248104 354822
rect 248052 354758 248104 354764
rect 248512 354816 248564 354822
rect 248512 354758 248564 354764
rect 224328 348894 224710 348922
rect 225432 348894 225814 348922
rect 226536 348894 226826 348922
rect 227732 348894 227930 348922
rect 228744 348894 229034 348922
rect 229848 348894 230138 348922
rect 230676 348894 231150 348922
rect 231872 348894 232254 348922
rect 233252 348894 233358 348922
rect 234080 348894 234370 348922
rect 235184 348894 235474 348922
rect 236196 348894 236578 348922
rect 237392 348894 237682 348922
rect 238312 348894 238694 348922
rect 239416 348894 239798 348922
rect 240520 348894 240902 348922
rect 241716 348894 241914 348922
rect 242912 348894 243018 348922
rect 243832 348894 244122 348922
rect 244936 348894 245226 348922
rect 245856 348894 246238 348922
rect 247052 348894 247342 348922
rect 248524 348786 248552 354758
rect 249168 348922 249196 357870
rect 250272 348922 250300 358142
rect 249168 348894 249458 348922
rect 250272 348894 250562 348922
rect 186332 348758 186990 348786
rect 189106 348758 189488 348786
rect 213946 348758 214052 348786
rect 223606 348758 223712 348786
rect 248446 348758 248552 348786
rect 251192 348786 251220 358142
rect 252572 348922 252600 358142
rect 253998 357898 254026 358156
rect 254872 358142 255208 358170
rect 256068 358142 256404 358170
rect 257356 358142 257692 358170
rect 258552 358142 258888 358170
rect 259564 358142 260084 358170
rect 261036 358142 261280 358170
rect 262232 358142 262568 358170
rect 263612 358142 263764 358170
rect 264624 358142 264960 358170
rect 265912 358142 266248 358170
rect 267108 358142 267444 358170
rect 268304 358142 268640 358170
rect 269500 358142 269836 358170
rect 270512 358142 271124 358170
rect 271892 358142 272320 358170
rect 273272 358142 273516 358170
rect 274744 358142 274804 358170
rect 275664 358142 276000 358170
rect 276216 358142 277196 358170
rect 277412 358142 278392 358170
rect 278792 358142 279680 358170
rect 280172 358142 280876 358170
rect 281736 358142 282072 358170
rect 253998 357870 254072 357898
rect 254044 355994 254072 357870
rect 253860 355966 254072 355994
rect 252572 348894 252770 348922
rect 253860 348786 253888 355966
rect 254872 355162 254900 358142
rect 256068 355706 256096 358142
rect 255320 355700 255372 355706
rect 255320 355642 255372 355648
rect 256056 355700 256108 355706
rect 256056 355642 256108 355648
rect 254124 355156 254176 355162
rect 254124 355098 254176 355104
rect 254860 355156 254912 355162
rect 254860 355098 254912 355104
rect 251192 348758 251666 348786
rect 253782 348758 253888 348786
rect 254136 348786 254164 355098
rect 255332 348786 255360 355642
rect 257356 355434 257384 358142
rect 258552 356046 258580 358142
rect 258080 356040 258132 356046
rect 258080 355982 258132 355988
rect 258540 356040 258592 356046
rect 259564 355994 259592 358142
rect 258540 355982 258592 355988
rect 256700 355428 256752 355434
rect 256700 355370 256752 355376
rect 257344 355428 257396 355434
rect 257344 355370 257396 355376
rect 256712 348922 256740 355370
rect 258092 349058 258120 355982
rect 259380 355966 259592 355994
rect 258092 349030 258212 349058
rect 256712 348894 257002 348922
rect 258184 348786 258212 349030
rect 259380 348786 259408 355966
rect 261036 354754 261064 358142
rect 262232 356046 262260 358142
rect 263612 356046 263640 358142
rect 261576 356040 261628 356046
rect 261576 355982 261628 355988
rect 262220 356040 262272 356046
rect 262220 355982 262272 355988
rect 262680 356040 262732 356046
rect 262680 355982 262732 355988
rect 263600 356040 263652 356046
rect 263600 355982 263652 355988
rect 260564 354748 260616 354754
rect 260564 354690 260616 354696
rect 261024 354748 261076 354754
rect 261024 354690 261076 354696
rect 260576 348786 260604 354690
rect 261588 348786 261616 355982
rect 262692 348786 262720 355982
rect 264624 355570 264652 358142
rect 263416 355564 263468 355570
rect 263416 355506 263468 355512
rect 264612 355564 264664 355570
rect 264612 355506 264664 355512
rect 263428 348922 263456 355506
rect 265912 355298 265940 358142
rect 267108 355434 267136 358142
rect 266084 355428 266136 355434
rect 266084 355370 266136 355376
rect 267096 355428 267148 355434
rect 267096 355370 267148 355376
rect 264888 355292 264940 355298
rect 264888 355234 264940 355240
rect 265900 355292 265952 355298
rect 265900 355234 265952 355240
rect 263428 348894 263534 348922
rect 264900 348786 264928 355234
rect 266096 348786 266124 355370
rect 268200 355156 268252 355162
rect 268200 355098 268252 355104
rect 267096 354748 267148 354754
rect 267096 354690 267148 354696
rect 267108 348786 267136 354690
rect 268212 348786 268240 355098
rect 268304 354754 268332 358142
rect 269500 355162 269528 358142
rect 269488 355156 269540 355162
rect 269488 355098 269540 355104
rect 268292 354748 268344 354754
rect 268292 354690 268344 354696
rect 270512 351490 270540 358142
rect 271328 351552 271380 351558
rect 271328 351494 271380 351500
rect 269028 351484 269080 351490
rect 269028 351426 269080 351432
rect 270500 351484 270552 351490
rect 270500 351426 270552 351432
rect 269040 348786 269068 351426
rect 270224 351416 270276 351422
rect 270224 351358 270276 351364
rect 270236 348786 270264 351358
rect 271340 348786 271368 351494
rect 271892 351422 271920 358142
rect 273272 351558 273300 358142
rect 274640 356448 274692 356454
rect 274640 356390 274692 356396
rect 273260 351552 273312 351558
rect 273260 351494 273312 351500
rect 274652 351490 274680 356390
rect 273076 351484 273128 351490
rect 273076 351426 273128 351432
rect 274640 351484 274692 351490
rect 274640 351426 274692 351432
rect 271880 351416 271932 351422
rect 271880 351358 271932 351364
rect 272432 350940 272484 350946
rect 272432 350882 272484 350888
rect 272444 348786 272472 350882
rect 273088 348922 273116 351426
rect 274548 351416 274600 351422
rect 274548 351358 274600 351364
rect 273088 348894 273194 348922
rect 274560 348786 274588 351358
rect 274744 350946 274772 358142
rect 275664 356454 275692 358142
rect 275652 356448 275704 356454
rect 275652 356390 275704 356396
rect 275744 351892 275796 351898
rect 275744 351834 275796 351840
rect 274732 350940 274784 350946
rect 274732 350882 274784 350888
rect 275756 348786 275784 351834
rect 276216 351422 276244 358142
rect 277412 351898 277440 358142
rect 277400 351892 277452 351898
rect 277400 351834 277452 351840
rect 278688 351484 278740 351490
rect 278688 351426 278740 351432
rect 276204 351416 276256 351422
rect 276204 351358 276256 351364
rect 277768 351416 277820 351422
rect 277768 351358 277820 351364
rect 276664 351348 276716 351354
rect 276664 351290 276716 351296
rect 276676 348786 276704 351290
rect 277780 348786 277808 351358
rect 278700 348786 278728 351426
rect 278792 351354 278820 358142
rect 280172 351422 280200 358142
rect 281736 355842 281764 358142
rect 281448 355836 281500 355842
rect 281448 355778 281500 355784
rect 281724 355836 281776 355842
rect 281724 355778 281776 355784
rect 281460 351490 281488 355778
rect 281448 351484 281500 351490
rect 281448 351426 281500 351432
rect 280160 351416 280212 351422
rect 280160 351358 280212 351364
rect 278780 351348 278832 351354
rect 278780 351290 278832 351296
rect 254136 348758 254886 348786
rect 255332 348758 255990 348786
rect 258106 348758 258212 348786
rect 259210 348758 259408 348786
rect 260314 348758 260604 348786
rect 261326 348758 261616 348786
rect 262430 348758 262720 348786
rect 264546 348758 264928 348786
rect 265650 348758 266124 348786
rect 266754 348758 267136 348786
rect 267858 348758 268240 348786
rect 268870 348758 269068 348786
rect 269974 348758 270264 348786
rect 271078 348758 271368 348786
rect 272090 348758 272472 348786
rect 274298 348758 274588 348786
rect 275402 348758 275784 348786
rect 276414 348758 276704 348786
rect 277518 348758 277808 348786
rect 278622 348758 278728 348786
rect 282196 336025 282224 360130
rect 282182 336016 282238 336025
rect 282182 335951 282238 335960
rect 21364 323536 21416 323542
rect 21364 323478 21416 323484
rect 22192 323536 22244 323542
rect 22192 323478 22244 323484
rect 22008 320204 22060 320210
rect 22008 320146 22060 320152
rect 20628 318776 20680 318782
rect 20628 318718 20680 318724
rect 20640 315588 20668 318718
rect 22020 315602 22048 320146
rect 22112 319462 22140 322932
rect 22204 321638 22232 323478
rect 22192 321632 22244 321638
rect 22192 321574 22244 321580
rect 22100 319456 22152 319462
rect 22100 319398 22152 319404
rect 23124 318782 23152 322932
rect 23296 320476 23348 320482
rect 23296 320418 23348 320424
rect 23112 318776 23164 318782
rect 23112 318718 23164 318724
rect 23308 315602 23336 320418
rect 24228 320210 24256 322932
rect 24768 320884 24820 320890
rect 24768 320826 24820 320832
rect 24216 320204 24268 320210
rect 24216 320146 24268 320152
rect 24780 315602 24808 320826
rect 25332 320482 25360 322932
rect 26344 320890 26372 322932
rect 26884 321564 26936 321570
rect 26884 321506 26936 321512
rect 26332 320884 26384 320890
rect 26332 320826 26384 320832
rect 25320 320476 25372 320482
rect 25320 320418 25372 320424
rect 25320 320340 25372 320346
rect 25320 320282 25372 320288
rect 21758 315574 22048 315602
rect 22954 315574 23336 315602
rect 24596 315574 24808 315602
rect 25332 315588 25360 320282
rect 26516 320204 26568 320210
rect 26516 320146 26568 320152
rect 26528 315588 26556 320146
rect 24596 315466 24624 315574
rect 24150 315438 24624 315466
rect 26896 315382 26924 321506
rect 27448 320346 27476 322932
rect 27436 320340 27488 320346
rect 27436 320282 27488 320288
rect 27712 320272 27764 320278
rect 27712 320214 27764 320220
rect 27724 315588 27752 320214
rect 28552 320210 28580 322932
rect 29656 320278 29684 322932
rect 29644 320272 29696 320278
rect 29644 320214 29696 320220
rect 30288 320272 30340 320278
rect 30288 320214 30340 320220
rect 28540 320204 28592 320210
rect 28540 320146 28592 320152
rect 28908 320204 28960 320210
rect 28908 320146 28960 320152
rect 28920 315588 28948 320146
rect 30300 315602 30328 320214
rect 30668 320210 30696 322932
rect 31772 320278 31800 322932
rect 31760 320272 31812 320278
rect 31760 320214 31812 320220
rect 32876 320210 32904 322932
rect 33692 320272 33744 320278
rect 33692 320214 33744 320220
rect 30656 320204 30708 320210
rect 30656 320146 30708 320152
rect 31668 320204 31720 320210
rect 31668 320146 31720 320152
rect 32864 320204 32916 320210
rect 32864 320146 32916 320152
rect 33048 320204 33100 320210
rect 33048 320146 33100 320152
rect 31680 315602 31708 320146
rect 30130 315574 30328 315602
rect 31326 315574 31708 315602
rect 33060 315466 33088 320146
rect 33704 315588 33732 320214
rect 33888 320210 33916 322932
rect 34888 320884 34940 320890
rect 34888 320826 34940 320832
rect 33876 320204 33928 320210
rect 33876 320146 33928 320152
rect 34900 315588 34928 320826
rect 34992 320278 35020 322932
rect 35912 322918 36110 322946
rect 35808 320884 35860 320890
rect 35912 320872 35940 322918
rect 35860 320844 35940 320872
rect 35808 320826 35860 320832
rect 34980 320272 35032 320278
rect 34980 320214 35032 320220
rect 37200 320210 37228 322932
rect 38212 320210 38240 322932
rect 39316 320210 39344 322932
rect 40052 322918 40434 322946
rect 40052 320226 40080 322918
rect 41432 320226 41460 322932
rect 35900 320204 35952 320210
rect 35900 320146 35952 320152
rect 37188 320204 37240 320210
rect 37188 320146 37240 320152
rect 37280 320204 37332 320210
rect 37280 320146 37332 320152
rect 38200 320204 38252 320210
rect 38200 320146 38252 320152
rect 38568 320204 38620 320210
rect 38568 320146 38620 320152
rect 39304 320204 39356 320210
rect 39304 320146 39356 320152
rect 39960 320198 40080 320226
rect 41340 320198 41460 320226
rect 42536 320210 42564 322932
rect 43640 320210 43668 322932
rect 44192 322918 44758 322946
rect 45664 322918 45770 322946
rect 46584 322918 46874 322946
rect 42524 320204 42576 320210
rect 35912 315602 35940 320146
rect 35912 315574 36110 315602
rect 37292 315588 37320 320146
rect 38580 315602 38608 320146
rect 39960 315602 39988 320198
rect 38502 315574 38608 315602
rect 39698 315574 39988 315602
rect 41340 315466 41368 320198
rect 42524 320146 42576 320152
rect 42800 320204 42852 320210
rect 42800 320146 42852 320152
rect 43628 320204 43680 320210
rect 43628 320146 43680 320152
rect 41420 320136 41472 320142
rect 41420 320078 41472 320084
rect 32522 315438 33088 315466
rect 40894 315438 41368 315466
rect 41432 315466 41460 320078
rect 42812 315602 42840 320146
rect 44192 315602 44220 322918
rect 42812 315574 43286 315602
rect 44192 315574 44482 315602
rect 45664 315588 45692 322918
rect 46584 315602 46612 322918
rect 47964 320210 47992 322932
rect 48332 322918 48990 322946
rect 49712 322918 50094 322946
rect 51092 322918 51198 322946
rect 52302 322918 52408 322946
rect 53314 322918 53788 322946
rect 46940 320204 46992 320210
rect 46940 320146 46992 320152
rect 47952 320204 48004 320210
rect 47952 320146 48004 320152
rect 46584 315574 46874 315602
rect 46952 315466 46980 320146
rect 48332 315466 48360 322918
rect 49712 315466 49740 322918
rect 51092 315466 51120 322918
rect 52380 320226 52408 322918
rect 53760 320226 53788 322918
rect 54404 320890 54432 322932
rect 55522 322918 56088 322946
rect 54392 320884 54444 320890
rect 54392 320826 54444 320832
rect 55312 320884 55364 320890
rect 55312 320826 55364 320832
rect 52380 320198 52500 320226
rect 53760 320198 53880 320226
rect 52472 315602 52500 320198
rect 53852 315602 53880 320198
rect 55324 315602 55352 320826
rect 52472 315574 52854 315602
rect 53852 315574 54050 315602
rect 55246 315574 55352 315602
rect 56060 315602 56088 322918
rect 56520 320226 56548 322932
rect 57638 322918 57928 322946
rect 58742 322918 59308 322946
rect 57900 320226 57928 322918
rect 59280 320226 59308 322918
rect 56520 320198 56640 320226
rect 57900 320198 58020 320226
rect 59280 320198 59400 320226
rect 59832 320210 59860 322932
rect 60844 320210 60872 322932
rect 61948 320278 61976 322932
rect 61936 320272 61988 320278
rect 61936 320214 61988 320220
rect 63052 320210 63080 322932
rect 64064 320890 64092 322932
rect 64052 320884 64104 320890
rect 64052 320826 64104 320832
rect 64880 320884 64932 320890
rect 64880 320826 64932 320832
rect 63500 320272 63552 320278
rect 63500 320214 63552 320220
rect 56060 315574 56442 315602
rect 56612 315466 56640 320198
rect 57992 315466 58020 320198
rect 59372 315466 59400 320198
rect 59820 320204 59872 320210
rect 59820 320146 59872 320152
rect 60740 320204 60792 320210
rect 60740 320146 60792 320152
rect 60832 320204 60884 320210
rect 60832 320146 60884 320152
rect 62120 320204 62172 320210
rect 62120 320146 62172 320152
rect 63040 320204 63092 320210
rect 63040 320146 63092 320152
rect 60752 315466 60780 320146
rect 62132 315602 62160 320146
rect 63512 315602 63540 320214
rect 64328 320204 64380 320210
rect 64328 320146 64380 320152
rect 64340 315602 64368 320146
rect 64892 315738 64920 320826
rect 65168 320210 65196 322932
rect 66272 320346 66300 322932
rect 66260 320340 66312 320346
rect 66260 320282 66312 320288
rect 67376 320210 67404 322932
rect 67640 320340 67692 320346
rect 67640 320282 67692 320288
rect 65156 320204 65208 320210
rect 65156 320146 65208 320152
rect 66260 320204 66312 320210
rect 66260 320146 66312 320152
rect 67364 320204 67416 320210
rect 67364 320146 67416 320152
rect 64892 315710 65564 315738
rect 62132 315574 62422 315602
rect 63512 315574 63618 315602
rect 64340 315574 64814 315602
rect 65536 315466 65564 315710
rect 66272 315466 66300 320146
rect 67652 315466 67680 320282
rect 68388 320278 68416 322932
rect 68376 320272 68428 320278
rect 68376 320214 68428 320220
rect 69492 320210 69520 322932
rect 70596 320278 70624 322932
rect 71608 320346 71636 322932
rect 72712 320890 72740 322932
rect 72700 320884 72752 320890
rect 72700 320826 72752 320832
rect 73816 320822 73844 322932
rect 74540 320884 74592 320890
rect 74540 320826 74592 320832
rect 73804 320816 73856 320822
rect 73804 320758 73856 320764
rect 71596 320340 71648 320346
rect 71596 320282 71648 320288
rect 73896 320340 73948 320346
rect 73896 320282 73948 320288
rect 70400 320272 70452 320278
rect 70400 320214 70452 320220
rect 70584 320272 70636 320278
rect 70584 320214 70636 320220
rect 73252 320272 73304 320278
rect 73252 320214 73304 320220
rect 69020 320204 69072 320210
rect 69020 320146 69072 320152
rect 69480 320204 69532 320210
rect 69480 320146 69532 320152
rect 69032 315466 69060 320146
rect 70412 315602 70440 320214
rect 71780 320204 71832 320210
rect 71780 320146 71832 320152
rect 71792 315602 71820 320146
rect 73264 315602 73292 320214
rect 70412 315574 70794 315602
rect 71792 315574 71990 315602
rect 73186 315574 73292 315602
rect 73908 315602 73936 320282
rect 73908 315574 74382 315602
rect 74552 315466 74580 320826
rect 74920 320210 74948 322932
rect 75932 320958 75960 322932
rect 75920 320952 75972 320958
rect 75920 320894 75972 320900
rect 75920 320816 75972 320822
rect 75920 320758 75972 320764
rect 74908 320204 74960 320210
rect 74908 320146 74960 320152
rect 75932 315466 75960 320758
rect 77036 320278 77064 322932
rect 78140 320414 78168 322932
rect 78680 320952 78732 320958
rect 78680 320894 78732 320900
rect 78128 320408 78180 320414
rect 78128 320350 78180 320356
rect 77024 320272 77076 320278
rect 77024 320214 77076 320220
rect 77300 320204 77352 320210
rect 77300 320146 77352 320152
rect 77312 315466 77340 320146
rect 78692 315602 78720 320894
rect 79152 320210 79180 322932
rect 80256 320346 80284 322932
rect 81256 320408 81308 320414
rect 81256 320350 81308 320356
rect 80244 320340 80296 320346
rect 80244 320282 80296 320288
rect 79968 320272 80020 320278
rect 79968 320214 80020 320220
rect 79140 320204 79192 320210
rect 79140 320146 79192 320152
rect 79980 318730 80008 320214
rect 81268 318730 81296 320350
rect 81360 320278 81388 322932
rect 82464 320890 82492 322932
rect 82452 320884 82504 320890
rect 82452 320826 82504 320832
rect 83476 320754 83504 322932
rect 83464 320748 83516 320754
rect 83464 320690 83516 320696
rect 83004 320340 83056 320346
rect 83004 320282 83056 320288
rect 81348 320272 81400 320278
rect 81348 320214 81400 320220
rect 82820 320272 82872 320278
rect 82820 320214 82872 320220
rect 81624 320204 81676 320210
rect 81624 320146 81676 320152
rect 79980 318702 80376 318730
rect 81268 318702 81572 318730
rect 78692 315574 79166 315602
rect 80348 315588 80376 318702
rect 81544 315588 81572 318702
rect 81636 315738 81664 320146
rect 82832 317558 82860 320214
rect 82820 317552 82872 317558
rect 82820 317494 82872 317500
rect 83016 317370 83044 320282
rect 84580 320210 84608 322932
rect 85684 320890 85712 322932
rect 85120 320884 85172 320890
rect 85120 320826 85172 320832
rect 85672 320884 85724 320890
rect 85672 320826 85724 320832
rect 84568 320204 84620 320210
rect 84568 320146 84620 320152
rect 85132 318442 85160 320826
rect 85672 320748 85724 320754
rect 85672 320690 85724 320696
rect 85120 318436 85172 318442
rect 85120 318378 85172 318384
rect 85684 318374 85712 320690
rect 86696 320346 86724 322932
rect 86684 320340 86736 320346
rect 86684 320282 86736 320288
rect 87800 320210 87828 322932
rect 88904 320414 88932 322932
rect 89628 320884 89680 320890
rect 89628 320826 89680 320832
rect 88892 320408 88944 320414
rect 88892 320350 88944 320356
rect 87696 320204 87748 320210
rect 87696 320146 87748 320152
rect 87788 320204 87840 320210
rect 87788 320146 87840 320152
rect 86316 318436 86368 318442
rect 86316 318378 86368 318384
rect 85672 318368 85724 318374
rect 85672 318310 85724 318316
rect 85120 317552 85172 317558
rect 85120 317494 85172 317500
rect 82832 317342 83044 317370
rect 81636 315710 82308 315738
rect 82280 315466 82308 315710
rect 82832 315466 82860 317342
rect 85132 315588 85160 317494
rect 86328 315588 86356 318378
rect 87512 318368 87564 318374
rect 87512 318310 87564 318316
rect 87524 315588 87552 318310
rect 87708 318238 87736 320146
rect 89640 318730 89668 320826
rect 90008 320278 90036 322932
rect 91020 320482 91048 322932
rect 92124 321094 92152 322932
rect 92112 321088 92164 321094
rect 92112 321030 92164 321036
rect 93228 320958 93256 322932
rect 93216 320952 93268 320958
rect 93216 320894 93268 320900
rect 91008 320476 91060 320482
rect 91008 320418 91060 320424
rect 94240 320414 94268 322932
rect 95240 320476 95292 320482
rect 95240 320418 95292 320424
rect 92388 320408 92440 320414
rect 92388 320350 92440 320356
rect 94228 320408 94280 320414
rect 94228 320350 94280 320356
rect 91100 320340 91152 320346
rect 91100 320282 91152 320288
rect 89996 320272 90048 320278
rect 89996 320214 90048 320220
rect 90180 320204 90232 320210
rect 90180 320146 90232 320152
rect 90192 318782 90220 320146
rect 90180 318776 90232 318782
rect 89640 318702 89944 318730
rect 90180 318718 90232 318724
rect 87696 318232 87748 318238
rect 87696 318174 87748 318180
rect 88708 318232 88760 318238
rect 88708 318174 88760 318180
rect 88720 315588 88748 318174
rect 89916 315588 89944 318702
rect 91112 315588 91140 320282
rect 92296 318776 92348 318782
rect 92296 318718 92348 318724
rect 92308 315588 92336 318718
rect 92400 318578 92428 320350
rect 92756 320272 92808 320278
rect 92756 320214 92808 320220
rect 92388 318572 92440 318578
rect 92388 318514 92440 318520
rect 92768 317490 92796 320214
rect 93492 318572 93544 318578
rect 93492 318514 93544 318520
rect 92756 317484 92808 317490
rect 92756 317426 92808 317432
rect 93504 315588 93532 318514
rect 94688 317484 94740 317490
rect 94688 317426 94740 317432
rect 94700 315588 94728 317426
rect 95252 315466 95280 320418
rect 95344 320210 95372 322932
rect 96448 320278 96476 322932
rect 96620 321088 96672 321094
rect 96620 321030 96672 321036
rect 96436 320272 96488 320278
rect 96436 320214 96488 320220
rect 95332 320204 95384 320210
rect 95332 320146 95384 320152
rect 96632 315466 96660 321030
rect 97552 320346 97580 322932
rect 98000 320952 98052 320958
rect 98000 320894 98052 320900
rect 97540 320340 97592 320346
rect 97540 320282 97592 320288
rect 98012 315602 98040 320894
rect 98564 320618 98592 322932
rect 98552 320612 98604 320618
rect 98552 320554 98604 320560
rect 99668 320482 99696 322932
rect 100772 321230 100800 322932
rect 100760 321224 100812 321230
rect 100760 321166 100812 321172
rect 101784 321026 101812 322932
rect 101772 321020 101824 321026
rect 101772 320962 101824 320968
rect 102888 320958 102916 322932
rect 102876 320952 102928 320958
rect 102876 320894 102928 320900
rect 103520 320612 103572 320618
rect 103520 320554 103572 320560
rect 99656 320476 99708 320482
rect 99656 320418 99708 320424
rect 99564 320408 99616 320414
rect 99564 320350 99616 320356
rect 98736 320204 98788 320210
rect 98736 320146 98788 320152
rect 98748 318578 98776 320146
rect 98736 318572 98788 318578
rect 98736 318514 98788 318520
rect 99576 315602 99604 320350
rect 102140 320340 102192 320346
rect 102140 320282 102192 320288
rect 100760 320272 100812 320278
rect 100760 320214 100812 320220
rect 100668 318572 100720 318578
rect 100668 318514 100720 318520
rect 98012 315574 98302 315602
rect 99498 315574 99604 315602
rect 100680 315588 100708 318514
rect 100772 315466 100800 320214
rect 102152 315466 102180 320282
rect 103532 315466 103560 320554
rect 103992 320346 104020 322932
rect 104900 320476 104952 320482
rect 104900 320418 104952 320424
rect 103980 320340 104032 320346
rect 103980 320282 104032 320288
rect 104912 315466 104940 320418
rect 105096 320278 105124 322932
rect 106108 320890 106136 322932
rect 106280 321224 106332 321230
rect 106280 321166 106332 321172
rect 106096 320884 106148 320890
rect 106096 320826 106148 320832
rect 105084 320272 105136 320278
rect 105084 320214 105136 320220
rect 106292 315602 106320 321166
rect 106372 321020 106424 321026
rect 106372 320962 106424 320968
rect 106384 318578 106412 320962
rect 107212 320210 107240 322932
rect 108316 321094 108344 322932
rect 108304 321088 108356 321094
rect 108304 321030 108356 321036
rect 109328 321026 109356 322932
rect 109316 321020 109368 321026
rect 109316 320962 109368 320968
rect 108948 320952 109000 320958
rect 108948 320894 109000 320900
rect 107200 320204 107252 320210
rect 107200 320146 107252 320152
rect 108960 318730 108988 320894
rect 110432 320822 110460 322932
rect 111536 321162 111564 322932
rect 112654 322918 113128 322946
rect 111524 321156 111576 321162
rect 111524 321098 111576 321104
rect 110420 320816 110472 320822
rect 110420 320758 110472 320764
rect 109776 320340 109828 320346
rect 109776 320282 109828 320288
rect 108960 318702 109080 318730
rect 106372 318572 106424 318578
rect 106372 318514 106424 318520
rect 107844 318572 107896 318578
rect 107844 318514 107896 318520
rect 106292 315574 106674 315602
rect 107856 315588 107884 318514
rect 109052 315588 109080 318702
rect 109788 315602 109816 320282
rect 110420 320272 110472 320278
rect 110420 320214 110472 320220
rect 110432 316010 110460 320214
rect 112444 320204 112496 320210
rect 112444 320146 112496 320152
rect 110432 315982 111012 316010
rect 109788 315574 110262 315602
rect 110984 315466 111012 315982
rect 41432 315438 42090 315466
rect 46952 315438 48070 315466
rect 48332 315438 49266 315466
rect 49712 315438 50462 315466
rect 51092 315438 51658 315466
rect 56612 315438 57638 315466
rect 57992 315438 58834 315466
rect 59372 315438 60030 315466
rect 60752 315438 61226 315466
rect 65536 315438 66010 315466
rect 66272 315438 67206 315466
rect 67652 315438 68402 315466
rect 69032 315438 69598 315466
rect 74552 315438 75578 315466
rect 75932 315438 76774 315466
rect 77312 315438 77970 315466
rect 82280 315438 82754 315466
rect 82832 315438 83950 315466
rect 95252 315438 95910 315466
rect 96632 315438 97106 315466
rect 100772 315438 101890 315466
rect 102152 315438 103086 315466
rect 103532 315438 104282 315466
rect 104912 315438 105478 315466
rect 110984 315438 111458 315466
rect 26884 315376 26936 315382
rect 26884 315318 26936 315324
rect 111800 315376 111852 315382
rect 111800 315318 111852 315324
rect 15844 315308 15896 315314
rect 15844 315250 15896 315256
rect 111812 313682 111840 315318
rect 111800 313676 111852 313682
rect 111800 313618 111852 313624
rect 15844 294024 15896 294030
rect 15844 293966 15896 293972
rect 15856 227050 15884 293966
rect 17132 276004 17184 276010
rect 17132 275946 17184 275952
rect 17144 274961 17172 275946
rect 17130 274952 17186 274961
rect 17130 274887 17186 274896
rect 15844 227044 15896 227050
rect 15844 226986 15896 226992
rect 14464 225616 14516 225622
rect 14464 225558 14516 225564
rect 112456 224262 112484 320146
rect 113100 224534 113128 322918
rect 113652 319462 113680 322932
rect 113824 320816 113876 320822
rect 113824 320758 113876 320764
rect 113180 319456 113232 319462
rect 113180 319398 113232 319404
rect 113640 319456 113692 319462
rect 113640 319398 113692 319404
rect 113192 295361 113220 319398
rect 113548 313676 113600 313682
rect 113548 313618 113600 313624
rect 113560 311642 113588 313618
rect 113548 311636 113600 311642
rect 113548 311578 113600 311584
rect 113178 295352 113234 295361
rect 113178 295287 113234 295296
rect 113836 224602 113864 320758
rect 114756 320210 114784 322932
rect 115204 321088 115256 321094
rect 115204 321030 115256 321036
rect 114744 320204 114796 320210
rect 114744 320146 114796 320152
rect 113914 254552 113970 254561
rect 113914 254487 113970 254496
rect 113928 235958 113956 254487
rect 113916 235952 113968 235958
rect 113916 235894 113968 235900
rect 115216 224874 115244 321030
rect 115860 320958 115888 322932
rect 116886 322918 117268 322946
rect 117990 322918 118648 322946
rect 115848 320952 115900 320958
rect 115848 320894 115900 320900
rect 115848 320204 115900 320210
rect 115848 320146 115900 320152
rect 115204 224868 115256 224874
rect 115204 224810 115256 224816
rect 115860 224670 115888 320146
rect 116584 311636 116636 311642
rect 116584 311578 116636 311584
rect 115848 224664 115900 224670
rect 115848 224606 115900 224612
rect 113824 224596 113876 224602
rect 113824 224538 113876 224544
rect 113088 224528 113140 224534
rect 113088 224470 113140 224476
rect 112444 224256 112496 224262
rect 112444 224198 112496 224204
rect 13084 222896 13136 222902
rect 13084 222838 13136 222844
rect 116398 221232 116454 221241
rect 116398 221167 116454 221176
rect 116412 220930 116440 221167
rect 55220 220924 55272 220930
rect 55220 220866 55272 220872
rect 116400 220924 116452 220930
rect 116400 220866 116452 220872
rect 11704 220108 11756 220114
rect 11704 220050 11756 220056
rect 55232 219708 55260 220866
rect 116122 220008 116178 220017
rect 116122 219943 116178 219952
rect 116136 219502 116164 219943
rect 116124 219496 116176 219502
rect 116124 219438 116176 219444
rect 104808 219428 104860 219434
rect 104808 219370 104860 219376
rect 104820 219337 104848 219370
rect 104806 219328 104862 219337
rect 104806 219263 104862 219272
rect 116398 218920 116454 218929
rect 116398 218855 116454 218864
rect 116412 218074 116440 218855
rect 116400 218068 116452 218074
rect 116400 218010 116452 218016
rect 104808 218000 104860 218006
rect 104806 217968 104808 217977
rect 104860 217968 104862 217977
rect 104806 217903 104862 217912
rect 116398 217696 116454 217705
rect 116398 217631 116454 217640
rect 116412 216714 116440 217631
rect 116400 216708 116452 216714
rect 116400 216650 116452 216656
rect 104808 216640 104860 216646
rect 104806 216608 104808 216617
rect 104860 216608 104862 216617
rect 104806 216543 104862 216552
rect 115938 216608 115994 216617
rect 115938 216543 115994 216552
rect 115952 215966 115980 216543
rect 104808 215960 104860 215966
rect 104808 215902 104860 215908
rect 115940 215960 115992 215966
rect 115940 215902 115992 215908
rect 104820 215665 104848 215902
rect 104806 215656 104862 215665
rect 104806 215591 104862 215600
rect 116398 215384 116454 215393
rect 116398 215319 116400 215328
rect 116452 215319 116454 215328
rect 116400 215290 116452 215296
rect 104808 215280 104860 215286
rect 104808 215222 104860 215228
rect 104820 214713 104848 215222
rect 104806 214704 104862 214713
rect 104806 214639 104862 214648
rect 116398 214160 116454 214169
rect 116398 214095 116454 214104
rect 116412 213994 116440 214095
rect 116400 213988 116452 213994
rect 116400 213930 116452 213936
rect 104808 213920 104860 213926
rect 104808 213862 104860 213868
rect 104820 213489 104848 213862
rect 104806 213480 104862 213489
rect 104806 213415 104862 213424
rect 115938 213072 115994 213081
rect 115938 213007 115994 213016
rect 115952 212566 115980 213007
rect 115940 212560 115992 212566
rect 115940 212502 115992 212508
rect 104440 212492 104492 212498
rect 104440 212434 104492 212440
rect 104452 212129 104480 212434
rect 104438 212120 104494 212129
rect 104438 212055 104494 212064
rect 116306 211848 116362 211857
rect 116306 211783 116362 211792
rect 116320 211206 116348 211783
rect 116308 211200 116360 211206
rect 116308 211142 116360 211148
rect 104808 211132 104860 211138
rect 104808 211074 104860 211080
rect 104820 210905 104848 211074
rect 104806 210896 104862 210905
rect 104806 210831 104862 210840
rect 116306 210760 116362 210769
rect 116306 210695 116362 210704
rect 116320 209846 116348 210695
rect 116308 209840 116360 209846
rect 116308 209782 116360 209788
rect 104808 209772 104860 209778
rect 104808 209714 104860 209720
rect 104820 209545 104848 209714
rect 104806 209536 104862 209545
rect 104806 209471 104862 209480
rect 116030 209536 116086 209545
rect 116030 209471 116086 209480
rect 116044 208418 116072 209471
rect 116032 208412 116084 208418
rect 116032 208354 116084 208360
rect 104808 208344 104860 208350
rect 104808 208286 104860 208292
rect 115938 208312 115994 208321
rect 104820 208185 104848 208286
rect 115938 208247 115994 208256
rect 104806 208176 104862 208185
rect 104806 208111 104862 208120
rect 113088 207120 113140 207126
rect 113088 207062 113140 207068
rect 104806 206952 104862 206961
rect 104806 206887 104808 206896
rect 104860 206887 104862 206896
rect 104808 206858 104860 206864
rect 113100 206854 113128 207062
rect 115952 207058 115980 208247
rect 116030 207224 116086 207233
rect 116030 207159 116086 207168
rect 116044 207126 116072 207159
rect 116032 207120 116084 207126
rect 116032 207062 116084 207068
rect 115940 207052 115992 207058
rect 115940 206994 115992 207000
rect 104716 206848 104768 206854
rect 104716 206790 104768 206796
rect 113088 206848 113140 206854
rect 113088 206790 113140 206796
rect 104728 206281 104756 206790
rect 104714 206272 104770 206281
rect 104714 206207 104770 206216
rect 115938 206000 115994 206009
rect 115938 205935 115994 205944
rect 115952 205698 115980 205935
rect 115940 205692 115992 205698
rect 115940 205634 115992 205640
rect 104808 205624 104860 205630
rect 104808 205566 104860 205572
rect 104820 205057 104848 205566
rect 104806 205048 104862 205057
rect 104806 204983 104862 204992
rect 116398 204912 116454 204921
rect 116398 204847 116454 204856
rect 116412 204338 116440 204847
rect 116400 204332 116452 204338
rect 116400 204274 116452 204280
rect 104808 204264 104860 204270
rect 104808 204206 104860 204212
rect 104820 203697 104848 204206
rect 104806 203688 104862 203697
rect 104806 203623 104862 203632
rect 116306 203688 116362 203697
rect 116306 203623 116362 203632
rect 116320 202910 116348 203623
rect 116308 202904 116360 202910
rect 116308 202846 116360 202852
rect 104808 202836 104860 202842
rect 104808 202778 104860 202784
rect 104820 202473 104848 202778
rect 104806 202464 104862 202473
rect 104806 202399 104862 202408
rect 116122 202464 116178 202473
rect 116122 202399 116178 202408
rect 116136 201550 116164 202399
rect 116124 201544 116176 201550
rect 116124 201486 116176 201492
rect 104808 201476 104860 201482
rect 104808 201418 104860 201424
rect 104820 201113 104848 201418
rect 116122 201376 116178 201385
rect 116122 201311 116178 201320
rect 104806 201104 104862 201113
rect 104806 201039 104862 201048
rect 116136 200258 116164 201311
rect 116124 200252 116176 200258
rect 116124 200194 116176 200200
rect 113272 200184 113324 200190
rect 115940 200184 115992 200190
rect 113272 200126 113324 200132
rect 115938 200152 115940 200161
rect 115992 200152 115994 200161
rect 104808 200116 104860 200122
rect 104808 200058 104860 200064
rect 104820 199889 104848 200058
rect 104806 199880 104862 199889
rect 104806 199815 104862 199824
rect 113180 198756 113232 198762
rect 113180 198698 113232 198704
rect 104808 198688 104860 198694
rect 104808 198630 104860 198636
rect 104820 198529 104848 198630
rect 104806 198520 104862 198529
rect 104806 198455 104862 198464
rect 113192 197418 113220 198698
rect 113284 198694 113312 200126
rect 115938 200087 115994 200096
rect 116398 199064 116454 199073
rect 116398 198999 116454 199008
rect 116412 198762 116440 198999
rect 116400 198756 116452 198762
rect 116400 198698 116452 198704
rect 113272 198688 113324 198694
rect 113272 198630 113324 198636
rect 116398 197840 116454 197849
rect 116398 197775 116454 197784
rect 113100 197390 113220 197418
rect 116412 197402 116440 197775
rect 116400 197396 116452 197402
rect 113100 197334 113128 197390
rect 116400 197338 116452 197344
rect 104808 197328 104860 197334
rect 104806 197296 104808 197305
rect 113088 197328 113140 197334
rect 104860 197296 104862 197305
rect 104532 197260 104584 197266
rect 113088 197270 113140 197276
rect 104806 197231 104862 197240
rect 104532 197202 104584 197208
rect 104544 196625 104572 197202
rect 116398 196752 116454 196761
rect 116398 196687 116454 196696
rect 104530 196616 104586 196625
rect 104530 196551 104586 196560
rect 116412 196042 116440 196687
rect 116400 196036 116452 196042
rect 116400 195978 116452 195984
rect 104808 195968 104860 195974
rect 104808 195910 104860 195916
rect 104820 195401 104848 195910
rect 115938 195528 115994 195537
rect 115938 195463 115994 195472
rect 104806 195392 104862 195401
rect 104806 195327 104862 195336
rect 115952 194614 115980 195463
rect 115940 194608 115992 194614
rect 115940 194550 115992 194556
rect 104808 194540 104860 194546
rect 104808 194482 104860 194488
rect 104820 194041 104848 194482
rect 116122 194304 116178 194313
rect 116122 194239 116178 194248
rect 104806 194032 104862 194041
rect 104806 193967 104862 193976
rect 116136 193254 116164 194239
rect 116124 193248 116176 193254
rect 116124 193190 116176 193196
rect 116398 193216 116454 193225
rect 104440 193180 104492 193186
rect 116398 193151 116454 193160
rect 104440 193122 104492 193128
rect 104452 192817 104480 193122
rect 104438 192808 104494 192817
rect 104438 192743 104494 192752
rect 116412 192030 116440 193151
rect 113180 192024 113232 192030
rect 116400 192024 116452 192030
rect 113180 191966 113232 191972
rect 116030 191992 116086 192001
rect 113192 191826 113220 191966
rect 113272 191956 113324 191962
rect 116400 191966 116452 191972
rect 116030 191927 116032 191936
rect 113272 191898 113324 191904
rect 116084 191927 116086 191936
rect 116032 191898 116084 191904
rect 104808 191820 104860 191826
rect 104808 191762 104860 191768
rect 113180 191820 113232 191826
rect 113180 191762 113232 191768
rect 104820 191457 104848 191762
rect 104806 191448 104862 191457
rect 104806 191383 104862 191392
rect 113284 190466 113312 191898
rect 116490 190904 116546 190913
rect 116490 190839 116546 190848
rect 116504 190670 116532 190839
rect 113364 190664 113416 190670
rect 113364 190606 113416 190612
rect 116492 190664 116544 190670
rect 116492 190606 116544 190612
rect 104716 190460 104768 190466
rect 104716 190402 104768 190408
rect 113272 190460 113324 190466
rect 113272 190402 113324 190408
rect 104728 190233 104756 190402
rect 104714 190224 104770 190233
rect 104714 190159 104770 190168
rect 113376 189038 113404 190606
rect 116398 189680 116454 189689
rect 116398 189615 116454 189624
rect 116412 189106 116440 189615
rect 114192 189100 114244 189106
rect 114192 189042 114244 189048
rect 116400 189100 116452 189106
rect 116400 189042 116452 189048
rect 104808 189032 104860 189038
rect 104808 188974 104860 188980
rect 113364 189032 113416 189038
rect 113364 188974 113416 188980
rect 104820 188873 104848 188974
rect 104806 188864 104862 188873
rect 104806 188799 104862 188808
rect 113180 187740 113232 187746
rect 113180 187682 113232 187688
rect 104808 187672 104860 187678
rect 104808 187614 104860 187620
rect 104820 187513 104848 187614
rect 104806 187504 104862 187513
rect 104806 187439 104862 187448
rect 113192 186402 113220 187682
rect 114204 187678 114232 189042
rect 116214 188456 116270 188465
rect 116214 188391 116270 188400
rect 116228 187746 116256 188391
rect 116216 187740 116268 187746
rect 116216 187682 116268 187688
rect 114192 187672 114244 187678
rect 114192 187614 114244 187620
rect 116306 187368 116362 187377
rect 116306 187303 116362 187312
rect 113100 186374 113220 186402
rect 116320 186386 116348 187303
rect 116308 186380 116360 186386
rect 113100 186318 113128 186374
rect 116308 186322 116360 186328
rect 104808 186312 104860 186318
rect 104806 186280 104808 186289
rect 113088 186312 113140 186318
rect 104860 186280 104862 186289
rect 104532 186244 104584 186250
rect 113088 186254 113140 186260
rect 104806 186215 104862 186224
rect 104532 186186 104584 186192
rect 104544 185609 104572 186186
rect 116030 186144 116086 186153
rect 116030 186079 116086 186088
rect 104530 185600 104586 185609
rect 104530 185535 104586 185544
rect 114468 185020 114520 185026
rect 114468 184962 114520 184968
rect 104808 184884 104860 184890
rect 104808 184826 104860 184832
rect 104820 184385 104848 184826
rect 104806 184376 104862 184385
rect 104806 184311 104862 184320
rect 114376 183592 114428 183598
rect 114376 183534 114428 183540
rect 104808 183524 104860 183530
rect 104808 183466 104860 183472
rect 104820 183025 104848 183466
rect 104806 183016 104862 183025
rect 104806 182951 104862 182960
rect 113180 182232 113232 182238
rect 113180 182174 113232 182180
rect 104808 182164 104860 182170
rect 104808 182106 104860 182112
rect 104820 181801 104848 182106
rect 104806 181792 104862 181801
rect 104806 181727 104862 181736
rect 113192 180810 113220 182174
rect 114388 182170 114416 183534
rect 114480 183530 114508 184962
rect 116044 184958 116072 186079
rect 116398 185056 116454 185065
rect 116398 184991 116400 185000
rect 116452 184991 116454 185000
rect 116400 184962 116452 184968
rect 116032 184952 116084 184958
rect 116032 184894 116084 184900
rect 116398 183832 116454 183841
rect 116398 183767 116454 183776
rect 116412 183598 116440 183767
rect 116400 183592 116452 183598
rect 116400 183534 116452 183540
rect 114468 183524 114520 183530
rect 114468 183466 114520 183472
rect 115938 182608 115994 182617
rect 115938 182543 115994 182552
rect 115952 182238 115980 182543
rect 115940 182232 115992 182238
rect 115940 182174 115992 182180
rect 114376 182164 114428 182170
rect 114376 182106 114428 182112
rect 115938 181520 115994 181529
rect 115938 181455 115994 181464
rect 115952 181150 115980 181455
rect 113272 181144 113324 181150
rect 113272 181086 113324 181092
rect 115940 181144 115992 181150
rect 115940 181086 115992 181092
rect 104808 180804 104860 180810
rect 104808 180746 104860 180752
rect 113180 180804 113232 180810
rect 113180 180746 113232 180752
rect 104820 180441 104848 180746
rect 104806 180432 104862 180441
rect 104806 180367 104862 180376
rect 113284 179382 113312 181086
rect 116398 180296 116454 180305
rect 116398 180231 116454 180240
rect 116412 179450 116440 180231
rect 113916 179444 113968 179450
rect 113916 179386 113968 179392
rect 116400 179444 116452 179450
rect 116400 179386 116452 179392
rect 104808 179376 104860 179382
rect 104808 179318 104860 179324
rect 113272 179376 113324 179382
rect 113272 179318 113324 179324
rect 104820 179081 104848 179318
rect 104806 179072 104862 179081
rect 104806 179007 104862 179016
rect 113928 178022 113956 179386
rect 115938 179208 115994 179217
rect 115938 179143 115994 179152
rect 115952 178090 115980 179143
rect 114192 178084 114244 178090
rect 114192 178026 114244 178032
rect 115940 178084 115992 178090
rect 115940 178026 115992 178032
rect 104164 178016 104216 178022
rect 104164 177958 104216 177964
rect 113916 178016 113968 178022
rect 113916 177958 113968 177964
rect 104176 177857 104204 177958
rect 104162 177848 104218 177857
rect 104162 177783 104218 177792
rect 113916 176792 113968 176798
rect 113916 176734 113968 176740
rect 104164 176656 104216 176662
rect 104164 176598 104216 176604
rect 104176 176497 104204 176598
rect 104162 176488 104218 176497
rect 104162 176423 104218 176432
rect 104440 175228 104492 175234
rect 104440 175170 104492 175176
rect 104452 174729 104480 175170
rect 113928 175166 113956 176734
rect 114204 176662 114232 178026
rect 115938 177984 115994 177993
rect 115938 177919 115994 177928
rect 115952 176798 115980 177919
rect 116398 176896 116454 176905
rect 116398 176831 116454 176840
rect 115940 176792 115992 176798
rect 115940 176734 115992 176740
rect 116412 176730 116440 176831
rect 114468 176724 114520 176730
rect 114468 176666 114520 176672
rect 116400 176724 116452 176730
rect 116400 176666 116452 176672
rect 114192 176656 114244 176662
rect 114192 176598 114244 176604
rect 114284 175296 114336 175302
rect 114284 175238 114336 175244
rect 104808 175160 104860 175166
rect 104806 175128 104808 175137
rect 113916 175160 113968 175166
rect 104860 175128 104862 175137
rect 113916 175102 113968 175108
rect 104806 175063 104862 175072
rect 104438 174720 104494 174729
rect 104438 174655 104494 174664
rect 114296 173874 114324 175238
rect 114480 175234 114508 176666
rect 116398 175672 116454 175681
rect 116398 175607 116454 175616
rect 116412 175302 116440 175607
rect 116400 175296 116452 175302
rect 116400 175238 116452 175244
rect 114468 175228 114520 175234
rect 114468 175170 114520 175176
rect 115938 174448 115994 174457
rect 115938 174383 115994 174392
rect 115952 173942 115980 174383
rect 114376 173936 114428 173942
rect 114376 173878 114428 173884
rect 115940 173936 115992 173942
rect 115940 173878 115992 173884
rect 104808 173868 104860 173874
rect 104808 173810 104860 173816
rect 114284 173868 114336 173874
rect 114284 173810 114336 173816
rect 104820 173369 104848 173810
rect 104806 173360 104862 173369
rect 104806 173295 104862 173304
rect 113180 172576 113232 172582
rect 113180 172518 113232 172524
rect 104440 172508 104492 172514
rect 104440 172450 104492 172456
rect 104452 172145 104480 172450
rect 104438 172136 104494 172145
rect 104438 172071 104494 172080
rect 113192 171086 113220 172518
rect 114388 172514 114416 173878
rect 116398 173360 116454 173369
rect 116398 173295 116454 173304
rect 116412 172582 116440 173295
rect 116400 172576 116452 172582
rect 116400 172518 116452 172524
rect 114376 172508 114428 172514
rect 114376 172450 114428 172456
rect 116122 172136 116178 172145
rect 116122 172071 116178 172080
rect 116136 171630 116164 172071
rect 113272 171624 113324 171630
rect 113272 171566 113324 171572
rect 116124 171624 116176 171630
rect 116124 171566 116176 171572
rect 104808 171080 104860 171086
rect 104808 171022 104860 171028
rect 113180 171080 113232 171086
rect 113180 171022 113232 171028
rect 104820 170785 104848 171022
rect 104806 170776 104862 170785
rect 104806 170711 104862 170720
rect 104256 169788 104308 169794
rect 104256 169730 104308 169736
rect 104164 168360 104216 168366
rect 104164 168302 104216 168308
rect 104176 168201 104204 168302
rect 104162 168192 104218 168201
rect 104162 168127 104218 168136
rect 104268 166977 104296 169730
rect 113284 169726 113312 171566
rect 116306 171048 116362 171057
rect 116306 170983 116362 170992
rect 116320 169862 116348 170983
rect 113916 169856 113968 169862
rect 113916 169798 113968 169804
rect 116308 169856 116360 169862
rect 116308 169798 116360 169804
rect 116398 169824 116454 169833
rect 104808 169720 104860 169726
rect 104808 169662 104860 169668
rect 113272 169720 113324 169726
rect 113272 169662 113324 169668
rect 104820 169425 104848 169662
rect 104806 169416 104862 169425
rect 104806 169351 104862 169360
rect 104808 168428 104860 168434
rect 104808 168370 104860 168376
rect 104254 166968 104310 166977
rect 104254 166903 104310 166912
rect 104820 165617 104848 168370
rect 113928 168366 113956 169798
rect 116398 169759 116400 169768
rect 116452 169759 116454 169768
rect 116400 169730 116452 169736
rect 116398 168600 116454 168609
rect 116398 168535 116454 168544
rect 116412 168434 116440 168535
rect 116400 168428 116452 168434
rect 116400 168370 116452 168376
rect 113916 168360 113968 168366
rect 113916 168302 113968 168308
rect 115938 167512 115994 167521
rect 115938 167447 115994 167456
rect 115952 167074 115980 167447
rect 114468 167068 114520 167074
rect 114468 167010 114520 167016
rect 115940 167068 115992 167074
rect 115940 167010 115992 167016
rect 113824 165640 113876 165646
rect 104806 165608 104862 165617
rect 104624 165572 104676 165578
rect 113824 165582 113876 165588
rect 104806 165543 104862 165552
rect 104624 165514 104676 165520
rect 104636 164937 104664 165514
rect 104622 164928 104678 164937
rect 104622 164863 104678 164872
rect 113836 164218 113864 165582
rect 114480 165578 114508 167010
rect 115938 166288 115994 166297
rect 115938 166223 115994 166232
rect 115952 165646 115980 166223
rect 115940 165640 115992 165646
rect 115940 165582 115992 165588
rect 114468 165572 114520 165578
rect 114468 165514 114520 165520
rect 116122 165200 116178 165209
rect 116122 165135 116178 165144
rect 116136 164286 116164 165135
rect 114468 164280 114520 164286
rect 114468 164222 114520 164228
rect 116124 164280 116176 164286
rect 116124 164222 116176 164228
rect 104808 164212 104860 164218
rect 104808 164154 104860 164160
rect 113824 164212 113876 164218
rect 113824 164154 113876 164160
rect 104820 163713 104848 164154
rect 104806 163704 104862 163713
rect 104806 163639 104862 163648
rect 113180 162920 113232 162926
rect 113180 162862 113232 162868
rect 104808 162852 104860 162858
rect 104808 162794 104860 162800
rect 104820 162353 104848 162794
rect 104806 162344 104862 162353
rect 104806 162279 104862 162288
rect 103704 161492 103756 161498
rect 103704 161434 103756 161440
rect 103716 158681 103744 161434
rect 113192 161430 113220 162862
rect 114480 162858 114508 164222
rect 116398 163976 116454 163985
rect 116398 163911 116454 163920
rect 116412 162926 116440 163911
rect 116400 162920 116452 162926
rect 116400 162862 116452 162868
rect 114468 162852 114520 162858
rect 114468 162794 114520 162800
rect 116214 162752 116270 162761
rect 116214 162687 116270 162696
rect 116228 162042 116256 162687
rect 113272 162036 113324 162042
rect 113272 161978 113324 161984
rect 116216 162036 116268 162042
rect 116216 161978 116268 161984
rect 104808 161424 104860 161430
rect 104808 161366 104860 161372
rect 113180 161424 113232 161430
rect 113180 161366 113232 161372
rect 104820 160993 104848 161366
rect 104806 160984 104862 160993
rect 104806 160919 104862 160928
rect 104256 160132 104308 160138
rect 104256 160074 104308 160080
rect 103702 158672 103758 158681
rect 103702 158607 103758 158616
rect 104268 157321 104296 160074
rect 113284 160070 113312 161978
rect 116398 161664 116454 161673
rect 116398 161599 116454 161608
rect 116412 161498 116440 161599
rect 116400 161492 116452 161498
rect 116400 161434 116452 161440
rect 116398 160440 116454 160449
rect 116398 160375 116454 160384
rect 116412 160138 116440 160375
rect 116400 160132 116452 160138
rect 116400 160074 116452 160080
rect 104808 160064 104860 160070
rect 104808 160006 104860 160012
rect 113272 160064 113324 160070
rect 113272 160006 113324 160012
rect 104820 159769 104848 160006
rect 104806 159760 104862 159769
rect 104806 159695 104862 159704
rect 116398 159352 116454 159361
rect 116398 159287 116454 159296
rect 116412 158778 116440 159287
rect 104808 158772 104860 158778
rect 104808 158714 104860 158720
rect 116400 158772 116452 158778
rect 116400 158714 116452 158720
rect 104348 157412 104400 157418
rect 104348 157354 104400 157360
rect 104254 157312 104310 157321
rect 104254 157247 104310 157256
rect 104164 154624 104216 154630
rect 104164 154566 104216 154572
rect 103796 153264 103848 153270
rect 103796 153206 103848 153212
rect 103704 151836 103756 151842
rect 103704 151778 103756 151784
rect 103716 149025 103744 151778
rect 103808 150385 103836 153206
rect 104176 151609 104204 154566
rect 104360 154465 104388 157354
rect 104820 155961 104848 158714
rect 116398 158128 116454 158137
rect 116398 158063 116454 158072
rect 116412 157418 116440 158063
rect 116400 157412 116452 157418
rect 116400 157354 116452 157360
rect 116030 157040 116086 157049
rect 116030 156975 116086 156984
rect 116044 155990 116072 156975
rect 114284 155984 114336 155990
rect 104806 155952 104862 155961
rect 114284 155926 114336 155932
rect 116032 155984 116084 155990
rect 116032 155926 116084 155932
rect 104806 155887 104862 155896
rect 113456 154692 113508 154698
rect 113456 154634 113508 154640
rect 104624 154556 104676 154562
rect 104624 154498 104676 154504
rect 104346 154456 104402 154465
rect 104346 154391 104402 154400
rect 104636 153921 104664 154498
rect 104622 153912 104678 153921
rect 104622 153847 104678 153856
rect 113468 153202 113496 154634
rect 114296 154562 114324 155926
rect 116030 155816 116086 155825
rect 116030 155751 116086 155760
rect 116044 154698 116072 155751
rect 116032 154692 116084 154698
rect 116032 154634 116084 154640
rect 116400 154624 116452 154630
rect 116398 154592 116400 154601
rect 116452 154592 116454 154601
rect 114284 154556 114336 154562
rect 116398 154527 116454 154536
rect 114284 154498 114336 154504
rect 115938 153504 115994 153513
rect 115938 153439 115994 153448
rect 115952 153270 115980 153439
rect 115940 153264 115992 153270
rect 115940 153206 115992 153212
rect 104808 153196 104860 153202
rect 104808 153138 104860 153144
rect 113456 153196 113508 153202
rect 113456 153138 113508 153144
rect 104820 152697 104848 153138
rect 104806 152688 104862 152697
rect 104806 152623 104862 152632
rect 116398 152280 116454 152289
rect 116398 152215 116454 152224
rect 116412 151842 116440 152215
rect 116400 151836 116452 151842
rect 116400 151778 116452 151784
rect 104162 151600 104218 151609
rect 104162 151535 104218 151544
rect 116398 151192 116454 151201
rect 116398 151127 116454 151136
rect 116412 150482 116440 151127
rect 104348 150476 104400 150482
rect 104348 150418 104400 150424
rect 116400 150476 116452 150482
rect 116400 150418 116452 150424
rect 103794 150376 103850 150385
rect 103794 150311 103850 150320
rect 103702 149016 103758 149025
rect 103702 148951 103758 148960
rect 104360 147665 104388 150418
rect 116398 149968 116454 149977
rect 116398 149903 116454 149912
rect 116412 149122 116440 149903
rect 104440 149116 104492 149122
rect 104440 149058 104492 149064
rect 116400 149116 116452 149122
rect 116400 149058 116452 149064
rect 104346 147656 104402 147665
rect 104346 147591 104402 147600
rect 104164 146328 104216 146334
rect 104452 146305 104480 149058
rect 116398 148744 116454 148753
rect 116398 148679 116454 148688
rect 116412 147694 116440 148679
rect 104808 147688 104860 147694
rect 116400 147688 116452 147694
rect 104808 147630 104860 147636
rect 115938 147656 115994 147665
rect 104164 146270 104216 146276
rect 104438 146296 104494 146305
rect 103520 143608 103572 143614
rect 103520 143550 103572 143556
rect 103532 140593 103560 143550
rect 104176 143041 104204 146270
rect 104438 146231 104494 146240
rect 104532 144968 104584 144974
rect 104532 144910 104584 144916
rect 104162 143032 104218 143041
rect 104162 142967 104218 142976
rect 103704 142180 103756 142186
rect 103704 142122 103756 142128
rect 103518 140584 103574 140593
rect 103518 140519 103574 140528
rect 103716 139369 103744 142122
rect 104544 141817 104572 144910
rect 104624 144900 104676 144906
rect 104624 144842 104676 144848
rect 104636 144265 104664 144842
rect 104820 144809 104848 147630
rect 116400 147630 116452 147636
rect 115938 147591 115994 147600
rect 115952 146402 115980 147591
rect 116398 146432 116454 146441
rect 113640 146396 113692 146402
rect 113640 146338 113692 146344
rect 115940 146396 115992 146402
rect 116398 146367 116454 146376
rect 115940 146338 115992 146344
rect 113652 144906 113680 146338
rect 116412 146334 116440 146367
rect 116400 146328 116452 146334
rect 116400 146270 116452 146276
rect 116030 145344 116086 145353
rect 116030 145279 116086 145288
rect 116044 144974 116072 145279
rect 116032 144968 116084 144974
rect 116032 144910 116084 144916
rect 113640 144900 113692 144906
rect 113640 144842 113692 144848
rect 104806 144800 104862 144809
rect 104806 144735 104862 144744
rect 104622 144256 104678 144265
rect 104622 144191 104678 144200
rect 116398 144120 116454 144129
rect 116398 144055 116454 144064
rect 116412 143614 116440 144055
rect 116400 143608 116452 143614
rect 116400 143550 116452 143556
rect 116398 142896 116454 142905
rect 116398 142831 116454 142840
rect 116412 142186 116440 142831
rect 116400 142180 116452 142186
rect 116400 142122 116452 142128
rect 104530 141808 104586 141817
rect 104530 141743 104586 141752
rect 116398 141808 116454 141817
rect 116398 141743 116454 141752
rect 116412 140826 116440 141743
rect 104348 140820 104400 140826
rect 104348 140762 104400 140768
rect 116400 140820 116452 140826
rect 116400 140762 116452 140768
rect 103702 139360 103758 139369
rect 103702 139295 103758 139304
rect 104360 138009 104388 140762
rect 116398 140584 116454 140593
rect 116398 140519 116454 140528
rect 113548 139528 113600 139534
rect 116308 139528 116360 139534
rect 113548 139470 113600 139476
rect 116306 139496 116308 139505
rect 116360 139496 116362 139505
rect 104808 139460 104860 139466
rect 104808 139402 104860 139408
rect 104346 138000 104402 138009
rect 104346 137935 104402 137944
rect 104716 136672 104768 136678
rect 104820 136649 104848 139402
rect 104716 136614 104768 136620
rect 104806 136640 104862 136649
rect 104348 135312 104400 135318
rect 104348 135254 104400 135260
rect 104360 132025 104388 135254
rect 104728 133249 104756 136614
rect 104806 136575 104862 136584
rect 113560 135250 113588 139470
rect 116412 139466 116440 140519
rect 116306 139431 116362 139440
rect 116400 139460 116452 139466
rect 116400 139402 116452 139408
rect 115846 138272 115902 138281
rect 115846 138207 115902 138216
rect 104808 135244 104860 135250
rect 104808 135186 104860 135192
rect 113548 135244 113600 135250
rect 113548 135186 113600 135192
rect 104820 135153 104848 135186
rect 104806 135144 104862 135153
rect 104806 135079 104862 135088
rect 109868 133952 109920 133958
rect 109868 133894 109920 133900
rect 104808 133884 104860 133890
rect 104808 133826 104860 133832
rect 104820 133793 104848 133826
rect 104806 133784 104862 133793
rect 104806 133719 104862 133728
rect 104714 133240 104770 133249
rect 104714 133175 104770 133184
rect 104346 132016 104402 132025
rect 104346 131951 104402 131960
rect 109880 130762 109908 133894
rect 115860 133890 115888 138207
rect 116398 137184 116454 137193
rect 116398 137119 116454 137128
rect 116412 136678 116440 137119
rect 116400 136672 116452 136678
rect 116400 136614 116452 136620
rect 115938 135960 115994 135969
rect 115938 135895 115994 135904
rect 115952 135318 115980 135895
rect 115940 135312 115992 135318
rect 115940 135254 115992 135260
rect 116398 134736 116454 134745
rect 116398 134671 116454 134680
rect 116412 133958 116440 134671
rect 116400 133952 116452 133958
rect 116400 133894 116452 133900
rect 115848 133884 115900 133890
rect 115848 133826 115900 133832
rect 114560 132932 114612 132938
rect 114560 132874 114612 132880
rect 113732 131164 113784 131170
rect 113732 131106 113784 131112
rect 103980 130756 104032 130762
rect 103980 130698 104032 130704
rect 109868 130756 109920 130762
rect 109868 130698 109920 130704
rect 103992 130665 104020 130698
rect 103978 130656 104034 130665
rect 103978 130591 104034 130600
rect 100760 130416 100812 130422
rect 100760 130358 100812 130364
rect 32232 125089 32260 127228
rect 78232 125526 78260 127228
rect 100772 125526 100800 130358
rect 104808 129736 104860 129742
rect 104808 129678 104860 129684
rect 104820 129305 104848 129678
rect 104806 129296 104862 129305
rect 104806 129231 104862 129240
rect 113744 128246 113772 131106
rect 114572 129742 114600 132874
rect 116122 132424 116178 132433
rect 116122 132359 116178 132368
rect 116136 131170 116164 132359
rect 116398 131336 116454 131345
rect 116398 131271 116454 131280
rect 116124 131164 116176 131170
rect 116124 131106 116176 131112
rect 116412 130422 116440 131271
rect 116400 130416 116452 130422
rect 116400 130358 116452 130364
rect 114560 129736 114612 129742
rect 114560 129678 114612 129684
rect 116400 129328 116452 129334
rect 116400 129270 116452 129276
rect 116412 128897 116440 129270
rect 116398 128888 116454 128897
rect 116398 128823 116454 128832
rect 116400 128308 116452 128314
rect 116400 128250 116452 128256
rect 104808 128240 104860 128246
rect 104808 128182 104860 128188
rect 113732 128240 113784 128246
rect 113732 128182 113784 128188
rect 104820 128081 104848 128182
rect 104806 128072 104862 128081
rect 104806 128007 104862 128016
rect 116412 127809 116440 128250
rect 116398 127800 116454 127809
rect 116398 127735 116454 127744
rect 116400 126948 116452 126954
rect 116400 126890 116452 126896
rect 116412 126585 116440 126890
rect 116398 126576 116454 126585
rect 116398 126511 116454 126520
rect 116400 125588 116452 125594
rect 116400 125530 116452 125536
rect 78220 125520 78272 125526
rect 78220 125462 78272 125468
rect 100760 125520 100812 125526
rect 116412 125497 116440 125530
rect 100760 125462 100812 125468
rect 116398 125488 116454 125497
rect 116398 125423 116454 125432
rect 32218 125080 32274 125089
rect 32218 125015 32274 125024
rect 116596 123049 116624 311578
rect 117240 236706 117268 322918
rect 117964 321156 118016 321162
rect 117964 321098 118016 321104
rect 117228 236700 117280 236706
rect 117228 236642 117280 236648
rect 117976 224738 118004 321098
rect 117964 224732 118016 224738
rect 117964 224674 118016 224680
rect 118620 224466 118648 322918
rect 119080 320210 119108 322932
rect 119344 321020 119396 321026
rect 119344 320962 119396 320968
rect 119068 320204 119120 320210
rect 119068 320146 119120 320152
rect 119356 224942 119384 320962
rect 120184 320210 120212 322932
rect 121210 322918 121408 322946
rect 122314 322918 122788 322946
rect 123418 322918 124168 322946
rect 119988 320204 120040 320210
rect 119988 320146 120040 320152
rect 120172 320204 120224 320210
rect 120172 320146 120224 320152
rect 121276 320204 121328 320210
rect 121276 320146 121328 320152
rect 119344 224936 119396 224942
rect 119344 224878 119396 224884
rect 120000 224806 120028 320146
rect 121288 227050 121316 320146
rect 120080 227044 120132 227050
rect 120080 226986 120132 226992
rect 121276 227044 121328 227050
rect 121276 226986 121328 226992
rect 119988 224800 120040 224806
rect 119988 224742 120040 224748
rect 118608 224460 118660 224466
rect 118608 224402 118660 224408
rect 120092 221748 120120 226986
rect 121380 224398 121408 322918
rect 121552 320884 121604 320890
rect 121552 320826 121604 320832
rect 121368 224392 121420 224398
rect 121368 224334 121420 224340
rect 121564 221626 121592 320826
rect 122760 224330 122788 322918
rect 122748 224324 122800 224330
rect 122748 224266 122800 224272
rect 123208 224256 123260 224262
rect 123208 224198 123260 224204
rect 123220 221748 123248 224198
rect 124140 224058 124168 322918
rect 124416 320210 124444 322932
rect 125428 322918 125534 322946
rect 126638 322918 126928 322946
rect 127742 322918 128308 322946
rect 124404 320204 124456 320210
rect 124404 320146 124456 320152
rect 125428 226658 125456 322918
rect 126244 320952 126296 320958
rect 126244 320894 126296 320900
rect 125508 320204 125560 320210
rect 125508 320146 125560 320152
rect 125244 226630 125456 226658
rect 124312 224868 124364 224874
rect 124312 224810 124364 224816
rect 124128 224052 124180 224058
rect 124128 223994 124180 224000
rect 124324 221748 124352 224810
rect 125244 224262 125272 226630
rect 125520 224942 125548 320146
rect 125416 224936 125468 224942
rect 125416 224878 125468 224884
rect 125508 224936 125560 224942
rect 125508 224878 125560 224884
rect 125232 224256 125284 224262
rect 125232 224198 125284 224204
rect 125428 221748 125456 224878
rect 126256 224806 126284 320894
rect 126152 224800 126204 224806
rect 126152 224742 126204 224748
rect 126244 224800 126296 224806
rect 126244 224742 126296 224748
rect 126164 224126 126192 224742
rect 126900 224602 126928 322918
rect 128280 224738 128308 322918
rect 128740 320210 128768 322932
rect 129844 320210 129872 322932
rect 130962 322918 131068 322946
rect 131974 322918 132448 322946
rect 128728 320204 128780 320210
rect 128728 320146 128780 320152
rect 129648 320204 129700 320210
rect 129648 320146 129700 320152
rect 129832 320204 129884 320210
rect 129832 320146 129884 320152
rect 130936 320204 130988 320210
rect 130936 320146 130988 320152
rect 128452 319456 128504 319462
rect 128452 319398 128504 319404
rect 127532 224732 127584 224738
rect 127532 224674 127584 224680
rect 128268 224732 128320 224738
rect 128268 224674 128320 224680
rect 126428 224596 126480 224602
rect 126428 224538 126480 224544
rect 126888 224596 126940 224602
rect 126888 224538 126940 224544
rect 126152 224120 126204 224126
rect 126152 224062 126204 224068
rect 126440 221748 126468 224538
rect 127544 221748 127572 224674
rect 128464 224618 128492 319398
rect 128464 224590 129228 224618
rect 128636 224528 128688 224534
rect 128636 224470 128688 224476
rect 128648 221748 128676 224470
rect 129200 221626 129228 224590
rect 129660 223990 129688 320146
rect 130948 224874 130976 320146
rect 130936 224868 130988 224874
rect 130936 224810 130988 224816
rect 130752 224664 130804 224670
rect 130752 224606 130804 224612
rect 129648 223984 129700 223990
rect 129648 223926 129700 223932
rect 130764 221748 130792 224606
rect 131040 224534 131068 322918
rect 131764 224800 131816 224806
rect 131764 224742 131816 224748
rect 131028 224528 131080 224534
rect 131028 224470 131080 224476
rect 131776 221748 131804 224742
rect 132420 224670 132448 322918
rect 133064 320210 133092 322932
rect 134168 320210 134196 322932
rect 135272 320210 135300 322932
rect 136298 322918 136588 322946
rect 137402 322918 137968 322946
rect 133052 320204 133104 320210
rect 133052 320146 133104 320152
rect 133788 320204 133840 320210
rect 133788 320146 133840 320152
rect 134156 320204 134208 320210
rect 134156 320146 134208 320152
rect 135168 320204 135220 320210
rect 135168 320146 135220 320152
rect 135260 320204 135312 320210
rect 135260 320146 135312 320152
rect 136456 320204 136508 320210
rect 136456 320146 136508 320152
rect 132500 236700 132552 236706
rect 132500 236642 132552 236648
rect 132408 224664 132460 224670
rect 132408 224606 132460 224612
rect 132512 221762 132540 236642
rect 133800 224942 133828 320146
rect 135180 227118 135208 320146
rect 135168 227112 135220 227118
rect 135168 227054 135220 227060
rect 136088 227044 136140 227050
rect 136088 226986 136140 226992
rect 133696 224936 133748 224942
rect 133696 224878 133748 224884
rect 133788 224936 133840 224942
rect 133788 224878 133840 224884
rect 133708 223922 133736 224878
rect 133972 224460 134024 224466
rect 133972 224402 134024 224408
rect 133696 223916 133748 223922
rect 133696 223858 133748 223864
rect 132512 221734 132894 221762
rect 133984 221748 134012 224402
rect 134984 224120 135036 224126
rect 134984 224062 135036 224068
rect 134996 221748 135024 224062
rect 136100 221748 136128 226986
rect 136468 224806 136496 320146
rect 136456 224800 136508 224806
rect 136456 224742 136508 224748
rect 136560 224466 136588 322918
rect 136548 224460 136600 224466
rect 136548 224402 136600 224408
rect 137940 224398 137968 322918
rect 138492 320210 138520 322932
rect 139504 320210 139532 322932
rect 140622 322918 140728 322946
rect 141726 322918 142108 322946
rect 142830 322918 143488 322946
rect 138480 320204 138532 320210
rect 138480 320146 138532 320152
rect 139308 320204 139360 320210
rect 139308 320146 139360 320152
rect 139492 320204 139544 320210
rect 139492 320146 139544 320152
rect 139320 228410 139348 320146
rect 140700 229770 140728 322918
rect 141424 320204 141476 320210
rect 141424 320146 141476 320152
rect 140688 229764 140740 229770
rect 140688 229706 140740 229712
rect 139308 228404 139360 228410
rect 139308 228346 139360 228352
rect 141436 226522 141464 320146
rect 141344 226494 141464 226522
rect 139400 224936 139452 224942
rect 139400 224878 139452 224884
rect 137192 224392 137244 224398
rect 137192 224334 137244 224340
rect 137928 224392 137980 224398
rect 137928 224334 137980 224340
rect 137204 221748 137232 224334
rect 138204 224324 138256 224330
rect 138204 224266 138256 224272
rect 138216 221748 138244 224266
rect 139412 224194 139440 224878
rect 139308 224188 139360 224194
rect 139308 224130 139360 224136
rect 139400 224188 139452 224194
rect 139400 224130 139452 224136
rect 139320 221748 139348 224130
rect 141344 224058 141372 226494
rect 142080 224330 142108 322918
rect 143460 231130 143488 322918
rect 143828 320210 143856 322932
rect 144932 320210 144960 322932
rect 146036 320822 146064 322932
rect 147062 322918 147628 322946
rect 146024 320816 146076 320822
rect 146024 320758 146076 320764
rect 143816 320204 143868 320210
rect 143816 320146 143868 320152
rect 144828 320204 144880 320210
rect 144828 320146 144880 320152
rect 144920 320204 144972 320210
rect 144920 320146 144972 320152
rect 146208 320204 146260 320210
rect 146208 320146 146260 320152
rect 143448 231124 143500 231130
rect 143448 231066 143500 231072
rect 144840 224942 144868 320146
rect 146220 232558 146248 320146
rect 146208 232552 146260 232558
rect 146208 232494 146260 232500
rect 147600 227050 147628 322918
rect 148152 320210 148180 322932
rect 149256 320210 149284 322932
rect 148140 320204 148192 320210
rect 148140 320146 148192 320152
rect 148968 320204 149020 320210
rect 148968 320146 149020 320152
rect 149244 320204 149296 320210
rect 149244 320146 149296 320152
rect 150256 320204 150308 320210
rect 150256 320146 150308 320152
rect 147588 227044 147640 227050
rect 147588 226986 147640 226992
rect 144828 224936 144880 224942
rect 144828 224878 144880 224884
rect 145748 224868 145800 224874
rect 145748 224810 145800 224816
rect 143540 224732 143592 224738
rect 143540 224674 143592 224680
rect 142528 224596 142580 224602
rect 142528 224538 142580 224544
rect 142068 224324 142120 224330
rect 142068 224266 142120 224272
rect 141424 224256 141476 224262
rect 141424 224198 141476 224204
rect 141332 224052 141384 224058
rect 141332 223994 141384 224000
rect 140320 223916 140372 223922
rect 140320 223858 140372 223864
rect 140332 221748 140360 223858
rect 141436 221748 141464 224198
rect 142540 221748 142568 224538
rect 143552 221748 143580 224674
rect 144644 224120 144696 224126
rect 144644 224062 144696 224068
rect 144656 221748 144684 224062
rect 145760 221748 145788 224810
rect 148980 224670 149008 320146
rect 149980 227112 150032 227118
rect 149980 227054 150032 227060
rect 147864 224664 147916 224670
rect 147864 224606 147916 224612
rect 148968 224664 149020 224670
rect 148968 224606 149020 224612
rect 146760 224528 146812 224534
rect 146760 224470 146812 224476
rect 146772 221748 146800 224470
rect 147876 221748 147904 224606
rect 148876 224188 148928 224194
rect 148876 224130 148928 224136
rect 148888 221748 148916 224130
rect 149992 221748 150020 227054
rect 150268 224602 150296 320146
rect 150256 224596 150308 224602
rect 150256 224538 150308 224544
rect 150360 224262 150388 322932
rect 151386 322918 151768 322946
rect 152490 322918 153148 322946
rect 151084 224800 151136 224806
rect 151084 224742 151136 224748
rect 150348 224256 150400 224262
rect 150348 224198 150400 224204
rect 151096 221748 151124 224742
rect 151740 224534 151768 322918
rect 152464 320816 152516 320822
rect 152464 320758 152516 320764
rect 152476 224874 152504 320758
rect 152464 224868 152516 224874
rect 152464 224810 152516 224816
rect 153120 224738 153148 322918
rect 153580 320210 153608 322932
rect 154684 320210 154712 322932
rect 155710 322918 155816 322946
rect 156814 322918 157288 322946
rect 153568 320204 153620 320210
rect 153568 320146 153620 320152
rect 154488 320204 154540 320210
rect 154488 320146 154540 320152
rect 154672 320204 154724 320210
rect 154672 320146 154724 320152
rect 154304 228404 154356 228410
rect 154304 228346 154356 228352
rect 153108 224732 153160 224738
rect 153108 224674 153160 224680
rect 151728 224528 151780 224534
rect 151728 224470 151780 224476
rect 152096 224460 152148 224466
rect 152096 224402 152148 224408
rect 152108 221748 152136 224402
rect 153200 224392 153252 224398
rect 153200 224334 153252 224340
rect 153212 221748 153240 224334
rect 154316 221748 154344 228346
rect 154500 224806 154528 320146
rect 155788 228410 155816 322918
rect 155868 320204 155920 320210
rect 155868 320146 155920 320152
rect 155776 228404 155828 228410
rect 155776 228346 155828 228352
rect 154488 224800 154540 224806
rect 154488 224742 154540 224748
rect 155880 224466 155908 320146
rect 155960 229764 156012 229770
rect 155960 229706 156012 229712
rect 155868 224460 155920 224466
rect 155868 224402 155920 224408
rect 155316 224052 155368 224058
rect 155316 223994 155368 224000
rect 155328 221748 155356 223994
rect 155972 221762 156000 229706
rect 157260 224126 157288 322918
rect 157904 320210 157932 322932
rect 158916 320210 158944 322932
rect 159928 322918 160034 322946
rect 161138 322918 161428 322946
rect 162242 322918 162808 322946
rect 157892 320204 157944 320210
rect 157892 320146 157944 320152
rect 158628 320204 158680 320210
rect 158628 320146 158680 320152
rect 158904 320204 158956 320210
rect 158904 320146 158956 320152
rect 157524 231124 157576 231130
rect 157524 231066 157576 231072
rect 157432 224324 157484 224330
rect 157432 224266 157484 224272
rect 157248 224120 157300 224126
rect 157248 224062 157300 224068
rect 155972 221734 156446 221762
rect 157444 221748 157472 224266
rect 157536 221626 157564 231066
rect 158640 224194 158668 320146
rect 159928 229770 159956 322918
rect 160008 320204 160060 320210
rect 160008 320146 160060 320152
rect 159916 229764 159968 229770
rect 159916 229706 159968 229712
rect 160020 224942 160048 320146
rect 160100 232552 160152 232558
rect 160100 232494 160152 232500
rect 159640 224936 159692 224942
rect 159640 224878 159692 224884
rect 160008 224936 160060 224942
rect 160008 224878 160060 224884
rect 158628 224188 158680 224194
rect 158628 224130 158680 224136
rect 159652 221748 159680 224878
rect 160112 221626 160140 232494
rect 161400 224330 161428 322918
rect 162780 227118 162808 322918
rect 163240 320278 163268 322932
rect 163228 320272 163280 320278
rect 163228 320214 163280 320220
rect 164344 320210 164372 322932
rect 165462 322918 165568 322946
rect 166474 322918 166948 322946
rect 167578 322918 168328 322946
rect 164332 320204 164384 320210
rect 164332 320146 164384 320152
rect 165436 320204 165488 320210
rect 165436 320146 165488 320152
rect 162768 227112 162820 227118
rect 162768 227054 162820 227060
rect 162860 227044 162912 227050
rect 162860 226986 162912 226992
rect 161756 224868 161808 224874
rect 161756 224810 161808 224816
rect 161388 224324 161440 224330
rect 161388 224266 161440 224272
rect 161768 221748 161796 224810
rect 162872 221748 162900 226986
rect 163872 224664 163924 224670
rect 163872 224606 163924 224612
rect 163884 221748 163912 224606
rect 165448 224602 165476 320146
rect 164976 224596 165028 224602
rect 164976 224538 165028 224544
rect 165436 224596 165488 224602
rect 165436 224538 165488 224544
rect 164988 221748 165016 224538
rect 165540 224398 165568 322918
rect 166920 231130 166948 322918
rect 167644 320272 167696 320278
rect 167644 320214 167696 320220
rect 166908 231124 166960 231130
rect 166908 231066 166960 231072
rect 167092 224528 167144 224534
rect 167092 224470 167144 224476
rect 165528 224392 165580 224398
rect 165528 224334 165580 224340
rect 166080 224256 166132 224262
rect 166080 224198 166132 224204
rect 166092 221748 166120 224198
rect 167104 221748 167132 224470
rect 167656 224058 167684 320214
rect 168196 224732 168248 224738
rect 168196 224674 168248 224680
rect 167644 224052 167696 224058
rect 167644 223994 167696 224000
rect 168208 221748 168236 224674
rect 168300 224534 168328 322918
rect 168668 320210 168696 322932
rect 169772 320210 169800 322932
rect 170798 322918 171088 322946
rect 171902 322918 172468 322946
rect 168656 320204 168708 320210
rect 168656 320146 168708 320152
rect 169668 320204 169720 320210
rect 169668 320146 169720 320152
rect 169760 320204 169812 320210
rect 169760 320146 169812 320152
rect 170956 320204 171008 320210
rect 170956 320146 171008 320152
rect 169680 224874 169708 320146
rect 169668 224868 169720 224874
rect 169668 224810 169720 224816
rect 169208 224800 169260 224806
rect 169208 224742 169260 224748
rect 168288 224528 168340 224534
rect 168288 224470 168340 224476
rect 169220 221748 169248 224742
rect 170968 224466 170996 320146
rect 170312 224460 170364 224466
rect 170312 224402 170364 224408
rect 170956 224460 171008 224466
rect 170956 224402 171008 224408
rect 170324 221748 170352 224402
rect 171060 224262 171088 322918
rect 171416 228404 171468 228410
rect 171416 228346 171468 228352
rect 171048 224256 171100 224262
rect 171048 224198 171100 224204
rect 171428 221748 171456 228346
rect 172440 224806 172468 322918
rect 172992 320210 173020 322932
rect 174004 320210 174032 322932
rect 172980 320204 173032 320210
rect 172980 320146 173032 320152
rect 173808 320204 173860 320210
rect 173808 320146 173860 320152
rect 173992 320204 174044 320210
rect 173992 320146 174044 320152
rect 172428 224800 172480 224806
rect 172428 224742 172480 224748
rect 173820 224194 173848 320146
rect 175108 228410 175136 322932
rect 176226 322918 176608 322946
rect 177330 322918 177988 322946
rect 175188 320204 175240 320210
rect 175188 320146 175240 320152
rect 175096 228404 175148 228410
rect 175096 228346 175148 228352
rect 174636 224936 174688 224942
rect 174636 224878 174688 224884
rect 173532 224188 173584 224194
rect 173532 224130 173584 224136
rect 173808 224188 173860 224194
rect 173808 224130 173860 224136
rect 172428 224120 172480 224126
rect 172428 224062 172480 224068
rect 172440 221748 172468 224062
rect 173544 221748 173572 224130
rect 174648 221748 174676 224878
rect 175200 224738 175228 320146
rect 175280 229764 175332 229770
rect 175280 229706 175332 229712
rect 175188 224732 175240 224738
rect 175188 224674 175240 224680
rect 175292 221762 175320 229706
rect 176580 224942 176608 322918
rect 177764 227112 177816 227118
rect 177764 227054 177816 227060
rect 176568 224936 176620 224942
rect 176568 224878 176620 224884
rect 176752 224324 176804 224330
rect 176752 224266 176804 224272
rect 175292 221734 175674 221762
rect 176764 221748 176792 224266
rect 177776 221748 177804 227054
rect 177960 224670 177988 322918
rect 178328 320210 178356 322932
rect 179432 320210 179460 322932
rect 180550 322918 180748 322946
rect 178316 320204 178368 320210
rect 178316 320146 178368 320152
rect 179328 320204 179380 320210
rect 179328 320146 179380 320152
rect 179420 320204 179472 320210
rect 179420 320146 179472 320152
rect 180616 320204 180668 320210
rect 180616 320146 180668 320152
rect 177948 224664 178000 224670
rect 177948 224606 178000 224612
rect 179340 224126 179368 320146
rect 180628 235278 180656 320146
rect 180616 235272 180668 235278
rect 180616 235214 180668 235220
rect 179972 224596 180024 224602
rect 179972 224538 180024 224544
rect 179328 224120 179380 224126
rect 179328 224062 179380 224068
rect 178868 224052 178920 224058
rect 178868 223994 178920 224000
rect 178880 221748 178908 223994
rect 179984 221748 180012 224538
rect 180720 224330 180748 322918
rect 181548 320278 181576 322932
rect 181536 320272 181588 320278
rect 181536 320214 181588 320220
rect 182652 320210 182680 322932
rect 183756 320210 183784 322932
rect 184860 320346 184888 322932
rect 185886 322918 186268 322946
rect 186990 322918 187648 322946
rect 188094 322918 188476 322946
rect 184848 320340 184900 320346
rect 184848 320282 184900 320288
rect 184204 320272 184256 320278
rect 184204 320214 184256 320220
rect 182640 320204 182692 320210
rect 182640 320146 182692 320152
rect 183468 320204 183520 320210
rect 183468 320146 183520 320152
rect 183744 320204 183796 320210
rect 183744 320146 183796 320152
rect 180892 231124 180944 231130
rect 180892 231066 180944 231072
rect 180904 224482 180932 231066
rect 183480 224534 183508 320146
rect 184216 224874 184244 320214
rect 184848 320204 184900 320210
rect 184848 320146 184900 320152
rect 183836 224868 183888 224874
rect 183836 224810 183888 224816
rect 184204 224868 184256 224874
rect 184204 224810 184256 224816
rect 183192 224528 183244 224534
rect 180904 224454 181668 224482
rect 183192 224470 183244 224476
rect 183468 224528 183520 224534
rect 183468 224470 183520 224476
rect 180984 224392 181036 224398
rect 180984 224334 181036 224340
rect 180708 224324 180760 224330
rect 180708 224266 180760 224272
rect 180996 221748 181024 224334
rect 181640 221626 181668 224454
rect 183204 221748 183232 224470
rect 183848 221762 183876 224810
rect 184020 224732 184072 224738
rect 184020 224674 184072 224680
rect 184032 224058 184060 224674
rect 184860 224602 184888 320146
rect 185584 315308 185636 315314
rect 185584 315250 185636 315256
rect 185596 274961 185624 315250
rect 185582 274952 185638 274961
rect 185582 274887 185638 274896
rect 184848 224596 184900 224602
rect 184848 224538 184900 224544
rect 186240 224466 186268 322918
rect 186964 320340 187016 320346
rect 186964 320282 187016 320288
rect 186976 224806 187004 320282
rect 186964 224800 187016 224806
rect 186964 224742 187016 224748
rect 187424 224732 187476 224738
rect 187424 224674 187476 224680
rect 185308 224460 185360 224466
rect 185308 224402 185360 224408
rect 186228 224460 186280 224466
rect 186228 224402 186280 224408
rect 184020 224052 184072 224058
rect 184020 223994 184072 224000
rect 183848 221734 184230 221762
rect 185320 221748 185348 224402
rect 186320 224256 186372 224262
rect 186320 224198 186372 224204
rect 186332 221748 186360 224198
rect 187436 221748 187464 224674
rect 187620 224398 187648 322918
rect 187608 224392 187660 224398
rect 187608 224334 187660 224340
rect 188448 224262 188476 322918
rect 189092 320385 189120 322932
rect 189078 320376 189134 320385
rect 189078 320311 189134 320320
rect 190196 320249 190224 322932
rect 191300 320249 191328 322932
rect 192404 320249 192432 322932
rect 193416 320385 193444 322932
rect 193402 320376 193458 320385
rect 193402 320311 193458 320320
rect 192484 320272 192536 320278
rect 190182 320240 190238 320249
rect 190182 320175 190238 320184
rect 191286 320240 191342 320249
rect 191286 320175 191342 320184
rect 192390 320240 192446 320249
rect 194520 320249 194548 322932
rect 192484 320214 192536 320220
rect 194506 320240 194562 320249
rect 192390 320175 192446 320184
rect 192392 318776 192444 318782
rect 192392 318718 192444 318724
rect 191196 318300 191248 318306
rect 191196 318242 191248 318248
rect 190000 318096 190052 318102
rect 190000 318038 190052 318044
rect 188620 317484 188672 317490
rect 188620 317426 188672 317432
rect 188632 315602 188660 317426
rect 190012 315602 190040 318038
rect 191208 315602 191236 318242
rect 192404 315602 192432 318718
rect 192496 317490 192524 320214
rect 194506 320175 194562 320184
rect 195624 319462 195652 322932
rect 195980 320476 196032 320482
rect 195980 320418 196032 320424
rect 195612 319456 195664 319462
rect 195612 319398 195664 319404
rect 194508 318504 194560 318510
rect 194508 318446 194560 318452
rect 193588 317892 193640 317898
rect 193588 317834 193640 317840
rect 192484 317484 192536 317490
rect 192484 317426 192536 317432
rect 193600 315602 193628 317834
rect 194520 315602 194548 318446
rect 195888 318368 195940 318374
rect 195888 318310 195940 318316
rect 195900 315602 195928 318310
rect 195992 318306 196020 320418
rect 196636 320278 196664 322932
rect 197372 322918 197754 322946
rect 196624 320272 196676 320278
rect 197372 320226 197400 322918
rect 198740 320884 198792 320890
rect 198740 320826 198792 320832
rect 196624 320214 196676 320220
rect 197280 320198 197400 320226
rect 197452 320204 197504 320210
rect 195980 318300 196032 318306
rect 195980 318242 196032 318248
rect 197280 318102 197308 320198
rect 197452 320146 197504 320152
rect 197464 318782 197492 320146
rect 197452 318776 197504 318782
rect 197452 318718 197504 318724
rect 198752 318510 198780 320826
rect 198844 320482 198872 322932
rect 198832 320476 198884 320482
rect 198832 320418 198884 320424
rect 198832 320340 198884 320346
rect 198832 320282 198884 320288
rect 198740 318504 198792 318510
rect 198740 318446 198792 318452
rect 198372 318164 198424 318170
rect 198372 318106 198424 318112
rect 197268 318096 197320 318102
rect 197268 318038 197320 318044
rect 197176 317552 197228 317558
rect 197176 317494 197228 317500
rect 197188 315602 197216 317494
rect 198384 315602 198412 318106
rect 198844 317898 198872 320282
rect 199948 320210 199976 322932
rect 200960 320346 200988 322932
rect 202064 320890 202092 322932
rect 202052 320884 202104 320890
rect 202052 320826 202104 320832
rect 202880 320544 202932 320550
rect 202880 320486 202932 320492
rect 200948 320340 201000 320346
rect 200948 320282 201000 320288
rect 202144 320272 202196 320278
rect 202144 320214 202196 320220
rect 199936 320204 199988 320210
rect 199936 320146 199988 320152
rect 201132 320204 201184 320210
rect 201132 320146 201184 320152
rect 200764 318708 200816 318714
rect 200764 318650 200816 318656
rect 199568 318300 199620 318306
rect 199568 318242 199620 318248
rect 198832 317892 198884 317898
rect 198832 317834 198884 317840
rect 199580 315602 199608 318242
rect 200776 315602 200804 318650
rect 201144 318374 201172 320146
rect 201960 318776 202012 318782
rect 201960 318718 202012 318724
rect 201132 318368 201184 318374
rect 201132 318310 201184 318316
rect 201972 315602 202000 318718
rect 202156 317558 202184 320214
rect 202788 318640 202840 318646
rect 202788 318582 202840 318588
rect 202144 317552 202196 317558
rect 202144 317494 202196 317500
rect 188600 315574 188660 315602
rect 189704 315574 190040 315602
rect 190900 315574 191236 315602
rect 192096 315574 192432 315602
rect 193292 315574 193628 315602
rect 194488 315574 194548 315602
rect 195684 315574 195928 315602
rect 196880 315574 197216 315602
rect 198076 315574 198412 315602
rect 199272 315574 199608 315602
rect 200468 315574 200804 315602
rect 201664 315574 202000 315602
rect 202800 315602 202828 318582
rect 202892 318170 202920 320486
rect 203168 320210 203196 322932
rect 204180 320278 204208 322932
rect 204260 320612 204312 320618
rect 204260 320554 204312 320560
rect 204168 320272 204220 320278
rect 204168 320214 204220 320220
rect 203156 320204 203208 320210
rect 203156 320146 203208 320152
rect 204168 318368 204220 318374
rect 204168 318310 204220 318316
rect 202880 318164 202932 318170
rect 202880 318106 202932 318112
rect 204180 315602 204208 318310
rect 204272 318306 204300 320554
rect 205284 320550 205312 322932
rect 206388 320618 206416 322932
rect 207032 322918 207506 322946
rect 208412 322918 208518 322946
rect 206376 320612 206428 320618
rect 206376 320554 206428 320560
rect 205272 320544 205324 320550
rect 205272 320486 205324 320492
rect 207032 320192 207060 322918
rect 208412 320770 208440 322918
rect 208320 320742 208440 320770
rect 206940 320164 207060 320192
rect 207112 320204 207164 320210
rect 206940 318714 206968 320164
rect 207112 320146 207164 320152
rect 206928 318708 206980 318714
rect 206928 318650 206980 318656
rect 207124 318646 207152 320146
rect 208320 318782 208348 320742
rect 208400 320612 208452 320618
rect 208400 320554 208452 320560
rect 208308 318776 208360 318782
rect 208308 318718 208360 318724
rect 207112 318640 207164 318646
rect 207112 318582 207164 318588
rect 208412 318374 208440 320554
rect 209608 320210 209636 322932
rect 210712 320618 210740 322932
rect 211172 322918 211738 322946
rect 212552 322918 212842 322946
rect 210700 320612 210752 320618
rect 210700 320554 210752 320560
rect 211172 320226 211200 322918
rect 212552 320226 212580 322918
rect 213932 320226 213960 322932
rect 209596 320204 209648 320210
rect 209596 320146 209648 320152
rect 211080 320198 211200 320226
rect 212460 320198 212580 320226
rect 213840 320198 213960 320226
rect 209136 318504 209188 318510
rect 209136 318446 209188 318452
rect 208400 318368 208452 318374
rect 208400 318310 208452 318316
rect 204260 318300 204312 318306
rect 204260 318242 204312 318248
rect 207940 318232 207992 318238
rect 207940 318174 207992 318180
rect 206744 317620 206796 317626
rect 206744 317562 206796 317568
rect 205548 317552 205600 317558
rect 205548 317494 205600 317500
rect 205560 315602 205588 317494
rect 206756 315602 206784 317562
rect 207952 315602 207980 318174
rect 209148 315602 209176 318446
rect 210332 317756 210384 317762
rect 210332 317698 210384 317704
rect 210344 315602 210372 317698
rect 211080 317558 211108 320198
rect 211528 318776 211580 318782
rect 211528 318718 211580 318724
rect 211068 317552 211120 317558
rect 211068 317494 211120 317500
rect 211540 315602 211568 318718
rect 212460 317626 212488 320198
rect 213840 318238 213868 320198
rect 215036 318510 215064 322932
rect 215024 318504 215076 318510
rect 215024 318446 215076 318452
rect 213828 318232 213880 318238
rect 213828 318174 213880 318180
rect 213828 317960 213880 317966
rect 213828 317902 213880 317908
rect 212448 317620 212500 317626
rect 212448 317562 212500 317568
rect 212448 317484 212500 317490
rect 212448 317426 212500 317432
rect 212460 315602 212488 317426
rect 213840 315602 213868 317902
rect 216048 317762 216076 322932
rect 217152 318782 217180 322932
rect 218072 322918 218270 322946
rect 218072 320226 218100 322918
rect 217980 320198 218100 320226
rect 217140 318776 217192 318782
rect 217140 318718 217192 318724
rect 217508 318300 217560 318306
rect 217508 318242 217560 318248
rect 216036 317756 216088 317762
rect 216036 317698 216088 317704
rect 216312 317620 216364 317626
rect 216312 317562 216364 317568
rect 215116 317484 215168 317490
rect 215116 317426 215168 317432
rect 215128 315602 215156 317426
rect 216324 315602 216352 317562
rect 217520 315602 217548 318242
rect 217980 317558 218008 320198
rect 218704 318096 218756 318102
rect 218704 318038 218756 318044
rect 217968 317552 218020 317558
rect 217968 317494 218020 317500
rect 218716 315602 218744 318038
rect 219268 317966 219296 322932
rect 219900 320204 219952 320210
rect 219900 320146 219952 320152
rect 219256 317960 219308 317966
rect 219256 317902 219308 317908
rect 219912 315602 219940 320146
rect 220372 317490 220400 322932
rect 220636 318708 220688 318714
rect 220636 318650 220688 318656
rect 220360 317484 220412 317490
rect 220360 317426 220412 317432
rect 202800 315574 202860 315602
rect 204056 315574 204208 315602
rect 205252 315574 205588 315602
rect 206448 315574 206784 315602
rect 207644 315574 207980 315602
rect 208840 315574 209176 315602
rect 210036 315574 210372 315602
rect 211232 315574 211568 315602
rect 212428 315574 212488 315602
rect 213624 315574 213868 315602
rect 214820 315574 215156 315602
rect 216016 315574 216352 315602
rect 217212 315574 217548 315602
rect 218408 315574 218744 315602
rect 219604 315574 219940 315602
rect 220648 315602 220676 318650
rect 221476 317626 221504 322932
rect 222580 318306 222608 322932
rect 223488 318776 223540 318782
rect 223488 318718 223540 318724
rect 222568 318300 222620 318306
rect 222568 318242 222620 318248
rect 222016 317960 222068 317966
rect 222016 317902 222068 317908
rect 221464 317620 221516 317626
rect 221464 317562 221516 317568
rect 222028 315602 222056 317902
rect 223500 315602 223528 318718
rect 223592 318102 223620 322932
rect 224696 320210 224724 322932
rect 224684 320204 224736 320210
rect 224684 320146 224736 320152
rect 224868 320204 224920 320210
rect 224868 320146 224920 320152
rect 223580 318096 223632 318102
rect 223580 318038 223632 318044
rect 220648 315574 220800 315602
rect 221996 315574 222056 315602
rect 223192 315574 223528 315602
rect 224880 315466 224908 320146
rect 225800 318714 225828 322932
rect 226248 320680 226300 320686
rect 226248 320622 226300 320628
rect 225788 318708 225840 318714
rect 225788 318650 225840 318656
rect 226260 315602 226288 320622
rect 226812 317966 226840 322932
rect 227076 320816 227128 320822
rect 227076 320758 227128 320764
rect 226800 317960 226852 317966
rect 226800 317902 226852 317908
rect 227088 315602 227116 320758
rect 227916 318782 227944 322932
rect 228272 321088 228324 321094
rect 228272 321030 228324 321036
rect 227904 318776 227956 318782
rect 227904 318718 227956 318724
rect 228284 315602 228312 321030
rect 229020 320210 229048 322932
rect 230124 320686 230152 322932
rect 231136 320822 231164 322932
rect 231768 321156 231820 321162
rect 231768 321098 231820 321104
rect 231124 320816 231176 320822
rect 231124 320758 231176 320764
rect 230112 320680 230164 320686
rect 230112 320622 230164 320628
rect 229284 320340 229336 320346
rect 229284 320282 229336 320288
rect 229008 320204 229060 320210
rect 229008 320146 229060 320152
rect 229296 315602 229324 320282
rect 230296 320204 230348 320210
rect 230296 320146 230348 320152
rect 226076 315574 226288 315602
rect 226780 315574 227116 315602
rect 227976 315574 228312 315602
rect 229172 315574 229324 315602
rect 230308 315602 230336 320146
rect 231780 315602 231808 321098
rect 232240 321094 232268 322932
rect 232228 321088 232280 321094
rect 232228 321030 232280 321036
rect 233344 320346 233372 322932
rect 233332 320340 233384 320346
rect 233332 320282 233384 320288
rect 233148 320272 233200 320278
rect 233148 320214 233200 320220
rect 233160 315602 233188 320214
rect 234356 320210 234384 322932
rect 235460 321162 235488 322932
rect 235448 321156 235500 321162
rect 235448 321098 235500 321104
rect 235448 320476 235500 320482
rect 235448 320418 235500 320424
rect 234344 320204 234396 320210
rect 234344 320146 234396 320152
rect 234528 320204 234580 320210
rect 234528 320146 234580 320152
rect 230308 315574 230368 315602
rect 231564 315574 231808 315602
rect 232760 315574 233188 315602
rect 226076 315466 226104 315574
rect 234540 315466 234568 320146
rect 235460 315602 235488 320418
rect 236564 320278 236592 322932
rect 236644 320408 236696 320414
rect 236644 320350 236696 320356
rect 236552 320272 236604 320278
rect 236552 320214 236604 320220
rect 236656 315602 236684 320350
rect 237668 320210 237696 322932
rect 238680 320482 238708 322932
rect 238668 320476 238720 320482
rect 238668 320418 238720 320424
rect 239784 320414 239812 322932
rect 239772 320408 239824 320414
rect 239772 320350 239824 320356
rect 238668 320340 238720 320346
rect 238668 320282 238720 320288
rect 237840 320272 237892 320278
rect 237840 320214 237892 320220
rect 237656 320204 237708 320210
rect 237656 320146 237708 320152
rect 237852 315602 237880 320214
rect 235152 315574 235488 315602
rect 236348 315574 236684 315602
rect 237544 315574 237880 315602
rect 238680 315602 238708 320282
rect 240888 320278 240916 322932
rect 241900 320346 241928 322932
rect 241888 320340 241940 320346
rect 241888 320282 241940 320288
rect 242624 320340 242676 320346
rect 242624 320282 242676 320288
rect 240876 320272 240928 320278
rect 240876 320214 240928 320220
rect 241428 320272 241480 320278
rect 241428 320214 241480 320220
rect 240048 320204 240100 320210
rect 240048 320146 240100 320152
rect 240060 315602 240088 320146
rect 241440 315602 241468 320214
rect 242636 315602 242664 320282
rect 243004 320210 243032 322932
rect 244108 320278 244136 322932
rect 245212 320346 245240 322932
rect 246120 320816 246172 320822
rect 246120 320758 246172 320764
rect 245200 320340 245252 320346
rect 245200 320282 245252 320288
rect 244096 320272 244148 320278
rect 244096 320214 244148 320220
rect 245016 320272 245068 320278
rect 245016 320214 245068 320220
rect 242992 320204 243044 320210
rect 242992 320146 243044 320152
rect 243820 320204 243872 320210
rect 243820 320146 243872 320152
rect 243832 315602 243860 320146
rect 245028 315602 245056 320214
rect 246132 318458 246160 320758
rect 246224 320210 246252 322932
rect 247328 320278 247356 322932
rect 247408 320884 247460 320890
rect 247408 320826 247460 320832
rect 247316 320272 247368 320278
rect 247316 320214 247368 320220
rect 246212 320204 246264 320210
rect 246212 320146 246264 320152
rect 246132 318430 246252 318458
rect 246224 315602 246252 318430
rect 247420 315602 247448 320826
rect 248432 320822 248460 322932
rect 249444 320890 249472 322932
rect 249432 320884 249484 320890
rect 249432 320826 249484 320832
rect 248420 320816 248472 320822
rect 248420 320758 248472 320764
rect 250548 320754 250576 322932
rect 248328 320748 248380 320754
rect 248328 320690 248380 320696
rect 250536 320748 250588 320754
rect 250536 320690 250588 320696
rect 248340 315602 248368 320690
rect 251088 320272 251140 320278
rect 251088 320214 251140 320220
rect 249708 320204 249760 320210
rect 249708 320146 249760 320152
rect 249720 315602 249748 320146
rect 251100 315602 251128 320214
rect 251652 320210 251680 322932
rect 252756 320278 252784 322932
rect 253388 320340 253440 320346
rect 253388 320282 253440 320288
rect 252744 320272 252796 320278
rect 252744 320214 252796 320220
rect 251640 320204 251692 320210
rect 251640 320146 251692 320152
rect 252468 320204 252520 320210
rect 252468 320146 252520 320152
rect 238680 315574 238740 315602
rect 239936 315574 240088 315602
rect 241132 315574 241468 315602
rect 242328 315574 242664 315602
rect 243524 315574 243860 315602
rect 244720 315574 245056 315602
rect 245916 315574 246252 315602
rect 247112 315574 247448 315602
rect 248308 315574 248368 315602
rect 249504 315574 249748 315602
rect 250700 315574 251128 315602
rect 252480 315466 252508 320146
rect 253400 315602 253428 320282
rect 253768 320210 253796 322932
rect 254872 320346 254900 322932
rect 254860 320340 254912 320346
rect 254860 320282 254912 320288
rect 255976 320278 256004 322932
rect 256516 320816 256568 320822
rect 256516 320758 256568 320764
rect 254584 320272 254636 320278
rect 254584 320214 254636 320220
rect 255964 320272 256016 320278
rect 255964 320214 256016 320220
rect 253756 320204 253808 320210
rect 253756 320146 253808 320152
rect 254596 315602 254624 320214
rect 255780 320204 255832 320210
rect 255780 320146 255832 320152
rect 255792 315602 255820 320146
rect 253092 315574 253428 315602
rect 254288 315574 254624 315602
rect 255484 315574 255820 315602
rect 256528 315602 256556 320758
rect 256988 320210 257016 322932
rect 258092 320822 258120 322932
rect 258080 320816 258132 320822
rect 258080 320758 258132 320764
rect 259196 320278 259224 322932
rect 257988 320272 258040 320278
rect 257988 320214 258040 320220
rect 259184 320272 259236 320278
rect 259184 320214 259236 320220
rect 256976 320204 257028 320210
rect 256976 320146 257028 320152
rect 258000 315602 258028 320214
rect 260300 320210 260328 322932
rect 260852 322918 261326 322946
rect 262232 322918 262430 322946
rect 259368 320204 259420 320210
rect 259368 320146 259420 320152
rect 260288 320204 260340 320210
rect 260852 320192 260880 322918
rect 262232 320192 262260 322918
rect 263520 320210 263548 322932
rect 264532 320210 264560 322932
rect 264992 322918 265650 322946
rect 266372 322918 266754 322946
rect 267752 322918 267858 322946
rect 260288 320146 260340 320152
rect 260760 320164 260880 320192
rect 262140 320164 262260 320192
rect 263508 320204 263560 320210
rect 259380 315602 259408 320146
rect 256528 315574 256680 315602
rect 257876 315574 258028 315602
rect 259072 315574 259408 315602
rect 260760 315466 260788 320164
rect 262140 315466 262168 320164
rect 263508 320146 263560 320152
rect 263600 320204 263652 320210
rect 263600 320146 263652 320152
rect 264520 320204 264572 320210
rect 264520 320146 264572 320152
rect 262220 320068 262272 320074
rect 262220 320010 262272 320016
rect 262232 315602 262260 320010
rect 263612 315602 263640 320146
rect 264992 315602 265020 322918
rect 266372 320192 266400 322918
rect 267752 320872 267780 322918
rect 266280 320164 266400 320192
rect 267660 320844 267780 320872
rect 266280 315602 266308 320164
rect 267660 315602 267688 320844
rect 268856 320210 268884 322932
rect 269960 320210 269988 322932
rect 270512 322918 271078 322946
rect 271892 322918 272090 322946
rect 267740 320204 267792 320210
rect 267740 320146 267792 320152
rect 268844 320204 268896 320210
rect 268844 320146 268896 320152
rect 269120 320204 269172 320210
rect 269120 320146 269172 320152
rect 269948 320204 270000 320210
rect 269948 320146 270000 320152
rect 262232 315574 262660 315602
rect 263612 315574 263856 315602
rect 264992 315574 265052 315602
rect 266248 315574 266308 315602
rect 267444 315574 267688 315602
rect 224388 315438 224908 315466
rect 225584 315438 226104 315466
rect 233956 315438 234568 315466
rect 251896 315438 252508 315466
rect 260268 315438 260788 315466
rect 261464 315438 262168 315466
rect 267752 315466 267780 320146
rect 269132 315466 269160 320146
rect 270512 315466 270540 322918
rect 271892 315602 271920 322918
rect 273180 320226 273208 322932
rect 273180 320198 273392 320226
rect 273364 315602 273392 320198
rect 274284 315602 274312 322932
rect 275388 315602 275416 322932
rect 276032 322918 276414 322946
rect 277412 322918 277518 322946
rect 278622 322918 278728 322946
rect 276032 315738 276060 322918
rect 277412 315738 277440 322918
rect 278700 320226 278728 322918
rect 278700 320198 278820 320226
rect 276032 315710 276520 315738
rect 277412 315710 277716 315738
rect 271892 315574 272228 315602
rect 273364 315574 273424 315602
rect 274284 315574 274620 315602
rect 275388 315574 275816 315602
rect 276492 315466 276520 315710
rect 277688 315466 277716 315710
rect 278792 315466 278820 320198
rect 280160 319456 280212 319462
rect 280160 319398 280212 319404
rect 267752 315438 268640 315466
rect 269132 315438 269836 315466
rect 270512 315438 271032 315466
rect 276492 315438 277012 315466
rect 277688 315438 278208 315466
rect 278792 315438 279404 315466
rect 280172 295905 280200 319398
rect 282196 305658 282224 335951
rect 282288 322153 282316 700266
rect 283944 698290 283972 703446
rect 332520 700602 332548 703520
rect 348804 700641 348832 703520
rect 348790 700632 348846 700641
rect 287704 700596 287756 700602
rect 287704 700538 287756 700544
rect 332508 700596 332560 700602
rect 348790 700567 348846 700576
rect 332508 700538 332560 700544
rect 283288 698284 283340 698290
rect 283288 698226 283340 698232
rect 283932 698284 283984 698290
rect 283932 698226 283984 698232
rect 283300 694142 283328 698226
rect 283104 694136 283156 694142
rect 283104 694078 283156 694084
rect 283288 694136 283340 694142
rect 283288 694078 283340 694084
rect 283116 684554 283144 694078
rect 283012 684548 283064 684554
rect 283012 684490 283064 684496
rect 283104 684548 283156 684554
rect 283104 684490 283156 684496
rect 283024 684457 283052 684490
rect 283010 684448 283066 684457
rect 283010 684383 283066 684392
rect 283102 678872 283158 678881
rect 283102 678807 283158 678816
rect 283116 666602 283144 678807
rect 283104 666596 283156 666602
rect 283104 666538 283156 666544
rect 283380 666596 283432 666602
rect 283380 666538 283432 666544
rect 283392 661774 283420 666538
rect 283104 661768 283156 661774
rect 283104 661710 283156 661716
rect 283380 661768 283432 661774
rect 283380 661710 283432 661716
rect 283116 656946 283144 661710
rect 283104 656940 283156 656946
rect 283104 656882 283156 656888
rect 283196 656940 283248 656946
rect 283196 656882 283248 656888
rect 283208 647290 283236 656882
rect 283104 647284 283156 647290
rect 283104 647226 283156 647232
rect 283196 647284 283248 647290
rect 283196 647226 283248 647232
rect 283116 640422 283144 647226
rect 283104 640416 283156 640422
rect 283104 640358 283156 640364
rect 283196 640416 283248 640422
rect 283196 640358 283248 640364
rect 283208 630698 283236 640358
rect 282920 630692 282972 630698
rect 282920 630634 282972 630640
rect 283196 630692 283248 630698
rect 283196 630634 283248 630640
rect 282932 625954 282960 630634
rect 282932 625926 283236 625954
rect 283012 621716 283064 621722
rect 283012 621658 283064 621664
rect 282920 611380 282972 611386
rect 282920 611322 282972 611328
rect 282932 592006 282960 611322
rect 282920 592000 282972 592006
rect 282920 591942 282972 591948
rect 283024 585993 283052 621658
rect 283208 621058 283236 625926
rect 283208 621030 283328 621058
rect 283300 611386 283328 621030
rect 284300 618928 284352 618934
rect 284300 618870 284352 618876
rect 283288 611380 283340 611386
rect 283288 611322 283340 611328
rect 283196 592000 283248 592006
rect 283196 591942 283248 591948
rect 283010 585984 283066 585993
rect 283010 585919 283066 585928
rect 283208 582486 283236 591942
rect 283196 582480 283248 582486
rect 283196 582422 283248 582428
rect 283196 582344 283248 582350
rect 283196 582286 283248 582292
rect 283208 572762 283236 582286
rect 283196 572756 283248 572762
rect 283196 572698 283248 572704
rect 283196 572620 283248 572626
rect 283196 572562 283248 572568
rect 283208 568585 283236 572562
rect 283194 568576 283250 568585
rect 283194 568511 283250 568520
rect 283378 568576 283434 568585
rect 283378 568511 283434 568520
rect 283392 558958 283420 568511
rect 283196 558952 283248 558958
rect 283196 558894 283248 558900
rect 283380 558952 283432 558958
rect 283380 558894 283432 558900
rect 283208 553450 283236 558894
rect 283196 553444 283248 553450
rect 283196 553386 283248 553392
rect 283288 553308 283340 553314
rect 283288 553250 283340 553256
rect 283300 543862 283328 553250
rect 283288 543856 283340 543862
rect 283288 543798 283340 543804
rect 283104 543720 283156 543726
rect 283104 543662 283156 543668
rect 282828 528012 282880 528018
rect 282828 527954 282880 527960
rect 282840 527542 282868 527954
rect 282828 527536 282880 527542
rect 282828 527478 282880 527484
rect 283116 527134 283144 543662
rect 282828 527128 282880 527134
rect 282828 527070 282880 527076
rect 283104 527128 283156 527134
rect 283104 527070 283156 527076
rect 282840 519330 282868 527070
rect 282840 519302 283052 519330
rect 283024 512038 283052 519302
rect 283012 512032 283064 512038
rect 282918 512000 282974 512009
rect 283104 512032 283156 512038
rect 283012 511974 283064 511980
rect 283102 512000 283104 512009
rect 283156 512000 283158 512009
rect 282918 511935 282974 511944
rect 283102 511935 283158 511944
rect 282932 502382 282960 511935
rect 282920 502376 282972 502382
rect 282920 502318 282972 502324
rect 283196 502376 283248 502382
rect 283196 502318 283248 502324
rect 283208 495394 283236 502318
rect 283024 495366 283236 495394
rect 283024 485858 283052 495366
rect 283012 485852 283064 485858
rect 283012 485794 283064 485800
rect 283104 485784 283156 485790
rect 283104 485726 283156 485732
rect 283116 483002 283144 485726
rect 283104 482996 283156 483002
rect 283104 482938 283156 482944
rect 283288 482996 283340 483002
rect 283288 482938 283340 482944
rect 283300 473414 283328 482938
rect 283012 473408 283064 473414
rect 283012 473350 283064 473356
rect 283288 473408 283340 473414
rect 283288 473350 283340 473356
rect 283024 473278 283052 473350
rect 283012 473272 283064 473278
rect 283012 473214 283064 473220
rect 283196 473272 283248 473278
rect 283196 473214 283248 473220
rect 283208 454073 283236 473214
rect 282918 454064 282974 454073
rect 282918 453999 282974 454008
rect 283194 454064 283250 454073
rect 283194 453999 283250 454008
rect 282932 447166 282960 453999
rect 282920 447160 282972 447166
rect 282920 447102 282972 447108
rect 283012 447092 283064 447098
rect 283012 447034 283064 447040
rect 283024 444378 283052 447034
rect 282736 444372 282788 444378
rect 282736 444314 282788 444320
rect 283012 444372 283064 444378
rect 283012 444314 283064 444320
rect 282748 434761 282776 444314
rect 282734 434752 282790 434761
rect 282734 434687 282790 434696
rect 282918 434752 282974 434761
rect 282918 434687 282974 434696
rect 282932 427854 282960 434687
rect 282920 427848 282972 427854
rect 282920 427790 282972 427796
rect 283012 427780 283064 427786
rect 283012 427722 283064 427728
rect 283024 418146 283052 427722
rect 283024 418118 283144 418146
rect 283116 415410 283144 418118
rect 282920 415404 282972 415410
rect 282920 415346 282972 415352
rect 283104 415404 283156 415410
rect 283104 415346 283156 415352
rect 282932 405754 282960 415346
rect 282920 405748 282972 405754
rect 282920 405690 282972 405696
rect 283196 405748 283248 405754
rect 283196 405690 283248 405696
rect 283208 403617 283236 405690
rect 283194 403608 283250 403617
rect 283194 403543 283250 403552
rect 284312 369617 284340 618870
rect 284390 608832 284446 608841
rect 284390 608767 284446 608776
rect 284404 569906 284432 608767
rect 284392 569900 284444 569906
rect 284392 569842 284444 569848
rect 286324 569220 286376 569226
rect 286324 569162 286376 569168
rect 284390 392728 284446 392737
rect 284390 392663 284446 392672
rect 284404 377262 284432 392663
rect 284392 377256 284444 377262
rect 284392 377198 284444 377204
rect 284298 369608 284354 369617
rect 284298 369543 284354 369552
rect 282274 322144 282330 322153
rect 282274 322079 282330 322088
rect 282184 305652 282236 305658
rect 282184 305594 282236 305600
rect 280158 295896 280214 295905
rect 280158 295831 280214 295840
rect 282196 254017 282224 305594
rect 281538 254008 281594 254017
rect 281538 253943 281594 253952
rect 282182 254008 282238 254017
rect 282182 253943 282238 253952
rect 281552 235958 281580 253943
rect 281540 235952 281592 235958
rect 281540 235894 281592 235900
rect 194600 235272 194652 235278
rect 194600 235214 194652 235220
rect 235262 235240 235318 235249
rect 190644 228404 190696 228410
rect 190644 228346 190696 228352
rect 188436 224256 188488 224262
rect 188436 224198 188488 224204
rect 188528 224188 188580 224194
rect 188528 224130 188580 224136
rect 188540 221748 188568 224130
rect 189540 224052 189592 224058
rect 189540 223994 189592 224000
rect 189552 221748 189580 223994
rect 190656 221748 190684 228346
rect 191748 224936 191800 224942
rect 191748 224878 191800 224884
rect 191760 221748 191788 224878
rect 192760 224664 192812 224670
rect 192760 224606 192812 224612
rect 192772 221748 192800 224606
rect 193864 224120 193916 224126
rect 193864 224062 193916 224068
rect 193876 221748 193904 224062
rect 194612 221762 194640 235214
rect 235262 235175 235318 235184
rect 227628 232552 227680 232558
rect 227628 232494 227680 232500
rect 214748 231124 214800 231130
rect 214748 231066 214800 231072
rect 214564 229764 214616 229770
rect 214564 229706 214616 229712
rect 207754 224904 207810 224913
rect 197084 224868 197136 224874
rect 207754 224839 207810 224848
rect 197084 224810 197136 224816
rect 195980 224324 196032 224330
rect 195980 224266 196032 224272
rect 194612 221734 194902 221762
rect 195992 221748 196020 224266
rect 197096 221748 197124 224810
rect 200304 224800 200356 224806
rect 200304 224742 200356 224748
rect 199200 224596 199252 224602
rect 199200 224538 199252 224544
rect 198096 224528 198148 224534
rect 198096 224470 198148 224476
rect 198108 221748 198136 224470
rect 199212 221748 199240 224538
rect 200316 221748 200344 224742
rect 206650 224632 206706 224641
rect 206650 224567 206706 224576
rect 204534 224496 204590 224505
rect 201316 224460 201368 224466
rect 204534 224431 204590 224440
rect 201316 224402 201368 224408
rect 201328 221748 201356 224402
rect 202420 224392 202472 224398
rect 202420 224334 202472 224340
rect 202432 221748 202460 224334
rect 203432 224256 203484 224262
rect 203432 224198 203484 224204
rect 203444 221748 203472 224198
rect 204548 221748 204576 224431
rect 205638 224360 205694 224369
rect 205638 224295 205694 224304
rect 205652 221748 205680 224295
rect 206664 221748 206692 224567
rect 207768 221748 207796 224839
rect 208858 224768 208914 224777
rect 208858 224703 208914 224712
rect 208872 221748 208900 224703
rect 210976 224256 211028 224262
rect 209870 224224 209926 224233
rect 210976 224198 211028 224204
rect 209870 224159 209926 224168
rect 209884 221748 209912 224159
rect 210988 221748 211016 224198
rect 121564 221598 122222 221626
rect 129200 221598 129674 221626
rect 157536 221598 158562 221626
rect 160112 221598 160678 221626
rect 181640 221598 182114 221626
rect 120724 221536 120776 221542
rect 120776 221484 121118 221490
rect 120724 221478 121118 221484
rect 120736 221462 121118 221478
rect 116676 220108 116728 220114
rect 116676 220050 116728 220056
rect 116688 130121 116716 220050
rect 214380 213852 214432 213858
rect 214380 213794 214432 213800
rect 214392 212673 214420 213794
rect 214378 212664 214434 212673
rect 214378 212599 214434 212608
rect 214196 211132 214248 211138
rect 214196 211074 214248 211080
rect 214208 210361 214236 211074
rect 214194 210352 214250 210361
rect 214194 210287 214250 210296
rect 214196 209704 214248 209710
rect 214196 209646 214248 209652
rect 214208 208865 214236 209646
rect 214194 208856 214250 208865
rect 214194 208791 214250 208800
rect 214288 208276 214340 208282
rect 214288 208218 214340 208224
rect 214300 207233 214328 208218
rect 214286 207224 214342 207233
rect 214286 207159 214342 207168
rect 214380 206916 214432 206922
rect 214380 206858 214432 206864
rect 214392 205737 214420 206858
rect 214378 205728 214434 205737
rect 214378 205663 214434 205672
rect 214288 202836 214340 202842
rect 214288 202778 214340 202784
rect 214300 201793 214328 202778
rect 214286 201784 214342 201793
rect 214286 201719 214342 201728
rect 214380 201476 214432 201482
rect 214380 201418 214432 201424
rect 214392 200977 214420 201418
rect 214378 200968 214434 200977
rect 214378 200903 214434 200912
rect 214104 200116 214156 200122
rect 214104 200058 214156 200064
rect 214116 199345 214144 200058
rect 214102 199336 214158 199345
rect 214102 199271 214158 199280
rect 214104 198620 214156 198626
rect 214104 198562 214156 198568
rect 214116 197849 214144 198562
rect 214102 197840 214158 197849
rect 214102 197775 214158 197784
rect 214380 197328 214432 197334
rect 214380 197270 214432 197276
rect 214392 196217 214420 197270
rect 214378 196208 214434 196217
rect 214378 196143 214434 196152
rect 214288 191820 214340 191826
rect 214288 191762 214340 191768
rect 214300 190777 214328 191762
rect 214286 190768 214342 190777
rect 214286 190703 214342 190712
rect 214380 190460 214432 190466
rect 214380 190402 214432 190408
rect 214392 189281 214420 190402
rect 214378 189272 214434 189281
rect 214378 189207 214434 189216
rect 214012 189032 214064 189038
rect 214012 188974 214064 188980
rect 214024 188465 214052 188974
rect 214010 188456 214066 188465
rect 214010 188391 214066 188400
rect 214472 185700 214524 185706
rect 214472 185642 214524 185648
rect 213920 185564 213972 185570
rect 213920 185506 213972 185512
rect 213932 185337 213960 185506
rect 213918 185328 213974 185337
rect 213918 185263 213974 185272
rect 214196 184816 214248 184822
rect 214196 184758 214248 184764
rect 214208 183705 214236 184758
rect 214484 184521 214512 185642
rect 214470 184512 214526 184521
rect 214470 184447 214526 184456
rect 214194 183696 214250 183705
rect 214194 183631 214250 183640
rect 214196 182164 214248 182170
rect 214196 182106 214248 182112
rect 214208 181393 214236 182106
rect 214194 181384 214250 181393
rect 214194 181319 214250 181328
rect 214012 180804 214064 180810
rect 214012 180746 214064 180752
rect 214024 179761 214052 180746
rect 214102 180568 214158 180577
rect 214102 180503 214158 180512
rect 214116 179790 214144 180503
rect 214104 179784 214156 179790
rect 214010 179752 214066 179761
rect 214104 179726 214156 179732
rect 214010 179687 214066 179696
rect 213920 179240 213972 179246
rect 213920 179182 213972 179188
rect 213932 179081 213960 179182
rect 213918 179072 213974 179081
rect 213918 179007 213974 179016
rect 214104 178628 214156 178634
rect 214104 178570 214156 178576
rect 214116 178265 214144 178570
rect 214102 178256 214158 178265
rect 214102 178191 214158 178200
rect 214104 175228 214156 175234
rect 214104 175170 214156 175176
rect 214116 174321 214144 175170
rect 214102 174312 214158 174321
rect 214102 174247 214158 174256
rect 214288 173868 214340 173874
rect 214288 173810 214340 173816
rect 214300 172825 214328 173810
rect 214286 172816 214342 172825
rect 214286 172751 214342 172760
rect 214288 172508 214340 172514
rect 214288 172450 214340 172456
rect 214300 172009 214328 172450
rect 214286 172000 214342 172009
rect 214286 171935 214342 171944
rect 213920 168088 213972 168094
rect 213918 168056 213920 168065
rect 213972 168056 213974 168065
rect 213918 167991 213974 168000
rect 214288 167612 214340 167618
rect 214288 167554 214340 167560
rect 214300 167249 214328 167554
rect 214286 167240 214342 167249
rect 214286 167175 214342 167184
rect 214380 166864 214432 166870
rect 214380 166806 214432 166812
rect 214392 165753 214420 166806
rect 214378 165744 214434 165753
rect 214378 165679 214434 165688
rect 214104 165572 214156 165578
rect 214104 165514 214156 165520
rect 214116 164937 214144 165514
rect 214102 164928 214158 164937
rect 214102 164863 214158 164872
rect 214380 164212 214432 164218
rect 214380 164154 214432 164160
rect 214392 163305 214420 164154
rect 214378 163296 214434 163305
rect 214378 163231 214434 163240
rect 214288 162852 214340 162858
rect 214288 162794 214340 162800
rect 214300 161809 214328 162794
rect 214286 161800 214342 161809
rect 214286 161735 214342 161744
rect 214378 155544 214434 155553
rect 214378 155479 214434 155488
rect 214392 154698 214420 155479
rect 214380 154692 214432 154698
rect 214380 154634 214432 154640
rect 214010 152416 214066 152425
rect 214010 152351 214066 152360
rect 214024 151910 214052 152351
rect 214012 151904 214064 151910
rect 214012 151846 214064 151852
rect 214378 151600 214434 151609
rect 214378 151535 214434 151544
rect 214392 150550 214420 151535
rect 214380 150544 214432 150550
rect 214380 150486 214432 150492
rect 214378 149968 214434 149977
rect 214378 149903 214434 149912
rect 214392 149258 214420 149903
rect 214380 149252 214432 149258
rect 214380 149194 214432 149200
rect 214470 144528 214526 144537
rect 214470 144463 214526 144472
rect 214484 143614 214512 144463
rect 214472 143608 214524 143614
rect 214472 143550 214524 143556
rect 214378 139904 214434 139913
rect 214378 139839 214434 139848
rect 214392 139534 214420 139839
rect 214380 139528 214432 139534
rect 214380 139470 214432 139476
rect 214470 139088 214526 139097
rect 214470 139023 214526 139032
rect 214484 138038 214512 139023
rect 214472 138032 214524 138038
rect 214472 137974 214524 137980
rect 214286 137456 214342 137465
rect 214286 137391 214342 137400
rect 214300 136678 214328 137391
rect 214288 136672 214340 136678
rect 214288 136614 214340 136620
rect 214194 135960 214250 135969
rect 214194 135895 214250 135904
rect 214208 135318 214236 135895
rect 214196 135312 214248 135318
rect 214196 135254 214248 135260
rect 117134 133648 117190 133657
rect 117134 133583 117190 133592
rect 117148 132938 117176 133583
rect 117136 132932 117188 132938
rect 117136 132874 117188 132880
rect 214010 132832 214066 132841
rect 214010 132767 214066 132776
rect 214024 132598 214052 132767
rect 214012 132592 214064 132598
rect 214012 132534 214064 132540
rect 214378 132016 214434 132025
rect 214378 131951 214434 131960
rect 214392 131170 214420 131951
rect 214380 131164 214432 131170
rect 214380 131106 214432 131112
rect 214194 130384 214250 130393
rect 214194 130319 214250 130328
rect 116674 130112 116730 130121
rect 116674 130047 116730 130056
rect 214208 129810 214236 130319
rect 214196 129804 214248 129810
rect 214196 129746 214248 129752
rect 214194 129704 214250 129713
rect 214194 129639 214250 129648
rect 214208 129062 214236 129639
rect 214196 129056 214248 129062
rect 214196 128998 214248 129004
rect 214010 128888 214066 128897
rect 214010 128823 214066 128832
rect 214024 128382 214052 128823
rect 214012 128376 214064 128382
rect 214012 128318 214064 128324
rect 116582 123040 116638 123049
rect 116582 122975 116638 122984
rect 116398 121952 116454 121961
rect 116398 121887 116454 121896
rect 116412 121514 116440 121887
rect 50988 121508 51040 121514
rect 50988 121450 51040 121456
rect 116400 121508 116452 121514
rect 116400 121450 116452 121456
rect 51000 99362 51028 121450
rect 116398 120728 116454 120737
rect 116398 120663 116454 120672
rect 116412 120154 116440 120663
rect 100024 120148 100076 120154
rect 100024 120090 100076 120096
rect 116400 120148 116452 120154
rect 116400 120090 116452 120096
rect 94780 118720 94832 118726
rect 94780 118662 94832 118668
rect 94688 117360 94740 117366
rect 94688 117302 94740 117308
rect 94596 116000 94648 116006
rect 94596 115942 94648 115948
rect 94504 114572 94556 114578
rect 94504 114514 94556 114520
rect 50646 99334 51028 99362
rect 94516 94489 94544 114514
rect 94608 95441 94636 115942
rect 94700 97209 94728 117302
rect 94792 98025 94820 118662
rect 94872 116068 94924 116074
rect 94872 116010 94924 116016
rect 94778 98016 94834 98025
rect 94778 97951 94834 97960
rect 94686 97200 94742 97209
rect 94686 97135 94742 97144
rect 94884 96257 94912 116010
rect 95884 113212 95936 113218
rect 95884 113154 95936 113160
rect 94964 109064 95016 109070
rect 94964 109006 95016 109012
rect 94870 96248 94926 96257
rect 94870 96183 94926 96192
rect 94594 95432 94650 95441
rect 94594 95367 94650 95376
rect 94688 95260 94740 95266
rect 94688 95202 94740 95208
rect 94502 94480 94558 94489
rect 94502 94415 94558 94424
rect 94596 93900 94648 93906
rect 94596 93842 94648 93848
rect 94412 93356 94464 93362
rect 94412 93298 94464 93304
rect 94424 92721 94452 93298
rect 94410 92712 94466 92721
rect 94410 92647 94466 92656
rect 94412 87916 94464 87922
rect 94412 87858 94464 87864
rect 94424 87281 94452 87858
rect 94410 87272 94466 87281
rect 94410 87207 94466 87216
rect 94504 86760 94556 86766
rect 94504 86702 94556 86708
rect 94516 86465 94544 86702
rect 94502 86456 94558 86465
rect 94502 86391 94558 86400
rect 94044 86216 94096 86222
rect 94044 86158 94096 86164
rect 94056 83745 94084 86158
rect 94042 83736 94098 83745
rect 94042 83671 94098 83680
rect 94228 83428 94280 83434
rect 94228 83370 94280 83376
rect 94240 82929 94268 83370
rect 94226 82920 94282 82929
rect 94226 82855 94282 82864
rect 94412 81388 94464 81394
rect 94412 81330 94464 81336
rect 94424 81025 94452 81330
rect 94410 81016 94466 81025
rect 94410 80951 94466 80960
rect 94412 78668 94464 78674
rect 94412 78610 94464 78616
rect 94228 77988 94280 77994
rect 94228 77930 94280 77936
rect 94044 76900 94096 76906
rect 94044 76842 94096 76848
rect 94056 73001 94084 76842
rect 94240 76537 94268 77930
rect 94424 77489 94452 78610
rect 94608 78441 94636 93842
rect 94700 80209 94728 95202
rect 94872 93696 94924 93702
rect 94872 93638 94924 93644
rect 94884 93537 94912 93638
rect 94870 93528 94926 93537
rect 94870 93463 94926 93472
rect 94976 90953 95004 109006
rect 95148 99000 95200 99006
rect 95146 98968 95148 98977
rect 95200 98968 95202 98977
rect 95146 98903 95202 98912
rect 95896 93702 95924 113154
rect 98644 111852 98696 111858
rect 98644 111794 98696 111800
rect 97264 107704 97316 107710
rect 97264 107646 97316 107652
rect 95976 102196 96028 102202
rect 95976 102138 96028 102144
rect 95884 93696 95936 93702
rect 95884 93638 95936 93644
rect 95148 92472 95200 92478
rect 95148 92414 95200 92420
rect 95160 91769 95188 92414
rect 95146 91760 95202 91769
rect 95146 91695 95202 91704
rect 95056 91044 95108 91050
rect 95056 90986 95108 90992
rect 94962 90944 95018 90953
rect 94962 90879 95018 90888
rect 95068 90001 95096 90986
rect 95054 89992 95110 90001
rect 95054 89927 95110 89936
rect 95148 89344 95200 89350
rect 95148 89286 95200 89292
rect 95160 89185 95188 89286
rect 95146 89176 95202 89185
rect 95146 89111 95202 89120
rect 95148 88256 95200 88262
rect 95146 88224 95148 88233
rect 95200 88224 95202 88233
rect 95146 88159 95202 88168
rect 95988 85542 96016 102138
rect 96068 96688 96120 96694
rect 96068 96630 96120 96636
rect 94872 85536 94924 85542
rect 94870 85504 94872 85513
rect 95976 85536 96028 85542
rect 94924 85504 94926 85513
rect 95976 85478 96028 85484
rect 94870 85439 94926 85448
rect 95148 84856 95200 84862
rect 95148 84798 95200 84804
rect 95160 84697 95188 84798
rect 95146 84688 95202 84697
rect 95146 84623 95202 84632
rect 95884 82884 95936 82890
rect 95884 82826 95936 82832
rect 95148 82816 95200 82822
rect 95148 82758 95200 82764
rect 95160 81977 95188 82758
rect 95146 81968 95202 81977
rect 95146 81903 95202 81912
rect 94964 81456 95016 81462
rect 94964 81398 95016 81404
rect 94686 80200 94742 80209
rect 94686 80135 94742 80144
rect 94594 78432 94650 78441
rect 94594 78367 94650 78376
rect 94410 77480 94466 77489
rect 94410 77415 94466 77424
rect 94226 76528 94282 76537
rect 94226 76463 94282 76472
rect 94596 75744 94648 75750
rect 94594 75712 94596 75721
rect 94648 75712 94650 75721
rect 94594 75647 94650 75656
rect 94976 74769 95004 81398
rect 95240 80708 95292 80714
rect 95240 80650 95292 80656
rect 95146 79248 95202 79257
rect 95252 79234 95280 80650
rect 95202 79206 95280 79234
rect 95146 79183 95202 79192
rect 94962 74760 95018 74769
rect 94962 74695 95018 74704
rect 94596 74588 94648 74594
rect 94596 74530 94648 74536
rect 94042 72992 94098 73001
rect 94042 72927 94098 72936
rect 94412 72684 94464 72690
rect 94412 72626 94464 72632
rect 94424 72185 94452 72626
rect 94410 72176 94466 72185
rect 94410 72111 94466 72120
rect 94228 71732 94280 71738
rect 94228 71674 94280 71680
rect 94240 71233 94268 71674
rect 94226 71224 94282 71233
rect 94226 71159 94282 71168
rect 94504 70440 94556 70446
rect 94504 70382 94556 70388
rect 94044 68604 94096 68610
rect 94044 68546 94096 68552
rect 94056 68513 94084 68546
rect 94042 68504 94098 68513
rect 94042 68439 94098 68448
rect 94412 66020 94464 66026
rect 94412 65962 94464 65968
rect 94136 65952 94188 65958
rect 94134 65920 94136 65929
rect 94188 65920 94190 65929
rect 94134 65855 94190 65864
rect 94424 64977 94452 65962
rect 94410 64968 94466 64977
rect 94410 64903 94466 64912
rect 94320 61804 94372 61810
rect 94320 61746 94372 61752
rect 94332 61441 94360 61746
rect 94318 61432 94374 61441
rect 94318 61367 94374 61376
rect 94516 60489 94544 70382
rect 94608 64025 94636 74530
rect 95148 74248 95200 74254
rect 95148 74190 95200 74196
rect 95160 73953 95188 74190
rect 95146 73944 95202 73953
rect 95146 73879 95202 73888
rect 94780 71800 94832 71806
rect 94780 71742 94832 71748
rect 94688 67652 94740 67658
rect 94688 67594 94740 67600
rect 94594 64016 94650 64025
rect 94594 63951 94650 63960
rect 94596 62144 94648 62150
rect 94596 62086 94648 62092
rect 94502 60480 94558 60489
rect 94502 60415 94558 60424
rect 94320 59900 94372 59906
rect 94320 59842 94372 59848
rect 94332 59537 94360 59842
rect 94318 59528 94374 59537
rect 94318 59463 94374 59472
rect 94412 57928 94464 57934
rect 94412 57870 94464 57876
rect 94424 57769 94452 57870
rect 94410 57760 94466 57769
rect 94410 57695 94466 57704
rect 94044 55344 94096 55350
rect 94044 55286 94096 55292
rect 94056 49745 94084 55286
rect 94136 55276 94188 55282
rect 94136 55218 94188 55224
rect 94042 49736 94098 49745
rect 94042 49671 94098 49680
rect 94148 48929 94176 55218
rect 94608 55185 94636 62086
rect 94700 58721 94728 67594
rect 94792 62257 94820 71742
rect 95056 70508 95108 70514
rect 95056 70450 95108 70456
rect 94872 70304 94924 70310
rect 94870 70272 94872 70281
rect 94924 70272 94926 70281
rect 94870 70207 94926 70216
rect 95068 69465 95096 70450
rect 95896 70310 95924 82826
rect 96080 81394 96108 96630
rect 97276 89350 97304 107646
rect 97356 104916 97408 104922
rect 97356 104858 97408 104864
rect 97264 89344 97316 89350
rect 97264 89286 97316 89292
rect 97368 87922 97396 104858
rect 98656 93362 98684 111794
rect 98736 100768 98788 100774
rect 98736 100710 98788 100716
rect 98644 93356 98696 93362
rect 98644 93298 98696 93304
rect 97448 89752 97500 89758
rect 97448 89694 97500 89700
rect 97356 87916 97408 87922
rect 97356 87858 97408 87864
rect 96068 81388 96120 81394
rect 96068 81330 96120 81336
rect 97264 80096 97316 80102
rect 97264 80038 97316 80044
rect 96068 79348 96120 79354
rect 96068 79290 96120 79296
rect 95976 75948 96028 75954
rect 95976 75890 96028 75896
rect 95884 70304 95936 70310
rect 95884 70246 95936 70252
rect 95148 69896 95200 69902
rect 95148 69838 95200 69844
rect 95054 69456 95110 69465
rect 95054 69391 95110 69400
rect 95160 67697 95188 69838
rect 95146 67688 95202 67697
rect 95146 67623 95202 67632
rect 95148 67516 95200 67522
rect 95148 67458 95200 67464
rect 95160 66745 95188 67458
rect 95146 66736 95202 66745
rect 95146 66671 95202 66680
rect 95988 66026 96016 75890
rect 96080 71738 96108 79290
rect 96620 73840 96672 73846
rect 96620 73782 96672 73788
rect 96068 71732 96120 71738
rect 96068 71674 96120 71680
rect 96068 69080 96120 69086
rect 96068 69022 96120 69028
rect 95976 66020 96028 66026
rect 95976 65962 96028 65968
rect 94872 64932 94924 64938
rect 94872 64874 94924 64880
rect 94778 62248 94834 62257
rect 94778 62183 94834 62192
rect 94780 60784 94832 60790
rect 94780 60726 94832 60732
rect 94686 58712 94742 58721
rect 94686 58647 94742 58656
rect 94594 55176 94650 55185
rect 94594 55111 94650 55120
rect 94596 54732 94648 54738
rect 94596 54674 94648 54680
rect 94608 54233 94636 54674
rect 94594 54224 94650 54233
rect 94594 54159 94650 54168
rect 94792 53281 94820 60726
rect 94884 56953 94912 64874
rect 95240 63572 95292 63578
rect 95240 63514 95292 63520
rect 95148 63232 95200 63238
rect 95146 63200 95148 63209
rect 95200 63200 95202 63209
rect 95146 63135 95202 63144
rect 94964 57996 95016 58002
rect 94964 57938 95016 57944
rect 94870 56944 94926 56953
rect 94870 56879 94926 56888
rect 94872 53848 94924 53854
rect 94872 53790 94924 53796
rect 94778 53272 94834 53281
rect 94778 53207 94834 53216
rect 94780 52488 94832 52494
rect 94780 52430 94832 52436
rect 94134 48920 94190 48929
rect 94134 48855 94190 48864
rect 94412 48340 94464 48346
rect 94412 48282 94464 48288
rect 94136 46980 94188 46986
rect 94136 46922 94188 46928
rect 93952 45620 94004 45626
rect 93952 45562 94004 45568
rect 93964 41721 93992 45562
rect 94148 42537 94176 46922
rect 94424 44441 94452 48282
rect 94792 47025 94820 52430
rect 94884 47977 94912 53790
rect 94976 51513 95004 57938
rect 95252 56794 95280 63514
rect 96080 59906 96108 69022
rect 96632 67522 96660 73782
rect 97276 68610 97304 80038
rect 97460 75750 97488 89694
rect 97540 88392 97592 88398
rect 97540 88334 97592 88340
rect 97552 81462 97580 88334
rect 98644 87032 98696 87038
rect 98644 86974 98696 86980
rect 97540 81456 97592 81462
rect 97540 81398 97592 81404
rect 97448 75744 97500 75750
rect 97448 75686 97500 75692
rect 98656 74254 98684 86974
rect 98748 86222 98776 100710
rect 100036 99006 100064 120090
rect 214196 120080 214248 120086
rect 214196 120022 214248 120028
rect 116398 119640 116454 119649
rect 116398 119575 116454 119584
rect 116412 118726 116440 119575
rect 214208 119513 214236 120022
rect 214194 119504 214250 119513
rect 214194 119439 214250 119448
rect 116400 118720 116452 118726
rect 116400 118662 116452 118668
rect 214288 118652 214340 118658
rect 214288 118594 214340 118600
rect 116398 118416 116454 118425
rect 116398 118351 116454 118360
rect 116412 117366 116440 118351
rect 214300 117881 214328 118594
rect 214286 117872 214342 117881
rect 214286 117807 214342 117816
rect 116400 117360 116452 117366
rect 116400 117302 116452 117308
rect 116306 117192 116362 117201
rect 116306 117127 116362 117136
rect 116320 116074 116348 117127
rect 116398 116104 116454 116113
rect 116308 116068 116360 116074
rect 116398 116039 116454 116048
rect 116308 116010 116360 116016
rect 116412 116006 116440 116039
rect 116400 116000 116452 116006
rect 116400 115942 116452 115948
rect 116398 114880 116454 114889
rect 116398 114815 116454 114824
rect 116412 114578 116440 114815
rect 116400 114572 116452 114578
rect 116400 114514 116452 114520
rect 214012 114436 214064 114442
rect 214012 114378 214064 114384
rect 214024 113937 214052 114378
rect 214010 113928 214066 113937
rect 214010 113863 214066 113872
rect 116398 113792 116454 113801
rect 116398 113727 116454 113736
rect 116412 113218 116440 113727
rect 116400 113212 116452 113218
rect 116400 113154 116452 113160
rect 214380 113144 214432 113150
rect 214380 113086 214432 113092
rect 116398 112568 116454 112577
rect 116398 112503 116454 112512
rect 116412 111858 116440 112503
rect 214392 112441 214420 113086
rect 214378 112432 214434 112441
rect 214378 112367 214434 112376
rect 116400 111852 116452 111858
rect 116400 111794 116452 111800
rect 116398 111480 116454 111489
rect 116398 111415 116454 111424
rect 116412 110498 116440 111415
rect 104164 110492 104216 110498
rect 104164 110434 104216 110440
rect 116400 110492 116452 110498
rect 116400 110434 116452 110440
rect 101404 106344 101456 106350
rect 101404 106286 101456 106292
rect 100116 99408 100168 99414
rect 100116 99350 100168 99356
rect 100024 99000 100076 99006
rect 100024 98942 100076 98948
rect 98828 93152 98880 93158
rect 98828 93094 98880 93100
rect 98736 86216 98788 86222
rect 98736 86158 98788 86164
rect 98840 84862 98868 93094
rect 98828 84856 98880 84862
rect 98828 84798 98880 84804
rect 100024 84856 100076 84862
rect 100024 84798 100076 84804
rect 98736 81456 98788 81462
rect 98736 81398 98788 81404
rect 98644 74248 98696 74254
rect 98644 74190 98696 74196
rect 98748 70514 98776 81398
rect 98828 73228 98880 73234
rect 98828 73170 98880 73176
rect 98736 70508 98788 70514
rect 98736 70450 98788 70456
rect 97264 68604 97316 68610
rect 97264 68546 97316 68552
rect 96620 67516 96672 67522
rect 96620 67458 96672 67464
rect 97264 66292 97316 66298
rect 97264 66234 97316 66240
rect 96160 60036 96212 60042
rect 96160 59978 96212 59984
rect 96068 59900 96120 59906
rect 96068 59842 96120 59848
rect 95160 56766 95280 56794
rect 95160 56001 95188 56766
rect 95240 56636 95292 56642
rect 95240 56578 95292 56584
rect 95146 55992 95202 56001
rect 95146 55927 95202 55936
rect 95146 52456 95202 52465
rect 95146 52391 95148 52400
rect 95200 52391 95202 52400
rect 95148 52362 95200 52368
rect 94962 51504 95018 51513
rect 94962 51439 95018 51448
rect 95056 51128 95108 51134
rect 95056 51070 95108 51076
rect 94964 48408 95016 48414
rect 94964 48350 95016 48356
rect 94870 47968 94926 47977
rect 94870 47903 94926 47912
rect 94778 47016 94834 47025
rect 94778 46951 94834 46960
rect 94410 44432 94466 44441
rect 94410 44367 94466 44376
rect 94976 43489 95004 48350
rect 95068 46209 95096 51070
rect 95146 50688 95202 50697
rect 95252 50674 95280 56578
rect 96172 54738 96200 59978
rect 97276 57934 97304 66234
rect 98840 63238 98868 73170
rect 100036 72690 100064 84798
rect 100128 83434 100156 99350
rect 101416 88262 101444 106286
rect 102784 103556 102836 103562
rect 102784 103498 102836 103504
rect 101496 92540 101548 92546
rect 101496 92482 101548 92488
rect 101404 88256 101456 88262
rect 101404 88198 101456 88204
rect 100116 83428 100168 83434
rect 100116 83370 100168 83376
rect 101508 78674 101536 92482
rect 102796 86766 102824 103498
rect 104176 92478 104204 110434
rect 214472 110356 214524 110362
rect 214472 110298 214524 110304
rect 116398 110256 116454 110265
rect 116398 110191 116454 110200
rect 116412 109070 116440 110191
rect 214484 109313 214512 110298
rect 214470 109304 214526 109313
rect 214470 109239 214526 109248
rect 116400 109064 116452 109070
rect 116306 109032 116362 109041
rect 116400 109006 116452 109012
rect 116306 108967 116362 108976
rect 116320 107778 116348 108967
rect 116398 107944 116454 107953
rect 116398 107879 116454 107888
rect 105544 107772 105596 107778
rect 105544 107714 105596 107720
rect 116308 107772 116360 107778
rect 116308 107714 116360 107720
rect 104164 92472 104216 92478
rect 104164 92414 104216 92420
rect 104256 91112 104308 91118
rect 104256 91054 104308 91060
rect 102784 86760 102836 86766
rect 102784 86702 102836 86708
rect 102876 85604 102928 85610
rect 102876 85546 102928 85552
rect 102784 78736 102836 78742
rect 102784 78678 102836 78684
rect 101496 78668 101548 78674
rect 101496 78610 101548 78616
rect 101404 77308 101456 77314
rect 101404 77250 101456 77256
rect 100024 72684 100076 72690
rect 100024 72626 100076 72632
rect 100024 70508 100076 70514
rect 100024 70450 100076 70456
rect 98828 63232 98880 63238
rect 98828 63174 98880 63180
rect 100036 61810 100064 70450
rect 101416 65958 101444 77250
rect 102796 69902 102824 78678
rect 102888 76906 102916 85546
rect 104268 77994 104296 91054
rect 105556 91050 105584 107714
rect 116412 107710 116440 107879
rect 116400 107704 116452 107710
rect 116400 107646 116452 107652
rect 214196 107636 214248 107642
rect 214196 107578 214248 107584
rect 214208 107001 214236 107578
rect 214194 106992 214250 107001
rect 214194 106927 214250 106936
rect 116398 106720 116454 106729
rect 116398 106655 116454 106664
rect 116412 106350 116440 106655
rect 116400 106344 116452 106350
rect 116400 106286 116452 106292
rect 214380 106208 214432 106214
rect 214380 106150 214432 106156
rect 116398 105632 116454 105641
rect 116398 105567 116454 105576
rect 116412 104922 116440 105567
rect 214392 105369 214420 106150
rect 214378 105360 214434 105369
rect 214378 105295 214434 105304
rect 116400 104916 116452 104922
rect 116400 104858 116452 104864
rect 214380 104780 214432 104786
rect 214380 104722 214432 104728
rect 116398 104408 116454 104417
rect 116398 104343 116454 104352
rect 116412 103562 116440 104343
rect 214392 103873 214420 104722
rect 214378 103864 214434 103873
rect 214378 103799 214434 103808
rect 116400 103556 116452 103562
rect 116400 103498 116452 103504
rect 116306 103184 116362 103193
rect 116306 103119 116362 103128
rect 116320 102202 116348 103119
rect 116308 102196 116360 102202
rect 116308 102138 116360 102144
rect 116674 102096 116730 102105
rect 116674 102031 116730 102040
rect 116398 100872 116454 100881
rect 116398 100807 116454 100816
rect 116412 100774 116440 100807
rect 116400 100768 116452 100774
rect 116400 100710 116452 100716
rect 116398 99784 116454 99793
rect 116398 99719 116454 99728
rect 116412 99414 116440 99719
rect 116400 99408 116452 99414
rect 116400 99350 116452 99356
rect 116398 98560 116454 98569
rect 116398 98495 116454 98504
rect 116412 98054 116440 98495
rect 106924 98048 106976 98054
rect 106924 97990 106976 97996
rect 116400 98048 116452 98054
rect 116400 97990 116452 97996
rect 105544 91044 105596 91050
rect 105544 90986 105596 90992
rect 106936 82822 106964 97990
rect 116398 97336 116454 97345
rect 116398 97271 116454 97280
rect 116412 96694 116440 97271
rect 116400 96688 116452 96694
rect 116400 96630 116452 96636
rect 116306 96248 116362 96257
rect 116306 96183 116362 96192
rect 116320 95266 116348 96183
rect 116308 95260 116360 95266
rect 116308 95202 116360 95208
rect 116582 95024 116638 95033
rect 116582 94959 116638 94968
rect 116398 93936 116454 93945
rect 116398 93871 116400 93880
rect 116452 93871 116454 93880
rect 116400 93842 116452 93848
rect 116398 92712 116454 92721
rect 116398 92647 116454 92656
rect 116412 92546 116440 92647
rect 116400 92540 116452 92546
rect 116400 92482 116452 92488
rect 116398 91624 116454 91633
rect 116398 91559 116454 91568
rect 116412 91118 116440 91559
rect 116400 91112 116452 91118
rect 116400 91054 116452 91060
rect 116398 90400 116454 90409
rect 116398 90335 116454 90344
rect 116412 89758 116440 90335
rect 116400 89752 116452 89758
rect 116400 89694 116452 89700
rect 115938 89176 115994 89185
rect 115938 89111 115994 89120
rect 115952 88398 115980 89111
rect 115940 88392 115992 88398
rect 115940 88334 115992 88340
rect 116398 88088 116454 88097
rect 116398 88023 116454 88032
rect 116412 87038 116440 88023
rect 116400 87032 116452 87038
rect 116400 86974 116452 86980
rect 116122 86864 116178 86873
rect 116122 86799 116178 86808
rect 116136 85610 116164 86799
rect 116398 85776 116454 85785
rect 116398 85711 116454 85720
rect 116124 85604 116176 85610
rect 116124 85546 116176 85552
rect 116412 84862 116440 85711
rect 116400 84856 116452 84862
rect 116400 84798 116452 84804
rect 116398 83328 116454 83337
rect 116398 83263 116454 83272
rect 116412 82890 116440 83263
rect 116400 82884 116452 82890
rect 116400 82826 116452 82832
rect 106924 82816 106976 82822
rect 106924 82758 106976 82764
rect 115938 82240 115994 82249
rect 115938 82175 115994 82184
rect 115952 81462 115980 82175
rect 115940 81456 115992 81462
rect 115940 81398 115992 81404
rect 116398 81016 116454 81025
rect 116398 80951 116454 80960
rect 116412 80102 116440 80951
rect 116596 80714 116624 94959
rect 116688 93158 116716 102031
rect 214472 100700 214524 100706
rect 214472 100642 214524 100648
rect 214484 99929 214512 100642
rect 214470 99920 214526 99929
rect 214470 99855 214526 99864
rect 214576 99634 214604 229706
rect 214656 227044 214708 227050
rect 214656 226986 214708 226992
rect 214300 99606 214604 99634
rect 214104 97980 214156 97986
rect 214104 97922 214156 97928
rect 214116 97481 214144 97922
rect 214102 97472 214158 97481
rect 214102 97407 214158 97416
rect 214300 95985 214328 99606
rect 214668 99498 214696 226986
rect 214760 157865 214788 231066
rect 214932 228404 214984 228410
rect 214932 228346 214984 228352
rect 214840 182232 214892 182238
rect 214840 182174 214892 182180
rect 214852 170377 214880 182174
rect 214838 170368 214894 170377
rect 214838 170303 214894 170312
rect 214944 166274 214972 228346
rect 227640 221377 227668 232494
rect 229744 223644 229796 223650
rect 229744 223586 229796 223592
rect 215114 221368 215170 221377
rect 215114 221303 215170 221312
rect 227626 221368 227682 221377
rect 227626 221303 227682 221312
rect 215128 220862 215156 221303
rect 215116 220856 215168 220862
rect 226340 220856 226392 220862
rect 215116 220798 215168 220804
rect 226338 220824 226340 220833
rect 226392 220824 226394 220833
rect 226338 220759 226394 220768
rect 215206 220552 215262 220561
rect 215206 220487 215262 220496
rect 215116 220176 215168 220182
rect 215116 220118 215168 220124
rect 215128 219745 215156 220118
rect 215220 220114 215248 220487
rect 226432 220176 226484 220182
rect 226338 220144 226394 220153
rect 215208 220108 215260 220114
rect 226432 220118 226484 220124
rect 226338 220079 226340 220088
rect 215208 220050 215260 220056
rect 226392 220079 226394 220088
rect 226340 220050 226392 220056
rect 215114 219736 215170 219745
rect 215114 219671 215170 219680
rect 226444 219609 226472 220118
rect 226430 219600 226486 219609
rect 226430 219535 226486 219544
rect 226338 219056 226394 219065
rect 226338 218991 226394 219000
rect 215114 218920 215170 218929
rect 215114 218855 215170 218864
rect 215128 218822 215156 218855
rect 226352 218822 226380 218991
rect 215116 218816 215168 218822
rect 215116 218758 215168 218764
rect 226340 218816 226392 218822
rect 226340 218758 226392 218764
rect 215208 218748 215260 218754
rect 215208 218690 215260 218696
rect 226432 218748 226484 218754
rect 226432 218690 226484 218696
rect 215220 218249 215248 218690
rect 226444 218385 226472 218690
rect 226430 218376 226486 218385
rect 226430 218311 226486 218320
rect 215206 218240 215262 218249
rect 215206 218175 215262 218184
rect 226338 217832 226394 217841
rect 226338 217767 226394 217776
rect 215114 217424 215170 217433
rect 215114 217359 215170 217368
rect 215128 217326 215156 217359
rect 226352 217326 226380 217767
rect 215116 217320 215168 217326
rect 215116 217262 215168 217268
rect 226340 217320 226392 217326
rect 226340 217262 226392 217268
rect 226430 217288 226486 217297
rect 226430 217223 226486 217232
rect 226444 216646 226472 217223
rect 215116 216640 215168 216646
rect 215114 216608 215116 216617
rect 226432 216640 226484 216646
rect 215168 216608 215170 216617
rect 215114 216543 215170 216552
rect 226338 216608 226394 216617
rect 226432 216582 226484 216588
rect 226338 216543 226394 216552
rect 226352 215966 226380 216543
rect 226430 216064 226486 216073
rect 226430 215999 226486 216008
rect 215116 215960 215168 215966
rect 215116 215902 215168 215908
rect 226340 215960 226392 215966
rect 226340 215902 226392 215908
rect 215128 215801 215156 215902
rect 215114 215792 215170 215801
rect 215114 215727 215170 215736
rect 226338 215520 226394 215529
rect 226338 215455 226394 215464
rect 215116 215280 215168 215286
rect 215116 215222 215168 215228
rect 215128 215121 215156 215222
rect 226352 215218 226380 215455
rect 226444 215286 226472 215999
rect 226432 215280 226484 215286
rect 226432 215222 226484 215228
rect 215208 215212 215260 215218
rect 215208 215154 215260 215160
rect 226340 215212 226392 215218
rect 226340 215154 226392 215160
rect 215114 215112 215170 215121
rect 215114 215047 215170 215056
rect 215220 214305 215248 215154
rect 226430 214840 226486 214849
rect 226430 214775 226486 214784
rect 215206 214296 215262 214305
rect 215206 214231 215262 214240
rect 226338 214296 226394 214305
rect 226338 214231 226394 214240
rect 215116 213920 215168 213926
rect 215116 213862 215168 213868
rect 215128 213489 215156 213862
rect 226352 213858 226380 214231
rect 226444 213926 226472 214775
rect 226432 213920 226484 213926
rect 226432 213862 226484 213868
rect 226340 213852 226392 213858
rect 226340 213794 226392 213800
rect 226430 213616 226486 213625
rect 226430 213551 226486 213560
rect 215114 213480 215170 213489
rect 215114 213415 215170 213424
rect 226338 213072 226394 213081
rect 226338 213007 226394 213016
rect 215116 212492 215168 212498
rect 215116 212434 215168 212440
rect 215128 211993 215156 212434
rect 226352 212430 226380 213007
rect 226444 212498 226472 213551
rect 226522 212528 226578 212537
rect 226432 212492 226484 212498
rect 226522 212463 226578 212472
rect 226432 212434 226484 212440
rect 215208 212424 215260 212430
rect 215208 212366 215260 212372
rect 226340 212424 226392 212430
rect 226340 212366 226392 212372
rect 215114 211984 215170 211993
rect 215114 211919 215170 211928
rect 215220 211177 215248 212366
rect 226154 211848 226210 211857
rect 226154 211783 226210 211792
rect 215206 211168 215262 211177
rect 215206 211103 215262 211112
rect 226062 210760 226118 210769
rect 226062 210695 226118 210704
rect 225970 210080 226026 210089
rect 225970 210015 226026 210024
rect 215116 209772 215168 209778
rect 215116 209714 215168 209720
rect 215128 209545 215156 209714
rect 215114 209536 215170 209545
rect 215114 209471 215170 209480
rect 215116 208344 215168 208350
rect 215116 208286 215168 208292
rect 215128 208049 215156 208286
rect 225984 208282 226012 210015
rect 226076 208350 226104 210695
rect 226168 209778 226196 211783
rect 226246 211304 226302 211313
rect 226246 211239 226302 211248
rect 226156 209772 226208 209778
rect 226156 209714 226208 209720
rect 226260 209710 226288 211239
rect 226536 211138 226564 212463
rect 226524 211132 226576 211138
rect 226524 211074 226576 211080
rect 226248 209704 226300 209710
rect 226248 209646 226300 209652
rect 226154 209536 226210 209545
rect 226154 209471 226210 209480
rect 226064 208344 226116 208350
rect 226064 208286 226116 208292
rect 225972 208276 226024 208282
rect 225972 208218 226024 208224
rect 226168 208162 226196 209471
rect 226246 208992 226302 209001
rect 226246 208927 226302 208936
rect 226076 208134 226196 208162
rect 215114 208040 215170 208049
rect 215114 207975 215170 207984
rect 225878 207768 225934 207777
rect 225878 207703 225934 207712
rect 215116 206984 215168 206990
rect 215116 206926 215168 206932
rect 215128 206417 215156 206926
rect 225786 206544 225842 206553
rect 225786 206479 225842 206488
rect 215114 206408 215170 206417
rect 215114 206343 215170 206352
rect 215116 205624 215168 205630
rect 215116 205566 215168 205572
rect 215128 204921 215156 205566
rect 225602 205320 225658 205329
rect 225602 205255 225658 205264
rect 215114 204912 215170 204921
rect 215114 204847 215170 204856
rect 215208 204264 215260 204270
rect 215208 204206 215260 204212
rect 215116 204196 215168 204202
rect 215116 204138 215168 204144
rect 215128 204105 215156 204138
rect 215114 204096 215170 204105
rect 215114 204031 215170 204040
rect 215220 203289 215248 204206
rect 215206 203280 215262 203289
rect 215206 203215 215262 203224
rect 215116 202768 215168 202774
rect 215116 202710 215168 202716
rect 215128 202473 215156 202710
rect 215114 202464 215170 202473
rect 215114 202399 215170 202408
rect 225616 201482 225644 205255
rect 225694 203008 225750 203017
rect 225694 202943 225750 202952
rect 225604 201476 225656 201482
rect 225604 201418 225656 201424
rect 215116 201408 215168 201414
rect 215116 201350 215168 201356
rect 215128 200161 215156 201350
rect 215114 200152 215170 200161
rect 215114 200087 215170 200096
rect 224040 198824 224092 198830
rect 224040 198766 224092 198772
rect 215116 198688 215168 198694
rect 215114 198656 215116 198665
rect 215168 198656 215170 198665
rect 215114 198591 215170 198600
rect 223948 197464 224000 197470
rect 223948 197406 224000 197412
rect 215116 197260 215168 197266
rect 215116 197202 215168 197208
rect 215128 197033 215156 197202
rect 215114 197024 215170 197033
rect 215114 196959 215170 196968
rect 215208 195968 215260 195974
rect 215208 195910 215260 195916
rect 215116 195900 215168 195906
rect 215116 195842 215168 195848
rect 215128 195537 215156 195842
rect 215114 195528 215170 195537
rect 215114 195463 215170 195472
rect 215220 194721 215248 195910
rect 215206 194712 215262 194721
rect 215206 194647 215262 194656
rect 215116 194540 215168 194546
rect 215116 194482 215168 194488
rect 215128 193905 215156 194482
rect 215114 193896 215170 193905
rect 215114 193831 215170 193840
rect 220268 193316 220320 193322
rect 220268 193258 220320 193264
rect 215944 193248 215996 193254
rect 215944 193190 215996 193196
rect 215116 193180 215168 193186
rect 215116 193122 215168 193128
rect 215128 193089 215156 193122
rect 215208 193112 215260 193118
rect 215114 193080 215170 193089
rect 215208 193054 215260 193060
rect 215114 193015 215170 193024
rect 215220 192409 215248 193054
rect 215206 192400 215262 192409
rect 215206 192335 215262 192344
rect 215116 191752 215168 191758
rect 215116 191694 215168 191700
rect 215128 191593 215156 191694
rect 215114 191584 215170 191593
rect 215114 191519 215170 191528
rect 215300 191140 215352 191146
rect 215300 191082 215352 191088
rect 215116 190392 215168 190398
rect 215116 190334 215168 190340
rect 215128 189961 215156 190334
rect 215114 189952 215170 189961
rect 215114 189887 215170 189896
rect 215206 187640 215262 187649
rect 215116 187604 215168 187610
rect 215312 187626 215340 191082
rect 215262 187598 215340 187626
rect 215206 187575 215262 187584
rect 215116 187546 215168 187552
rect 215128 186017 215156 187546
rect 215208 187196 215260 187202
rect 215208 187138 215260 187144
rect 215220 186833 215248 187138
rect 215206 186824 215262 186833
rect 215206 186759 215262 186768
rect 215114 186008 215170 186017
rect 215114 185943 215170 185952
rect 215300 185632 215352 185638
rect 215300 185574 215352 185580
rect 215024 183592 215076 183598
rect 215024 183534 215076 183540
rect 215036 177698 215064 183534
rect 215114 182880 215170 182889
rect 215114 182815 215170 182824
rect 215128 182578 215156 182815
rect 215116 182572 215168 182578
rect 215116 182514 215168 182520
rect 215206 182200 215262 182209
rect 215312 182186 215340 185574
rect 215956 185570 215984 193190
rect 218152 191888 218204 191894
rect 218152 191830 218204 191836
rect 218060 189780 218112 189786
rect 218060 189722 218112 189728
rect 216036 187740 216088 187746
rect 216036 187682 216088 187688
rect 215944 185564 215996 185570
rect 215944 185506 215996 185512
rect 215262 182158 215340 182186
rect 215206 182135 215262 182144
rect 216048 179246 216076 187682
rect 218072 187202 218100 189722
rect 218060 187196 218112 187202
rect 218060 187138 218112 187144
rect 218164 184822 218192 191830
rect 220084 189100 220136 189106
rect 220084 189042 220136 189048
rect 218796 186516 218848 186522
rect 218796 186458 218848 186464
rect 218152 184816 218204 184822
rect 218152 184758 218204 184764
rect 216036 179240 216088 179246
rect 216036 179182 216088 179188
rect 215944 178696 215996 178702
rect 215944 178638 215996 178644
rect 215036 177670 215248 177698
rect 215024 177540 215076 177546
rect 215024 177482 215076 177488
rect 215036 177449 215064 177482
rect 215022 177440 215078 177449
rect 215022 177375 215078 177384
rect 215116 176656 215168 176662
rect 215114 176624 215116 176633
rect 215168 176624 215170 176633
rect 215114 176559 215170 176568
rect 215116 176180 215168 176186
rect 215116 176122 215168 176128
rect 215128 175953 215156 176122
rect 215114 175944 215170 175953
rect 215114 175879 215170 175888
rect 215116 175160 215168 175166
rect 215114 175128 215116 175137
rect 215168 175128 215170 175137
rect 215114 175063 215170 175072
rect 215220 173505 215248 177670
rect 215206 173496 215262 173505
rect 215206 173431 215262 173440
rect 215024 172032 215076 172038
rect 215024 171974 215076 171980
rect 215036 171193 215064 171974
rect 215022 171184 215078 171193
rect 215022 171119 215078 171128
rect 215116 169720 215168 169726
rect 215116 169662 215168 169668
rect 215128 169561 215156 169662
rect 215114 169552 215170 169561
rect 215114 169487 215170 169496
rect 215114 168872 215170 168881
rect 215114 168807 215170 168816
rect 215128 168638 215156 168807
rect 215116 168632 215168 168638
rect 215116 168574 215168 168580
rect 215956 168094 215984 178638
rect 218808 177546 218836 186458
rect 218888 181484 218940 181490
rect 218888 181426 218940 181432
rect 218796 177540 218848 177546
rect 218796 177482 218848 177488
rect 218704 176724 218756 176730
rect 218704 176666 218756 176672
rect 215944 168088 215996 168094
rect 215944 168030 215996 168036
rect 215300 167680 215352 167686
rect 215300 167622 215352 167628
rect 215206 166424 215262 166433
rect 215312 166410 215340 167622
rect 215262 166382 215340 166410
rect 215206 166359 215262 166368
rect 214852 166246 214972 166274
rect 214852 158681 214880 166246
rect 217232 165844 217284 165850
rect 217232 165786 217284 165792
rect 214932 164144 214984 164150
rect 214930 164112 214932 164121
rect 214984 164112 214986 164121
rect 214930 164047 214986 164056
rect 217244 163402 217272 165786
rect 218716 164150 218744 176666
rect 218900 172038 218928 181426
rect 220096 179790 220124 189042
rect 220280 187610 220308 193258
rect 223960 191758 223988 197406
rect 224052 193186 224080 198766
rect 224132 198756 224184 198762
rect 224132 198698 224184 198704
rect 224040 193180 224092 193186
rect 224040 193122 224092 193128
rect 224144 193118 224172 198698
rect 225708 198626 225736 202943
rect 225800 202774 225828 206479
rect 225892 204202 225920 207703
rect 225970 207224 226026 207233
rect 225970 207159 226026 207168
rect 225984 204270 226012 207159
rect 226076 206990 226104 208134
rect 226154 208040 226210 208049
rect 226154 207975 226210 207984
rect 226064 206984 226116 206990
rect 226064 206926 226116 206932
rect 226062 206000 226118 206009
rect 226062 205935 226118 205944
rect 225972 204264 226024 204270
rect 225972 204206 226024 204212
rect 225880 204196 225932 204202
rect 225880 204138 225932 204144
rect 225970 203552 226026 203561
rect 225970 203487 226026 203496
rect 225788 202768 225840 202774
rect 225788 202710 225840 202716
rect 225878 202464 225934 202473
rect 225878 202399 225934 202408
rect 225786 200016 225842 200025
rect 225786 199951 225842 199960
rect 225696 198620 225748 198626
rect 225696 198562 225748 198568
rect 224316 197396 224368 197402
rect 224316 197338 224368 197344
rect 224224 196104 224276 196110
rect 224224 196046 224276 196052
rect 224132 193112 224184 193118
rect 224132 193054 224184 193060
rect 223948 191752 224000 191758
rect 223948 191694 224000 191700
rect 221464 190936 221516 190942
rect 221464 190878 221516 190884
rect 220268 187604 220320 187610
rect 220268 187546 220320 187552
rect 220176 186380 220228 186386
rect 220176 186322 220228 186328
rect 220084 179784 220136 179790
rect 220084 179726 220136 179732
rect 220084 178084 220136 178090
rect 220084 178026 220136 178032
rect 218888 172032 218940 172038
rect 218888 171974 218940 171980
rect 220096 166870 220124 178026
rect 220188 176186 220216 186322
rect 221476 182578 221504 190878
rect 222844 190528 222896 190534
rect 222844 190470 222896 190476
rect 221648 187808 221700 187814
rect 221648 187750 221700 187756
rect 221464 182572 221516 182578
rect 221464 182514 221516 182520
rect 221556 180940 221608 180946
rect 221556 180882 221608 180888
rect 221464 179512 221516 179518
rect 221464 179454 221516 179460
rect 220176 176180 220228 176186
rect 220176 176122 220228 176128
rect 220268 175636 220320 175642
rect 220268 175578 220320 175584
rect 220084 166864 220136 166870
rect 220084 166806 220136 166812
rect 220280 165850 220308 175578
rect 221476 167618 221504 179454
rect 221568 168638 221596 180882
rect 221660 178634 221688 187750
rect 222856 182170 222884 190470
rect 224236 190398 224264 196046
rect 224328 191826 224356 197338
rect 224592 196036 224644 196042
rect 224592 195978 224644 195984
rect 224408 194608 224460 194614
rect 224408 194550 224460 194556
rect 224316 191820 224368 191826
rect 224316 191762 224368 191768
rect 224224 190392 224276 190398
rect 224224 190334 224276 190340
rect 224420 189038 224448 194550
rect 224604 190466 224632 195978
rect 225800 194546 225828 199951
rect 225892 197266 225920 202399
rect 225984 198694 226012 203487
rect 226076 202842 226104 205935
rect 226168 205630 226196 207975
rect 226260 206922 226288 208927
rect 226248 206916 226300 206922
rect 226248 206858 226300 206864
rect 226156 205624 226208 205630
rect 226156 205566 226208 205572
rect 226154 204776 226210 204785
rect 226154 204711 226210 204720
rect 226064 202836 226116 202842
rect 226064 202778 226116 202784
rect 226168 201906 226196 204711
rect 226246 204232 226302 204241
rect 226246 204167 226302 204176
rect 226076 201878 226196 201906
rect 226076 201414 226104 201878
rect 226154 201784 226210 201793
rect 226154 201719 226210 201728
rect 226064 201408 226116 201414
rect 226064 201350 226116 201356
rect 226062 200696 226118 200705
rect 226062 200631 226118 200640
rect 225972 198688 226024 198694
rect 225972 198630 226024 198636
rect 225880 197260 225932 197266
rect 225880 197202 225932 197208
rect 226076 195974 226104 200631
rect 226168 197334 226196 201719
rect 226260 200122 226288 204167
rect 226338 201240 226394 201249
rect 226338 201175 226394 201184
rect 226248 200116 226300 200122
rect 226248 200058 226300 200064
rect 226352 200002 226380 201175
rect 226260 199974 226380 200002
rect 226156 197328 226208 197334
rect 226156 197270 226208 197276
rect 226064 195968 226116 195974
rect 226064 195910 226116 195916
rect 226260 195906 226288 199974
rect 226430 199472 226486 199481
rect 226430 199407 226486 199416
rect 226338 198928 226394 198937
rect 226338 198863 226394 198872
rect 226352 198762 226380 198863
rect 226444 198830 226472 199407
rect 226432 198824 226484 198830
rect 226432 198766 226484 198772
rect 226340 198756 226392 198762
rect 226340 198698 226392 198704
rect 226430 198248 226486 198257
rect 226430 198183 226486 198192
rect 226338 197704 226394 197713
rect 226338 197639 226394 197648
rect 226352 197402 226380 197639
rect 226444 197470 226472 198183
rect 226432 197464 226484 197470
rect 226432 197406 226484 197412
rect 226340 197396 226392 197402
rect 226340 197338 226392 197344
rect 226614 197024 226670 197033
rect 226614 196959 226670 196968
rect 226628 196110 226656 196959
rect 226706 196480 226762 196489
rect 226706 196415 226762 196424
rect 226616 196104 226668 196110
rect 226616 196046 226668 196052
rect 226720 196042 226748 196415
rect 226708 196036 226760 196042
rect 226708 195978 226760 195984
rect 226338 195936 226394 195945
rect 226248 195900 226300 195906
rect 226338 195871 226394 195880
rect 226248 195842 226300 195848
rect 226352 194614 226380 195871
rect 226614 195256 226670 195265
rect 226614 195191 226670 195200
rect 226340 194608 226392 194614
rect 226340 194550 226392 194556
rect 225788 194540 225840 194546
rect 225788 194482 225840 194488
rect 226430 194168 226486 194177
rect 226430 194103 226486 194112
rect 226338 193488 226394 193497
rect 226338 193423 226394 193432
rect 226352 193254 226380 193423
rect 226444 193322 226472 194103
rect 226432 193316 226484 193322
rect 226432 193258 226484 193264
rect 226340 193248 226392 193254
rect 226340 193190 226392 193196
rect 226430 192944 226486 192953
rect 226430 192879 226486 192888
rect 226338 192400 226394 192409
rect 226338 192335 226394 192344
rect 224868 191956 224920 191962
rect 224868 191898 224920 191904
rect 224592 190460 224644 190466
rect 224592 190402 224644 190408
rect 224408 189032 224460 189038
rect 224408 188974 224460 188980
rect 224880 185706 224908 191898
rect 226352 191894 226380 192335
rect 226444 191962 226472 192879
rect 226432 191956 226484 191962
rect 226432 191898 226484 191904
rect 226340 191888 226392 191894
rect 226340 191830 226392 191836
rect 226338 191720 226394 191729
rect 226338 191655 226394 191664
rect 226352 190942 226380 191655
rect 226522 191176 226578 191185
rect 226628 191146 226656 195191
rect 226982 194712 227038 194721
rect 226982 194647 227038 194656
rect 226522 191111 226578 191120
rect 226616 191140 226668 191146
rect 226340 190936 226392 190942
rect 226340 190878 226392 190884
rect 226340 190528 226392 190534
rect 226338 190496 226340 190505
rect 226392 190496 226394 190505
rect 226338 190431 226394 190440
rect 226338 189952 226394 189961
rect 226338 189887 226394 189896
rect 225786 189408 225842 189417
rect 225786 189343 225842 189352
rect 225602 186960 225658 186969
rect 225602 186895 225658 186904
rect 224868 185700 224920 185706
rect 224868 185642 224920 185648
rect 224224 184952 224276 184958
rect 224224 184894 224276 184900
rect 222936 182300 222988 182306
rect 222936 182242 222988 182248
rect 222844 182164 222896 182170
rect 222844 182106 222896 182112
rect 221648 178628 221700 178634
rect 221648 178570 221700 178576
rect 222844 175296 222896 175302
rect 222844 175238 222896 175244
rect 221556 168632 221608 168638
rect 221556 168574 221608 168580
rect 221464 167612 221516 167618
rect 221464 167554 221516 167560
rect 220268 165844 220320 165850
rect 220268 165786 220320 165792
rect 218704 164144 218756 164150
rect 218704 164086 218756 164092
rect 214932 163396 214984 163402
rect 214932 163338 214984 163344
rect 217232 163396 217284 163402
rect 217232 163338 217284 163344
rect 214944 160177 214972 163338
rect 222856 162790 222884 175238
rect 222948 172514 222976 182242
rect 224236 175166 224264 184894
rect 224316 183660 224368 183666
rect 224316 183602 224368 183608
rect 224224 175160 224276 175166
rect 224224 175102 224276 175108
rect 224328 173874 224356 183602
rect 224960 178016 225012 178022
rect 224960 177958 225012 177964
rect 224972 175234 225000 177958
rect 225616 176662 225644 186895
rect 225800 180810 225828 189343
rect 226352 189106 226380 189887
rect 226340 189100 226392 189106
rect 226340 189042 226392 189048
rect 226338 188728 226394 188737
rect 226338 188663 226394 188672
rect 226352 187746 226380 188663
rect 226430 188184 226486 188193
rect 226430 188119 226486 188128
rect 226444 187814 226472 188119
rect 226432 187808 226484 187814
rect 226432 187750 226484 187756
rect 226340 187740 226392 187746
rect 226340 187682 226392 187688
rect 226338 187640 226394 187649
rect 226338 187575 226394 187584
rect 226352 186522 226380 187575
rect 226340 186516 226392 186522
rect 226340 186458 226392 186464
rect 226338 186416 226394 186425
rect 226338 186351 226340 186360
rect 226392 186351 226394 186360
rect 226340 186322 226392 186328
rect 226338 185872 226394 185881
rect 226338 185807 226394 185816
rect 226352 184958 226380 185807
rect 226536 185638 226564 191111
rect 226616 191082 226668 191088
rect 226996 189786 227024 194647
rect 226984 189780 227036 189786
rect 226984 189722 227036 189728
rect 226524 185632 226576 185638
rect 226524 185574 226576 185580
rect 226982 185192 227038 185201
rect 226982 185127 227038 185136
rect 226340 184952 226392 184958
rect 226340 184894 226392 184900
rect 226338 184648 226394 184657
rect 226338 184583 226394 184592
rect 226352 183598 226380 184583
rect 226522 184104 226578 184113
rect 226522 184039 226578 184048
rect 226536 183666 226564 184039
rect 226524 183660 226576 183666
rect 226524 183602 226576 183608
rect 226340 183592 226392 183598
rect 226340 183534 226392 183540
rect 226522 183424 226578 183433
rect 226522 183359 226578 183368
rect 226430 182880 226486 182889
rect 226430 182815 226486 182824
rect 226340 182232 226392 182238
rect 226338 182200 226340 182209
rect 226392 182200 226394 182209
rect 226338 182135 226394 182144
rect 226444 181490 226472 182815
rect 226536 182306 226564 183359
rect 226524 182300 226576 182306
rect 226524 182242 226576 182248
rect 226432 181484 226484 181490
rect 226432 181426 226484 181432
rect 226338 181112 226394 181121
rect 226338 181047 226394 181056
rect 226352 180946 226380 181047
rect 226340 180940 226392 180946
rect 226340 180882 226392 180888
rect 225788 180804 225840 180810
rect 225788 180746 225840 180752
rect 226338 180432 226394 180441
rect 226338 180367 226394 180376
rect 225696 179444 225748 179450
rect 225696 179386 225748 179392
rect 225604 176656 225656 176662
rect 225604 176598 225656 176604
rect 224960 175228 225012 175234
rect 224960 175170 225012 175176
rect 225604 173936 225656 173942
rect 225604 173878 225656 173884
rect 224316 173868 224368 173874
rect 224316 173810 224368 173816
rect 224316 173324 224368 173330
rect 224316 173266 224368 173272
rect 222936 172508 222988 172514
rect 222936 172450 222988 172456
rect 224328 165578 224356 173266
rect 224316 165572 224368 165578
rect 224316 165514 224368 165520
rect 225616 164218 225644 173878
rect 225708 169726 225736 179386
rect 226352 178702 226380 180367
rect 226430 179888 226486 179897
rect 226430 179823 226486 179832
rect 226444 179518 226472 179823
rect 226432 179512 226484 179518
rect 226432 179454 226484 179460
rect 226340 178696 226392 178702
rect 226340 178638 226392 178644
rect 226430 178664 226486 178673
rect 226430 178599 226486 178608
rect 226444 178090 226472 178599
rect 226706 178120 226762 178129
rect 226432 178084 226484 178090
rect 226706 178055 226762 178064
rect 226432 178026 226484 178032
rect 226338 177576 226394 177585
rect 226338 177511 226394 177520
rect 226352 176730 226380 177511
rect 226340 176724 226392 176730
rect 226340 176666 226392 176672
rect 226720 173330 226748 178055
rect 226996 178022 227024 185127
rect 227168 184884 227220 184890
rect 227168 184826 227220 184832
rect 227074 179344 227130 179353
rect 227074 179279 227130 179288
rect 226984 178016 227036 178022
rect 226984 177958 227036 177964
rect 226982 175808 227038 175817
rect 226982 175743 227038 175752
rect 226708 173324 226760 173330
rect 226708 173266 226760 173272
rect 225696 169720 225748 169726
rect 225696 169662 225748 169668
rect 225604 164212 225656 164218
rect 225604 164154 225656 164160
rect 226996 162858 227024 175743
rect 227088 167686 227116 179279
rect 227180 175642 227208 184826
rect 227626 181656 227682 181665
rect 227626 181591 227682 181600
rect 227640 179450 227668 181591
rect 227628 179444 227680 179450
rect 227628 179386 227680 179392
rect 227350 176896 227406 176905
rect 227350 176831 227406 176840
rect 227168 175636 227220 175642
rect 227168 175578 227220 175584
rect 227364 173942 227392 176831
rect 227442 176352 227498 176361
rect 227442 176287 227498 176296
rect 227456 175302 227484 176287
rect 227444 175296 227496 175302
rect 227444 175238 227496 175244
rect 227352 173936 227404 173942
rect 227352 173878 227404 173884
rect 227076 167680 227128 167686
rect 227076 167622 227128 167628
rect 226984 162852 227036 162858
rect 226984 162794 227036 162800
rect 215116 162784 215168 162790
rect 215116 162726 215168 162732
rect 222844 162784 222896 162790
rect 222844 162726 222896 162732
rect 215128 162625 215156 162726
rect 215114 162616 215170 162625
rect 215114 162551 215170 162560
rect 229756 161430 229784 223586
rect 235276 222494 235304 235175
rect 286336 224262 286364 569162
rect 287716 228410 287744 700538
rect 397472 700534 397500 703520
rect 305644 700528 305696 700534
rect 305644 700470 305696 700476
rect 397460 700528 397512 700534
rect 397460 700470 397512 700476
rect 304264 556232 304316 556238
rect 304264 556174 304316 556180
rect 302148 528080 302200 528086
rect 302148 528022 302200 528028
rect 288532 527944 288584 527950
rect 288532 527886 288584 527892
rect 288544 527814 288572 527886
rect 302160 527882 302188 528022
rect 302240 528012 302292 528018
rect 302240 527954 302292 527960
rect 302424 528012 302476 528018
rect 302424 527954 302476 527960
rect 302252 527898 302280 527954
rect 302436 527898 302464 527954
rect 302148 527876 302200 527882
rect 302252 527870 302464 527898
rect 302148 527818 302200 527824
rect 288532 527808 288584 527814
rect 288532 527750 288584 527756
rect 289728 500268 289780 500274
rect 289728 500210 289780 500216
rect 289636 438932 289688 438938
rect 289636 438874 289688 438880
rect 288898 317112 288954 317121
rect 288898 317047 288954 317056
rect 288912 316742 288940 317047
rect 288900 316736 288952 316742
rect 288900 316678 288952 316684
rect 289648 308961 289676 438874
rect 289740 325281 289768 500210
rect 299388 496120 299440 496126
rect 299388 496062 299440 496068
rect 299400 495514 299428 496062
rect 298100 495508 298152 495514
rect 298100 495450 298152 495456
rect 299388 495508 299440 495514
rect 299388 495450 299440 495456
rect 292580 421592 292632 421598
rect 292580 421534 292632 421540
rect 292592 329338 292620 421534
rect 298112 329338 298140 495450
rect 292592 329310 292988 329338
rect 298112 329310 298508 329338
rect 292960 329066 292988 329310
rect 298480 329066 298508 329310
rect 292960 329038 293526 329066
rect 298480 329038 298954 329066
rect 304276 328273 304304 556174
rect 304356 415472 304408 415478
rect 304356 415414 304408 415420
rect 304262 328264 304318 328273
rect 304262 328199 304318 328208
rect 303620 327072 303672 327078
rect 303620 327014 303672 327020
rect 303632 326369 303660 327014
rect 303618 326360 303674 326369
rect 303618 326295 303674 326304
rect 303620 325644 303672 325650
rect 303620 325586 303672 325592
rect 289726 325272 289782 325281
rect 289726 325207 289782 325216
rect 303632 324465 303660 325586
rect 303618 324456 303674 324465
rect 303618 324391 303674 324400
rect 304368 322561 304396 415414
rect 304448 368552 304500 368558
rect 304448 368494 304500 368500
rect 304354 322552 304410 322561
rect 304354 322487 304410 322496
rect 303620 321632 303672 321638
rect 303620 321574 303672 321580
rect 303632 318753 303660 321574
rect 304460 320657 304488 368494
rect 304446 320648 304502 320657
rect 304446 320583 304502 320592
rect 303618 318744 303674 318753
rect 303618 318679 303674 318688
rect 304354 316976 304410 316985
rect 304354 316911 304410 316920
rect 304262 315072 304318 315081
rect 304262 315007 304318 315016
rect 303618 313168 303674 313177
rect 303618 313103 303674 313112
rect 303632 311914 303660 313103
rect 303620 311908 303672 311914
rect 303620 311850 303672 311856
rect 303618 311264 303674 311273
rect 303618 311199 303674 311208
rect 303632 310554 303660 311199
rect 303620 310548 303672 310554
rect 303620 310490 303672 310496
rect 303618 309360 303674 309369
rect 303618 309295 303674 309304
rect 303632 309194 303660 309295
rect 303620 309188 303672 309194
rect 303620 309130 303672 309136
rect 289634 308952 289690 308961
rect 289634 308887 289690 308896
rect 303618 307456 303674 307465
rect 303618 307391 303674 307400
rect 303632 306406 303660 307391
rect 303620 306400 303672 306406
rect 303620 306342 303672 306348
rect 300860 305652 300912 305658
rect 300860 305594 300912 305600
rect 300872 305561 300900 305594
rect 300858 305552 300914 305561
rect 300858 305487 300914 305496
rect 292592 302841 292620 304844
rect 296180 303618 296208 304844
rect 299492 304830 299782 304858
rect 296168 303612 296220 303618
rect 296168 303554 296220 303560
rect 292578 302832 292634 302841
rect 292578 302767 292634 302776
rect 299492 233918 299520 304830
rect 299480 233912 299532 233918
rect 299480 233854 299532 233860
rect 304276 229090 304304 315007
rect 304368 276010 304396 316911
rect 304356 276004 304408 276010
rect 304356 275946 304408 275952
rect 305656 231130 305684 700470
rect 413664 700466 413692 703520
rect 313924 700460 313976 700466
rect 313924 700402 313976 700408
rect 413652 700460 413704 700466
rect 413652 700402 413704 700408
rect 308404 700392 308456 700398
rect 308404 700334 308456 700340
rect 305644 231124 305696 231130
rect 305644 231066 305696 231072
rect 308416 229770 308444 700334
rect 309784 700324 309836 700330
rect 309784 700266 309836 700272
rect 309046 473920 309102 473929
rect 309046 473855 309102 473864
rect 309060 473385 309088 473855
rect 309046 473376 309102 473385
rect 309046 473311 309102 473320
rect 308404 229764 308456 229770
rect 308404 229706 308456 229712
rect 304264 229084 304316 229090
rect 304264 229026 304316 229032
rect 287704 228404 287756 228410
rect 287704 228346 287756 228352
rect 309796 227050 309824 700266
rect 312544 627224 312596 627230
rect 312544 627166 312596 627172
rect 312556 613465 312584 627166
rect 312542 613456 312598 613465
rect 312542 613391 312598 613400
rect 312544 552084 312596 552090
rect 312544 552026 312596 552032
rect 312556 462777 312584 552026
rect 312542 462768 312598 462777
rect 312542 462703 312598 462712
rect 313278 439648 313334 439657
rect 313278 439583 313334 439592
rect 313292 438938 313320 439583
rect 313280 438932 313332 438938
rect 313280 438874 313332 438880
rect 313936 232558 313964 700402
rect 462332 700398 462360 703520
rect 478524 700505 478552 703520
rect 478510 700496 478566 700505
rect 478510 700431 478566 700440
rect 462320 700392 462372 700398
rect 462320 700334 462372 700340
rect 527192 700330 527220 703520
rect 543476 700369 543504 703520
rect 543462 700360 543518 700369
rect 527180 700324 527232 700330
rect 543462 700295 543518 700304
rect 527180 700266 527232 700272
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 576124 696992 576176 696998
rect 576124 696934 576176 696940
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 453304 681760 453356 681766
rect 453304 681702 453356 681708
rect 453316 616826 453344 681702
rect 506018 663912 506074 663921
rect 506018 663847 506074 663856
rect 506032 662388 506060 663847
rect 553398 649632 553454 649641
rect 553398 649567 553454 649576
rect 551742 638208 551798 638217
rect 551742 638143 551798 638152
rect 551374 636984 551430 636993
rect 551204 636942 551374 636970
rect 456062 635216 456118 635225
rect 456062 635151 456118 635160
rect 453304 616820 453356 616826
rect 453304 616762 453356 616768
rect 455418 591696 455474 591705
rect 455418 591631 455474 591640
rect 316894 570030 317368 570058
rect 317340 536246 317368 570030
rect 318536 570030 318642 570058
rect 318536 569974 318564 570030
rect 318524 569968 318576 569974
rect 318524 569910 318576 569916
rect 318708 569968 318760 569974
rect 318708 569910 318760 569916
rect 317328 536240 317380 536246
rect 317328 536182 317380 536188
rect 318720 533730 318748 569910
rect 320376 567254 320404 570044
rect 322230 570030 322888 570058
rect 323978 570030 324268 570058
rect 320364 567248 320416 567254
rect 320364 567190 320416 567196
rect 321468 567248 321520 567254
rect 321468 567190 321520 567196
rect 318708 533724 318760 533730
rect 318708 533666 318760 533672
rect 321284 533588 321336 533594
rect 321284 533530 321336 533536
rect 320732 533520 320784 533526
rect 320732 533462 320784 533468
rect 319628 533452 319680 533458
rect 319628 533394 319680 533400
rect 318524 533384 318576 533390
rect 318524 533326 318576 533332
rect 318536 528850 318564 533326
rect 319640 528850 319668 533394
rect 320744 528850 320772 533462
rect 318228 528822 318564 528850
rect 319332 528822 319668 528850
rect 320436 528822 320772 528850
rect 321296 528714 321324 533530
rect 321480 532098 321508 567190
rect 322860 545766 322888 570030
rect 324136 552696 324188 552702
rect 324136 552638 324188 552644
rect 322848 545760 322900 545766
rect 322848 545702 322900 545708
rect 322848 533656 322900 533662
rect 322848 533598 322900 533604
rect 321468 532092 321520 532098
rect 321468 532034 321520 532040
rect 322860 528850 322888 533598
rect 322552 528822 322888 528850
rect 324148 528714 324176 552638
rect 324240 543046 324268 570030
rect 325804 568274 325832 570044
rect 327552 568410 327580 570044
rect 327540 568404 327592 568410
rect 327540 568346 327592 568352
rect 328276 568404 328328 568410
rect 328276 568346 328328 568352
rect 325792 568268 325844 568274
rect 325792 568210 325844 568216
rect 326988 567860 327040 567866
rect 326988 567802 327040 567808
rect 326896 544400 326948 544406
rect 326896 544342 326948 544348
rect 324228 543040 324280 543046
rect 324228 542982 324280 542988
rect 325608 541680 325660 541686
rect 325608 541622 325660 541628
rect 325620 531078 325648 541622
rect 325056 531072 325108 531078
rect 325056 531014 325108 531020
rect 325608 531072 325660 531078
rect 325608 531014 325660 531020
rect 325068 528850 325096 531014
rect 326068 530936 326120 530942
rect 326068 530878 326120 530884
rect 326080 528850 326108 530878
rect 326908 528850 326936 544342
rect 327000 530942 327028 567802
rect 328288 533798 328316 568346
rect 329392 568342 329420 570044
rect 331048 570030 331154 570058
rect 329380 568336 329432 568342
rect 329380 568278 329432 568284
rect 328368 567928 328420 567934
rect 328368 567870 328420 567876
rect 328276 533792 328328 533798
rect 328276 533734 328328 533740
rect 326988 530936 327040 530942
rect 326988 530878 327040 530884
rect 328380 528850 328408 567870
rect 329748 551336 329800 551342
rect 329748 551278 329800 551284
rect 329760 531078 329788 551278
rect 331048 533866 331076 570030
rect 332980 568410 333008 570044
rect 334742 570030 335216 570058
rect 332968 568404 333020 568410
rect 332968 568346 333020 568352
rect 332508 568064 332560 568070
rect 332508 568006 332560 568012
rect 331128 567996 331180 568002
rect 331128 567938 331180 567944
rect 331036 533860 331088 533866
rect 331036 533802 331088 533808
rect 331140 531078 331168 567938
rect 332416 549908 332468 549914
rect 332416 549850 332468 549856
rect 332428 531282 332456 549850
rect 331496 531276 331548 531282
rect 331496 531218 331548 531224
rect 332416 531276 332468 531282
rect 332416 531218 332468 531224
rect 329288 531072 329340 531078
rect 329288 531014 329340 531020
rect 329748 531072 329800 531078
rect 329748 531014 329800 531020
rect 330392 531072 330444 531078
rect 330392 531014 330444 531020
rect 331128 531072 331180 531078
rect 331128 531014 331180 531020
rect 329300 528850 329328 531014
rect 330404 528850 330432 531014
rect 331508 528850 331536 531218
rect 332520 528850 332548 568006
rect 333888 548548 333940 548554
rect 333888 548490 333940 548496
rect 324760 528822 325096 528850
rect 325772 528822 326108 528850
rect 326876 528822 326936 528850
rect 327980 528822 328408 528850
rect 328992 528822 329328 528850
rect 330096 528822 330432 528850
rect 331200 528822 331536 528850
rect 332304 528822 332548 528850
rect 333900 528714 333928 548490
rect 335188 533934 335216 570030
rect 336568 568478 336596 570044
rect 338316 568546 338344 570044
rect 340156 568546 340184 570044
rect 341918 570030 342208 570058
rect 338304 568540 338356 568546
rect 338304 568482 338356 568488
rect 339316 568540 339368 568546
rect 339316 568482 339368 568488
rect 340144 568540 340196 568546
rect 340144 568482 340196 568488
rect 336556 568472 336608 568478
rect 336556 568414 336608 568420
rect 336648 568200 336700 568206
rect 336648 568142 336700 568148
rect 335268 568132 335320 568138
rect 335268 568074 335320 568080
rect 335176 533928 335228 533934
rect 335176 533870 335228 533876
rect 335280 531282 335308 568074
rect 336556 547188 336608 547194
rect 336556 547130 336608 547136
rect 336568 531282 336596 547130
rect 334716 531276 334768 531282
rect 334716 531218 334768 531224
rect 335268 531276 335320 531282
rect 335268 531218 335320 531224
rect 335820 531276 335872 531282
rect 335820 531218 335872 531224
rect 336556 531276 336608 531282
rect 336556 531218 336608 531224
rect 334728 528850 334756 531218
rect 335832 528850 335860 531218
rect 336660 528850 336688 568142
rect 339328 534002 339356 568482
rect 339408 565140 339460 565146
rect 339408 565082 339460 565088
rect 339316 533996 339368 534002
rect 339316 533938 339368 533944
rect 337936 532024 337988 532030
rect 337936 531966 337988 531972
rect 337948 528850 337976 531966
rect 339420 528986 339448 565082
rect 342076 563712 342128 563718
rect 342076 563654 342128 563660
rect 340052 532160 340104 532166
rect 340052 532102 340104 532108
rect 339144 528958 339448 528986
rect 339144 528850 339172 528958
rect 340064 528850 340092 532102
rect 340144 531820 340196 531826
rect 340144 531762 340196 531768
rect 340156 530806 340184 531762
rect 342088 531282 342116 563654
rect 342180 534070 342208 570030
rect 343744 567798 343772 570044
rect 343732 567792 343784 567798
rect 343732 567734 343784 567740
rect 345492 567730 345520 570044
rect 347332 567730 347360 570044
rect 345480 567724 345532 567730
rect 345480 567666 345532 567672
rect 346308 567724 346360 567730
rect 346308 567666 346360 567672
rect 347320 567724 347372 567730
rect 347320 567666 347372 567672
rect 346216 562352 346268 562358
rect 346216 562294 346268 562300
rect 343548 540252 343600 540258
rect 343548 540194 343600 540200
rect 342168 534064 342220 534070
rect 342168 534006 342220 534012
rect 342168 532228 342220 532234
rect 342168 532170 342220 532176
rect 341156 531276 341208 531282
rect 341156 531218 341208 531224
rect 342076 531276 342128 531282
rect 342076 531218 342128 531224
rect 340144 530800 340196 530806
rect 340144 530742 340196 530748
rect 341168 528850 341196 531218
rect 342180 528850 342208 532170
rect 334420 528822 334756 528850
rect 335524 528822 335860 528850
rect 336536 528822 336688 528850
rect 337640 528822 337976 528850
rect 338744 528822 339172 528850
rect 339848 528822 340092 528850
rect 340860 528822 341196 528850
rect 341964 528822 342208 528850
rect 343560 528714 343588 540194
rect 344376 532296 344428 532302
rect 344376 532238 344428 532244
rect 343640 531752 343692 531758
rect 343640 531694 343692 531700
rect 343652 530874 343680 531694
rect 343640 530868 343692 530874
rect 343640 530810 343692 530816
rect 344388 528850 344416 532238
rect 346228 531282 346256 562294
rect 346320 533322 346348 567666
rect 347688 560992 347740 560998
rect 347688 560934 347740 560940
rect 346308 533316 346360 533322
rect 346308 533258 346360 533264
rect 346308 532364 346360 532370
rect 346308 532306 346360 532312
rect 345480 531276 345532 531282
rect 345480 531218 345532 531224
rect 346216 531276 346268 531282
rect 346216 531218 346268 531224
rect 345492 528850 345520 531218
rect 346320 528850 346348 532306
rect 347700 528850 347728 560934
rect 349080 533254 349108 570044
rect 350920 567662 350948 570044
rect 352682 570030 353248 570058
rect 350908 567656 350960 567662
rect 350908 567598 350960 567604
rect 350448 559564 350500 559570
rect 350448 559506 350500 559512
rect 349068 533248 349120 533254
rect 349068 533190 349120 533196
rect 348700 532432 348752 532438
rect 348700 532374 348752 532380
rect 348712 528850 348740 532374
rect 349068 531684 349120 531690
rect 349068 531626 349120 531632
rect 349080 530942 349108 531626
rect 350460 531282 350488 559506
rect 351736 558204 351788 558210
rect 351736 558146 351788 558152
rect 350908 532500 350960 532506
rect 350908 532442 350960 532448
rect 349804 531276 349856 531282
rect 349804 531218 349856 531224
rect 350448 531276 350500 531282
rect 350448 531218 350500 531224
rect 349068 530936 349120 530942
rect 349068 530878 349120 530884
rect 348884 530528 348936 530534
rect 348884 530470 348936 530476
rect 348896 529650 348924 530470
rect 348884 529644 348936 529650
rect 348884 529586 348936 529592
rect 349816 528850 349844 531218
rect 350920 528850 350948 532442
rect 351748 528850 351776 558146
rect 353220 537538 353248 570030
rect 354416 570030 354522 570058
rect 354416 569974 354444 570030
rect 354404 569968 354456 569974
rect 354404 569910 354456 569916
rect 354588 569968 354640 569974
rect 354588 569910 354640 569916
rect 354496 555484 354548 555490
rect 354496 555426 354548 555432
rect 353208 537532 353260 537538
rect 353208 537474 353260 537480
rect 353024 532568 353076 532574
rect 353024 532510 353076 532516
rect 351920 531616 351972 531622
rect 351920 531558 351972 531564
rect 351932 531010 351960 531558
rect 351920 531004 351972 531010
rect 351920 530946 351972 530952
rect 353036 528850 353064 532510
rect 354508 531282 354536 555426
rect 354600 533186 354628 569910
rect 356256 567254 356284 570044
rect 358110 570030 358768 570058
rect 359858 570030 360148 570058
rect 356244 567248 356296 567254
rect 356244 567190 356296 567196
rect 357348 567248 357400 567254
rect 357348 567190 357400 567196
rect 355876 566500 355928 566506
rect 355876 566442 355928 566448
rect 354588 533180 354640 533186
rect 354588 533122 354640 533128
rect 355232 532636 355284 532642
rect 355232 532578 355284 532584
rect 354036 531276 354088 531282
rect 354036 531218 354088 531224
rect 354496 531276 354548 531282
rect 354496 531218 354548 531224
rect 354048 528850 354076 531218
rect 355244 528850 355272 532578
rect 355888 529122 355916 566442
rect 357360 538898 357388 567190
rect 358636 554056 358688 554062
rect 358636 553998 358688 554004
rect 357348 538892 357400 538898
rect 357348 538834 357400 538840
rect 357256 532704 357308 532710
rect 357256 532646 357308 532652
rect 355888 529094 355962 529122
rect 344080 528822 344416 528850
rect 345184 528822 345520 528850
rect 346288 528822 346348 528850
rect 347392 528822 347728 528850
rect 348404 528822 348740 528850
rect 349508 528822 349844 528850
rect 350612 528822 350948 528850
rect 351624 528822 351776 528850
rect 352728 528822 353064 528850
rect 353832 528822 354076 528850
rect 354936 528822 355272 528850
rect 355934 528836 355962 529094
rect 357268 528850 357296 532646
rect 357348 531548 357400 531554
rect 357348 531490 357400 531496
rect 357360 531078 357388 531490
rect 357348 531072 357400 531078
rect 357348 531014 357400 531020
rect 357052 528822 357296 528850
rect 358648 528714 358676 553998
rect 358740 534886 358768 570030
rect 360120 540326 360148 570030
rect 361684 567594 361712 570044
rect 363432 567594 363460 570044
rect 365194 570030 365668 570058
rect 361672 567588 361724 567594
rect 361672 567530 361724 567536
rect 362868 567588 362920 567594
rect 362868 567530 362920 567536
rect 363420 567588 363472 567594
rect 363420 567530 363472 567536
rect 364248 567588 364300 567594
rect 364248 567530 364300 567536
rect 360108 540320 360160 540326
rect 360108 540262 360160 540268
rect 362880 534954 362908 567530
rect 364260 541754 364288 567530
rect 364248 541748 364300 541754
rect 364248 541690 364300 541696
rect 363788 536308 363840 536314
rect 363788 536250 363840 536256
rect 362868 534948 362920 534954
rect 362868 534890 362920 534896
rect 358728 534880 358780 534886
rect 358728 534822 358780 534828
rect 362776 534812 362828 534818
rect 362776 534754 362828 534760
rect 360568 534744 360620 534750
rect 360568 534686 360620 534692
rect 359464 531956 359516 531962
rect 359464 531898 359516 531904
rect 359476 528850 359504 531898
rect 360580 528850 360608 534686
rect 361488 531888 361540 531894
rect 361488 531830 361540 531836
rect 361500 528850 361528 531830
rect 362788 528850 362816 534754
rect 363800 528850 363828 536250
rect 364892 535152 364944 535158
rect 364892 535094 364944 535100
rect 364904 528850 364932 535094
rect 365640 535022 365668 570030
rect 366916 545828 366968 545834
rect 366916 545770 366968 545776
rect 365628 535016 365680 535022
rect 365628 534958 365680 534964
rect 366928 531282 366956 545770
rect 367020 543318 367048 570044
rect 368492 570030 368782 570058
rect 369872 570030 370622 570058
rect 371252 570030 372370 570058
rect 374012 570030 374210 570058
rect 375392 570030 375958 570058
rect 376772 570030 377798 570058
rect 368388 543788 368440 543794
rect 368388 543730 368440 543736
rect 367008 543312 367060 543318
rect 367008 543254 367060 543260
rect 367008 534948 367060 534954
rect 367008 534890 367060 534896
rect 365996 531276 366048 531282
rect 365996 531218 366048 531224
rect 366916 531276 366968 531282
rect 366916 531218 366968 531224
rect 366008 528850 366036 531218
rect 367020 528850 367048 534890
rect 368400 528850 368428 543730
rect 359168 528822 359504 528850
rect 360272 528822 360608 528850
rect 361376 528822 361528 528850
rect 362480 528822 362816 528850
rect 363492 528822 363828 528850
rect 364596 528822 364932 528850
rect 365700 528822 366036 528850
rect 366712 528822 367048 528850
rect 367816 528822 368428 528850
rect 368492 528850 368520 570030
rect 369872 543794 369900 570030
rect 369860 543788 369912 543794
rect 369860 543730 369912 543736
rect 369860 543312 369912 543318
rect 369860 543254 369912 543260
rect 369872 528850 369900 543254
rect 370688 535016 370740 535022
rect 370688 534958 370740 534964
rect 370700 528850 370728 534958
rect 371252 534954 371280 570030
rect 374012 545834 374040 570030
rect 374000 545828 374052 545834
rect 374000 545770 374052 545776
rect 371332 541748 371384 541754
rect 371332 541690 371384 541696
rect 371240 534948 371292 534954
rect 371240 534890 371292 534896
rect 371344 528850 371372 541690
rect 374000 540320 374052 540326
rect 374000 540262 374052 540268
rect 372896 535084 372948 535090
rect 372896 535026 372948 535032
rect 372908 528850 372936 535026
rect 374012 528850 374040 540262
rect 375392 535022 375420 570030
rect 375472 538892 375524 538898
rect 375472 538834 375524 538840
rect 375380 535016 375432 535022
rect 375380 534958 375432 534964
rect 375380 534880 375432 534886
rect 375380 534822 375432 534828
rect 375392 528850 375420 534822
rect 368492 528822 368920 528850
rect 369872 528822 370024 528850
rect 370700 528822 371036 528850
rect 371344 528822 372140 528850
rect 372908 528822 373244 528850
rect 374012 528822 374256 528850
rect 375360 528822 375420 528850
rect 321296 528686 321448 528714
rect 323656 528686 324176 528714
rect 333316 528686 333928 528714
rect 343068 528686 343588 528714
rect 358156 528686 358676 528714
rect 375484 528714 375512 538834
rect 376772 536314 376800 570030
rect 379532 568562 379560 570044
rect 381004 570030 381386 570058
rect 382292 570030 383134 570058
rect 383672 570030 384974 570058
rect 386432 570030 386722 570058
rect 387812 570030 388562 570058
rect 389192 570030 390310 570058
rect 392044 570030 392150 570058
rect 393332 570030 393898 570058
rect 394804 570030 395738 570058
rect 379532 568534 379652 568562
rect 379520 567656 379572 567662
rect 379520 567598 379572 567604
rect 378232 537532 378284 537538
rect 378232 537474 378284 537480
rect 376760 536308 376812 536314
rect 376760 536250 376812 536256
rect 377220 533180 377272 533186
rect 377220 533122 377272 533128
rect 377232 528850 377260 533122
rect 378244 528850 378272 537474
rect 379532 528850 379560 567598
rect 379624 534818 379652 568534
rect 380900 567724 380952 567730
rect 380900 567666 380952 567672
rect 379612 534812 379664 534818
rect 379612 534754 379664 534760
rect 380440 533248 380492 533254
rect 380440 533190 380492 533196
rect 380452 528850 380480 533190
rect 380912 528986 380940 567666
rect 381004 531894 381032 570030
rect 382292 534750 382320 570030
rect 382280 534744 382332 534750
rect 382280 534686 382332 534692
rect 382556 533316 382608 533322
rect 382556 533258 382608 533264
rect 380992 531888 381044 531894
rect 380992 531830 381044 531836
rect 380912 528958 381400 528986
rect 381372 528850 381400 528958
rect 382568 528850 382596 533258
rect 383672 531962 383700 570030
rect 385040 568540 385092 568546
rect 385040 568482 385092 568488
rect 383752 567792 383804 567798
rect 383752 567734 383804 567740
rect 383660 531956 383712 531962
rect 383660 531898 383712 531904
rect 383764 528850 383792 567734
rect 385052 534154 385080 568482
rect 386432 554062 386460 570030
rect 386420 554056 386472 554062
rect 386420 553998 386472 554004
rect 385052 534126 385540 534154
rect 385132 534064 385184 534070
rect 385132 534006 385184 534012
rect 385144 528850 385172 534006
rect 377232 528822 377568 528850
rect 378244 528822 378580 528850
rect 379532 528822 379684 528850
rect 380452 528822 380788 528850
rect 381372 528822 381800 528850
rect 382568 528822 382904 528850
rect 383764 528822 384008 528850
rect 385112 528822 385172 528850
rect 385406 528864 385462 528873
rect 385512 528850 385540 534126
rect 386880 533996 386932 534002
rect 386880 533938 386932 533944
rect 386892 528850 386920 533938
rect 387812 532710 387840 570030
rect 387892 568472 387944 568478
rect 387892 568414 387944 568420
rect 387800 532704 387852 532710
rect 387800 532646 387852 532652
rect 387338 528864 387394 528873
rect 385512 528822 386124 528850
rect 386892 528822 387228 528850
rect 385406 528799 385462 528808
rect 387904 528850 387932 568414
rect 389192 566506 389220 570030
rect 389364 568404 389416 568410
rect 389364 568346 389416 568352
rect 389180 566500 389232 566506
rect 389180 566442 389232 566448
rect 389180 533928 389232 533934
rect 389180 533870 389232 533876
rect 389192 528850 389220 533870
rect 389376 528986 389404 568346
rect 391940 568336 391992 568342
rect 391940 568278 391992 568284
rect 391204 533860 391256 533866
rect 391204 533802 391256 533808
rect 389376 528958 390140 528986
rect 390112 528850 390140 528958
rect 391216 528850 391244 533802
rect 391952 528986 391980 568278
rect 392044 532642 392072 570030
rect 393332 555490 393360 570030
rect 394700 568268 394752 568274
rect 394700 568210 394752 568216
rect 393320 555484 393372 555490
rect 393320 555426 393372 555432
rect 393320 533792 393372 533798
rect 393320 533734 393372 533740
rect 392032 532636 392084 532642
rect 392032 532578 392084 532584
rect 391952 528958 392256 528986
rect 392228 528850 392256 528958
rect 393332 528850 393360 533734
rect 394712 529122 394740 568210
rect 394804 532574 394832 570030
rect 397472 558210 397500 570044
rect 398852 570030 399326 570058
rect 400232 570030 401074 570058
rect 401612 570030 402914 570058
rect 404372 570030 404662 570058
rect 405752 570030 406502 570058
rect 407132 570030 408250 570058
rect 409892 570030 409998 570058
rect 411272 570030 411838 570058
rect 412652 570030 413586 570058
rect 397460 558204 397512 558210
rect 397460 558146 397512 558152
rect 396080 545760 396132 545766
rect 396080 545702 396132 545708
rect 394884 543040 394936 543046
rect 394884 542982 394936 542988
rect 394792 532568 394844 532574
rect 394792 532510 394844 532516
rect 394712 529094 394786 529122
rect 387904 528822 388332 528850
rect 389192 528822 389344 528850
rect 390112 528822 390448 528850
rect 391216 528822 391552 528850
rect 392228 528822 392656 528850
rect 393332 528822 393668 528850
rect 394758 528836 394786 529094
rect 394896 528986 394924 542982
rect 396092 528986 396120 545702
rect 398852 532506 398880 570030
rect 400232 559570 400260 570030
rect 400220 559564 400272 559570
rect 400220 559506 400272 559512
rect 400220 536240 400272 536246
rect 400220 536182 400272 536188
rect 398932 533724 398984 533730
rect 398932 533666 398984 533672
rect 398840 532500 398892 532506
rect 398840 532442 398892 532448
rect 397644 532092 397696 532098
rect 397644 532034 397696 532040
rect 394896 528958 395568 528986
rect 396092 528958 396580 528986
rect 395540 528850 395568 528958
rect 396552 528850 396580 528958
rect 397656 528850 397684 532034
rect 398838 529000 398894 529009
rect 398838 528935 398894 528944
rect 395540 528822 395876 528850
rect 396552 528822 396888 528850
rect 397656 528822 397992 528850
rect 387338 528799 387394 528808
rect 375484 528686 376464 528714
rect 315396 528556 315448 528562
rect 315396 528498 315448 528504
rect 319628 528556 319680 528562
rect 319628 528498 319680 528504
rect 315302 528456 315358 528465
rect 315302 528391 315358 528400
rect 315210 528320 315266 528329
rect 315210 528255 315212 528264
rect 315264 528255 315266 528264
rect 315212 528226 315264 528232
rect 315316 527882 315344 528391
rect 315408 528222 315436 528498
rect 318064 528488 318116 528494
rect 318064 528430 318116 528436
rect 315396 528216 315448 528222
rect 315396 528158 315448 528164
rect 318076 528154 318104 528430
rect 319640 528290 319668 528498
rect 322020 528488 322072 528494
rect 320086 528456 320142 528465
rect 322020 528430 322072 528436
rect 320086 528391 320142 528400
rect 319628 528284 319680 528290
rect 319628 528226 319680 528232
rect 320100 528222 320128 528391
rect 322032 528222 322060 528430
rect 324148 528426 324268 528442
rect 324136 528420 324280 528426
rect 324188 528414 324228 528420
rect 324136 528362 324188 528368
rect 324228 528362 324280 528368
rect 324226 528320 324282 528329
rect 323952 528284 324004 528290
rect 324226 528255 324228 528264
rect 323952 528226 324004 528232
rect 324280 528255 324282 528264
rect 324228 528226 324280 528232
rect 320088 528216 320140 528222
rect 320088 528158 320140 528164
rect 322020 528216 322072 528222
rect 322020 528158 322072 528164
rect 323964 528170 323992 528226
rect 385420 528222 385448 528799
rect 385682 528728 385738 528737
rect 385682 528663 385738 528672
rect 386234 528728 386290 528737
rect 386234 528663 386290 528672
rect 385696 528426 385724 528663
rect 385958 528592 386014 528601
rect 385958 528527 386014 528536
rect 385866 528456 385922 528465
rect 385684 528420 385736 528426
rect 385866 528391 385922 528400
rect 385684 528362 385736 528368
rect 385776 528352 385828 528358
rect 385774 528320 385776 528329
rect 385828 528320 385830 528329
rect 385774 528255 385830 528264
rect 385880 528222 385908 528391
rect 385972 528290 386000 528527
rect 386248 528426 386276 528663
rect 386510 528592 386566 528601
rect 386510 528527 386566 528536
rect 386418 528456 386474 528465
rect 386236 528420 386288 528426
rect 386418 528391 386474 528400
rect 386236 528362 386288 528368
rect 386328 528352 386380 528358
rect 386326 528320 386328 528329
rect 386380 528320 386382 528329
rect 385960 528284 386012 528290
rect 386326 528255 386382 528264
rect 385960 528226 386012 528232
rect 386432 528222 386460 528391
rect 386524 528290 386552 528527
rect 386512 528284 386564 528290
rect 386512 528226 386564 528232
rect 387352 528222 387380 528799
rect 398852 528766 398880 528935
rect 398944 528850 398972 533666
rect 399206 529000 399262 529009
rect 399206 528935 399262 528944
rect 398944 528822 399096 528850
rect 399220 528766 399248 528935
rect 400232 528850 400260 536182
rect 401612 532438 401640 570030
rect 404372 560998 404400 570030
rect 404360 560992 404412 560998
rect 404360 560934 404412 560940
rect 401968 536172 402020 536178
rect 401968 536114 402020 536120
rect 401600 532432 401652 532438
rect 401600 532374 401652 532380
rect 401508 532092 401560 532098
rect 401508 532034 401560 532040
rect 401520 528850 401548 532034
rect 400200 528822 400260 528850
rect 401212 528822 401548 528850
rect 401980 528850 402008 536114
rect 403164 536104 403216 536110
rect 403164 536046 403216 536052
rect 403176 528850 403204 536046
rect 404452 534676 404504 534682
rect 404452 534618 404504 534624
rect 404464 528850 404492 534618
rect 405752 532370 405780 570030
rect 407132 562358 407160 570030
rect 407120 562352 407172 562358
rect 407120 562294 407172 562300
rect 407396 534608 407448 534614
rect 407396 534550 407448 534556
rect 405740 532364 405792 532370
rect 405740 532306 405792 532312
rect 405188 529576 405240 529582
rect 405188 529518 405240 529524
rect 401980 528822 402316 528850
rect 403176 528822 403420 528850
rect 404432 528822 404492 528850
rect 405200 528850 405228 529518
rect 407408 528850 407436 534550
rect 408592 532840 408644 532846
rect 408592 532782 408644 532788
rect 408604 528850 408632 532782
rect 409892 532302 409920 570030
rect 411272 540258 411300 570030
rect 411260 540252 411312 540258
rect 411260 540194 411312 540200
rect 410616 534540 410668 534546
rect 410616 534482 410668 534488
rect 409880 532296 409932 532302
rect 409880 532238 409932 532244
rect 409880 530732 409932 530738
rect 409880 530674 409932 530680
rect 409892 528850 409920 530674
rect 405200 528822 405536 528850
rect 407408 528822 407744 528850
rect 408604 528822 408756 528850
rect 409860 528822 409920 528850
rect 410628 528850 410656 534482
rect 412652 532234 412680 570030
rect 415412 563718 415440 570044
rect 416792 570030 417174 570058
rect 418172 570030 419014 570058
rect 419552 570030 420762 570058
rect 415400 563712 415452 563718
rect 415400 563654 415452 563660
rect 412640 532228 412692 532234
rect 412640 532170 412692 532176
rect 416792 532166 416820 570030
rect 418172 565146 418200 570030
rect 418160 565140 418212 565146
rect 418160 565082 418212 565088
rect 417056 534472 417108 534478
rect 417056 534414 417108 534420
rect 416780 532160 416832 532166
rect 416780 532102 416832 532108
rect 412732 531480 412784 531486
rect 412732 531422 412784 531428
rect 411628 530664 411680 530670
rect 411628 530606 411680 530612
rect 411640 528850 411668 530606
rect 412744 528850 412772 531422
rect 414020 530596 414072 530602
rect 414020 530538 414072 530544
rect 414032 528850 414060 530538
rect 415952 530460 416004 530466
rect 415952 530402 416004 530408
rect 415964 528850 415992 530402
rect 417068 528850 417096 534414
rect 419552 532030 419580 570030
rect 422588 568206 422616 570044
rect 423692 570030 424350 570058
rect 422576 568200 422628 568206
rect 422576 568142 422628 568148
rect 423692 547194 423720 570030
rect 426176 568138 426204 570044
rect 427832 570030 427938 570058
rect 426164 568132 426216 568138
rect 426164 568074 426216 568080
rect 427832 548554 427860 570030
rect 429764 568070 429792 570044
rect 430592 570030 431526 570058
rect 429752 568064 429804 568070
rect 429752 568006 429804 568012
rect 430592 549914 430620 570030
rect 433352 568002 433380 570044
rect 434732 570030 435114 570058
rect 433340 567996 433392 568002
rect 433340 567938 433392 567944
rect 434732 551342 434760 570030
rect 436940 567934 436968 570044
rect 437492 570030 438702 570058
rect 436928 567928 436980 567934
rect 436928 567870 436980 567876
rect 434720 551336 434772 551342
rect 434720 551278 434772 551284
rect 430580 549908 430632 549914
rect 430580 549850 430632 549856
rect 427820 548548 427872 548554
rect 427820 548490 427872 548496
rect 423680 547188 423732 547194
rect 423680 547130 423732 547136
rect 437492 544406 437520 570030
rect 440528 567866 440556 570044
rect 441632 570030 442290 570058
rect 443012 570030 444130 570058
rect 445772 570030 445878 570058
rect 447152 570030 447718 570058
rect 448532 570030 449466 570058
rect 440516 567860 440568 567866
rect 440516 567802 440568 567808
rect 437480 544400 437532 544406
rect 437480 544342 437532 544348
rect 441632 541686 441660 570030
rect 443012 552702 443040 570030
rect 443000 552696 443052 552702
rect 443000 552638 443052 552644
rect 441620 541680 441672 541686
rect 441620 541622 441672 541628
rect 431040 537396 431092 537402
rect 431040 537338 431092 537344
rect 419632 534404 419684 534410
rect 419632 534346 419684 534352
rect 419540 532024 419592 532030
rect 419540 531966 419592 531972
rect 418252 530800 418304 530806
rect 418252 530742 418304 530748
rect 418264 528850 418292 530742
rect 419448 529984 419500 529990
rect 419448 529926 419500 529932
rect 419460 529446 419488 529926
rect 419448 529440 419500 529446
rect 419448 529382 419500 529388
rect 419644 528850 419672 534346
rect 423680 534336 423732 534342
rect 423680 534278 423732 534284
rect 422484 530936 422536 530942
rect 422484 530878 422536 530884
rect 420276 530868 420328 530874
rect 420276 530810 420328 530816
rect 410628 528822 410964 528850
rect 411640 528822 411976 528850
rect 412744 528822 413080 528850
rect 414032 528822 414184 528850
rect 415964 528822 416300 528850
rect 417068 528822 417404 528850
rect 418264 528822 418508 528850
rect 419520 528822 419672 528850
rect 420288 528850 420316 530810
rect 421380 529508 421432 529514
rect 421380 529450 421432 529456
rect 421392 528850 421420 529450
rect 422496 528850 422524 530878
rect 423692 528850 423720 534278
rect 425704 534268 425756 534274
rect 425704 534210 425756 534216
rect 424600 531004 424652 531010
rect 424600 530946 424652 530952
rect 424612 528850 424640 530946
rect 425716 528850 425744 534210
rect 430028 534200 430080 534206
rect 430028 534142 430080 534148
rect 427912 532772 427964 532778
rect 427912 532714 427964 532720
rect 426716 531072 426768 531078
rect 426716 531014 426768 531020
rect 426728 528850 426756 531014
rect 427924 528850 427952 532714
rect 429292 529984 429344 529990
rect 429292 529926 429344 529932
rect 429304 528850 429332 529926
rect 420288 528822 420624 528850
rect 421392 528822 421728 528850
rect 422496 528822 422832 528850
rect 423692 528822 423844 528850
rect 424612 528822 424948 528850
rect 425716 528822 426052 528850
rect 426728 528822 427064 528850
rect 427924 528822 428168 528850
rect 429272 528822 429332 528850
rect 430040 528850 430068 534142
rect 431052 528850 431080 537338
rect 433340 537328 433392 537334
rect 433340 537270 433392 537276
rect 432144 534132 432196 534138
rect 432144 534074 432196 534080
rect 432156 528850 432184 534074
rect 433352 528850 433380 537270
rect 437572 537260 437624 537266
rect 437572 537202 437624 537208
rect 435362 533080 435418 533089
rect 435362 533015 435418 533024
rect 435376 528850 435404 533015
rect 437584 528850 437612 537202
rect 439688 537192 439740 537198
rect 439688 537134 439740 537140
rect 438950 532944 439006 532953
rect 438950 532879 439006 532888
rect 438964 528850 438992 532879
rect 430040 528822 430376 528850
rect 431052 528822 431388 528850
rect 432156 528822 432492 528850
rect 433352 528822 433596 528850
rect 435376 528822 435712 528850
rect 437584 528822 437920 528850
rect 438932 528822 438992 528850
rect 439700 528850 439728 537134
rect 444380 537124 444432 537130
rect 444380 537066 444432 537072
rect 441804 536036 441856 536042
rect 441804 535978 441856 535984
rect 440792 529372 440844 529378
rect 440792 529314 440844 529320
rect 440804 528850 440832 529314
rect 441816 528850 441844 535978
rect 444392 528850 444420 537066
rect 445772 533662 445800 570030
rect 446128 537056 446180 537062
rect 446128 536998 446180 537004
rect 445760 533656 445812 533662
rect 445760 533598 445812 533604
rect 439700 528822 440036 528850
rect 440804 528822 441140 528850
rect 441816 528822 442152 528850
rect 444360 528822 444420 528850
rect 446140 528850 446168 536998
rect 447152 533594 447180 570030
rect 447140 533588 447192 533594
rect 447140 533530 447192 533536
rect 448532 533526 448560 570030
rect 448704 536988 448756 536994
rect 448704 536930 448756 536936
rect 448520 533520 448572 533526
rect 448520 533462 448572 533468
rect 447232 529304 447284 529310
rect 447232 529246 447284 529252
rect 447244 528850 447272 529246
rect 448716 528850 448744 536930
rect 450452 536920 450504 536926
rect 450452 536862 450504 536868
rect 449440 531412 449492 531418
rect 449440 531354 449492 531360
rect 446140 528822 446476 528850
rect 447244 528822 447580 528850
rect 448684 528822 448744 528850
rect 449452 528850 449480 531354
rect 450464 528850 450492 536862
rect 451292 533458 451320 570044
rect 452672 570030 453054 570058
rect 451280 533452 451332 533458
rect 451280 533394 451332 533400
rect 452672 533390 452700 570030
rect 454774 534440 454830 534449
rect 454774 534375 454830 534384
rect 452660 533384 452712 533390
rect 452660 533326 452712 533332
rect 454040 531344 454092 531350
rect 454040 531286 454092 531292
rect 451556 529236 451608 529242
rect 451556 529178 451608 529184
rect 451568 528850 451596 529178
rect 454052 528850 454080 531286
rect 449452 528822 449788 528850
rect 450464 528822 450800 528850
rect 451568 528822 451904 528850
rect 454020 528822 454080 528850
rect 454788 528850 454816 534375
rect 455432 532098 455460 591631
rect 456076 568546 456104 635151
rect 456800 616820 456852 616826
rect 456800 616762 456852 616768
rect 456812 616321 456840 616762
rect 456798 616312 456854 616321
rect 456798 616247 456854 616256
rect 551100 616208 551152 616214
rect 551100 616150 551152 616156
rect 551112 606558 551140 616150
rect 551100 606552 551152 606558
rect 551100 606494 551152 606500
rect 551100 596896 551152 596902
rect 551100 596838 551152 596844
rect 551112 587246 551140 596838
rect 551100 587240 551152 587246
rect 551100 587182 551152 587188
rect 551100 577584 551152 577590
rect 551100 577526 551152 577532
rect 551112 572694 551140 577526
rect 551100 572688 551152 572694
rect 551100 572630 551152 572636
rect 525708 570512 525760 570518
rect 525708 570454 525760 570460
rect 483046 570030 483704 570058
rect 483676 568546 483704 570030
rect 456064 568540 456116 568546
rect 456064 568482 456116 568488
rect 483664 568540 483716 568546
rect 483664 568482 483716 568488
rect 483676 556510 483704 568482
rect 483664 556504 483716 556510
rect 483664 556446 483716 556452
rect 485780 556504 485832 556510
rect 485780 556446 485832 556452
rect 485792 554062 485820 556446
rect 485780 554056 485832 554062
rect 485780 553998 485832 554004
rect 498200 554056 498252 554062
rect 498200 553998 498252 554004
rect 498212 551342 498240 553998
rect 498200 551336 498252 551342
rect 498200 551278 498252 551284
rect 504364 551336 504416 551342
rect 504364 551278 504416 551284
rect 483848 536852 483900 536858
rect 483848 536794 483900 536800
rect 456984 535968 457036 535974
rect 456984 535910 457036 535916
rect 455420 532092 455472 532098
rect 455420 532034 455472 532040
rect 455880 529168 455932 529174
rect 455880 529110 455932 529116
rect 455892 528850 455920 529110
rect 456996 528850 457024 535910
rect 459100 535900 459152 535906
rect 459100 535842 459152 535848
rect 458178 531720 458234 531729
rect 458178 531655 458234 531664
rect 458192 528850 458220 531655
rect 459112 528850 459140 535842
rect 468760 535832 468812 535838
rect 468760 535774 468812 535780
rect 464526 534304 464582 534313
rect 464526 534239 464582 534248
rect 461214 531584 461270 531593
rect 461214 531519 461270 531528
rect 460526 529100 460578 529106
rect 460526 529042 460578 529048
rect 454788 528822 455124 528850
rect 455892 528822 456228 528850
rect 456996 528822 457332 528850
rect 458192 528822 458344 528850
rect 459112 528822 459448 528850
rect 460538 528836 460566 529042
rect 461228 528850 461256 531519
rect 463792 530392 463844 530398
rect 463792 530334 463844 530340
rect 462642 529032 462694 529038
rect 462642 528974 462694 528980
rect 461228 528822 461564 528850
rect 462654 528836 462682 528974
rect 463804 528850 463832 530334
rect 463772 528822 463832 528850
rect 464540 528850 464568 534239
rect 466642 532808 466698 532817
rect 466642 532743 466698 532752
rect 465540 530324 465592 530330
rect 465540 530266 465592 530272
rect 465552 528850 465580 530266
rect 466656 528850 466684 532743
rect 467840 530256 467892 530262
rect 467840 530198 467892 530204
rect 467852 528850 467880 530198
rect 468772 528850 468800 535774
rect 470968 535764 471020 535770
rect 470968 535706 471020 535712
rect 469864 530188 469916 530194
rect 469864 530130 469916 530136
rect 469876 528850 469904 530130
rect 470980 528850 471008 535706
rect 473452 535696 473504 535702
rect 473452 535638 473504 535644
rect 472072 530120 472124 530126
rect 472072 530062 472124 530068
rect 472084 528850 472112 530062
rect 473464 528850 473492 535638
rect 475292 535628 475344 535634
rect 475292 535570 475344 535576
rect 474188 530052 474240 530058
rect 474188 529994 474240 530000
rect 464540 528822 464876 528850
rect 465552 528822 465888 528850
rect 466656 528822 466992 528850
rect 467852 528822 468096 528850
rect 468772 528822 469108 528850
rect 469876 528822 470212 528850
rect 470980 528822 471316 528850
rect 472084 528822 472420 528850
rect 473432 528822 473492 528850
rect 474200 528850 474228 529994
rect 475304 528850 475332 535570
rect 478880 535560 478932 535566
rect 478880 535502 478932 535508
rect 477500 531140 477552 531146
rect 477500 531082 477552 531088
rect 476304 528964 476356 528970
rect 476304 528906 476356 528912
rect 476316 528850 476344 528906
rect 477512 528850 477540 531082
rect 478892 528850 478920 535502
rect 483664 535492 483716 535498
rect 483664 535434 483716 535440
rect 481730 534168 481786 534177
rect 481730 534103 481786 534112
rect 480628 529644 480680 529650
rect 480628 529586 480680 529592
rect 474200 528822 474536 528850
rect 475304 528822 475640 528850
rect 476316 528822 476652 528850
rect 477512 528822 477756 528850
rect 478860 528822 478920 528850
rect 479616 528896 479668 528902
rect 480640 528850 480668 529586
rect 481744 528850 481772 534103
rect 483676 531282 483704 535434
rect 483664 531276 483716 531282
rect 483664 531218 483716 531224
rect 483860 528850 483888 536794
rect 501786 533488 501842 533497
rect 501786 533423 501842 533432
rect 499394 533352 499450 533361
rect 499394 533287 499450 533296
rect 498566 532400 498622 532409
rect 498566 532335 498622 532344
rect 496358 532128 496414 532137
rect 496358 532063 496414 532072
rect 484950 531448 485006 531457
rect 484950 531383 485006 531392
rect 484964 528850 484992 531383
rect 493046 531312 493102 531321
rect 487160 531276 487212 531282
rect 493046 531247 493102 531256
rect 487160 531218 487212 531224
rect 487172 528850 487200 531218
rect 492034 531176 492090 531185
rect 492034 531111 492090 531120
rect 490378 529952 490434 529961
rect 490378 529887 490434 529896
rect 490392 528850 490420 529887
rect 492048 528850 492076 531111
rect 493060 528850 493088 531247
rect 495346 530632 495402 530641
rect 495346 530567 495402 530576
rect 493782 529952 493838 529961
rect 493782 529887 493838 529896
rect 479668 528844 479964 528850
rect 479616 528838 479964 528844
rect 479628 528822 479964 528838
rect 480640 528822 480976 528850
rect 481744 528822 482080 528850
rect 483032 528834 483184 528850
rect 483020 528828 483184 528834
rect 483072 528822 483184 528828
rect 483860 528822 484196 528850
rect 484964 528822 485300 528850
rect 487172 528822 487508 528850
rect 490392 528822 490728 528850
rect 491740 528822 492076 528850
rect 492844 528822 493088 528850
rect 483020 528770 483072 528776
rect 398840 528760 398892 528766
rect 398840 528702 398892 528708
rect 399208 528760 399260 528766
rect 399208 528702 399260 528708
rect 486056 528760 486108 528766
rect 493796 528714 493824 529887
rect 495360 528850 495388 530567
rect 496372 528850 496400 532063
rect 497462 531992 497518 532001
rect 497462 531927 497518 531936
rect 497476 528850 497504 531927
rect 498580 528850 498608 532335
rect 499408 528850 499436 533287
rect 500682 532264 500738 532273
rect 500682 532199 500738 532208
rect 500696 528850 500724 532199
rect 501800 528850 501828 533423
rect 503628 533384 503680 533390
rect 503628 533326 503680 533332
rect 502890 532536 502946 532545
rect 502890 532471 502946 532480
rect 502904 528850 502932 532471
rect 503640 528850 503668 533326
rect 504376 532710 504404 551278
rect 520186 547088 520242 547097
rect 520186 547023 520242 547032
rect 518716 533860 518768 533866
rect 518716 533802 518768 533808
rect 516876 533792 516928 533798
rect 516876 533734 516928 533740
rect 514668 533724 514720 533730
rect 514668 533666 514720 533672
rect 512552 533656 512604 533662
rect 506110 533624 506166 533633
rect 512552 533598 512604 533604
rect 506110 533559 506166 533568
rect 510436 533588 510488 533594
rect 504364 532704 504416 532710
rect 504364 532646 504416 532652
rect 505008 530596 505060 530602
rect 505008 530538 505060 530544
rect 505020 528850 505048 530538
rect 506124 528850 506152 533559
rect 510436 533530 510488 533536
rect 508228 533452 508280 533458
rect 508228 533394 508280 533400
rect 507122 532672 507178 532681
rect 507122 532607 507178 532616
rect 507136 528850 507164 532607
rect 508240 528850 508268 533394
rect 508504 532704 508556 532710
rect 508504 532646 508556 532652
rect 495052 528822 495388 528850
rect 496064 528822 496400 528850
rect 497168 528822 497504 528850
rect 498272 528822 498608 528850
rect 499284 528822 499436 528850
rect 500388 528822 500724 528850
rect 501492 528822 501828 528850
rect 502596 528822 502932 528850
rect 503608 528822 503668 528850
rect 504712 528822 505048 528850
rect 505816 528822 506152 528850
rect 506828 528822 507164 528850
rect 507932 528822 508268 528850
rect 486108 528708 486404 528714
rect 486056 528702 486404 528708
rect 398932 528692 398984 528698
rect 398932 528634 398984 528640
rect 403624 528692 403676 528698
rect 486068 528686 486404 528702
rect 488368 528698 488520 528714
rect 488356 528692 488520 528698
rect 403624 528634 403676 528640
rect 488408 528686 488520 528692
rect 493796 528686 493948 528714
rect 488356 528634 488408 528640
rect 398838 528592 398894 528601
rect 398838 528527 398840 528536
rect 398892 528527 398894 528536
rect 398840 528498 398892 528504
rect 398944 528494 398972 528634
rect 403636 528494 403664 528634
rect 411260 528624 411312 528630
rect 403714 528592 403770 528601
rect 411444 528624 411496 528630
rect 411312 528584 411444 528612
rect 411260 528566 411312 528572
rect 411444 528566 411496 528572
rect 489276 528624 489328 528630
rect 489328 528572 489624 528578
rect 489276 528566 489624 528572
rect 489288 528550 489624 528566
rect 403714 528527 403770 528536
rect 403728 528494 403756 528527
rect 398932 528488 398984 528494
rect 398932 528430 398984 528436
rect 403624 528488 403676 528494
rect 403624 528430 403676 528436
rect 403716 528488 403768 528494
rect 408224 528488 408276 528494
rect 403716 528430 403768 528436
rect 406304 528426 406640 528442
rect 443368 528488 443420 528494
rect 408224 528430 408276 528436
rect 422298 528456 422354 528465
rect 406292 528420 406640 528426
rect 406344 528414 406640 528420
rect 406292 528362 406344 528368
rect 408236 528329 408264 528430
rect 422298 528391 422300 528400
rect 422352 528391 422354 528400
rect 431774 528456 431830 528465
rect 434732 528426 434852 528442
rect 443368 528430 443420 528436
rect 431774 528391 431830 528400
rect 431868 528420 431920 528426
rect 422300 528362 422352 528368
rect 414940 528352 414992 528358
rect 408222 528320 408278 528329
rect 422208 528352 422260 528358
rect 422206 528320 422208 528329
rect 422260 528320 422262 528329
rect 414992 528300 415288 528306
rect 414940 528294 415288 528300
rect 414952 528278 415288 528294
rect 408222 528255 408278 528264
rect 431788 528306 431816 528391
rect 431868 528362 431920 528368
rect 434720 528420 434864 528426
rect 434772 528414 434812 528420
rect 434720 528362 434772 528368
rect 434812 528362 434864 528368
rect 431880 528306 431908 528362
rect 431788 528278 431908 528306
rect 434272 528290 434608 528306
rect 434260 528284 434608 528290
rect 422206 528255 422262 528264
rect 434312 528278 434608 528284
rect 434260 528226 434312 528232
rect 443380 528222 443408 528430
rect 508516 528329 508544 532646
rect 509054 530768 509110 530777
rect 509054 530703 509110 530712
rect 509068 528850 509096 530703
rect 510448 528850 510476 533530
rect 511446 531856 511502 531865
rect 511446 531791 511502 531800
rect 511460 528850 511488 531791
rect 512564 528850 512592 533598
rect 513656 532024 513708 532030
rect 513656 531966 513708 531972
rect 513668 528850 513696 531966
rect 514680 528850 514708 533666
rect 515770 531720 515826 531729
rect 515770 531655 515826 531664
rect 515784 528850 515812 531655
rect 516888 528850 516916 533734
rect 517980 532092 518032 532098
rect 517980 532034 518032 532040
rect 517992 528850 518020 532034
rect 518728 528850 518756 533802
rect 520200 528850 520228 547023
rect 524328 538892 524380 538898
rect 524328 538834 524380 538840
rect 521200 532160 521252 532166
rect 521200 532102 521252 532108
rect 521212 528850 521240 532102
rect 524234 530904 524290 530913
rect 523316 530868 523368 530874
rect 524340 530874 524368 538834
rect 524234 530839 524290 530848
rect 524328 530868 524380 530874
rect 523316 530810 523368 530816
rect 522212 530664 522264 530670
rect 522212 530606 522264 530612
rect 522224 528850 522252 530606
rect 523328 528850 523356 530810
rect 524248 528850 524276 530839
rect 524328 530810 524380 530816
rect 525720 528986 525748 570454
rect 543648 570444 543700 570450
rect 543648 570386 543700 570392
rect 529032 567254 529060 570044
rect 529020 567248 529072 567254
rect 529020 567190 529072 567196
rect 530584 567248 530636 567254
rect 530584 567190 530636 567196
rect 528468 563712 528520 563718
rect 528468 563654 528520 563660
rect 527088 547188 527140 547194
rect 527088 547130 527140 547136
rect 527100 531282 527128 547130
rect 528480 531282 528508 563654
rect 529848 559564 529900 559570
rect 529848 559506 529900 559512
rect 526536 531276 526588 531282
rect 526536 531218 526588 531224
rect 527088 531276 527140 531282
rect 527088 531218 527140 531224
rect 527640 531276 527692 531282
rect 527640 531218 527692 531224
rect 528468 531276 528520 531282
rect 528468 531218 528520 531224
rect 525536 528958 525748 528986
rect 525536 528850 525564 528958
rect 526548 528850 526576 531218
rect 527652 528850 527680 531218
rect 528468 530732 528520 530738
rect 528468 530674 528520 530680
rect 528480 528850 528508 530674
rect 529860 528850 529888 559506
rect 530596 533526 530624 567190
rect 532608 565140 532660 565146
rect 532608 565082 532660 565088
rect 531228 547256 531280 547262
rect 531228 547198 531280 547204
rect 530584 533520 530636 533526
rect 530584 533462 530636 533468
rect 531240 531282 531268 547198
rect 532620 531282 532648 565082
rect 538128 562352 538180 562358
rect 538128 562294 538180 562300
rect 533988 560992 534040 560998
rect 533988 560934 534040 560940
rect 530860 531276 530912 531282
rect 530860 531218 530912 531224
rect 531228 531276 531280 531282
rect 531228 531218 531280 531224
rect 531964 531276 532016 531282
rect 531964 531218 532016 531224
rect 532608 531276 532660 531282
rect 532608 531218 532660 531224
rect 530872 528850 530900 531218
rect 531976 528850 532004 531218
rect 533068 530800 533120 530806
rect 533068 530742 533120 530748
rect 533080 528850 533108 530742
rect 534000 528850 534028 560934
rect 536748 551336 536800 551342
rect 536748 551278 536800 551284
rect 536760 531282 536788 551278
rect 536288 531276 536340 531282
rect 536288 531218 536340 531224
rect 536748 531276 536800 531282
rect 536748 531218 536800 531224
rect 535184 530868 535236 530874
rect 535184 530810 535236 530816
rect 535196 528850 535224 530810
rect 536300 528850 536328 531218
rect 537300 530936 537352 530942
rect 537300 530878 537352 530884
rect 537312 528850 537340 530878
rect 538140 528850 538168 562294
rect 540888 552696 540940 552702
rect 540888 552638 540940 552644
rect 539508 531004 539560 531010
rect 539508 530946 539560 530952
rect 539520 528850 539548 530946
rect 540900 528986 540928 552638
rect 543556 531140 543608 531146
rect 543556 531082 543608 531088
rect 541624 531072 541676 531078
rect 541624 531014 541676 531020
rect 540624 528958 540928 528986
rect 540624 528850 540652 528958
rect 541636 528850 541664 531014
rect 542728 530188 542780 530194
rect 542728 530130 542780 530136
rect 542740 528850 542768 530130
rect 543568 528850 543596 531082
rect 543660 530194 543688 570386
rect 547788 569968 547840 569974
rect 547788 569910 547840 569916
rect 544844 531344 544896 531350
rect 544844 531286 544896 531292
rect 543648 530188 543700 530194
rect 543648 530130 543700 530136
rect 544856 528850 544884 531286
rect 545580 531276 545632 531282
rect 545580 531218 545632 531224
rect 545592 530738 545620 531218
rect 545948 531072 546000 531078
rect 545948 531014 546000 531020
rect 545764 531004 545816 531010
rect 545764 530946 545816 530952
rect 545776 530874 545804 530946
rect 545672 530868 545724 530874
rect 545672 530810 545724 530816
rect 545764 530868 545816 530874
rect 545764 530810 545816 530816
rect 545684 530738 545712 530810
rect 545580 530732 545632 530738
rect 545580 530674 545632 530680
rect 545672 530732 545724 530738
rect 545672 530674 545724 530680
rect 545960 528850 545988 531014
rect 547800 530194 547828 569910
rect 549168 568608 549220 568614
rect 549168 568550 549220 568556
rect 549076 547732 549128 547738
rect 549076 547674 549128 547680
rect 549088 530194 549116 547674
rect 547052 530188 547104 530194
rect 547052 530130 547104 530136
rect 547788 530188 547840 530194
rect 547788 530130 547840 530136
rect 548156 530188 548208 530194
rect 548156 530130 548208 530136
rect 549076 530188 549128 530194
rect 549076 530130 549128 530136
rect 547064 528850 547092 530130
rect 548168 528850 548196 530130
rect 549180 528850 549208 568550
rect 551006 567760 551062 567769
rect 551006 567695 551062 567704
rect 551020 559201 551048 567695
rect 551100 563100 551152 563106
rect 551100 563042 551152 563048
rect 551006 559192 551062 559201
rect 551006 559127 551062 559136
rect 551112 558906 551140 563042
rect 551020 558878 551140 558906
rect 551020 553450 551048 558878
rect 551008 553444 551060 553450
rect 551008 553386 551060 553392
rect 551100 553376 551152 553382
rect 551100 553318 551152 553324
rect 551112 549302 551140 553318
rect 551008 549296 551060 549302
rect 551008 549238 551060 549244
rect 551100 549296 551152 549302
rect 551100 549238 551152 549244
rect 550548 547120 550600 547126
rect 550548 547062 550600 547068
rect 509036 528822 509096 528850
rect 510140 528822 510476 528850
rect 511152 528822 511488 528850
rect 512256 528822 512592 528850
rect 513360 528822 513696 528850
rect 514372 528822 514708 528850
rect 515476 528822 515812 528850
rect 516580 528822 516916 528850
rect 517684 528822 518020 528850
rect 518696 528822 518756 528850
rect 519800 528822 520228 528850
rect 520904 528822 521240 528850
rect 521916 528822 522252 528850
rect 523020 528822 523356 528850
rect 524124 528822 524276 528850
rect 525228 528822 525564 528850
rect 526240 528822 526576 528850
rect 527344 528822 527680 528850
rect 528448 528822 528508 528850
rect 529460 528822 529888 528850
rect 530564 528822 530900 528850
rect 531668 528822 532004 528850
rect 532772 528822 533108 528850
rect 533784 528822 534028 528850
rect 534888 528822 535224 528850
rect 535992 528822 536328 528850
rect 537004 528822 537340 528850
rect 538108 528822 538168 528850
rect 539212 528822 539548 528850
rect 540316 528822 540652 528850
rect 541328 528822 541664 528850
rect 542432 528822 542768 528850
rect 543536 528822 543596 528850
rect 544548 528822 544884 528850
rect 545652 528822 545988 528850
rect 546756 528822 547092 528850
rect 547860 528822 548196 528850
rect 548872 528822 549208 528850
rect 550560 528714 550588 547062
rect 551020 543810 551048 549238
rect 550928 543782 551048 543810
rect 550928 539617 550956 543782
rect 550730 539608 550786 539617
rect 550730 539543 550786 539552
rect 550914 539608 550970 539617
rect 550914 539543 550970 539552
rect 550744 532030 550772 539543
rect 551204 533730 551232 636942
rect 551374 636919 551430 636928
rect 551374 633584 551430 633593
rect 551296 633542 551374 633570
rect 551192 533724 551244 533730
rect 551192 533666 551244 533672
rect 551296 532098 551324 633542
rect 551374 633519 551430 633528
rect 551466 630864 551522 630873
rect 551466 630799 551522 630808
rect 551374 628416 551430 628425
rect 551374 628351 551430 628360
rect 551284 532092 551336 532098
rect 551284 532034 551336 532040
rect 550732 532024 550784 532030
rect 550732 531966 550784 531972
rect 551388 531298 551416 628351
rect 551480 628017 551508 630799
rect 551466 628008 551522 628017
rect 551466 627943 551522 627952
rect 551558 623792 551614 623801
rect 551558 623727 551614 623736
rect 551466 616312 551522 616321
rect 551466 616247 551522 616256
rect 551296 531270 551416 531298
rect 551296 530670 551324 531270
rect 551376 531140 551428 531146
rect 551376 531082 551428 531088
rect 551284 530664 551336 530670
rect 551284 530606 551336 530612
rect 551388 528850 551416 531082
rect 551480 530806 551508 616247
rect 551572 547194 551600 623727
rect 551650 618624 551706 618633
rect 551650 618559 551706 618568
rect 551664 547262 551692 618559
rect 551756 616214 551784 638143
rect 552018 621344 552074 621353
rect 552018 621279 552074 621288
rect 551834 616312 551890 616321
rect 551834 616247 551890 616256
rect 551744 616208 551796 616214
rect 551744 616150 551796 616156
rect 551848 612921 551876 616247
rect 551834 612912 551890 612921
rect 551834 612847 551890 612856
rect 551836 606552 551888 606558
rect 551836 606494 551888 606500
rect 551742 603120 551798 603129
rect 551742 603055 551798 603064
rect 551652 547256 551704 547262
rect 551652 547198 551704 547204
rect 551560 547188 551612 547194
rect 551560 547130 551612 547136
rect 551756 531350 551784 603055
rect 551848 596902 551876 606494
rect 551926 604344 551982 604353
rect 551926 604279 551982 604288
rect 551940 603090 551968 604279
rect 551928 603084 551980 603090
rect 551928 603026 551980 603032
rect 551836 596896 551888 596902
rect 551836 596838 551888 596844
rect 551836 596760 551888 596766
rect 551836 596702 551888 596708
rect 551848 588577 551876 596702
rect 551834 588568 551890 588577
rect 551834 588503 551890 588512
rect 551836 587240 551888 587246
rect 551836 587182 551888 587188
rect 551848 577590 551876 587182
rect 551836 577584 551888 577590
rect 551836 577526 551888 577532
rect 551836 572688 551888 572694
rect 551836 572630 551888 572636
rect 551848 563106 551876 572630
rect 551928 571260 551980 571266
rect 551928 571202 551980 571208
rect 551836 563100 551888 563106
rect 551836 563042 551888 563048
rect 551744 531344 551796 531350
rect 551744 531286 551796 531292
rect 551940 531146 551968 571202
rect 552032 531282 552060 621279
rect 552110 614408 552166 614417
rect 552110 614343 552166 614352
rect 552020 531276 552072 531282
rect 552020 531218 552072 531224
rect 551928 531140 551980 531146
rect 551928 531082 551980 531088
rect 551468 530800 551520 530806
rect 551468 530742 551520 530748
rect 552124 530738 552152 614343
rect 552202 611960 552258 611969
rect 552202 611895 552258 611904
rect 552216 530942 552244 611895
rect 552294 609512 552350 609521
rect 552294 609447 552350 609456
rect 552204 530936 552256 530942
rect 552204 530878 552256 530884
rect 552308 530874 552336 609447
rect 552386 607064 552442 607073
rect 552386 606999 552442 607008
rect 552400 531010 552428 606999
rect 552478 604616 552534 604625
rect 552478 604551 552534 604560
rect 552492 531214 552520 604551
rect 552664 603084 552716 603090
rect 552664 603026 552716 603032
rect 552570 602168 552626 602177
rect 552570 602103 552626 602112
rect 552480 531208 552532 531214
rect 552480 531150 552532 531156
rect 552584 531078 552612 602103
rect 552676 596766 552704 603026
rect 552938 600944 552994 600953
rect 552938 600879 552994 600888
rect 552754 599720 552810 599729
rect 552754 599655 552810 599664
rect 552664 596760 552716 596766
rect 552664 596702 552716 596708
rect 552662 594824 552718 594833
rect 552662 594759 552718 594768
rect 552572 531072 552624 531078
rect 552572 531014 552624 531020
rect 552388 531004 552440 531010
rect 552388 530946 552440 530952
rect 552296 530868 552348 530874
rect 552296 530810 552348 530816
rect 552112 530732 552164 530738
rect 552112 530674 552164 530680
rect 552676 528986 552704 594759
rect 552768 547738 552796 599655
rect 552846 597272 552902 597281
rect 552846 597207 552902 597216
rect 552756 547732 552808 547738
rect 552756 547674 552808 547680
rect 552860 547126 552888 597207
rect 552952 569974 552980 600879
rect 553030 598496 553086 598505
rect 553030 598431 553086 598440
rect 552940 569968 552992 569974
rect 552940 569910 552992 569916
rect 553044 568614 553072 598431
rect 553032 568608 553084 568614
rect 553032 568550 553084 568556
rect 552848 547120 552900 547126
rect 552848 547062 552900 547068
rect 553412 533390 553440 649567
rect 554410 648408 554466 648417
rect 554410 648343 554466 648352
rect 554424 647290 554452 648343
rect 554412 647284 554464 647290
rect 554412 647226 554464 647232
rect 556252 647284 556304 647290
rect 556252 647226 556304 647232
rect 553490 644736 553546 644745
rect 553490 644671 553546 644680
rect 553504 533458 553532 644671
rect 554042 643512 554098 643521
rect 554042 643447 554098 643456
rect 553582 642288 553638 642297
rect 553582 642223 553638 642232
rect 553596 533594 553624 642223
rect 553674 639976 553730 639985
rect 553674 639911 553730 639920
rect 553688 533662 553716 639911
rect 553766 635080 553822 635089
rect 553766 635015 553822 635024
rect 553780 533798 553808 635015
rect 553858 632632 553914 632641
rect 553858 632567 553914 632576
rect 553872 533866 553900 632567
rect 553950 630184 554006 630193
rect 553950 630119 554006 630128
rect 553860 533860 553912 533866
rect 553860 533802 553912 533808
rect 553768 533792 553820 533798
rect 553768 533734 553820 533740
rect 553676 533656 553728 533662
rect 553676 533598 553728 533604
rect 553584 533588 553636 533594
rect 553584 533530 553636 533536
rect 553492 533452 553544 533458
rect 553492 533394 553544 533400
rect 553400 533384 553452 533390
rect 553400 533326 553452 533332
rect 553964 532166 553992 630119
rect 554056 594017 554084 643447
rect 554870 627736 554926 627745
rect 554870 627671 554926 627680
rect 554226 625288 554282 625297
rect 554226 625223 554282 625232
rect 554134 610736 554190 610745
rect 554134 610671 554190 610680
rect 554148 610026 554176 610671
rect 554136 610020 554188 610026
rect 554136 609962 554188 609968
rect 554042 594008 554098 594017
rect 554042 593943 554098 593952
rect 554042 593736 554098 593745
rect 554042 593671 554098 593680
rect 553952 532160 554004 532166
rect 553952 532102 554004 532108
rect 554056 531282 554084 593671
rect 554134 592512 554190 592521
rect 554134 592447 554190 592456
rect 553216 531276 553268 531282
rect 553216 531218 553268 531224
rect 554044 531276 554096 531282
rect 554044 531218 554096 531224
rect 552492 528958 552704 528986
rect 552492 528850 552520 528958
rect 553228 528850 553256 531218
rect 551080 528822 551416 528850
rect 552092 528822 552520 528850
rect 553196 528822 553256 528850
rect 554148 528850 554176 592447
rect 554240 571826 554268 625223
rect 554778 617944 554834 617953
rect 554778 617879 554834 617888
rect 554410 605840 554466 605849
rect 554410 605775 554466 605784
rect 554318 588840 554374 588849
rect 554318 588775 554374 588784
rect 554332 587926 554360 588775
rect 554320 587920 554372 587926
rect 554320 587862 554372 587868
rect 554318 587616 554374 587625
rect 554318 587551 554374 587560
rect 554332 587042 554360 587551
rect 554320 587036 554372 587042
rect 554320 586978 554372 586984
rect 554320 585200 554372 585206
rect 554318 585168 554320 585177
rect 554372 585168 554374 585177
rect 554318 585103 554374 585112
rect 554318 583944 554374 583953
rect 554318 583879 554374 583888
rect 554332 583778 554360 583879
rect 554320 583772 554372 583778
rect 554320 583714 554372 583720
rect 554318 581496 554374 581505
rect 554318 581431 554374 581440
rect 554332 581058 554360 581431
rect 554320 581052 554372 581058
rect 554320 580994 554372 581000
rect 554318 580272 554374 580281
rect 554318 580207 554374 580216
rect 554332 579698 554360 580207
rect 554320 579692 554372 579698
rect 554320 579634 554372 579640
rect 554318 579048 554374 579057
rect 554318 578983 554374 578992
rect 554332 578270 554360 578983
rect 554320 578264 554372 578270
rect 554320 578206 554372 578212
rect 554318 577824 554374 577833
rect 554318 577759 554374 577768
rect 554332 576910 554360 577759
rect 554320 576904 554372 576910
rect 554320 576846 554372 576852
rect 554424 576722 554452 605775
rect 554594 596048 554650 596057
rect 554594 595983 554650 595992
rect 554502 591288 554558 591297
rect 554502 591223 554558 591232
rect 554516 590714 554544 591223
rect 554504 590708 554556 590714
rect 554504 590650 554556 590656
rect 554502 590064 554558 590073
rect 554502 589999 554558 590008
rect 554516 589354 554544 589999
rect 554504 589348 554556 589354
rect 554504 589290 554556 589296
rect 554502 586392 554558 586401
rect 554502 586327 554558 586336
rect 554516 585274 554544 586327
rect 554504 585268 554556 585274
rect 554504 585210 554556 585216
rect 554424 576694 554544 576722
rect 554410 576600 554466 576609
rect 554410 576535 554466 576544
rect 554424 575550 554452 576535
rect 554412 575544 554464 575550
rect 554412 575486 554464 575492
rect 554318 575376 554374 575385
rect 554318 575311 554374 575320
rect 554332 574190 554360 575311
rect 554320 574184 554372 574190
rect 554320 574126 554372 574132
rect 554410 574152 554466 574161
rect 554410 574087 554412 574096
rect 554464 574087 554466 574096
rect 554412 574058 554464 574064
rect 554410 572928 554466 572937
rect 554410 572863 554466 572872
rect 554424 572762 554452 572863
rect 554412 572756 554464 572762
rect 554412 572698 554464 572704
rect 554240 571798 554360 571826
rect 554226 571704 554282 571713
rect 554226 571639 554282 571648
rect 554240 571402 554268 571639
rect 554228 571396 554280 571402
rect 554228 571338 554280 571344
rect 554332 570722 554360 571798
rect 554320 570716 554372 570722
rect 554320 570658 554372 570664
rect 554410 570616 554466 570625
rect 554410 570551 554466 570560
rect 554424 569974 554452 570551
rect 554516 570450 554544 576694
rect 554608 571266 554636 595983
rect 554596 571260 554648 571266
rect 554596 571202 554648 571208
rect 554504 570444 554556 570450
rect 554504 570386 554556 570392
rect 554412 569968 554464 569974
rect 554412 569910 554464 569916
rect 554792 565146 554820 617879
rect 554780 565140 554832 565146
rect 554780 565082 554832 565088
rect 554884 538898 554912 627671
rect 555146 622840 555202 622849
rect 555146 622775 555202 622784
rect 555054 620392 555110 620401
rect 555054 620327 555110 620336
rect 554962 613184 555018 613193
rect 554962 613119 555018 613128
rect 554976 551342 555004 613119
rect 555068 559570 555096 620327
rect 555160 563718 555188 622775
rect 555330 615632 555386 615641
rect 555330 615567 555386 615576
rect 555238 608288 555294 608297
rect 555238 608223 555294 608232
rect 555148 563712 555200 563718
rect 555148 563654 555200 563660
rect 555056 559564 555108 559570
rect 555056 559506 555108 559512
rect 555252 552702 555280 608223
rect 555344 560998 555372 615567
rect 555516 610020 555568 610026
rect 555516 609962 555568 609968
rect 555422 582720 555478 582729
rect 555422 582655 555478 582664
rect 555332 560992 555384 560998
rect 555332 560934 555384 560940
rect 555240 552696 555292 552702
rect 555240 552638 555292 552644
rect 554964 551336 555016 551342
rect 554964 551278 555016 551284
rect 554872 538892 554924 538898
rect 554872 538834 554924 538840
rect 555436 530738 555464 582655
rect 555528 562358 555556 609962
rect 555608 590708 555660 590714
rect 555608 590650 555660 590656
rect 555516 562352 555568 562358
rect 555516 562294 555568 562300
rect 555424 530732 555476 530738
rect 555424 530674 555476 530680
rect 555620 528850 555648 590650
rect 556160 589348 556212 589354
rect 556160 589290 556212 589296
rect 554148 528822 554300 528850
rect 555404 528822 555648 528850
rect 556172 528850 556200 589290
rect 556264 530602 556292 647226
rect 557632 587920 557684 587926
rect 557632 587862 557684 587868
rect 556804 587036 556856 587042
rect 556804 586978 556856 586984
rect 556252 530596 556304 530602
rect 556252 530538 556304 530544
rect 556816 529990 556844 586978
rect 556804 529984 556856 529990
rect 556804 529926 556856 529932
rect 557644 528850 557672 587862
rect 558920 585268 558972 585274
rect 558920 585210 558972 585216
rect 558184 571396 558236 571402
rect 558184 571338 558236 571344
rect 558196 530602 558224 571338
rect 558184 530596 558236 530602
rect 558184 530538 558236 530544
rect 558276 529984 558328 529990
rect 558276 529926 558328 529932
rect 556172 528822 556416 528850
rect 557520 528822 557672 528850
rect 558288 528850 558316 529926
rect 558932 528986 558960 585210
rect 560300 585200 560352 585206
rect 560300 585142 560352 585148
rect 558932 528958 559328 528986
rect 559300 528850 559328 528958
rect 560312 528850 560340 585142
rect 561772 583772 561824 583778
rect 561772 583714 561824 583720
rect 560944 575544 560996 575550
rect 560944 575486 560996 575492
rect 560956 529990 560984 575486
rect 560944 529984 560996 529990
rect 560944 529926 560996 529932
rect 561784 529122 561812 583714
rect 563060 581052 563112 581058
rect 563060 580994 563112 581000
rect 562600 530732 562652 530738
rect 562600 530674 562652 530680
rect 561784 529094 561858 529122
rect 558288 528822 558624 528850
rect 559300 528822 559636 528850
rect 560312 528822 560740 528850
rect 561830 528836 561858 529094
rect 562612 528850 562640 530674
rect 563072 529666 563100 580994
rect 564440 579692 564492 579698
rect 564440 579634 564492 579640
rect 563072 529638 563652 529666
rect 563624 528850 563652 529638
rect 564452 528986 564480 579634
rect 565820 578264 565872 578270
rect 565820 578206 565872 578212
rect 564452 528958 564756 528986
rect 564728 528850 564756 528958
rect 565832 528850 565860 578206
rect 567292 576904 567344 576910
rect 567292 576846 567344 576852
rect 567304 528850 567332 576846
rect 568580 574184 568632 574190
rect 568580 574126 568632 574132
rect 567936 529984 567988 529990
rect 567936 529926 567988 529932
rect 562612 528822 562948 528850
rect 563624 528822 563960 528850
rect 564728 528822 565064 528850
rect 565832 528822 566168 528850
rect 567180 528822 567332 528850
rect 567948 528850 567976 529926
rect 567948 528822 568284 528850
rect 549976 528686 550588 528714
rect 568592 528714 568620 574126
rect 569960 574116 570012 574122
rect 569960 574058 570012 574064
rect 569972 528714 570000 574058
rect 571432 572756 571484 572762
rect 571432 572698 571484 572704
rect 571444 529122 571472 572698
rect 572720 569968 572772 569974
rect 572720 569910 572772 569916
rect 572260 530596 572312 530602
rect 572260 530538 572312 530544
rect 571444 529094 571518 529122
rect 571490 528836 571518 529094
rect 572272 528850 572300 530538
rect 572732 528986 572760 569910
rect 574376 533520 574428 533526
rect 574376 533462 574428 533468
rect 572732 528958 573220 528986
rect 572272 528822 572608 528850
rect 573192 528714 573220 528958
rect 574388 528850 574416 533462
rect 574388 528822 574724 528850
rect 568592 528686 569388 528714
rect 569972 528686 570492 528714
rect 573192 528686 573712 528714
rect 508502 528320 508558 528329
rect 508502 528255 508558 528264
rect 324136 528216 324188 528222
rect 323964 528164 324136 528170
rect 323964 528158 324188 528164
rect 385408 528216 385460 528222
rect 385408 528158 385460 528164
rect 385868 528216 385920 528222
rect 385868 528158 385920 528164
rect 386420 528216 386472 528222
rect 386420 528158 386472 528164
rect 387340 528216 387392 528222
rect 387340 528158 387392 528164
rect 436468 528216 436520 528222
rect 442816 528216 442868 528222
rect 436520 528164 436816 528170
rect 436468 528158 436816 528164
rect 443368 528216 443420 528222
rect 442868 528164 443256 528170
rect 442816 528158 443256 528164
rect 443368 528158 443420 528164
rect 444932 528216 444984 528222
rect 452752 528216 452804 528222
rect 444984 528164 445464 528170
rect 444932 528158 445464 528164
rect 452804 528164 453008 528170
rect 452752 528158 453008 528164
rect 318064 528148 318116 528154
rect 323964 528142 324176 528158
rect 436480 528142 436816 528158
rect 442828 528142 443256 528158
rect 444944 528142 445464 528158
rect 452764 528142 453008 528158
rect 318064 528090 318116 528096
rect 315304 527876 315356 527882
rect 315304 527818 315356 527824
rect 315946 515808 316002 515817
rect 315946 515743 316002 515752
rect 315960 473414 315988 515743
rect 416596 503056 416648 503062
rect 324332 502982 324760 503010
rect 416148 503004 416596 503010
rect 416148 502998 416648 503004
rect 418160 503056 418212 503062
rect 418804 503056 418856 503062
rect 418212 503004 418804 503010
rect 418160 502998 418856 503004
rect 420276 503056 420328 503062
rect 574008 503056 574060 503062
rect 420328 503004 420868 503010
rect 420276 502998 420868 503004
rect 412088 502988 412140 502994
rect 317892 502846 318228 502874
rect 318904 502846 319332 502874
rect 320284 502846 320436 502874
rect 321112 502846 321448 502874
rect 321572 502846 322552 502874
rect 323320 502846 323656 502874
rect 317892 500954 317920 502846
rect 317328 500948 317380 500954
rect 317328 500890 317380 500896
rect 317880 500948 317932 500954
rect 317880 500890 317932 500896
rect 317340 476882 317368 500890
rect 318904 499746 318932 502846
rect 320284 500834 320312 502846
rect 318720 499718 318932 499746
rect 320100 500806 320312 500834
rect 318720 476882 318748 499718
rect 320100 476882 320128 500806
rect 321112 500750 321140 502846
rect 320272 500744 320324 500750
rect 320272 500686 320324 500692
rect 321100 500744 321152 500750
rect 321100 500686 321152 500692
rect 316684 476876 316736 476882
rect 316684 476818 316736 476824
rect 317328 476876 317380 476882
rect 317328 476818 317380 476824
rect 317880 476876 317932 476882
rect 317880 476818 317932 476824
rect 318708 476876 318760 476882
rect 318708 476818 318760 476824
rect 319076 476876 319128 476882
rect 319076 476818 319128 476824
rect 320088 476876 320140 476882
rect 320088 476818 320140 476824
rect 316696 474164 316724 476818
rect 317892 474164 317920 476818
rect 319088 474164 319116 476818
rect 320284 474178 320312 500686
rect 320284 474150 320390 474178
rect 321572 474164 321600 502846
rect 323320 500410 323348 502846
rect 324332 500834 324360 502982
rect 412088 502930 412140 502936
rect 416148 502982 416636 502998
rect 418172 502982 418844 502998
rect 420288 502982 420868 502998
rect 325758 502602 325786 502860
rect 324240 500806 324360 500834
rect 325712 502574 325786 502602
rect 325896 502846 326876 502874
rect 327092 502846 327980 502874
rect 328472 502846 328992 502874
rect 329852 502846 330096 502874
rect 331200 502846 331352 502874
rect 322848 500404 322900 500410
rect 322848 500346 322900 500352
rect 323308 500404 323360 500410
rect 323308 500346 323360 500352
rect 322860 474178 322888 500346
rect 324240 474178 324268 500806
rect 325712 499610 325740 502574
rect 325620 499582 325740 499610
rect 325620 474178 325648 499582
rect 325896 476490 325924 502846
rect 327092 476626 327120 502846
rect 327092 476598 327396 476626
rect 325896 476462 326108 476490
rect 322782 474150 322888 474178
rect 323978 474150 324268 474178
rect 325266 474150 325648 474178
rect 326080 474178 326108 476462
rect 327368 474178 327396 476598
rect 328472 476490 328500 502846
rect 328472 476462 328684 476490
rect 328656 474178 328684 476462
rect 329852 474178 329880 502846
rect 326080 474150 326462 474178
rect 327368 474150 327658 474178
rect 328656 474150 328946 474178
rect 329852 474150 330142 474178
rect 331324 474164 331352 502846
rect 331416 502846 332304 502874
rect 332612 502846 333316 502874
rect 333992 502846 334420 502874
rect 335372 502846 335524 502874
rect 336536 502846 336688 502874
rect 337640 502846 338068 502874
rect 338744 502846 339448 502874
rect 339848 502846 340184 502874
rect 340860 502846 341196 502874
rect 341964 502846 342208 502874
rect 343068 502846 343220 502874
rect 344080 502846 344416 502874
rect 345184 502846 345520 502874
rect 346288 502846 346348 502874
rect 347392 502846 347728 502874
rect 348404 502846 349108 502874
rect 349508 502846 349844 502874
rect 350612 502846 350948 502874
rect 351624 502846 351776 502874
rect 352728 502846 353248 502874
rect 353832 502846 354168 502874
rect 354936 502846 355272 502874
rect 331416 476474 331444 502846
rect 332612 476882 332640 502846
rect 332600 476876 332652 476882
rect 332600 476818 332652 476824
rect 333796 476876 333848 476882
rect 333796 476818 333848 476824
rect 331404 476468 331456 476474
rect 331404 476410 331456 476416
rect 332508 476468 332560 476474
rect 332508 476410 332560 476416
rect 332520 474164 332548 476410
rect 333808 474164 333836 476818
rect 333992 476610 334020 502846
rect 335372 476882 335400 502846
rect 336660 476882 336688 502846
rect 335360 476876 335412 476882
rect 335360 476818 335412 476824
rect 336188 476876 336240 476882
rect 336188 476818 336240 476824
rect 336648 476876 336700 476882
rect 336648 476818 336700 476824
rect 337476 476876 337528 476882
rect 337476 476818 337528 476824
rect 333980 476604 334032 476610
rect 333980 476546 334032 476552
rect 334992 476604 335044 476610
rect 334992 476546 335044 476552
rect 335004 474164 335032 476546
rect 336200 474164 336228 476818
rect 337488 474164 337516 476818
rect 338040 476218 338068 502846
rect 339420 476218 339448 502846
rect 340156 500954 340184 502846
rect 341168 500954 341196 502846
rect 340144 500948 340196 500954
rect 340144 500890 340196 500896
rect 340788 500948 340840 500954
rect 340788 500890 340840 500896
rect 341156 500948 341208 500954
rect 341156 500890 341208 500896
rect 342076 500948 342128 500954
rect 342076 500890 342128 500896
rect 340800 476218 340828 500890
rect 342088 476218 342116 500890
rect 342180 476882 342208 502846
rect 343192 500954 343220 502846
rect 343180 500948 343232 500954
rect 343180 500890 343232 500896
rect 343732 500948 343784 500954
rect 343732 500890 343784 500896
rect 343744 476898 343772 500890
rect 344388 499866 344416 502846
rect 345492 500954 345520 502846
rect 345480 500948 345532 500954
rect 345480 500890 345532 500896
rect 346216 500948 346268 500954
rect 346216 500890 346268 500896
rect 344376 499860 344428 499866
rect 344376 499802 344428 499808
rect 344928 499860 344980 499866
rect 344928 499802 344980 499808
rect 344940 477494 344968 499802
rect 344928 477488 344980 477494
rect 344928 477430 344980 477436
rect 346032 477488 346084 477494
rect 346032 477430 346084 477436
rect 342168 476876 342220 476882
rect 342168 476818 342220 476824
rect 343548 476876 343600 476882
rect 343744 476870 344324 476898
rect 343548 476818 343600 476824
rect 338040 476190 338344 476218
rect 339420 476190 339540 476218
rect 340800 476190 340920 476218
rect 342088 476190 342300 476218
rect 338316 474178 338344 476190
rect 339512 474178 339540 476190
rect 340892 474178 340920 476190
rect 342272 474178 342300 476190
rect 338316 474150 338698 474178
rect 339512 474150 339894 474178
rect 340892 474150 341090 474178
rect 342272 474150 342378 474178
rect 343560 474164 343588 476818
rect 344296 474042 344324 476870
rect 346044 474164 346072 477430
rect 346228 476882 346256 500890
rect 346216 476876 346268 476882
rect 346216 476818 346268 476824
rect 346320 476338 346348 502846
rect 347228 476876 347280 476882
rect 347228 476818 347280 476824
rect 346308 476332 346360 476338
rect 346308 476274 346360 476280
rect 347240 474164 347268 476818
rect 347700 476406 347728 502846
rect 349080 476610 349108 502846
rect 349816 500954 349844 502846
rect 350920 500954 350948 502846
rect 349804 500948 349856 500954
rect 349804 500890 349856 500896
rect 350448 500948 350500 500954
rect 350448 500890 350500 500896
rect 350908 500948 350960 500954
rect 350908 500890 350960 500896
rect 350460 476882 350488 500890
rect 350448 476876 350500 476882
rect 350448 476818 350500 476824
rect 351748 476814 351776 502846
rect 351828 500948 351880 500954
rect 351828 500890 351880 500896
rect 351840 476950 351868 500890
rect 353220 477494 353248 502846
rect 354140 500954 354168 502846
rect 354128 500948 354180 500954
rect 354128 500890 354180 500896
rect 354588 500948 354640 500954
rect 354588 500890 354640 500896
rect 353208 477488 353260 477494
rect 353208 477430 353260 477436
rect 354600 477426 354628 500890
rect 355244 500818 355272 502846
rect 355934 502602 355962 502860
rect 357052 502846 357388 502874
rect 358156 502846 358768 502874
rect 359168 502846 359504 502874
rect 360272 502846 360608 502874
rect 361376 502846 361528 502874
rect 362480 502846 362908 502874
rect 363492 502846 363828 502874
rect 364596 502846 364932 502874
rect 365700 502846 366036 502874
rect 366712 502846 366956 502874
rect 367816 502846 368428 502874
rect 368920 502846 369256 502874
rect 370024 502846 370360 502874
rect 371036 502846 371188 502874
rect 372140 502846 372568 502874
rect 373244 502846 373948 502874
rect 374256 502846 374592 502874
rect 375360 502846 375696 502874
rect 376464 502846 376708 502874
rect 377568 502846 378088 502874
rect 378580 502846 378916 502874
rect 379684 502846 380020 502874
rect 380788 502846 380848 502874
rect 381800 502846 382228 502874
rect 382904 502846 383608 502874
rect 384008 502846 384344 502874
rect 385112 502846 385448 502874
rect 386124 502846 386276 502874
rect 387228 502846 387748 502874
rect 388332 502846 388668 502874
rect 389344 502846 389680 502874
rect 355888 502574 355962 502602
rect 355232 500812 355284 500818
rect 355232 500754 355284 500760
rect 355784 477488 355836 477494
rect 355784 477430 355836 477436
rect 354588 477420 354640 477426
rect 354588 477362 354640 477368
rect 351828 476944 351880 476950
rect 351828 476886 351880 476892
rect 353300 476944 353352 476950
rect 353300 476886 353352 476892
rect 352104 476876 352156 476882
rect 352104 476818 352156 476824
rect 351736 476808 351788 476814
rect 351736 476750 351788 476756
rect 349068 476604 349120 476610
rect 349068 476546 349120 476552
rect 350908 476604 350960 476610
rect 350908 476546 350960 476552
rect 347688 476400 347740 476406
rect 347688 476342 347740 476348
rect 349620 476400 349672 476406
rect 349620 476342 349672 476348
rect 348424 476332 348476 476338
rect 348424 476274 348476 476280
rect 348436 474164 348464 476274
rect 349632 474164 349660 476342
rect 350920 474164 350948 476546
rect 352116 474164 352144 476818
rect 353312 474164 353340 476886
rect 354588 476808 354640 476814
rect 354588 476750 354640 476756
rect 354600 474164 354628 476750
rect 355796 474164 355824 477430
rect 355888 476950 355916 502574
rect 355968 500812 356020 500818
rect 355968 500754 356020 500760
rect 355876 476944 355928 476950
rect 355876 476886 355928 476892
rect 355980 476882 356008 500754
rect 356980 477420 357032 477426
rect 356980 477362 357032 477368
rect 355968 476876 356020 476882
rect 355968 476818 356020 476824
rect 356992 474164 357020 477362
rect 357360 476610 357388 502846
rect 358740 476882 358768 502846
rect 359476 500954 359504 502846
rect 359464 500948 359516 500954
rect 359464 500890 359516 500896
rect 360108 500948 360160 500954
rect 360108 500890 360160 500896
rect 359464 476944 359516 476950
rect 359464 476886 359516 476892
rect 358176 476876 358228 476882
rect 358176 476818 358228 476824
rect 358728 476876 358780 476882
rect 358728 476818 358780 476824
rect 357348 476604 357400 476610
rect 357348 476546 357400 476552
rect 358188 474164 358216 476818
rect 359476 474164 359504 476886
rect 360120 476542 360148 500890
rect 360580 500682 360608 502846
rect 360568 500676 360620 500682
rect 360568 500618 360620 500624
rect 361396 500676 361448 500682
rect 361396 500618 361448 500624
rect 361408 476746 361436 500618
rect 361500 477018 361528 502846
rect 362880 477494 362908 502846
rect 363800 500546 363828 502846
rect 364904 500954 364932 502846
rect 366008 500954 366036 502846
rect 364892 500948 364944 500954
rect 364892 500890 364944 500896
rect 365628 500948 365680 500954
rect 365628 500890 365680 500896
rect 365996 500948 366048 500954
rect 365996 500890 366048 500896
rect 363788 500540 363840 500546
rect 363788 500482 363840 500488
rect 364248 500540 364300 500546
rect 364248 500482 364300 500488
rect 362868 477488 362920 477494
rect 362868 477430 362920 477436
rect 364260 477086 364288 500482
rect 364248 477080 364300 477086
rect 364248 477022 364300 477028
rect 361488 477012 361540 477018
rect 361488 476954 361540 476960
rect 365536 477012 365588 477018
rect 365536 476954 365588 476960
rect 361856 476876 361908 476882
rect 361856 476818 361908 476824
rect 361396 476740 361448 476746
rect 361396 476682 361448 476688
rect 360660 476604 360712 476610
rect 360660 476546 360712 476552
rect 360108 476536 360160 476542
rect 360108 476478 360160 476484
rect 360672 474164 360700 476546
rect 361868 474164 361896 476818
rect 364340 476740 364392 476746
rect 364340 476682 364392 476688
rect 363052 476536 363104 476542
rect 363052 476478 363104 476484
rect 363064 474164 363092 476478
rect 364352 474164 364380 476682
rect 365548 474164 365576 476954
rect 365640 476678 365668 500890
rect 366732 477488 366784 477494
rect 366732 477430 366784 477436
rect 365628 476672 365680 476678
rect 365628 476614 365680 476620
rect 366744 474164 366772 477430
rect 366928 476610 366956 502846
rect 367008 500948 367060 500954
rect 367008 500890 367060 500896
rect 366916 476604 366968 476610
rect 366916 476546 366968 476552
rect 367020 476406 367048 500890
rect 368020 477080 368072 477086
rect 368020 477022 368072 477028
rect 367008 476400 367060 476406
rect 367008 476342 367060 476348
rect 368032 474164 368060 477022
rect 368400 476950 368428 502846
rect 369228 500546 369256 502846
rect 370332 500682 370360 502846
rect 370320 500676 370372 500682
rect 370320 500618 370372 500624
rect 371056 500676 371108 500682
rect 371056 500618 371108 500624
rect 369216 500540 369268 500546
rect 369216 500482 369268 500488
rect 369768 500540 369820 500546
rect 369768 500482 369820 500488
rect 369780 477494 369808 500482
rect 369768 477488 369820 477494
rect 369768 477430 369820 477436
rect 368388 476944 368440 476950
rect 368388 476886 368440 476892
rect 371068 476882 371096 500618
rect 371056 476876 371108 476882
rect 371056 476818 371108 476824
rect 371160 476746 371188 502846
rect 372540 477018 372568 502846
rect 372528 477012 372580 477018
rect 372528 476954 372580 476960
rect 373920 476950 373948 502846
rect 374564 500002 374592 502846
rect 375668 500954 375696 502846
rect 375656 500948 375708 500954
rect 375656 500890 375708 500896
rect 376576 500948 376628 500954
rect 376576 500890 376628 500896
rect 374552 499996 374604 500002
rect 374552 499938 374604 499944
rect 375288 499996 375340 500002
rect 375288 499938 375340 499944
rect 374092 477488 374144 477494
rect 374092 477430 374144 477436
rect 372896 476944 372948 476950
rect 372896 476886 372948 476892
rect 373908 476944 373960 476950
rect 373908 476886 373960 476892
rect 371148 476740 371200 476746
rect 371148 476682 371200 476688
rect 369216 476672 369268 476678
rect 369216 476614 369268 476620
rect 369228 474164 369256 476614
rect 371608 476604 371660 476610
rect 371608 476546 371660 476552
rect 370412 476400 370464 476406
rect 370412 476342 370464 476348
rect 370424 474164 370452 476342
rect 371620 474164 371648 476546
rect 372908 474164 372936 476886
rect 374104 474164 374132 477430
rect 375300 477086 375328 499938
rect 375288 477080 375340 477086
rect 375288 477022 375340 477028
rect 376588 476882 376616 500890
rect 375288 476876 375340 476882
rect 375288 476818 375340 476824
rect 376576 476876 376628 476882
rect 376576 476818 376628 476824
rect 375300 474164 375328 476818
rect 376576 476740 376628 476746
rect 376576 476682 376628 476688
rect 376588 474164 376616 476682
rect 376680 476202 376708 502846
rect 377772 477012 377824 477018
rect 377772 476954 377824 476960
rect 376668 476196 376720 476202
rect 376668 476138 376720 476144
rect 377784 474164 377812 476954
rect 378060 476474 378088 502846
rect 378888 500002 378916 502846
rect 379992 500954 380020 502846
rect 379980 500948 380032 500954
rect 379980 500890 380032 500896
rect 380716 500948 380768 500954
rect 380716 500890 380768 500896
rect 378876 499996 378928 500002
rect 378876 499938 378928 499944
rect 379428 499996 379480 500002
rect 379428 499938 379480 499944
rect 378968 476944 379020 476950
rect 378968 476886 379020 476892
rect 378048 476468 378100 476474
rect 378048 476410 378100 476416
rect 378980 474164 379008 476886
rect 379440 476406 379468 499938
rect 380164 477080 380216 477086
rect 380164 477022 380216 477028
rect 379428 476400 379480 476406
rect 379428 476342 379480 476348
rect 380176 474164 380204 477022
rect 380728 476270 380756 500890
rect 380820 476950 380848 502846
rect 382200 477222 382228 502846
rect 382188 477216 382240 477222
rect 382188 477158 382240 477164
rect 380808 476944 380860 476950
rect 380808 476886 380860 476892
rect 381452 476876 381504 476882
rect 381452 476818 381504 476824
rect 380716 476264 380768 476270
rect 380716 476206 380768 476212
rect 381464 474164 381492 476818
rect 383580 476814 383608 502846
rect 384316 500954 384344 502846
rect 385420 500954 385448 502846
rect 384304 500948 384356 500954
rect 384304 500890 384356 500896
rect 384948 500948 385000 500954
rect 384948 500890 385000 500896
rect 385408 500948 385460 500954
rect 385408 500890 385460 500896
rect 383568 476808 383620 476814
rect 383568 476750 383620 476756
rect 383844 476468 383896 476474
rect 383844 476410 383896 476416
rect 382648 476196 382700 476202
rect 382648 476138 382700 476144
rect 382660 474164 382688 476138
rect 383856 474164 383884 476410
rect 384960 476202 384988 500890
rect 386248 477086 386276 502846
rect 386328 500948 386380 500954
rect 386328 500890 386380 500896
rect 386236 477080 386288 477086
rect 386236 477022 386288 477028
rect 386340 476882 386368 500890
rect 387524 476944 387576 476950
rect 387524 476886 387576 476892
rect 386328 476876 386380 476882
rect 386328 476818 386380 476824
rect 385132 476400 385184 476406
rect 385132 476342 385184 476348
rect 384948 476196 385000 476202
rect 384948 476138 385000 476144
rect 385144 474164 385172 476342
rect 386328 476264 386380 476270
rect 386328 476206 386380 476212
rect 386340 474164 386368 476206
rect 387536 474164 387564 476886
rect 387720 476474 387748 502846
rect 388640 499934 388668 502846
rect 389652 500002 389680 502846
rect 390434 502602 390462 502860
rect 391552 502846 391888 502874
rect 392656 502846 393268 502874
rect 393668 502846 394004 502874
rect 394772 502846 395108 502874
rect 395876 502846 396028 502874
rect 396888 502846 397408 502874
rect 397992 502846 398328 502874
rect 399096 502846 399432 502874
rect 400200 502846 400536 502874
rect 401212 502846 401456 502874
rect 403420 502846 403756 502874
rect 404432 502846 404768 502874
rect 409860 502846 409920 502874
rect 390388 502574 390462 502602
rect 389640 499996 389692 500002
rect 389640 499938 389692 499944
rect 388628 499928 388680 499934
rect 388628 499870 388680 499876
rect 389088 499928 389140 499934
rect 389088 499870 389140 499876
rect 388720 477216 388772 477222
rect 388720 477158 388772 477164
rect 387708 476468 387760 476474
rect 387708 476410 387760 476416
rect 388732 474164 388760 477158
rect 389100 476950 389128 499870
rect 389088 476944 389140 476950
rect 389088 476886 389140 476892
rect 390388 476814 390416 502574
rect 390468 499996 390520 500002
rect 390468 499938 390520 499944
rect 390480 477358 390508 499938
rect 390468 477352 390520 477358
rect 390468 477294 390520 477300
rect 391860 477222 391888 502846
rect 391848 477216 391900 477222
rect 391848 477158 391900 477164
rect 393240 477154 393268 502846
rect 393976 500002 394004 502846
rect 395080 500002 395108 502846
rect 393964 499996 394016 500002
rect 393964 499938 394016 499944
rect 394608 499996 394660 500002
rect 394608 499938 394660 499944
rect 395068 499996 395120 500002
rect 395068 499938 395120 499944
rect 395896 499996 395948 500002
rect 395896 499938 395948 499944
rect 393228 477148 393280 477154
rect 393228 477090 393280 477096
rect 392492 477080 392544 477086
rect 392492 477022 392544 477028
rect 392504 476882 392532 477022
rect 392400 476876 392452 476882
rect 392400 476818 392452 476824
rect 392492 476876 392544 476882
rect 392492 476818 392544 476824
rect 393688 476876 393740 476882
rect 393688 476818 393740 476824
rect 390008 476808 390060 476814
rect 390008 476750 390060 476756
rect 390376 476808 390428 476814
rect 390376 476750 390428 476756
rect 390020 474164 390048 476750
rect 391204 476196 391256 476202
rect 391204 476138 391256 476144
rect 391216 474164 391244 476138
rect 392412 474164 392440 476818
rect 393700 474164 393728 476818
rect 394620 476746 394648 499938
rect 395908 477086 395936 499938
rect 395896 477080 395948 477086
rect 395896 477022 395948 477028
rect 396000 477018 396028 502846
rect 397276 477352 397328 477358
rect 397276 477294 397328 477300
rect 395988 477012 396040 477018
rect 395988 476954 396040 476960
rect 396080 476944 396132 476950
rect 396080 476886 396132 476892
rect 394608 476740 394660 476746
rect 394608 476682 394660 476688
rect 394884 476468 394936 476474
rect 394884 476410 394936 476416
rect 394896 474164 394924 476410
rect 396092 474164 396120 476886
rect 397288 474164 397316 477294
rect 397380 476950 397408 502846
rect 398300 500410 398328 502846
rect 398288 500404 398340 500410
rect 398288 500346 398340 500352
rect 398748 500404 398800 500410
rect 398748 500346 398800 500352
rect 397368 476944 397420 476950
rect 397368 476886 397420 476892
rect 398760 476882 398788 500346
rect 399404 500002 399432 502846
rect 400508 500954 400536 502846
rect 400496 500948 400548 500954
rect 400496 500890 400548 500896
rect 399392 499996 399444 500002
rect 399392 499938 399444 499944
rect 400128 499996 400180 500002
rect 400128 499938 400180 499944
rect 400140 477222 400168 499938
rect 399760 477216 399812 477222
rect 399760 477158 399812 477164
rect 400128 477216 400180 477222
rect 400128 477158 400180 477164
rect 398748 476876 398800 476882
rect 398748 476818 398800 476824
rect 398564 476808 398616 476814
rect 398564 476750 398616 476756
rect 398576 474164 398604 476750
rect 399772 474164 399800 477158
rect 400956 477148 401008 477154
rect 400956 477090 401008 477096
rect 400968 474164 400996 477090
rect 401428 476814 401456 502846
rect 401508 500948 401560 500954
rect 401508 500890 401560 500896
rect 401520 477154 401548 500890
rect 403728 500886 403756 502846
rect 404740 500954 404768 502846
rect 404728 500948 404780 500954
rect 404728 500890 404780 500896
rect 409892 500886 409920 502846
rect 411640 502846 411976 502874
rect 411640 500954 411668 502846
rect 411628 500948 411680 500954
rect 411628 500890 411680 500896
rect 403716 500880 403768 500886
rect 403716 500822 403768 500828
rect 409880 500880 409932 500886
rect 409880 500822 409932 500828
rect 408316 477216 408368 477222
rect 408316 477158 408368 477164
rect 401508 477148 401560 477154
rect 401508 477090 401560 477096
rect 403440 477080 403492 477086
rect 403440 477022 403492 477028
rect 401416 476808 401468 476814
rect 401416 476750 401468 476756
rect 402244 476740 402296 476746
rect 402244 476682 402296 476688
rect 402256 474164 402284 476682
rect 403452 474164 403480 477022
rect 404636 477012 404688 477018
rect 404636 476954 404688 476960
rect 404648 474164 404676 476954
rect 405832 476944 405884 476950
rect 405832 476886 405884 476892
rect 405844 474164 405872 476886
rect 407120 476876 407172 476882
rect 407120 476818 407172 476824
rect 407132 474164 407160 476818
rect 408328 474164 408356 477158
rect 409512 477148 409564 477154
rect 409512 477090 409564 477096
rect 409524 474164 409552 477090
rect 410708 476808 410760 476814
rect 410708 476750 410760 476756
rect 410720 474164 410748 476750
rect 344296 474014 344770 474042
rect 389822 473920 389878 473929
rect 389822 473855 389878 473864
rect 389836 473657 389864 473855
rect 408590 473784 408646 473793
rect 408420 473742 408590 473770
rect 408420 473657 408448 473742
rect 408590 473719 408646 473728
rect 389822 473648 389878 473657
rect 389822 473583 389878 473592
rect 408406 473648 408462 473657
rect 408406 473583 408462 473592
rect 314660 473408 314712 473414
rect 314660 473350 314712 473356
rect 315948 473408 316000 473414
rect 315948 473350 316000 473356
rect 314672 439657 314700 473350
rect 314658 439648 314714 439657
rect 314658 439583 314714 439592
rect 338118 428768 338174 428777
rect 338118 428703 338174 428712
rect 336004 311908 336056 311914
rect 336004 311850 336056 311856
rect 313924 232552 313976 232558
rect 313924 232494 313976 232500
rect 309784 227044 309836 227050
rect 309784 226986 309836 226992
rect 286324 224256 286376 224262
rect 286324 224198 286376 224204
rect 283380 223644 283432 223650
rect 283380 223586 283432 223592
rect 231124 222488 231176 222494
rect 231124 222430 231176 222436
rect 235264 222488 235316 222494
rect 235264 222430 235316 222436
rect 230848 184884 230900 184890
rect 230848 184826 230900 184832
rect 230860 184770 230888 184826
rect 231136 184770 231164 222430
rect 283392 221612 283420 223586
rect 230860 184742 231164 184770
rect 336016 182170 336044 311850
rect 338132 198665 338160 428703
rect 338394 428632 338450 428641
rect 338394 428567 338450 428576
rect 338118 198656 338174 198665
rect 338118 198591 338174 198600
rect 336004 182164 336056 182170
rect 336004 182106 336056 182112
rect 283392 173913 283420 175508
rect 283378 173904 283434 173913
rect 283378 173839 283434 173848
rect 283392 173233 283420 173839
rect 232226 173224 232282 173233
rect 232226 173159 232282 173168
rect 283378 173224 283434 173233
rect 283378 173159 283434 173168
rect 232240 167006 232268 173159
rect 232228 167000 232280 167006
rect 232228 166942 232280 166948
rect 232596 167000 232648 167006
rect 232596 166942 232648 166948
rect 232608 164218 232636 166942
rect 232320 164212 232372 164218
rect 232320 164154 232372 164160
rect 232596 164212 232648 164218
rect 232596 164154 232648 164160
rect 215116 161424 215168 161430
rect 215116 161366 215168 161372
rect 229744 161424 229796 161430
rect 229744 161366 229796 161372
rect 215128 160993 215156 161366
rect 215114 160984 215170 160993
rect 215114 160919 215170 160928
rect 214930 160168 214986 160177
rect 214930 160103 214986 160112
rect 214838 158672 214894 158681
rect 214838 158607 214894 158616
rect 214746 157856 214802 157865
rect 214746 157791 214802 157800
rect 215114 157040 215170 157049
rect 215114 156975 215170 156984
rect 214746 156360 214802 156369
rect 214746 156295 214802 156304
rect 214760 149054 214788 156295
rect 215128 155990 215156 156975
rect 215116 155984 215168 155990
rect 215116 155926 215168 155932
rect 224684 155984 224736 155990
rect 224684 155926 224736 155932
rect 215114 154728 215170 154737
rect 215114 154663 215170 154672
rect 224592 154692 224644 154698
rect 215128 154630 215156 154663
rect 224592 154634 224644 154640
rect 215116 154624 215168 154630
rect 215116 154566 215168 154572
rect 215206 153912 215262 153921
rect 215206 153847 215262 153856
rect 215220 153338 215248 153847
rect 215208 153332 215260 153338
rect 215208 153274 215260 153280
rect 215116 153264 215168 153270
rect 215114 153232 215116 153241
rect 215168 153232 215170 153241
rect 215114 153167 215170 153176
rect 224500 151904 224552 151910
rect 224500 151846 224552 151852
rect 218704 151836 218756 151842
rect 218704 151778 218756 151784
rect 215114 150784 215170 150793
rect 215114 150719 215170 150728
rect 215128 150482 215156 150719
rect 216680 150544 216732 150550
rect 216680 150486 216732 150492
rect 215116 150476 215168 150482
rect 215116 150418 215168 150424
rect 215114 149288 215170 149297
rect 215114 149223 215170 149232
rect 215128 149122 215156 149223
rect 215116 149116 215168 149122
rect 215116 149058 215168 149064
rect 214748 149048 214800 149054
rect 214748 148990 214800 148996
rect 215114 148472 215170 148481
rect 215114 148407 215170 148416
rect 215128 147694 215156 148407
rect 215116 147688 215168 147694
rect 214838 147656 214894 147665
rect 215116 147630 215168 147636
rect 214838 147591 214894 147600
rect 214852 146334 214880 147591
rect 215206 146840 215262 146849
rect 215206 146775 215262 146784
rect 215220 146402 215248 146775
rect 215208 146396 215260 146402
rect 215208 146338 215260 146344
rect 214840 146328 214892 146334
rect 214840 146270 214892 146276
rect 216692 146266 216720 150486
rect 216864 149252 216916 149258
rect 216864 149194 216916 149200
rect 216772 147688 216824 147694
rect 216772 147630 216824 147636
rect 216680 146260 216732 146266
rect 216680 146202 216732 146208
rect 215022 146160 215078 146169
rect 215022 146095 215078 146104
rect 215036 144974 215064 146095
rect 215206 145344 215262 145353
rect 215206 145279 215262 145288
rect 215220 145042 215248 145279
rect 215208 145036 215260 145042
rect 215208 144978 215260 144984
rect 215024 144968 215076 144974
rect 215024 144910 215076 144916
rect 215206 143712 215262 143721
rect 215206 143647 215208 143656
rect 215260 143647 215262 143656
rect 216680 143676 216732 143682
rect 215208 143618 215260 143624
rect 216680 143618 216732 143624
rect 215114 143032 215170 143041
rect 215114 142967 215170 142976
rect 215128 142186 215156 142967
rect 215208 142248 215260 142254
rect 215206 142216 215208 142225
rect 215260 142216 215262 142225
rect 215116 142180 215168 142186
rect 215206 142151 215262 142160
rect 215116 142122 215168 142128
rect 215114 141400 215170 141409
rect 215114 141335 215170 141344
rect 215128 140826 215156 141335
rect 215116 140820 215168 140826
rect 215116 140762 215168 140768
rect 215114 140584 215170 140593
rect 215114 140519 215170 140528
rect 215128 139466 215156 140519
rect 215116 139460 215168 139466
rect 215116 139402 215168 139408
rect 216692 139398 216720 143618
rect 216784 143546 216812 147630
rect 216876 144906 216904 149194
rect 217692 146396 217744 146402
rect 217692 146338 217744 146344
rect 217416 145036 217468 145042
rect 217416 144978 217468 144984
rect 216864 144900 216916 144906
rect 216864 144842 216916 144848
rect 216772 143540 216824 143546
rect 216772 143482 216824 143488
rect 216772 142248 216824 142254
rect 216772 142190 216824 142196
rect 216680 139392 216732 139398
rect 216680 139334 216732 139340
rect 215114 138272 215170 138281
rect 215114 138207 215170 138216
rect 215128 138106 215156 138207
rect 215116 138100 215168 138106
rect 215116 138042 215168 138048
rect 216784 137970 216812 142190
rect 217428 140758 217456 144978
rect 217704 142118 217732 146338
rect 217692 142112 217744 142118
rect 217692 142054 217744 142060
rect 217416 140752 217468 140758
rect 217416 140694 217468 140700
rect 216772 137964 216824 137970
rect 216772 137906 216824 137912
rect 215114 136776 215170 136785
rect 215114 136711 215116 136720
rect 215168 136711 215170 136720
rect 215116 136682 215168 136688
rect 215206 135144 215262 135153
rect 215206 135079 215262 135088
rect 215114 134328 215170 134337
rect 215114 134263 215170 134272
rect 215128 134026 215156 134263
rect 215116 134020 215168 134026
rect 215116 133962 215168 133968
rect 215220 133958 215248 135079
rect 215208 133952 215260 133958
rect 215208 133894 215260 133900
rect 215114 133512 215170 133521
rect 215114 133447 215170 133456
rect 215128 132530 215156 133447
rect 215116 132524 215168 132530
rect 215116 132466 215168 132472
rect 215116 131232 215168 131238
rect 215114 131200 215116 131209
rect 215168 131200 215170 131209
rect 215114 131135 215170 131144
rect 215114 128072 215170 128081
rect 215114 128007 215170 128016
rect 215128 127634 215156 128007
rect 215116 127628 215168 127634
rect 215116 127570 215168 127576
rect 215114 127256 215170 127265
rect 215114 127191 215170 127200
rect 215128 127022 215156 127191
rect 215116 127016 215168 127022
rect 215116 126958 215168 126964
rect 215114 126576 215170 126585
rect 215114 126511 215170 126520
rect 215128 126274 215156 126511
rect 215116 126268 215168 126274
rect 215116 126210 215168 126216
rect 215114 125760 215170 125769
rect 215114 125695 215170 125704
rect 215128 125662 215156 125695
rect 215116 125656 215168 125662
rect 215116 125598 215168 125604
rect 215114 124944 215170 124953
rect 215114 124879 215116 124888
rect 215168 124879 215170 124888
rect 215116 124850 215168 124856
rect 215116 124160 215168 124166
rect 215114 124128 215116 124137
rect 215168 124128 215170 124137
rect 215114 124063 215170 124072
rect 215116 123480 215168 123486
rect 215114 123448 215116 123457
rect 215168 123448 215170 123457
rect 215114 123383 215170 123392
rect 215116 122800 215168 122806
rect 215116 122742 215168 122748
rect 215128 122641 215156 122742
rect 215114 122632 215170 122641
rect 215114 122567 215170 122576
rect 215116 122120 215168 122126
rect 215116 122062 215168 122068
rect 215128 121825 215156 122062
rect 215114 121816 215170 121825
rect 215114 121751 215170 121760
rect 215116 121440 215168 121446
rect 215116 121382 215168 121388
rect 215128 121009 215156 121382
rect 215114 121000 215170 121009
rect 215114 120935 215170 120944
rect 215116 120760 215168 120766
rect 215116 120702 215168 120708
rect 215128 120329 215156 120702
rect 215114 120320 215170 120329
rect 215114 120255 215170 120264
rect 215114 118688 215170 118697
rect 215114 118623 215170 118632
rect 215128 118590 215156 118623
rect 215116 118584 215168 118590
rect 215116 118526 215168 118532
rect 215208 117292 215260 117298
rect 215208 117234 215260 117240
rect 215116 117224 215168 117230
rect 215116 117166 215168 117172
rect 215128 117065 215156 117166
rect 215114 117056 215170 117065
rect 215114 116991 215170 117000
rect 215220 116385 215248 117234
rect 215206 116376 215262 116385
rect 215206 116311 215262 116320
rect 215208 115932 215260 115938
rect 215208 115874 215260 115880
rect 215116 115864 215168 115870
rect 215116 115806 215168 115812
rect 215128 115569 215156 115806
rect 215114 115560 215170 115569
rect 215114 115495 215170 115504
rect 215220 114753 215248 115874
rect 215206 114744 215262 114753
rect 215206 114679 215262 114688
rect 215116 114504 215168 114510
rect 215116 114446 215168 114452
rect 215128 113257 215156 114446
rect 215114 113248 215170 113257
rect 215114 113183 215170 113192
rect 215208 111784 215260 111790
rect 215208 111726 215260 111732
rect 215116 111716 215168 111722
rect 215116 111658 215168 111664
rect 215128 111625 215156 111658
rect 215114 111616 215170 111625
rect 215114 111551 215170 111560
rect 215220 110809 215248 111726
rect 215206 110800 215262 110809
rect 215206 110735 215262 110744
rect 215116 110424 215168 110430
rect 215116 110366 215168 110372
rect 215128 110129 215156 110366
rect 215114 110120 215170 110129
rect 215114 110055 215170 110064
rect 215208 108996 215260 109002
rect 215208 108938 215260 108944
rect 215116 108928 215168 108934
rect 215116 108870 215168 108876
rect 215128 108497 215156 108870
rect 215114 108488 215170 108497
rect 215114 108423 215170 108432
rect 215220 107681 215248 108938
rect 215206 107672 215262 107681
rect 215206 107607 215262 107616
rect 215116 106276 215168 106282
rect 215116 106218 215168 106224
rect 215128 106185 215156 106218
rect 215114 106176 215170 106185
rect 215114 106111 215170 106120
rect 215116 104848 215168 104854
rect 215116 104790 215168 104796
rect 215128 104553 215156 104790
rect 215114 104544 215170 104553
rect 215114 104479 215170 104488
rect 215116 103488 215168 103494
rect 215116 103430 215168 103436
rect 215128 102241 215156 103430
rect 215208 103420 215260 103426
rect 215208 103362 215260 103368
rect 215220 103057 215248 103362
rect 215206 103048 215262 103057
rect 215206 102983 215262 102992
rect 215114 102232 215170 102241
rect 215114 102167 215170 102176
rect 215116 102128 215168 102134
rect 215116 102070 215168 102076
rect 215128 101425 215156 102070
rect 215114 101416 215170 101425
rect 215114 101351 215170 101360
rect 215116 100632 215168 100638
rect 215114 100600 215116 100609
rect 215168 100600 215170 100609
rect 215114 100535 215170 100544
rect 214668 99470 214788 99498
rect 214656 99340 214708 99346
rect 214656 99282 214708 99288
rect 214668 98297 214696 99282
rect 214654 98288 214710 98297
rect 214654 98223 214710 98232
rect 214564 97028 214616 97034
rect 214564 96970 214616 96976
rect 214576 96801 214604 96970
rect 214562 96792 214618 96801
rect 214562 96727 214618 96736
rect 214286 95976 214342 95985
rect 214286 95911 214342 95920
rect 214760 95169 214788 99470
rect 215116 99272 215168 99278
rect 215116 99214 215168 99220
rect 215128 99113 215156 99214
rect 215114 99104 215170 99113
rect 215114 99039 215170 99048
rect 218716 97034 218744 151778
rect 224040 150476 224092 150482
rect 224040 150418 224092 150424
rect 224052 144838 224080 150418
rect 224224 149116 224276 149122
rect 224224 149058 224276 149064
rect 224040 144832 224092 144838
rect 224040 144774 224092 144780
rect 224236 143478 224264 149058
rect 224512 146198 224540 151846
rect 224604 148986 224632 154634
rect 224696 150414 224724 155926
rect 225604 154624 225656 154630
rect 232332 154601 232360 164154
rect 225604 154566 225656 154572
rect 232318 154592 232374 154601
rect 224868 153332 224920 153338
rect 224868 153274 224920 153280
rect 224776 153264 224828 153270
rect 224776 153206 224828 153212
rect 224684 150408 224736 150414
rect 224684 150350 224736 150356
rect 224592 148980 224644 148986
rect 224592 148922 224644 148928
rect 224788 147558 224816 153206
rect 224880 147626 224908 153274
rect 225616 147665 225644 154566
rect 232318 154527 232374 154536
rect 232502 154592 232558 154601
rect 232502 154527 232558 154536
rect 227444 150408 227496 150414
rect 227444 150350 227496 150356
rect 227456 149433 227484 150350
rect 232516 149734 232544 154527
rect 286140 151836 286192 151842
rect 286140 151778 286192 151784
rect 232136 149728 232188 149734
rect 232136 149670 232188 149676
rect 232504 149728 232556 149734
rect 232504 149670 232556 149676
rect 227442 149424 227498 149433
rect 227442 149359 227498 149368
rect 227444 149048 227496 149054
rect 227444 148990 227496 148996
rect 227456 148889 227484 148990
rect 227536 148980 227588 148986
rect 227536 148922 227588 148928
rect 227442 148880 227498 148889
rect 227442 148815 227498 148824
rect 227548 148209 227576 148922
rect 227534 148200 227590 148209
rect 227534 148135 227590 148144
rect 225602 147656 225658 147665
rect 224868 147620 224920 147626
rect 225602 147591 225658 147600
rect 226708 147620 226760 147626
rect 224868 147562 224920 147568
rect 226708 147562 226760 147568
rect 224776 147552 224828 147558
rect 224776 147494 224828 147500
rect 226524 147552 226576 147558
rect 226524 147494 226576 147500
rect 226536 146441 226564 147494
rect 226720 146985 226748 147562
rect 226706 146976 226762 146985
rect 226706 146911 226762 146920
rect 226522 146432 226578 146441
rect 226522 146367 226578 146376
rect 227628 146328 227680 146334
rect 227628 146270 227680 146276
rect 226708 146260 226760 146266
rect 226708 146202 226760 146208
rect 224500 146192 224552 146198
rect 224500 146134 224552 146140
rect 226720 145217 226748 146202
rect 227444 146192 227496 146198
rect 227444 146134 227496 146140
rect 227456 145897 227484 146134
rect 227442 145888 227498 145897
rect 227442 145823 227498 145832
rect 226706 145208 226762 145217
rect 226706 145143 226762 145152
rect 227260 144968 227312 144974
rect 227260 144910 227312 144916
rect 226524 144900 226576 144906
rect 226524 144842 226576 144848
rect 226536 143993 226564 144842
rect 226522 143984 226578 143993
rect 226522 143919 226578 143928
rect 226892 143540 226944 143546
rect 226892 143482 226944 143488
rect 224224 143472 224276 143478
rect 224224 143414 224276 143420
rect 226904 142905 226932 143482
rect 226890 142896 226946 142905
rect 226890 142831 226946 142840
rect 226708 142112 226760 142118
rect 226708 142054 226760 142060
rect 226720 141681 226748 142054
rect 226706 141672 226762 141681
rect 226706 141607 226762 141616
rect 227272 141001 227300 144910
rect 227444 144832 227496 144838
rect 227444 144774 227496 144780
rect 227456 144673 227484 144774
rect 227442 144664 227498 144673
rect 227442 144599 227498 144608
rect 227536 143608 227588 143614
rect 227536 143550 227588 143556
rect 227444 143472 227496 143478
rect 227442 143440 227444 143449
rect 227496 143440 227498 143449
rect 227442 143375 227498 143384
rect 227352 142180 227404 142186
rect 227352 142122 227404 142128
rect 227258 140992 227314 141001
rect 227258 140927 227314 140936
rect 226708 140820 226760 140826
rect 226708 140762 226760 140768
rect 226616 139528 226668 139534
rect 226616 139470 226668 139476
rect 226524 139460 226576 139466
rect 226524 139402 226576 139408
rect 226432 138032 226484 138038
rect 226432 137974 226484 137980
rect 226444 135697 226472 137974
rect 226536 136785 226564 139402
rect 226522 136776 226578 136785
rect 226522 136711 226578 136720
rect 226628 136241 226656 139470
rect 226720 137465 226748 140762
rect 227076 140752 227128 140758
rect 227076 140694 227128 140700
rect 227088 140457 227116 140694
rect 227074 140448 227130 140457
rect 227074 140383 227130 140392
rect 227364 138689 227392 142122
rect 227548 139777 227576 143550
rect 227640 142225 227668 146270
rect 227626 142216 227682 142225
rect 227626 142151 227682 142160
rect 227534 139768 227590 139777
rect 227534 139703 227590 139712
rect 227444 139392 227496 139398
rect 227444 139334 227496 139340
rect 227456 139233 227484 139334
rect 227442 139224 227498 139233
rect 227442 139159 227498 139168
rect 227350 138680 227406 138689
rect 227350 138615 227406 138624
rect 226800 138100 226852 138106
rect 226800 138042 226852 138048
rect 226706 137456 226762 137465
rect 226706 137391 226762 137400
rect 226614 136232 226670 136241
rect 226614 136167 226670 136176
rect 226430 135688 226486 135697
rect 226430 135623 226486 135632
rect 226524 135312 226576 135318
rect 226524 135254 226576 135260
rect 226536 133249 226564 135254
rect 226812 135017 226840 138042
rect 227442 138000 227498 138009
rect 227442 137935 227444 137944
rect 227496 137935 227498 137944
rect 227444 137906 227496 137912
rect 227260 136740 227312 136746
rect 227260 136682 227312 136688
rect 226798 135008 226854 135017
rect 226798 134943 226854 134952
rect 226708 134020 226760 134026
rect 226708 133962 226760 133968
rect 226522 133240 226578 133249
rect 226522 133175 226578 133184
rect 226720 132025 226748 133962
rect 227272 133793 227300 136682
rect 227444 136672 227496 136678
rect 227444 136614 227496 136620
rect 227456 134473 227484 136614
rect 227442 134464 227498 134473
rect 227442 134399 227498 134408
rect 227536 133952 227588 133958
rect 227536 133894 227588 133900
rect 227258 133784 227314 133793
rect 227258 133719 227314 133728
rect 227352 132592 227404 132598
rect 227548 132569 227576 133894
rect 227352 132534 227404 132540
rect 227534 132560 227590 132569
rect 226706 132016 226762 132025
rect 226706 131951 226762 131960
rect 226524 131232 226576 131238
rect 226524 131174 226576 131180
rect 226536 129577 226564 131174
rect 227076 131164 227128 131170
rect 227076 131106 227128 131112
rect 227088 130257 227116 131106
rect 227364 130801 227392 132534
rect 227444 132524 227496 132530
rect 227534 132495 227590 132504
rect 227444 132466 227496 132472
rect 227456 131481 227484 132466
rect 227442 131472 227498 131481
rect 227442 131407 227498 131416
rect 227350 130792 227406 130801
rect 227350 130727 227406 130736
rect 227074 130248 227130 130257
rect 227074 130183 227130 130192
rect 227536 129804 227588 129810
rect 227536 129746 227588 129752
rect 226522 129568 226578 129577
rect 226522 129503 226578 129512
rect 227444 129056 227496 129062
rect 227548 129033 227576 129746
rect 227444 128998 227496 129004
rect 227534 129024 227590 129033
rect 227456 128489 227484 128998
rect 227534 128959 227590 128968
rect 232148 128602 232176 149670
rect 286152 149668 286180 151778
rect 232056 128574 232176 128602
rect 227442 128480 227498 128489
rect 227442 128415 227498 128424
rect 226340 128376 226392 128382
rect 226340 128318 226392 128324
rect 226352 127809 226380 128318
rect 226338 127800 226394 127809
rect 226338 127735 226394 127744
rect 227444 127628 227496 127634
rect 227444 127570 227496 127576
rect 227456 127265 227484 127570
rect 227442 127256 227498 127265
rect 227442 127191 227498 127200
rect 227444 127016 227496 127022
rect 227444 126958 227496 126964
rect 227456 126585 227484 126958
rect 227442 126576 227498 126585
rect 227442 126511 227498 126520
rect 227444 126268 227496 126274
rect 227444 126210 227496 126216
rect 227456 126041 227484 126210
rect 227442 126032 227498 126041
rect 227442 125967 227498 125976
rect 227444 125656 227496 125662
rect 227444 125598 227496 125604
rect 227456 125361 227484 125598
rect 227442 125352 227498 125361
rect 227442 125287 227498 125296
rect 227260 124908 227312 124914
rect 227260 124850 227312 124856
rect 227272 124817 227300 124850
rect 227258 124808 227314 124817
rect 227258 124743 227314 124752
rect 227258 124264 227314 124273
rect 227258 124199 227314 124208
rect 227272 124166 227300 124199
rect 227260 124160 227312 124166
rect 227260 124102 227312 124108
rect 227258 123584 227314 123593
rect 227258 123519 227314 123528
rect 227272 123486 227300 123519
rect 227260 123480 227312 123486
rect 227260 123422 227312 123428
rect 227442 123040 227498 123049
rect 227442 122975 227498 122984
rect 227456 122806 227484 122975
rect 227444 122800 227496 122806
rect 227444 122742 227496 122748
rect 227442 122360 227498 122369
rect 227442 122295 227498 122304
rect 227456 122126 227484 122295
rect 227444 122120 227496 122126
rect 227444 122062 227496 122068
rect 227442 121816 227498 121825
rect 227442 121751 227498 121760
rect 227456 121446 227484 121751
rect 227444 121440 227496 121446
rect 227444 121382 227496 121388
rect 227442 121272 227498 121281
rect 227442 121207 227498 121216
rect 227456 120766 227484 121207
rect 227444 120760 227496 120766
rect 227444 120702 227496 120708
rect 227442 120592 227498 120601
rect 227442 120527 227498 120536
rect 227456 120086 227484 120527
rect 227444 120080 227496 120086
rect 226430 120048 226486 120057
rect 227444 120022 227496 120028
rect 226430 119983 226486 119992
rect 226338 119368 226394 119377
rect 226338 119303 226394 119312
rect 226246 118824 226302 118833
rect 226246 118759 226302 118768
rect 226154 117600 226210 117609
rect 226154 117535 226210 117544
rect 226168 115870 226196 117535
rect 226260 117230 226288 118759
rect 226352 118658 226380 119303
rect 226340 118652 226392 118658
rect 226340 118594 226392 118600
rect 226444 118590 226472 119983
rect 226432 118584 226484 118590
rect 226432 118526 226484 118532
rect 227442 118144 227498 118153
rect 227442 118079 227498 118088
rect 227456 117298 227484 118079
rect 227444 117292 227496 117298
rect 227444 117234 227496 117240
rect 226248 117224 226300 117230
rect 226248 117166 226300 117172
rect 227442 117056 227498 117065
rect 227442 116991 227498 117000
rect 226246 116376 226302 116385
rect 226246 116311 226302 116320
rect 226156 115864 226208 115870
rect 226156 115806 226208 115812
rect 226154 115152 226210 115161
rect 226154 115087 226210 115096
rect 226062 114608 226118 114617
rect 226062 114543 226118 114552
rect 225970 113384 226026 113393
rect 225970 113319 226026 113328
rect 225786 112160 225842 112169
rect 225786 112095 225842 112104
rect 225694 110392 225750 110401
rect 225694 110327 225750 110336
rect 225602 109168 225658 109177
rect 225602 109103 225658 109112
rect 224776 104916 224828 104922
rect 224776 104858 224828 104864
rect 224788 99278 224816 104858
rect 225616 104854 225644 109103
rect 225708 106282 225736 110327
rect 225800 108934 225828 112095
rect 225984 110430 226012 113319
rect 226076 111722 226104 114543
rect 226168 113150 226196 115087
rect 226260 114442 226288 116311
rect 227456 115938 227484 116991
rect 227444 115932 227496 115938
rect 227444 115874 227496 115880
rect 227074 115832 227130 115841
rect 232056 115818 232084 128574
rect 232056 115790 232176 115818
rect 227074 115767 227130 115776
rect 227088 114510 227116 115767
rect 227076 114504 227128 114510
rect 227076 114446 227128 114452
rect 226248 114436 226300 114442
rect 226248 114378 226300 114384
rect 226246 114064 226302 114073
rect 226246 113999 226302 114008
rect 226156 113144 226208 113150
rect 226156 113086 226208 113092
rect 226154 112840 226210 112849
rect 226154 112775 226210 112784
rect 226064 111716 226116 111722
rect 226064 111658 226116 111664
rect 226062 110936 226118 110945
rect 226062 110871 226118 110880
rect 225972 110424 226024 110430
rect 225972 110366 226024 110372
rect 225788 108928 225840 108934
rect 225788 108870 225840 108876
rect 225786 107944 225842 107953
rect 225786 107879 225842 107888
rect 225696 106276 225748 106282
rect 225696 106218 225748 106224
rect 225604 104848 225656 104854
rect 225604 104790 225656 104796
rect 224868 103692 224920 103698
rect 224868 103634 224920 103640
rect 224776 99272 224828 99278
rect 224776 99214 224828 99220
rect 224880 97986 224908 103634
rect 225800 103426 225828 107879
rect 226076 107642 226104 110871
rect 226168 110362 226196 112775
rect 226260 111790 226288 113999
rect 226248 111784 226300 111790
rect 226248 111726 226300 111732
rect 226246 111616 226302 111625
rect 226246 111551 226302 111560
rect 226156 110356 226208 110362
rect 226156 110298 226208 110304
rect 226154 109848 226210 109857
rect 226154 109783 226210 109792
rect 226064 107636 226116 107642
rect 226064 107578 226116 107584
rect 226062 107400 226118 107409
rect 226062 107335 226118 107344
rect 225878 106856 225934 106865
rect 225878 106791 225934 106800
rect 225788 103420 225840 103426
rect 225788 103362 225840 103368
rect 225892 102134 225920 106791
rect 225970 106176 226026 106185
rect 225970 106111 226026 106120
rect 225880 102128 225932 102134
rect 225880 102070 225932 102076
rect 225984 100638 226012 106111
rect 226076 103494 226104 107335
rect 226168 106214 226196 109783
rect 226260 109002 226288 111551
rect 226248 108996 226300 109002
rect 226248 108938 226300 108944
rect 226246 108624 226302 108633
rect 226246 108559 226302 108568
rect 226156 106208 226208 106214
rect 226156 106150 226208 106156
rect 226154 105632 226210 105641
rect 226154 105567 226210 105576
rect 226064 103488 226116 103494
rect 226064 103430 226116 103436
rect 226168 100706 226196 105567
rect 226260 104786 226288 108559
rect 227442 104952 227498 104961
rect 227442 104887 227444 104896
rect 227496 104887 227498 104896
rect 227444 104858 227496 104864
rect 226248 104780 226300 104786
rect 226248 104722 226300 104728
rect 226246 104408 226302 104417
rect 226246 104343 226302 104352
rect 226156 100700 226208 100706
rect 226156 100642 226208 100648
rect 225972 100632 226024 100638
rect 225972 100574 226024 100580
rect 226260 99346 226288 104343
rect 227442 103864 227498 103873
rect 227442 103799 227498 103808
rect 227456 103698 227484 103799
rect 227444 103692 227496 103698
rect 227444 103634 227496 103640
rect 232148 100706 232176 115790
rect 258092 100706 258120 103564
rect 314212 102134 314240 103564
rect 338408 102134 338436 428567
rect 343638 428496 343694 428505
rect 343638 428431 343694 428440
rect 341524 310548 341576 310554
rect 341524 310490 341576 310496
rect 340144 309188 340196 309194
rect 340144 309130 340196 309136
rect 314200 102128 314252 102134
rect 314200 102070 314252 102076
rect 338396 102128 338448 102134
rect 338396 102070 338448 102076
rect 232136 100700 232188 100706
rect 232136 100642 232188 100648
rect 258080 100700 258132 100706
rect 258080 100642 258132 100648
rect 232148 99346 232176 100642
rect 226248 99340 226300 99346
rect 226248 99282 226300 99288
rect 232136 99340 232188 99346
rect 232136 99282 232188 99288
rect 232504 99340 232556 99346
rect 232504 99282 232556 99288
rect 224868 97980 224920 97986
rect 224868 97922 224920 97928
rect 218704 97028 218756 97034
rect 218704 96970 218756 96976
rect 215116 95192 215168 95198
rect 214746 95160 214802 95169
rect 215116 95134 215168 95140
rect 214746 95095 214802 95104
rect 215128 94353 215156 95134
rect 215114 94344 215170 94353
rect 215114 94279 215170 94288
rect 215208 93832 215260 93838
rect 215208 93774 215260 93780
rect 215116 93764 215168 93770
rect 215116 93706 215168 93712
rect 215128 93673 215156 93706
rect 215114 93664 215170 93673
rect 215114 93599 215170 93608
rect 116676 93152 116728 93158
rect 116676 93094 116728 93100
rect 215220 92857 215248 93774
rect 215206 92848 215262 92857
rect 215206 92783 215262 92792
rect 214562 92032 214618 92041
rect 214562 91967 214618 91976
rect 214470 90536 214526 90545
rect 214470 90471 214526 90480
rect 214484 89758 214512 90471
rect 214472 89752 214524 89758
rect 214472 89694 214524 89700
rect 214102 88904 214158 88913
rect 214102 88839 214158 88848
rect 214116 88398 214144 88839
rect 214104 88392 214156 88398
rect 214104 88334 214156 88340
rect 117042 84552 117098 84561
rect 117042 84487 117098 84496
rect 116584 80708 116636 80714
rect 116584 80650 116636 80656
rect 116400 80096 116452 80102
rect 116400 80038 116452 80044
rect 116398 79928 116454 79937
rect 116398 79863 116454 79872
rect 116412 78742 116440 79863
rect 117056 79354 117084 84487
rect 214194 82648 214250 82657
rect 214194 82583 214250 82592
rect 214208 81462 214236 82583
rect 214196 81456 214248 81462
rect 214196 81398 214248 81404
rect 214576 81394 214604 91967
rect 214746 91216 214802 91225
rect 214746 91151 214802 91160
rect 214654 84960 214710 84969
rect 214654 84895 214710 84904
rect 214564 81388 214616 81394
rect 214564 81330 214616 81336
rect 214010 81016 214066 81025
rect 214010 80951 214066 80960
rect 214024 80102 214052 80951
rect 214012 80096 214064 80102
rect 214012 80038 214064 80044
rect 117044 79348 117096 79354
rect 117044 79290 117096 79296
rect 116400 78736 116452 78742
rect 116400 78678 116452 78684
rect 116582 78704 116638 78713
rect 116582 78639 116638 78648
rect 214562 78704 214618 78713
rect 214562 78639 214618 78648
rect 104256 77988 104308 77994
rect 104256 77930 104308 77936
rect 116398 77480 116454 77489
rect 116398 77415 116454 77424
rect 116412 77314 116440 77415
rect 116400 77308 116452 77314
rect 116400 77250 116452 77256
rect 102876 76900 102928 76906
rect 102876 76842 102928 76848
rect 116398 76392 116454 76401
rect 116398 76327 116454 76336
rect 116412 75954 116440 76327
rect 116400 75948 116452 75954
rect 116400 75890 116452 75896
rect 116398 75168 116454 75177
rect 116398 75103 116454 75112
rect 116412 74594 116440 75103
rect 116400 74588 116452 74594
rect 116400 74530 116452 74536
rect 116398 74080 116454 74089
rect 116398 74015 116454 74024
rect 116412 73234 116440 74015
rect 116596 73846 116624 78639
rect 214470 77208 214526 77217
rect 214470 77143 214526 77152
rect 214286 74080 214342 74089
rect 214286 74015 214342 74024
rect 116584 73840 116636 73846
rect 116584 73782 116636 73788
rect 116400 73228 116452 73234
rect 116400 73170 116452 73176
rect 116398 72856 116454 72865
rect 116398 72791 116454 72800
rect 116412 71806 116440 72791
rect 116400 71800 116452 71806
rect 116306 71768 116362 71777
rect 116400 71742 116452 71748
rect 116306 71703 116362 71712
rect 116320 70514 116348 71703
rect 214102 71632 214158 71641
rect 214102 71567 214158 71576
rect 116398 70544 116454 70553
rect 116308 70508 116360 70514
rect 116398 70479 116454 70488
rect 116308 70450 116360 70456
rect 116412 70446 116440 70479
rect 214116 70446 214144 71567
rect 116400 70440 116452 70446
rect 116400 70382 116452 70388
rect 214104 70440 214156 70446
rect 214104 70382 214156 70388
rect 102784 69896 102836 69902
rect 102784 69838 102836 69844
rect 116398 69320 116454 69329
rect 116398 69255 116454 69264
rect 116412 69086 116440 69255
rect 116400 69080 116452 69086
rect 116400 69022 116452 69028
rect 116398 68232 116454 68241
rect 116398 68167 116454 68176
rect 116412 67658 116440 68167
rect 116400 67652 116452 67658
rect 116400 67594 116452 67600
rect 116398 67008 116454 67017
rect 116398 66943 116454 66952
rect 116412 66298 116440 66943
rect 116400 66292 116452 66298
rect 116400 66234 116452 66240
rect 214300 66230 214328 74015
rect 214484 69018 214512 77143
rect 214576 70378 214604 78639
rect 214668 75886 214696 84895
rect 214760 81326 214788 91151
rect 227352 89752 227404 89758
rect 215114 89720 215170 89729
rect 227352 89694 227404 89700
rect 215114 89655 215170 89664
rect 215128 88466 215156 89655
rect 215116 88460 215168 88466
rect 215116 88402 215168 88408
rect 221464 88460 221516 88466
rect 221464 88402 221516 88408
rect 215022 88088 215078 88097
rect 215022 88023 215078 88032
rect 215036 87106 215064 88023
rect 215114 87408 215170 87417
rect 215114 87343 215170 87352
rect 215024 87100 215076 87106
rect 215024 87042 215076 87048
rect 215128 87038 215156 87343
rect 218704 87100 218756 87106
rect 218704 87042 218756 87048
rect 215116 87032 215168 87038
rect 215116 86974 215168 86980
rect 215206 86592 215262 86601
rect 215206 86527 215262 86536
rect 215114 85776 215170 85785
rect 215114 85711 215170 85720
rect 215128 85610 215156 85711
rect 215116 85604 215168 85610
rect 215116 85546 215168 85552
rect 215220 85354 215248 86527
rect 215128 85326 215248 85354
rect 214838 83464 214894 83473
rect 214838 83399 214894 83408
rect 214748 81320 214800 81326
rect 214748 81262 214800 81268
rect 214746 77888 214802 77897
rect 214746 77823 214802 77832
rect 214760 77314 214788 77823
rect 214748 77308 214800 77314
rect 214748 77250 214800 77256
rect 214656 75880 214708 75886
rect 214656 75822 214708 75828
rect 214852 74526 214880 83399
rect 214930 81832 214986 81841
rect 214930 81767 214986 81776
rect 214840 74520 214892 74526
rect 214840 74462 214892 74468
rect 214840 73500 214892 73506
rect 214840 73442 214892 73448
rect 214654 72448 214710 72457
rect 214654 72383 214710 72392
rect 214564 70372 214616 70378
rect 214564 70314 214616 70320
rect 214472 69012 214524 69018
rect 214472 68954 214524 68960
rect 214288 66224 214340 66230
rect 213918 66192 213974 66201
rect 214288 66166 214340 66172
rect 213918 66127 213974 66136
rect 101404 65952 101456 65958
rect 101404 65894 101456 65900
rect 116398 65920 116454 65929
rect 116398 65855 116454 65864
rect 116412 64938 116440 65855
rect 213932 65210 213960 66127
rect 214010 65376 214066 65385
rect 214010 65311 214066 65320
rect 213920 65204 213972 65210
rect 213920 65146 213972 65152
rect 214024 64938 214052 65311
rect 116400 64932 116452 64938
rect 116400 64874 116452 64880
rect 214012 64932 214064 64938
rect 214012 64874 214064 64880
rect 214668 64734 214696 72383
rect 214852 67590 214880 73442
rect 214944 73166 214972 81767
rect 215128 80730 215156 85326
rect 215206 84280 215262 84289
rect 215206 84215 215208 84224
rect 215260 84215 215262 84224
rect 215208 84186 215260 84192
rect 215944 82884 215996 82890
rect 215944 82826 215996 82832
rect 215128 80702 215248 80730
rect 215022 80336 215078 80345
rect 215022 80271 215078 80280
rect 214932 73160 214984 73166
rect 214932 73102 214984 73108
rect 215036 71738 215064 80271
rect 215114 79520 215170 79529
rect 215114 79455 215170 79464
rect 215128 78810 215156 79455
rect 215116 78804 215168 78810
rect 215116 78746 215168 78752
rect 215220 77246 215248 80702
rect 215208 77240 215260 77246
rect 215208 77182 215260 77188
rect 215206 76392 215262 76401
rect 215206 76327 215262 76336
rect 215220 75954 215248 76327
rect 215208 75948 215260 75954
rect 215208 75890 215260 75896
rect 215114 75576 215170 75585
rect 215114 75511 215170 75520
rect 215128 73506 215156 75511
rect 215206 74760 215262 74769
rect 215206 74695 215262 74704
rect 215220 74662 215248 74695
rect 215208 74656 215260 74662
rect 215208 74598 215260 74604
rect 215116 73500 215168 73506
rect 215116 73442 215168 73448
rect 215116 73364 215168 73370
rect 215116 73306 215168 73312
rect 215128 73273 215156 73306
rect 215114 73264 215170 73273
rect 215114 73199 215170 73208
rect 215024 71732 215076 71738
rect 215024 71674 215076 71680
rect 215114 70952 215170 70961
rect 215114 70887 215170 70896
rect 215128 70514 215156 70887
rect 215116 70508 215168 70514
rect 215116 70450 215168 70456
rect 214930 70136 214986 70145
rect 214930 70071 214986 70080
rect 214944 69154 214972 70071
rect 215114 69320 215170 69329
rect 215114 69255 215170 69264
rect 214932 69148 214984 69154
rect 214932 69090 214984 69096
rect 215128 69086 215156 69255
rect 215116 69080 215168 69086
rect 215116 69022 215168 69028
rect 215206 68504 215262 68513
rect 215206 68439 215262 68448
rect 215114 67824 215170 67833
rect 215114 67759 215170 67768
rect 215128 67658 215156 67759
rect 215220 67726 215248 68439
rect 215208 67720 215260 67726
rect 215208 67662 215260 67668
rect 215116 67652 215168 67658
rect 215116 67594 215168 67600
rect 214840 67584 214892 67590
rect 214840 67526 214892 67532
rect 215114 67008 215170 67017
rect 215114 66943 215170 66952
rect 215128 66298 215156 66943
rect 215116 66292 215168 66298
rect 215116 66234 215168 66240
rect 214656 64728 214708 64734
rect 115938 64696 115994 64705
rect 214656 64670 214708 64676
rect 115938 64631 115994 64640
rect 115952 63578 115980 64631
rect 214102 64560 214158 64569
rect 214102 64495 214158 64504
rect 214116 63646 214144 64495
rect 215114 63880 215170 63889
rect 215114 63815 215170 63824
rect 214104 63640 214156 63646
rect 214104 63582 214156 63588
rect 215128 63578 215156 63815
rect 115940 63572 115992 63578
rect 115940 63514 115992 63520
rect 215116 63572 215168 63578
rect 215116 63514 215168 63520
rect 116398 63472 116454 63481
rect 116398 63407 116454 63416
rect 116412 62150 116440 63407
rect 214378 63064 214434 63073
rect 214378 62999 214434 63008
rect 116490 62384 116546 62393
rect 116490 62319 116546 62328
rect 116400 62144 116452 62150
rect 116400 62086 116452 62092
rect 100024 61804 100076 61810
rect 100024 61746 100076 61752
rect 116398 61160 116454 61169
rect 116398 61095 116454 61104
rect 116412 60790 116440 61095
rect 116400 60784 116452 60790
rect 116400 60726 116452 60732
rect 116398 60072 116454 60081
rect 116504 60042 116532 62319
rect 214392 62218 214420 62999
rect 215114 62248 215170 62257
rect 214380 62212 214432 62218
rect 215114 62183 215170 62192
rect 214380 62154 214432 62160
rect 215128 62150 215156 62183
rect 215116 62144 215168 62150
rect 215116 62086 215168 62092
rect 214746 61432 214802 61441
rect 214746 61367 214802 61376
rect 214760 60858 214788 61367
rect 214748 60852 214800 60858
rect 214748 60794 214800 60800
rect 215116 60784 215168 60790
rect 215114 60752 215116 60761
rect 215168 60752 215170 60761
rect 215114 60687 215170 60696
rect 116398 60007 116454 60016
rect 116492 60036 116544 60042
rect 116412 59430 116440 60007
rect 116492 59978 116544 59984
rect 214378 59936 214434 59945
rect 214378 59871 214434 59880
rect 214392 59430 214420 59871
rect 97356 59424 97408 59430
rect 97356 59366 97408 59372
rect 116400 59424 116452 59430
rect 116400 59366 116452 59372
rect 214380 59424 214432 59430
rect 214380 59366 214432 59372
rect 97264 57928 97316 57934
rect 97264 57870 97316 57876
rect 96160 54732 96212 54738
rect 96160 54674 96212 54680
rect 97368 52426 97396 59366
rect 214286 59120 214342 59129
rect 214286 59055 214342 59064
rect 116398 58848 116454 58857
rect 116398 58783 116454 58792
rect 116412 58002 116440 58783
rect 214300 58070 214328 59055
rect 214378 58304 214434 58313
rect 214378 58239 214434 58248
rect 214288 58064 214340 58070
rect 214288 58006 214340 58012
rect 214392 58002 214420 58239
rect 116400 57996 116452 58002
rect 116400 57938 116452 57944
rect 214380 57996 214432 58002
rect 214380 57938 214432 57944
rect 116306 57624 116362 57633
rect 116306 57559 116362 57568
rect 213918 57624 213974 57633
rect 213918 57559 213974 57568
rect 116320 56642 116348 57559
rect 213932 56710 213960 57559
rect 214010 56808 214066 56817
rect 214010 56743 214066 56752
rect 213920 56704 213972 56710
rect 213920 56646 213972 56652
rect 214024 56642 214052 56743
rect 116308 56636 116360 56642
rect 116308 56578 116360 56584
rect 214012 56636 214064 56642
rect 214012 56578 214064 56584
rect 116306 56536 116362 56545
rect 116306 56471 116362 56480
rect 116320 55350 116348 56471
rect 215114 55992 215170 56001
rect 215114 55927 215170 55936
rect 116308 55344 116360 55350
rect 116308 55286 116360 55292
rect 116398 55312 116454 55321
rect 215128 55282 215156 55927
rect 116398 55247 116400 55256
rect 116452 55247 116454 55256
rect 215116 55276 215168 55282
rect 116400 55218 116452 55224
rect 215116 55218 215168 55224
rect 214746 55176 214802 55185
rect 214746 55111 214802 55120
rect 116398 54224 116454 54233
rect 116398 54159 116454 54168
rect 116412 53854 116440 54159
rect 214760 53922 214788 55111
rect 215114 54496 215170 54505
rect 215114 54431 215170 54440
rect 214748 53916 214800 53922
rect 214748 53858 214800 53864
rect 215128 53854 215156 54431
rect 116400 53848 116452 53854
rect 116400 53790 116452 53796
rect 215116 53848 215168 53854
rect 215116 53790 215168 53796
rect 214746 53680 214802 53689
rect 214746 53615 214802 53624
rect 116398 53000 116454 53009
rect 116398 52935 116454 52944
rect 116412 52494 116440 52935
rect 214760 52494 214788 53615
rect 215114 52864 215170 52873
rect 215114 52799 215170 52808
rect 215128 52562 215156 52799
rect 215116 52556 215168 52562
rect 215116 52498 215168 52504
rect 116400 52488 116452 52494
rect 116400 52430 116452 52436
rect 214748 52488 214800 52494
rect 214748 52430 214800 52436
rect 97356 52420 97408 52426
rect 97356 52362 97408 52368
rect 214562 52048 214618 52057
rect 214562 51983 214618 51992
rect 115938 51912 115994 51921
rect 115938 51847 115994 51856
rect 115952 51134 115980 51847
rect 214576 51134 214604 51983
rect 215114 51368 215170 51377
rect 215114 51303 215170 51312
rect 215128 51202 215156 51303
rect 215116 51196 215168 51202
rect 215116 51138 215168 51144
rect 115940 51128 115992 51134
rect 115940 51070 115992 51076
rect 214564 51128 214616 51134
rect 214564 51070 214616 51076
rect 95202 50646 95280 50674
rect 116398 50688 116454 50697
rect 95146 50623 95202 50632
rect 116398 50623 116454 50632
rect 116412 49774 116440 50623
rect 214378 50552 214434 50561
rect 214378 50487 214434 50496
rect 214392 49842 214420 50487
rect 214380 49836 214432 49842
rect 214380 49778 214432 49784
rect 95148 49768 95200 49774
rect 95148 49710 95200 49716
rect 116400 49768 116452 49774
rect 215116 49768 215168 49774
rect 116400 49710 116452 49716
rect 215114 49736 215116 49745
rect 215168 49736 215170 49745
rect 95054 46200 95110 46209
rect 95054 46135 95110 46144
rect 95160 45257 95188 49710
rect 215114 49671 215170 49680
rect 116398 49464 116454 49473
rect 116398 49399 116454 49408
rect 116124 48408 116176 48414
rect 116122 48376 116124 48385
rect 116176 48376 116178 48385
rect 116412 48346 116440 49399
rect 215114 48920 215170 48929
rect 215114 48855 215170 48864
rect 215128 48346 215156 48855
rect 116122 48311 116178 48320
rect 116400 48340 116452 48346
rect 116400 48282 116452 48288
rect 215116 48340 215168 48346
rect 215116 48282 215168 48288
rect 214746 48104 214802 48113
rect 214746 48039 214802 48048
rect 214010 47424 214066 47433
rect 214010 47359 214066 47368
rect 116398 47152 116454 47161
rect 116398 47087 116454 47096
rect 116412 46986 116440 47087
rect 214024 46986 214052 47359
rect 214760 47054 214788 48039
rect 214748 47048 214800 47054
rect 214748 46990 214800 46996
rect 116400 46980 116452 46986
rect 116400 46922 116452 46928
rect 214012 46980 214064 46986
rect 214012 46922 214064 46928
rect 215206 46608 215262 46617
rect 215206 46543 215262 46552
rect 116398 46064 116454 46073
rect 116398 45999 116454 46008
rect 116412 45626 116440 45999
rect 215114 45792 215170 45801
rect 215114 45727 215170 45736
rect 215128 45694 215156 45727
rect 215116 45688 215168 45694
rect 215116 45630 215168 45636
rect 215220 45626 215248 46543
rect 116400 45620 116452 45626
rect 116400 45562 116452 45568
rect 215208 45620 215260 45626
rect 215208 45562 215260 45568
rect 95146 45248 95202 45257
rect 95146 45183 95202 45192
rect 214470 44976 214526 44985
rect 214470 44911 214526 44920
rect 116398 44840 116454 44849
rect 116398 44775 116454 44784
rect 116412 44198 116440 44775
rect 214484 44198 214512 44911
rect 215114 44296 215170 44305
rect 215114 44231 215116 44240
rect 215168 44231 215170 44240
rect 215116 44202 215168 44208
rect 95056 44192 95108 44198
rect 95056 44134 95108 44140
rect 116400 44192 116452 44198
rect 116400 44134 116452 44140
rect 214472 44192 214524 44198
rect 214472 44134 214524 44140
rect 94962 43480 95018 43489
rect 94962 43415 95018 43424
rect 94596 42832 94648 42838
rect 94596 42774 94648 42780
rect 94134 42528 94190 42537
rect 94134 42463 94190 42472
rect 93950 41712 94006 41721
rect 93950 41647 94006 41656
rect 94504 40180 94556 40186
rect 94504 40122 94556 40128
rect 94516 38185 94544 40122
rect 94608 39953 94636 42774
rect 95068 40769 95096 44134
rect 115938 43616 115994 43625
rect 115938 43551 115994 43560
rect 115952 42838 115980 43551
rect 214378 43480 214434 43489
rect 214378 43415 214434 43424
rect 214392 42838 214420 43415
rect 115940 42832 115992 42838
rect 115940 42774 115992 42780
rect 214380 42832 214432 42838
rect 214380 42774 214432 42780
rect 214102 42664 214158 42673
rect 214102 42599 214158 42608
rect 116398 42528 116454 42537
rect 116398 42463 116454 42472
rect 116412 41478 116440 42463
rect 214116 41478 214144 42599
rect 215114 41848 215170 41857
rect 215114 41783 215170 41792
rect 215128 41546 215156 41783
rect 215116 41540 215168 41546
rect 215116 41482 215168 41488
rect 95148 41472 95200 41478
rect 95148 41414 95200 41420
rect 116400 41472 116452 41478
rect 116400 41414 116452 41420
rect 214104 41472 214156 41478
rect 214104 41414 214156 41420
rect 95054 40760 95110 40769
rect 95054 40695 95110 40704
rect 95056 40112 95108 40118
rect 95056 40054 95108 40060
rect 94594 39944 94650 39953
rect 94594 39879 94650 39888
rect 94596 38684 94648 38690
rect 94596 38626 94648 38632
rect 94502 38176 94558 38185
rect 94502 38111 94558 38120
rect 93860 37324 93912 37330
rect 93860 37266 93912 37272
rect 93872 35465 93900 37266
rect 94608 36281 94636 38626
rect 95068 37233 95096 40054
rect 95160 39001 95188 41414
rect 116306 41304 116362 41313
rect 116306 41239 116362 41248
rect 116320 40186 116348 41239
rect 214654 41168 214710 41177
rect 214654 41103 214710 41112
rect 116398 40216 116454 40225
rect 116308 40180 116360 40186
rect 116398 40151 116454 40160
rect 116308 40122 116360 40128
rect 116412 40118 116440 40151
rect 214668 40118 214696 41103
rect 215114 40352 215170 40361
rect 215114 40287 215170 40296
rect 215128 40186 215156 40287
rect 215116 40180 215168 40186
rect 215116 40122 215168 40128
rect 116400 40112 116452 40118
rect 116400 40054 116452 40060
rect 214656 40112 214708 40118
rect 214656 40054 214708 40060
rect 214470 39536 214526 39545
rect 214470 39471 214526 39480
rect 95146 38992 95202 39001
rect 95146 38927 95202 38936
rect 116398 38992 116454 39001
rect 116398 38927 116454 38936
rect 116412 38690 116440 38927
rect 214484 38758 214512 39471
rect 214472 38752 214524 38758
rect 214472 38694 214524 38700
rect 215114 38720 215170 38729
rect 116400 38684 116452 38690
rect 215114 38655 215116 38664
rect 116400 38626 116452 38632
rect 215168 38655 215170 38664
rect 215116 38626 215168 38632
rect 215114 38040 215170 38049
rect 215114 37975 215170 37984
rect 116398 37768 116454 37777
rect 116398 37703 116454 37712
rect 116412 37330 116440 37703
rect 215128 37330 215156 37975
rect 116400 37324 116452 37330
rect 116400 37266 116452 37272
rect 215116 37324 215168 37330
rect 215116 37266 215168 37272
rect 95054 37224 95110 37233
rect 95054 37159 95110 37168
rect 215114 37224 215170 37233
rect 215114 37159 215170 37168
rect 116398 36680 116454 36689
rect 116398 36615 116454 36624
rect 94594 36272 94650 36281
rect 94594 36207 94650 36216
rect 116412 35970 116440 36615
rect 214562 36408 214618 36417
rect 214562 36343 214618 36352
rect 214576 36038 214604 36343
rect 214564 36032 214616 36038
rect 214564 35974 214616 35980
rect 215128 35970 215156 37159
rect 93952 35964 94004 35970
rect 93952 35906 94004 35912
rect 116400 35964 116452 35970
rect 116400 35906 116452 35912
rect 215116 35964 215168 35970
rect 215116 35906 215168 35912
rect 93858 35456 93914 35465
rect 93858 35391 93914 35400
rect 93964 34513 93992 35906
rect 214654 35592 214710 35601
rect 214654 35527 214710 35536
rect 116398 35456 116454 35465
rect 116398 35391 116454 35400
rect 116412 34542 116440 35391
rect 214668 34542 214696 35527
rect 215114 34912 215170 34921
rect 215114 34847 215170 34856
rect 215128 34610 215156 34847
rect 215116 34604 215168 34610
rect 215116 34546 215168 34552
rect 95148 34536 95200 34542
rect 93950 34504 94006 34513
rect 95148 34478 95200 34484
rect 116400 34536 116452 34542
rect 116400 34478 116452 34484
rect 214656 34536 214708 34542
rect 214656 34478 214708 34484
rect 93950 34439 94006 34448
rect 95160 33697 95188 34478
rect 116306 34368 116362 34377
rect 116306 34303 116362 34312
rect 95146 33688 95202 33697
rect 95146 33623 95202 33632
rect 116320 33182 116348 34303
rect 214562 34096 214618 34105
rect 214562 34031 214618 34040
rect 214576 33182 214604 34031
rect 215114 33280 215170 33289
rect 215114 33215 215116 33224
rect 215168 33215 215170 33224
rect 215116 33186 215168 33192
rect 95148 33176 95200 33182
rect 95148 33118 95200 33124
rect 116308 33176 116360 33182
rect 214564 33176 214616 33182
rect 116308 33118 116360 33124
rect 116398 33144 116454 33153
rect 95160 32745 95188 33118
rect 214564 33118 214616 33124
rect 116398 33079 116454 33088
rect 95146 32736 95202 32745
rect 95146 32671 95202 32680
rect 116412 32434 116440 33079
rect 215956 32570 215984 82826
rect 216128 80096 216180 80102
rect 216128 80038 216180 80044
rect 216036 74656 216088 74662
rect 216036 74598 216088 74604
rect 216048 67522 216076 74598
rect 216140 73098 216168 80038
rect 218716 78674 218744 87042
rect 221476 80034 221504 88402
rect 222844 88392 222896 88398
rect 222844 88334 222896 88340
rect 221464 80028 221516 80034
rect 221464 79970 221516 79976
rect 221556 78804 221608 78810
rect 221556 78746 221608 78752
rect 218704 78668 218756 78674
rect 218704 78610 218756 78616
rect 218796 77308 218848 77314
rect 218796 77250 218848 77256
rect 218060 75948 218112 75954
rect 218060 75890 218112 75896
rect 216128 73092 216180 73098
rect 216128 73034 216180 73040
rect 218072 68950 218100 75890
rect 218808 70310 218836 77250
rect 220728 73364 220780 73370
rect 220728 73306 220780 73312
rect 218796 70304 218848 70310
rect 218796 70246 218848 70252
rect 218060 68944 218112 68950
rect 218060 68886 218112 68892
rect 216036 67516 216088 67522
rect 216036 67458 216088 67464
rect 220740 66162 220768 73306
rect 221568 71670 221596 78746
rect 222856 78606 222884 88334
rect 224224 87032 224276 87038
rect 224224 86974 224276 86980
rect 222844 78600 222896 78606
rect 222844 78542 222896 78548
rect 224236 77178 224264 86974
rect 225604 85604 225656 85610
rect 225604 85546 225656 85552
rect 224224 77172 224276 77178
rect 224224 77114 224276 77120
rect 225616 75857 225644 85546
rect 227076 84244 227128 84250
rect 227076 84186 227128 84192
rect 225602 75848 225658 75857
rect 225602 75783 225658 75792
rect 227088 74633 227116 84186
rect 227168 81456 227220 81462
rect 227168 81398 227220 81404
rect 227074 74624 227130 74633
rect 227074 74559 227130 74568
rect 227180 73273 227208 81398
rect 227364 79801 227392 89694
rect 232516 86970 232544 99282
rect 340156 88330 340184 309130
rect 341536 135250 341564 310490
rect 341524 135244 341576 135250
rect 341524 135186 341576 135192
rect 343652 126721 343680 428431
rect 411996 225616 412048 225622
rect 411996 225558 412048 225564
rect 411904 222896 411956 222902
rect 411904 222838 411956 222844
rect 343638 126712 343694 126721
rect 343638 126647 343694 126656
rect 340144 88324 340196 88330
rect 340144 88266 340196 88272
rect 232320 86964 232372 86970
rect 232320 86906 232372 86912
rect 232504 86964 232556 86970
rect 232504 86906 232556 86912
rect 227444 81388 227496 81394
rect 227444 81330 227496 81336
rect 227456 81161 227484 81330
rect 227536 81320 227588 81326
rect 227536 81262 227588 81268
rect 227442 81152 227498 81161
rect 227442 81087 227498 81096
rect 227548 80481 227576 81262
rect 227534 80472 227590 80481
rect 227534 80407 227590 80416
rect 232332 80102 232360 86906
rect 320824 83564 320876 83570
rect 320824 83506 320876 83512
rect 284484 83496 284536 83502
rect 284484 83438 284536 83444
rect 248144 82884 248196 82890
rect 248144 82826 248196 82832
rect 248156 81396 248184 82826
rect 284496 81396 284524 83438
rect 320836 81396 320864 83506
rect 232320 80096 232372 80102
rect 232320 80038 232372 80044
rect 227444 80028 227496 80034
rect 227444 79970 227496 79976
rect 227350 79792 227406 79801
rect 227350 79727 227406 79736
rect 227456 79121 227484 79970
rect 232320 79960 232372 79966
rect 232320 79902 232372 79908
rect 227442 79112 227498 79121
rect 227442 79047 227498 79056
rect 227536 78668 227588 78674
rect 227536 78610 227588 78616
rect 227444 78600 227496 78606
rect 227442 78568 227444 78577
rect 227496 78568 227498 78577
rect 227442 78503 227498 78512
rect 227548 77897 227576 78610
rect 227534 77888 227590 77897
rect 227534 77823 227590 77832
rect 227536 77240 227588 77246
rect 227442 77208 227498 77217
rect 227536 77182 227588 77188
rect 227442 77143 227444 77152
rect 227496 77143 227498 77152
rect 227444 77114 227496 77120
rect 227548 76537 227576 77182
rect 227534 76528 227590 76537
rect 227534 76463 227590 76472
rect 227444 75880 227496 75886
rect 227444 75822 227496 75828
rect 227456 75313 227484 75822
rect 227442 75304 227498 75313
rect 227442 75239 227498 75248
rect 227444 74520 227496 74526
rect 227444 74462 227496 74468
rect 227456 73953 227484 74462
rect 227442 73944 227498 73953
rect 227442 73879 227498 73888
rect 227166 73264 227222 73273
rect 227166 73199 227222 73208
rect 227444 73160 227496 73166
rect 227444 73102 227496 73108
rect 227456 72729 227484 73102
rect 227536 73092 227588 73098
rect 227536 73034 227588 73040
rect 227442 72720 227498 72729
rect 227442 72655 227498 72664
rect 227548 72049 227576 73034
rect 227534 72040 227590 72049
rect 227534 71975 227590 71984
rect 227444 71732 227496 71738
rect 227444 71674 227496 71680
rect 221556 71664 221608 71670
rect 221556 71606 221608 71612
rect 227456 71369 227484 71674
rect 227536 71664 227588 71670
rect 227536 71606 227588 71612
rect 227442 71360 227498 71369
rect 227442 71295 227498 71304
rect 227548 70689 227576 71606
rect 227534 70680 227590 70689
rect 227534 70615 227590 70624
rect 224132 70508 224184 70514
rect 224132 70450 224184 70456
rect 220728 66156 220780 66162
rect 220728 66098 220780 66104
rect 216864 65204 216916 65210
rect 216864 65146 216916 65152
rect 216680 62212 216732 62218
rect 216680 62154 216732 62160
rect 216692 57934 216720 62154
rect 216772 60852 216824 60858
rect 216772 60794 216824 60800
rect 216680 57928 216732 57934
rect 216680 57870 216732 57876
rect 216680 56636 216732 56642
rect 216680 56578 216732 56584
rect 216692 52426 216720 56578
rect 216784 56574 216812 60794
rect 216876 60722 216904 65146
rect 224144 64258 224172 70450
rect 224868 70440 224920 70446
rect 224868 70382 224920 70388
rect 224408 69148 224460 69154
rect 224408 69090 224460 69096
rect 224224 67720 224276 67726
rect 224224 67662 224276 67668
rect 224132 64252 224184 64258
rect 224132 64194 224184 64200
rect 216956 63640 217008 63646
rect 216956 63582 217008 63588
rect 216864 60716 216916 60722
rect 216864 60658 216916 60664
rect 216968 59362 216996 63582
rect 224132 62144 224184 62150
rect 224132 62086 224184 62092
rect 217324 59424 217376 59430
rect 217324 59366 217376 59372
rect 216956 59356 217008 59362
rect 216956 59298 217008 59304
rect 216864 56704 216916 56710
rect 216864 56646 216916 56652
rect 216772 56568 216824 56574
rect 216772 56510 216824 56516
rect 216680 52420 216732 52426
rect 216680 52362 216732 52368
rect 216876 52358 216904 56646
rect 217336 55214 217364 59366
rect 217692 58064 217744 58070
rect 217692 58006 217744 58012
rect 217324 55208 217376 55214
rect 217324 55150 217376 55156
rect 217704 53718 217732 58006
rect 217784 57996 217836 58002
rect 217784 57938 217836 57944
rect 217796 53786 217824 57938
rect 224144 56506 224172 62086
rect 224236 62014 224264 67662
rect 224316 63572 224368 63578
rect 224316 63514 224368 63520
rect 224224 62008 224276 62014
rect 224224 61950 224276 61956
rect 224328 57866 224356 63514
rect 224420 63442 224448 69090
rect 224592 69080 224644 69086
rect 224592 69022 224644 69028
rect 224500 64932 224552 64938
rect 224500 64874 224552 64880
rect 224408 63436 224460 63442
rect 224408 63378 224460 63384
rect 224408 60784 224460 60790
rect 224408 60726 224460 60732
rect 224316 57860 224368 57866
rect 224316 57802 224368 57808
rect 224132 56500 224184 56506
rect 224132 56442 224184 56448
rect 224420 55214 224448 60726
rect 224512 59294 224540 64874
rect 224604 63510 224632 69022
rect 224776 67652 224828 67658
rect 224776 67594 224828 67600
rect 224684 66292 224736 66298
rect 224684 66234 224736 66240
rect 224592 63504 224644 63510
rect 224592 63446 224644 63452
rect 224696 60654 224724 66234
rect 224788 62082 224816 67594
rect 224880 64530 224908 70382
rect 227444 70372 227496 70378
rect 227444 70314 227496 70320
rect 226524 70304 226576 70310
rect 226524 70246 226576 70252
rect 226536 69465 226564 70246
rect 227456 70009 227484 70314
rect 232332 70258 232360 79902
rect 232240 70230 232360 70258
rect 227442 70000 227498 70009
rect 227442 69935 227498 69944
rect 226522 69456 226578 69465
rect 226522 69391 226578 69400
rect 227444 69012 227496 69018
rect 227444 68954 227496 68960
rect 227456 68785 227484 68954
rect 227536 68944 227588 68950
rect 227536 68886 227588 68892
rect 227442 68776 227498 68785
rect 227442 68711 227498 68720
rect 227548 68105 227576 68886
rect 227534 68096 227590 68105
rect 227534 68031 227590 68040
rect 227444 67584 227496 67590
rect 227444 67526 227496 67532
rect 227456 67425 227484 67526
rect 227536 67516 227588 67522
rect 227536 67458 227588 67464
rect 227442 67416 227498 67425
rect 227442 67351 227498 67360
rect 227548 66881 227576 67458
rect 227534 66872 227590 66881
rect 227534 66807 227590 66816
rect 227444 66224 227496 66230
rect 227442 66192 227444 66201
rect 227496 66192 227498 66201
rect 227442 66127 227498 66136
rect 227536 66156 227588 66162
rect 227536 66098 227588 66104
rect 227548 65521 227576 66098
rect 227534 65512 227590 65521
rect 227534 65447 227590 65456
rect 227258 64832 227314 64841
rect 227258 64767 227314 64776
rect 227272 64734 227300 64767
rect 227260 64728 227312 64734
rect 227260 64670 227312 64676
rect 224868 64524 224920 64530
rect 224868 64466 224920 64472
rect 227444 64524 227496 64530
rect 227444 64466 227496 64472
rect 227456 64161 227484 64466
rect 227536 64252 227588 64258
rect 227536 64194 227588 64200
rect 227442 64152 227498 64161
rect 227442 64087 227498 64096
rect 227548 63617 227576 64194
rect 227534 63608 227590 63617
rect 227534 63543 227590 63552
rect 227076 63504 227128 63510
rect 227076 63446 227128 63452
rect 227088 62257 227116 63446
rect 227444 63436 227496 63442
rect 227444 63378 227496 63384
rect 227456 62937 227484 63378
rect 227442 62928 227498 62937
rect 227442 62863 227498 62872
rect 227074 62248 227130 62257
rect 227074 62183 227130 62192
rect 224776 62076 224828 62082
rect 224776 62018 224828 62024
rect 226708 62076 226760 62082
rect 226708 62018 226760 62024
rect 226720 61033 226748 62018
rect 227444 62008 227496 62014
rect 227444 61950 227496 61956
rect 227456 61577 227484 61950
rect 227442 61568 227498 61577
rect 227442 61503 227498 61512
rect 226706 61024 226762 61033
rect 226706 60959 226762 60968
rect 227536 60716 227588 60722
rect 227536 60658 227588 60664
rect 224684 60648 224736 60654
rect 224684 60590 224736 60596
rect 227444 60648 227496 60654
rect 227444 60590 227496 60596
rect 227456 60353 227484 60590
rect 227442 60344 227498 60353
rect 227442 60279 227498 60288
rect 227548 59673 227576 60658
rect 232240 60602 232268 70230
rect 232240 60574 232360 60602
rect 227534 59664 227590 59673
rect 227534 59599 227590 59608
rect 227536 59356 227588 59362
rect 227536 59298 227588 59304
rect 224500 59288 224552 59294
rect 224500 59230 224552 59236
rect 227444 59288 227496 59294
rect 227444 59230 227496 59236
rect 227456 58993 227484 59230
rect 227442 58984 227498 58993
rect 227442 58919 227498 58928
rect 227548 58313 227576 59298
rect 227534 58304 227590 58313
rect 227534 58239 227590 58248
rect 227444 57928 227496 57934
rect 232332 57882 232360 60574
rect 227444 57870 227496 57876
rect 227260 57860 227312 57866
rect 227260 57802 227312 57808
rect 227272 57769 227300 57802
rect 227258 57760 227314 57769
rect 227258 57695 227314 57704
rect 227456 57089 227484 57870
rect 232240 57854 232360 57882
rect 227442 57080 227498 57089
rect 227442 57015 227498 57024
rect 227444 56568 227496 56574
rect 227444 56510 227496 56516
rect 227260 56500 227312 56506
rect 227260 56442 227312 56448
rect 227272 56409 227300 56442
rect 227258 56400 227314 56409
rect 227258 56335 227314 56344
rect 227456 55729 227484 56510
rect 227442 55720 227498 55729
rect 227442 55655 227498 55664
rect 227536 55276 227588 55282
rect 227536 55218 227588 55224
rect 224408 55208 224460 55214
rect 227444 55208 227496 55214
rect 224408 55150 224460 55156
rect 227442 55176 227444 55185
rect 227496 55176 227498 55185
rect 227442 55111 227498 55120
rect 226524 55072 226576 55078
rect 226524 55014 226576 55020
rect 226536 54505 226564 55014
rect 226522 54496 226578 54505
rect 226522 54431 226578 54440
rect 226524 53916 226576 53922
rect 226524 53858 226576 53864
rect 217784 53780 217836 53786
rect 217784 53722 217836 53728
rect 217692 53712 217744 53718
rect 217692 53654 217744 53660
rect 216864 52352 216916 52358
rect 216864 52294 216916 52300
rect 226340 51128 226392 51134
rect 226340 51070 226392 51076
rect 226352 47977 226380 51070
rect 226536 50561 226564 53858
rect 226984 53848 227036 53854
rect 226984 53790 227036 53796
rect 227258 53816 227314 53825
rect 226800 52556 226852 52562
rect 226800 52498 226852 52504
rect 226708 52488 226760 52494
rect 226708 52430 226760 52436
rect 226616 51196 226668 51202
rect 226616 51138 226668 51144
rect 226522 50552 226578 50561
rect 226522 50487 226578 50496
rect 226338 47968 226394 47977
rect 226338 47903 226394 47912
rect 226628 47297 226656 51138
rect 226720 49337 226748 52430
rect 226706 49328 226762 49337
rect 226706 49263 226762 49272
rect 226812 48657 226840 52498
rect 226996 49881 227024 53790
rect 227258 53751 227314 53760
rect 227444 53780 227496 53786
rect 227272 53718 227300 53751
rect 227444 53722 227496 53728
rect 227260 53712 227312 53718
rect 227260 53654 227312 53660
rect 227456 53145 227484 53722
rect 227442 53136 227498 53145
rect 227442 53071 227498 53080
rect 227258 52456 227314 52465
rect 227258 52391 227314 52400
rect 227444 52420 227496 52426
rect 227272 52358 227300 52391
rect 227444 52362 227496 52368
rect 227260 52352 227312 52358
rect 227260 52294 227312 52300
rect 227456 51921 227484 52362
rect 227442 51912 227498 51921
rect 227442 51847 227498 51856
rect 227548 51241 227576 55218
rect 227534 51232 227590 51241
rect 227534 51167 227590 51176
rect 232240 51082 232268 57854
rect 232240 51054 232360 51082
rect 226982 49872 227038 49881
rect 226982 49807 227038 49816
rect 227352 49836 227404 49842
rect 227352 49778 227404 49784
rect 227076 49768 227128 49774
rect 227076 49710 227128 49716
rect 226798 48648 226854 48657
rect 226798 48583 226854 48592
rect 226614 47288 226670 47297
rect 226614 47223 226670 47232
rect 227088 46073 227116 49710
rect 227364 46617 227392 49778
rect 232332 48362 232360 51054
rect 227536 48340 227588 48346
rect 227536 48282 227588 48288
rect 232240 48334 232360 48362
rect 227444 47048 227496 47054
rect 227444 46990 227496 46996
rect 227350 46608 227406 46617
rect 227350 46543 227406 46552
rect 227074 46064 227130 46073
rect 227074 45999 227130 46008
rect 226708 45688 226760 45694
rect 226708 45630 226760 45636
rect 226432 42832 226484 42838
rect 226720 42809 226748 45630
rect 227076 45620 227128 45626
rect 227076 45562 227128 45568
rect 227088 43489 227116 45562
rect 227456 44713 227484 46990
rect 227548 45393 227576 48282
rect 227628 46980 227680 46986
rect 227628 46922 227680 46928
rect 227534 45384 227590 45393
rect 227534 45319 227590 45328
rect 227442 44704 227498 44713
rect 227442 44639 227498 44648
rect 227352 44260 227404 44266
rect 227352 44202 227404 44208
rect 227074 43480 227130 43489
rect 227074 43415 227130 43424
rect 226432 42774 226484 42780
rect 226706 42800 226762 42809
rect 226340 41472 226392 41478
rect 226340 41414 226392 41420
rect 226352 40225 226380 41414
rect 226444 40769 226472 42774
rect 226706 42735 226762 42744
rect 226616 41540 226668 41546
rect 226616 41482 226668 41488
rect 226430 40760 226486 40769
rect 226430 40695 226486 40704
rect 226338 40216 226394 40225
rect 226338 40151 226394 40160
rect 226628 39545 226656 41482
rect 227364 41449 227392 44202
rect 227444 44192 227496 44198
rect 227444 44134 227496 44140
rect 227456 42129 227484 44134
rect 227640 44033 227668 46922
rect 227626 44024 227682 44033
rect 227626 43959 227682 43968
rect 227442 42120 227498 42129
rect 227442 42055 227498 42064
rect 227350 41440 227406 41449
rect 227350 41375 227406 41384
rect 232240 41290 232268 48334
rect 232240 41262 232360 41290
rect 226892 40180 226944 40186
rect 226892 40122 226944 40128
rect 226614 39536 226670 39545
rect 226614 39471 226670 39480
rect 226904 38185 226932 40122
rect 227076 40112 227128 40118
rect 227076 40054 227128 40060
rect 227088 38865 227116 40054
rect 227074 38856 227130 38865
rect 227074 38791 227130 38800
rect 227444 38752 227496 38758
rect 227444 38694 227496 38700
rect 226890 38176 226946 38185
rect 226890 38111 226946 38120
rect 227456 37641 227484 38694
rect 227536 38684 227588 38690
rect 227536 38626 227588 38632
rect 227442 37632 227498 37641
rect 227442 37567 227498 37576
rect 227444 37324 227496 37330
rect 227444 37266 227496 37272
rect 227456 36281 227484 37266
rect 227548 36961 227576 38626
rect 232332 38570 232360 41262
rect 231964 38542 232360 38570
rect 227534 36952 227590 36961
rect 227534 36887 227590 36896
rect 227442 36272 227498 36281
rect 227442 36207 227498 36216
rect 227536 36032 227588 36038
rect 227536 35974 227588 35980
rect 227444 35964 227496 35970
rect 227444 35906 227496 35912
rect 227456 35601 227484 35906
rect 227442 35592 227498 35601
rect 227442 35527 227498 35536
rect 227548 34921 227576 35974
rect 227534 34912 227590 34921
rect 227534 34847 227590 34856
rect 227352 34604 227404 34610
rect 227352 34546 227404 34552
rect 227364 33697 227392 34546
rect 227444 34536 227496 34542
rect 227444 34478 227496 34484
rect 227456 34377 227484 34478
rect 227442 34368 227498 34377
rect 227442 34303 227498 34312
rect 227350 33688 227406 33697
rect 227350 33623 227406 33632
rect 227536 33244 227588 33250
rect 227536 33186 227588 33192
rect 227444 33176 227496 33182
rect 227444 33118 227496 33124
rect 227456 33017 227484 33118
rect 227442 33008 227498 33017
rect 227442 32943 227498 32952
rect 213920 32564 213972 32570
rect 213920 32506 213972 32512
rect 215944 32564 215996 32570
rect 215944 32506 215996 32512
rect 95148 32428 95200 32434
rect 95148 32370 95200 32376
rect 116400 32428 116452 32434
rect 116400 32370 116452 32376
rect 95160 31929 95188 32370
rect 116398 32056 116454 32065
rect 116398 31991 116454 32000
rect 95146 31920 95202 31929
rect 95146 31855 95202 31864
rect 116412 31822 116440 31991
rect 71688 31816 71740 31822
rect 71346 31764 71688 31770
rect 71346 31758 71740 31764
rect 116400 31816 116452 31822
rect 213932 31793 213960 32506
rect 215114 32464 215170 32473
rect 215114 32399 215116 32408
rect 215168 32399 215170 32408
rect 227444 32428 227496 32434
rect 215116 32370 215168 32376
rect 227444 32370 227496 32376
rect 227456 31793 227484 32370
rect 227548 32337 227576 33186
rect 227534 32328 227590 32337
rect 227534 32263 227590 32272
rect 116400 31758 116452 31764
rect 213918 31784 213974 31793
rect 71346 31742 71728 31758
rect 213918 31719 213974 31728
rect 227442 31784 227498 31793
rect 227442 31719 227498 31728
rect 121748 31606 122590 31634
rect 128740 31606 129490 31634
rect 149532 31606 150374 31634
rect 156524 31606 157274 31634
rect 159100 31606 159850 31634
rect 161676 31606 162518 31634
rect 164344 31606 165094 31634
rect 172992 31606 173742 31634
rect 175568 31606 176410 31634
rect 178236 31606 178986 31634
rect 179892 31606 180734 31634
rect 192128 31606 192878 31634
rect 208780 31606 209346 31634
rect 29932 30326 29960 31484
rect 120000 30326 120028 31484
rect 120092 31470 120842 31498
rect 29920 30320 29972 30326
rect 32312 30320 32364 30326
rect 29920 30262 29972 30268
rect 32310 30288 32312 30297
rect 119988 30320 120040 30326
rect 32364 30288 32366 30297
rect 119988 30262 120040 30268
rect 32310 30223 32366 30232
rect 115848 30252 115900 30258
rect 115848 30194 115900 30200
rect 107568 30184 107620 30190
rect 107568 30126 107620 30132
rect 51724 30116 51776 30122
rect 51724 30058 51776 30064
rect 32404 29980 32456 29986
rect 32404 29922 32456 29928
rect 28264 29912 28316 29918
rect 28264 29854 28316 29860
rect 24124 29844 24176 29850
rect 24124 29786 24176 29792
rect 22744 29708 22796 29714
rect 22744 29650 22796 29656
rect 11704 26920 11756 26926
rect 11704 26862 11756 26868
rect 10968 19984 11020 19990
rect 10968 19926 11020 19932
rect 10980 3534 11008 19926
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 10508 3460 10560 3466
rect 10508 3402 10560 3408
rect 11256 480 11284 3470
rect 11716 3262 11744 26862
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 13636 7608 13688 7614
rect 13636 7550 13688 7556
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 11704 3256 11756 3262
rect 11704 3198 11756 3204
rect 12452 480 12480 4762
rect 13648 480 13676 7550
rect 17132 3936 17184 3942
rect 17132 3878 17184 3884
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 14844 480 14872 3402
rect 16040 480 16068 3538
rect 17144 3534 17172 3878
rect 17880 3534 17908 17206
rect 22008 13116 22060 13122
rect 22008 13058 22060 13064
rect 18328 7676 18380 7682
rect 18328 7618 18380 7624
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17236 480 17264 3470
rect 18340 480 18368 7618
rect 20720 3392 20772 3398
rect 20720 3334 20772 3340
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 19536 480 19564 3130
rect 20732 480 20760 3334
rect 22020 626 22048 13058
rect 22756 3194 22784 29650
rect 23112 8968 23164 8974
rect 23112 8910 23164 8916
rect 22744 3188 22796 3194
rect 22744 3130 22796 3136
rect 21928 598 22048 626
rect 21928 480 21956 598
rect 23124 480 23152 8910
rect 24136 3942 24164 29786
rect 25504 29640 25556 29646
rect 25504 29582 25556 29588
rect 24124 3936 24176 3942
rect 24124 3878 24176 3884
rect 25516 3670 25544 29582
rect 27528 11824 27580 11830
rect 27528 11766 27580 11772
rect 24308 3664 24360 3670
rect 24308 3606 24360 3612
rect 25504 3664 25556 3670
rect 25504 3606 25556 3612
rect 25596 3664 25648 3670
rect 25596 3606 25648 3612
rect 24320 480 24348 3606
rect 25504 3528 25556 3534
rect 25504 3470 25556 3476
rect 25516 480 25544 3470
rect 25608 3398 25636 3606
rect 25596 3392 25648 3398
rect 25596 3334 25648 3340
rect 27540 3058 27568 11766
rect 28276 3602 28304 29854
rect 31024 29776 31076 29782
rect 31024 29718 31076 29724
rect 30288 18624 30340 18630
rect 30288 18566 30340 18572
rect 28908 14476 28960 14482
rect 28908 14418 28960 14424
rect 28264 3596 28316 3602
rect 28264 3538 28316 3544
rect 28920 3194 28948 14418
rect 29092 3596 29144 3602
rect 29092 3538 29144 3544
rect 27896 3188 27948 3194
rect 27896 3130 27948 3136
rect 28908 3188 28960 3194
rect 28908 3130 28960 3136
rect 26700 3052 26752 3058
rect 26700 2994 26752 3000
rect 27528 3052 27580 3058
rect 27528 2994 27580 3000
rect 26712 480 26740 2994
rect 27908 480 27936 3130
rect 29104 480 29132 3538
rect 30300 480 30328 18566
rect 31036 3602 31064 29718
rect 31668 10396 31720 10402
rect 31668 10338 31720 10344
rect 31024 3596 31076 3602
rect 31024 3538 31076 3544
rect 31680 3482 31708 10338
rect 32416 3670 32444 29922
rect 50988 28348 51040 28354
rect 50988 28290 51040 28296
rect 48228 20052 48280 20058
rect 48228 19994 48280 20000
rect 38568 17332 38620 17338
rect 38568 17274 38620 17280
rect 34428 15904 34480 15910
rect 34428 15846 34480 15852
rect 32680 3936 32732 3942
rect 32680 3878 32732 3884
rect 32404 3664 32456 3670
rect 32404 3606 32456 3612
rect 31496 3454 31708 3482
rect 31496 480 31524 3454
rect 32692 480 32720 3878
rect 34440 3602 34468 15846
rect 34980 7744 35032 7750
rect 34980 7686 35032 7692
rect 33876 3596 33928 3602
rect 33876 3538 33928 3544
rect 34428 3596 34480 3602
rect 34428 3538 34480 3544
rect 33888 480 33916 3538
rect 34992 480 35020 7686
rect 37372 6316 37424 6322
rect 37372 6258 37424 6264
rect 36176 3664 36228 3670
rect 36176 3606 36228 3612
rect 36188 480 36216 3606
rect 37384 480 37412 6258
rect 38580 480 38608 17274
rect 42708 13184 42760 13190
rect 42708 13126 42760 13132
rect 40960 6384 41012 6390
rect 40960 6326 41012 6332
rect 39764 4004 39816 4010
rect 39764 3946 39816 3952
rect 39776 480 39804 3946
rect 40972 480 41000 6326
rect 42720 3602 42748 13126
rect 46848 11892 46900 11898
rect 46848 11834 46900 11840
rect 44548 6452 44600 6458
rect 44548 6394 44600 6400
rect 43352 3664 43404 3670
rect 43352 3606 43404 3612
rect 42156 3596 42208 3602
rect 42156 3538 42208 3544
rect 42708 3596 42760 3602
rect 42708 3538 42760 3544
rect 42168 480 42196 3538
rect 43364 480 43392 3606
rect 44560 480 44588 6394
rect 46860 3398 46888 11834
rect 46940 3732 46992 3738
rect 46940 3674 46992 3680
rect 45744 3392 45796 3398
rect 45744 3334 45796 3340
rect 46848 3392 46900 3398
rect 46848 3334 46900 3340
rect 45756 480 45784 3334
rect 46952 480 46980 3674
rect 48240 3482 48268 19994
rect 49332 6520 49384 6526
rect 49332 6462 49384 6468
rect 48148 3454 48268 3482
rect 48148 480 48176 3454
rect 49344 480 49372 6462
rect 51000 3398 51028 28290
rect 51736 3942 51764 30058
rect 57244 30048 57296 30054
rect 57244 29990 57296 29996
rect 56508 22772 56560 22778
rect 56508 22714 56560 22720
rect 52368 21412 52420 21418
rect 52368 21354 52420 21360
rect 51724 3936 51776 3942
rect 51724 3878 51776 3884
rect 52380 3398 52408 21354
rect 55128 15972 55180 15978
rect 55128 15914 55180 15920
rect 52828 6656 52880 6662
rect 52828 6598 52880 6604
rect 50528 3392 50580 3398
rect 50528 3334 50580 3340
rect 50988 3392 51040 3398
rect 50988 3334 51040 3340
rect 51632 3392 51684 3398
rect 51632 3334 51684 3340
rect 52368 3392 52420 3398
rect 52368 3334 52420 3340
rect 50540 480 50568 3334
rect 51644 480 51672 3334
rect 52840 480 52868 6598
rect 55140 3398 55168 15914
rect 56416 6588 56468 6594
rect 56416 6530 56468 6536
rect 54024 3392 54076 3398
rect 54024 3334 54076 3340
rect 55128 3392 55180 3398
rect 55128 3334 55180 3340
rect 55220 3392 55272 3398
rect 55220 3334 55272 3340
rect 54036 480 54064 3334
rect 55232 480 55260 3334
rect 56428 480 56456 6530
rect 56520 3398 56548 22714
rect 57256 4010 57284 29990
rect 61384 29504 61436 29510
rect 61384 29446 61436 29452
rect 59268 25560 59320 25566
rect 59268 25502 59320 25508
rect 57888 24132 57940 24138
rect 57888 24074 57940 24080
rect 57244 4004 57296 4010
rect 57244 3946 57296 3952
rect 56508 3392 56560 3398
rect 57900 3346 57928 24074
rect 59280 3398 59308 25502
rect 60004 6724 60056 6730
rect 60004 6666 60056 6672
rect 56508 3334 56560 3340
rect 57624 3318 57928 3346
rect 58808 3392 58860 3398
rect 58808 3334 58860 3340
rect 59268 3392 59320 3398
rect 59268 3334 59320 3340
rect 57624 480 57652 3318
rect 58820 480 58848 3334
rect 60016 480 60044 6666
rect 61396 3874 61424 29446
rect 69664 29436 69716 29442
rect 69664 29378 69716 29384
rect 62028 26988 62080 26994
rect 62028 26930 62080 26936
rect 61384 3868 61436 3874
rect 61384 3810 61436 3816
rect 62040 3398 62068 26930
rect 68928 25628 68980 25634
rect 68928 25570 68980 25576
rect 63408 24200 63460 24206
rect 63408 24142 63460 24148
rect 63420 3398 63448 24142
rect 64788 22840 64840 22846
rect 64788 22782 64840 22788
rect 63592 6792 63644 6798
rect 63592 6734 63644 6740
rect 61200 3392 61252 3398
rect 61200 3334 61252 3340
rect 62028 3392 62080 3398
rect 62028 3334 62080 3340
rect 62396 3392 62448 3398
rect 62396 3334 62448 3340
rect 63408 3392 63460 3398
rect 63408 3334 63460 3340
rect 61212 480 61240 3334
rect 62408 480 62436 3334
rect 63604 480 63632 6734
rect 64800 480 64828 22782
rect 66168 14680 66220 14686
rect 66168 14622 66220 14628
rect 66180 3482 66208 14622
rect 67180 6860 67232 6866
rect 67180 6802 67232 6808
rect 65996 3454 66208 3482
rect 65996 480 66024 3454
rect 67192 480 67220 6802
rect 68940 3398 68968 25570
rect 69480 9172 69532 9178
rect 69480 9114 69532 9120
rect 68284 3392 68336 3398
rect 68284 3334 68336 3340
rect 68928 3392 68980 3398
rect 68928 3334 68980 3340
rect 68296 480 68324 3334
rect 69492 480 69520 9114
rect 69676 3806 69704 29378
rect 107476 27056 107528 27062
rect 107476 26998 107528 27004
rect 85488 25696 85540 25702
rect 85488 25638 85540 25644
rect 82728 21548 82780 21554
rect 82728 21490 82780 21496
rect 72976 21480 73028 21486
rect 72976 21422 73028 21428
rect 70676 6112 70728 6118
rect 70676 6054 70728 6060
rect 69664 3800 69716 3806
rect 69664 3742 69716 3748
rect 70688 480 70716 6054
rect 72988 3398 73016 21422
rect 75828 20120 75880 20126
rect 75828 20062 75880 20068
rect 74264 6044 74316 6050
rect 74264 5986 74316 5992
rect 73068 4888 73120 4894
rect 73068 4830 73120 4836
rect 71872 3392 71924 3398
rect 71872 3334 71924 3340
rect 72976 3392 73028 3398
rect 72976 3334 73028 3340
rect 71884 480 71912 3334
rect 73080 480 73108 4830
rect 74276 480 74304 5986
rect 75840 3482 75868 20062
rect 79968 18692 80020 18698
rect 79968 18634 80020 18640
rect 77852 5976 77904 5982
rect 77852 5918 77904 5924
rect 76656 4956 76708 4962
rect 76656 4898 76708 4904
rect 75472 3454 75868 3482
rect 75472 480 75500 3454
rect 76668 480 76696 4898
rect 77864 480 77892 5918
rect 79980 3398 80008 18634
rect 80244 5024 80296 5030
rect 80244 4966 80296 4972
rect 79048 3392 79100 3398
rect 79048 3334 79100 3340
rect 79968 3392 80020 3398
rect 79968 3334 80020 3340
rect 79060 480 79088 3334
rect 80256 480 80284 4966
rect 82740 4146 82768 21490
rect 83832 5092 83884 5098
rect 83832 5034 83884 5040
rect 81440 4140 81492 4146
rect 81440 4082 81492 4088
rect 82728 4140 82780 4146
rect 82728 4082 82780 4088
rect 81452 480 81480 4082
rect 82636 3868 82688 3874
rect 82636 3810 82688 3816
rect 82648 480 82676 3810
rect 83844 480 83872 5034
rect 85500 4146 85528 25638
rect 96528 24268 96580 24274
rect 96528 24210 96580 24216
rect 89628 22908 89680 22914
rect 89628 22850 89680 22856
rect 86132 10464 86184 10470
rect 86132 10406 86184 10412
rect 84936 4140 84988 4146
rect 84936 4082 84988 4088
rect 85488 4140 85540 4146
rect 85488 4082 85540 4088
rect 84948 480 84976 4082
rect 86144 480 86172 10406
rect 87328 5228 87380 5234
rect 87328 5170 87380 5176
rect 87340 480 87368 5170
rect 89640 4146 89668 22850
rect 93768 14748 93820 14754
rect 93768 14690 93820 14696
rect 92112 7812 92164 7818
rect 92112 7754 92164 7760
rect 90916 5160 90968 5166
rect 90916 5102 90968 5108
rect 88524 4140 88576 4146
rect 88524 4082 88576 4088
rect 89628 4140 89680 4146
rect 89628 4082 89680 4088
rect 88536 480 88564 4082
rect 89812 3868 89864 3874
rect 89812 3810 89864 3816
rect 89824 3346 89852 3810
rect 89732 3318 89852 3346
rect 89732 480 89760 3318
rect 90928 480 90956 5102
rect 92124 480 92152 7754
rect 93780 4146 93808 14690
rect 94504 5296 94556 5302
rect 94504 5238 94556 5244
rect 93308 4140 93360 4146
rect 93308 4082 93360 4088
rect 93768 4140 93820 4146
rect 93768 4082 93820 4088
rect 93320 480 93348 4082
rect 94516 480 94544 5238
rect 96540 4146 96568 24210
rect 100668 21616 100720 21622
rect 100668 21558 100720 21564
rect 99288 7880 99340 7886
rect 99288 7822 99340 7828
rect 98092 5364 98144 5370
rect 98092 5306 98144 5312
rect 95700 4140 95752 4146
rect 95700 4082 95752 4088
rect 96528 4140 96580 4146
rect 96528 4082 96580 4088
rect 95712 480 95740 4082
rect 96896 3936 96948 3942
rect 96896 3878 96948 3884
rect 96908 480 96936 3878
rect 98104 480 98132 5306
rect 99300 480 99328 7822
rect 100680 4842 100708 21558
rect 102784 7948 102836 7954
rect 102784 7890 102836 7896
rect 101588 5432 101640 5438
rect 101588 5374 101640 5380
rect 100496 4814 100708 4842
rect 100496 480 100524 4814
rect 101600 480 101628 5374
rect 102796 480 102824 7890
rect 105176 4752 105228 4758
rect 105176 4694 105228 4700
rect 103520 4140 103572 4146
rect 103520 4082 103572 4088
rect 103532 3806 103560 4082
rect 103980 4004 104032 4010
rect 103980 3946 104032 3952
rect 103520 3800 103572 3806
rect 103520 3742 103572 3748
rect 103992 480 104020 3946
rect 105188 480 105216 4694
rect 107488 3398 107516 26998
rect 106372 3392 106424 3398
rect 106372 3334 106424 3340
rect 107476 3392 107528 3398
rect 107476 3334 107528 3340
rect 106384 480 106412 3334
rect 107580 480 107608 30126
rect 113088 28416 113140 28422
rect 113088 28358 113140 28364
rect 109960 8016 110012 8022
rect 109960 7958 110012 7964
rect 108764 5500 108816 5506
rect 108764 5442 108816 5448
rect 108776 480 108804 5442
rect 109972 480 110000 7958
rect 112996 4140 113048 4146
rect 112996 4082 113048 4088
rect 111156 4072 111208 4078
rect 111156 4014 111208 4020
rect 111168 480 111196 4014
rect 113008 3806 113036 4082
rect 112996 3800 113048 3806
rect 112996 3742 113048 3748
rect 113100 3398 113128 28358
rect 113548 8152 113600 8158
rect 113548 8094 113600 8100
rect 113180 3800 113232 3806
rect 113180 3742 113232 3748
rect 112352 3392 112404 3398
rect 112352 3334 112404 3340
rect 113088 3392 113140 3398
rect 113088 3334 113140 3340
rect 112364 480 112392 3334
rect 113192 3330 113220 3742
rect 113180 3324 113232 3330
rect 113180 3266 113232 3272
rect 113560 480 113588 8094
rect 115860 3398 115888 30194
rect 118608 29572 118660 29578
rect 118608 29514 118660 29520
rect 117228 27124 117280 27130
rect 117228 27066 117280 27072
rect 117136 8084 117188 8090
rect 117136 8026 117188 8032
rect 114744 3392 114796 3398
rect 114744 3334 114796 3340
rect 115848 3392 115900 3398
rect 115848 3334 115900 3340
rect 114756 480 114784 3334
rect 115940 2916 115992 2922
rect 115940 2858 115992 2864
rect 115952 480 115980 2858
rect 117148 480 117176 8026
rect 117240 2922 117268 27066
rect 118620 3482 118648 29514
rect 119988 20188 120040 20194
rect 119988 20130 120040 20136
rect 118252 3454 118648 3482
rect 117228 2916 117280 2922
rect 117228 2858 117280 2864
rect 118252 480 118280 3454
rect 120000 3398 120028 20130
rect 120092 10334 120120 31470
rect 121656 28286 121684 31484
rect 121644 28280 121696 28286
rect 121644 28222 121696 28228
rect 121748 26738 121776 31606
rect 123404 29510 123432 31484
rect 123392 29504 123444 29510
rect 123392 29446 123444 29452
rect 123484 29504 123536 29510
rect 123484 29446 123536 29452
rect 121564 26710 121776 26738
rect 121564 21978 121592 26710
rect 121564 21950 121684 21978
rect 120080 10328 120132 10334
rect 120080 10270 120132 10276
rect 121656 6186 121684 21950
rect 121644 6180 121696 6186
rect 121644 6122 121696 6128
rect 120632 4684 120684 4690
rect 120632 4626 120684 4632
rect 119436 3392 119488 3398
rect 119436 3334 119488 3340
rect 119988 3392 120040 3398
rect 119988 3334 120040 3340
rect 119448 480 119476 3334
rect 120644 480 120672 4626
rect 123024 4616 123076 4622
rect 123024 4558 123076 4564
rect 121828 4140 121880 4146
rect 121828 4082 121880 4088
rect 121840 480 121868 4082
rect 122748 3800 122800 3806
rect 122748 3742 122800 3748
rect 122760 3330 122788 3742
rect 122748 3324 122800 3330
rect 122748 3266 122800 3272
rect 123036 480 123064 4558
rect 123496 4146 123524 29446
rect 124324 29442 124352 31484
rect 124312 29436 124364 29442
rect 124312 29378 124364 29384
rect 125152 26926 125180 31484
rect 125612 31470 126086 31498
rect 126624 31470 126914 31498
rect 125508 28280 125560 28286
rect 125508 28222 125560 28228
rect 125140 26920 125192 26926
rect 125140 26862 125192 26868
rect 123484 4140 123536 4146
rect 123484 4082 123536 4088
rect 125520 3466 125548 28222
rect 125612 6254 125640 31470
rect 126244 29436 126296 29442
rect 126244 29378 126296 29384
rect 125876 26784 125928 26790
rect 125876 26726 125928 26732
rect 125888 19990 125916 26726
rect 125876 19984 125928 19990
rect 125876 19926 125928 19932
rect 125600 6248 125652 6254
rect 125600 6190 125652 6196
rect 124220 3460 124272 3466
rect 124220 3402 124272 3408
rect 125508 3460 125560 3466
rect 125508 3402 125560 3408
rect 124232 480 124260 3402
rect 126256 3398 126284 29378
rect 126624 26790 126652 31470
rect 127728 29850 127756 31484
rect 128372 31470 128662 31498
rect 127716 29844 127768 29850
rect 127716 29786 127768 29792
rect 126612 26784 126664 26790
rect 126612 26726 126664 26732
rect 126886 14512 126942 14521
rect 126886 14447 126942 14456
rect 125416 3392 125468 3398
rect 125416 3334 125468 3340
rect 126244 3392 126296 3398
rect 126900 3346 126928 14447
rect 127806 7576 127862 7585
rect 127806 7511 127862 7520
rect 126244 3334 126296 3340
rect 125428 480 125456 3334
rect 126624 3318 126928 3346
rect 126624 480 126652 3318
rect 127820 480 127848 7511
rect 128372 4826 128400 31470
rect 128740 28914 128768 31606
rect 128556 28886 128768 28914
rect 129844 31470 130410 31498
rect 128556 7614 128584 28886
rect 129648 18012 129700 18018
rect 129648 17954 129700 17960
rect 128544 7608 128596 7614
rect 128544 7550 128596 7556
rect 128360 4820 128412 4826
rect 128360 4762 128412 4768
rect 129660 3466 129688 17954
rect 129004 3460 129056 3466
rect 129004 3402 129056 3408
rect 129648 3460 129700 3466
rect 129648 3402 129700 3408
rect 129016 480 129044 3402
rect 129844 3330 129872 31470
rect 131224 29918 131252 31484
rect 131316 31470 132158 31498
rect 132604 31470 132986 31498
rect 131212 29912 131264 29918
rect 131212 29854 131264 29860
rect 131316 17270 131344 31470
rect 131304 17264 131356 17270
rect 131304 17206 131356 17212
rect 132408 16652 132460 16658
rect 132408 16594 132460 16600
rect 131026 15328 131082 15337
rect 131026 15263 131082 15272
rect 131040 3466 131068 15263
rect 132420 3466 132448 16594
rect 132604 7682 132632 31470
rect 133800 29714 133828 31484
rect 134720 29986 134748 31484
rect 135364 31470 135562 31498
rect 136192 31470 136482 31498
rect 134708 29980 134760 29986
rect 134708 29922 134760 29928
rect 133788 29708 133840 29714
rect 133788 29650 133840 29656
rect 135260 28892 135312 28898
rect 135260 28834 135312 28840
rect 133788 11756 133840 11762
rect 133788 11698 133840 11704
rect 132592 7676 132644 7682
rect 132592 7618 132644 7624
rect 132500 3800 132552 3806
rect 132500 3742 132552 3748
rect 130200 3460 130252 3466
rect 130200 3402 130252 3408
rect 131028 3460 131080 3466
rect 131028 3402 131080 3408
rect 131396 3460 131448 3466
rect 131396 3402 131448 3408
rect 132408 3460 132460 3466
rect 132408 3402 132460 3408
rect 129832 3324 129884 3330
rect 129832 3266 129884 3272
rect 130212 480 130240 3402
rect 131408 480 131436 3402
rect 132512 3330 132540 3742
rect 133800 3534 133828 11698
rect 135168 10328 135220 10334
rect 135168 10270 135220 10276
rect 132592 3528 132644 3534
rect 132592 3470 132644 3476
rect 133788 3528 133840 3534
rect 135180 3482 135208 10270
rect 135272 8974 135300 28834
rect 135364 13122 135392 31470
rect 136192 28898 136220 31470
rect 137296 29646 137324 31484
rect 137284 29640 137336 29646
rect 137284 29582 137336 29588
rect 136180 28892 136232 28898
rect 136180 28834 136232 28840
rect 138112 28892 138164 28898
rect 138112 28834 138164 28840
rect 135352 13116 135404 13122
rect 135352 13058 135404 13064
rect 136546 13016 136602 13025
rect 136546 12951 136602 12960
rect 135260 8968 135312 8974
rect 135260 8910 135312 8916
rect 136560 3534 136588 12951
rect 138124 11830 138152 28834
rect 138112 11824 138164 11830
rect 138112 11766 138164 11772
rect 137284 4140 137336 4146
rect 137284 4082 137336 4088
rect 133788 3470 133840 3476
rect 132500 3324 132552 3330
rect 132500 3266 132552 3272
rect 132604 480 132632 3470
rect 134904 3454 135208 3482
rect 136088 3528 136140 3534
rect 136088 3470 136140 3476
rect 136548 3528 136600 3534
rect 136548 3470 136600 3476
rect 133788 2100 133840 2106
rect 133788 2042 133840 2048
rect 133800 480 133828 2042
rect 134904 480 134932 3454
rect 136100 480 136128 3470
rect 137296 480 137324 4082
rect 138216 3398 138244 31484
rect 138768 31470 139058 31498
rect 139412 31470 139886 31498
rect 138768 28898 138796 31470
rect 138756 28892 138808 28898
rect 138756 28834 138808 28840
rect 139412 14482 139440 31470
rect 140792 29782 140820 31484
rect 140884 31470 141634 31498
rect 142264 31470 142554 31498
rect 140780 29776 140832 29782
rect 140780 29718 140832 29724
rect 140884 18630 140912 31470
rect 140872 18624 140924 18630
rect 140872 18566 140924 18572
rect 139400 14476 139452 14482
rect 139400 14418 139452 14424
rect 140688 13252 140740 13258
rect 140688 13194 140740 13200
rect 138478 8936 138534 8945
rect 138478 8871 138534 8880
rect 138204 3392 138256 3398
rect 138204 3334 138256 3340
rect 138492 480 138520 8871
rect 140700 3534 140728 13194
rect 142066 11656 142122 11665
rect 142066 11591 142122 11600
rect 139676 3528 139728 3534
rect 139676 3470 139728 3476
rect 140688 3528 140740 3534
rect 140688 3470 140740 3476
rect 139688 480 139716 3470
rect 140872 3392 140924 3398
rect 140872 3334 140924 3340
rect 140884 480 140912 3334
rect 142080 480 142108 11591
rect 142264 10402 142292 31470
rect 143368 30122 143396 31484
rect 143552 31470 144302 31498
rect 145024 31470 145130 31498
rect 143356 30116 143408 30122
rect 143356 30058 143408 30064
rect 142804 29028 142856 29034
rect 142804 28970 142856 28976
rect 142252 10396 142304 10402
rect 142252 10338 142304 10344
rect 142816 3602 142844 28970
rect 143552 15910 143580 31470
rect 143540 15904 143592 15910
rect 143540 15846 143592 15852
rect 143448 14476 143500 14482
rect 143448 14418 143500 14424
rect 142804 3596 142856 3602
rect 142804 3538 142856 3544
rect 143460 3346 143488 14418
rect 145024 7750 145052 31470
rect 146036 29034 146064 31484
rect 146312 31470 146878 31498
rect 147706 31470 147812 31498
rect 146024 29028 146076 29034
rect 146024 28970 146076 28976
rect 145012 7744 145064 7750
rect 145012 7686 145064 7692
rect 145654 7712 145710 7721
rect 145654 7647 145710 7656
rect 143276 3318 143488 3346
rect 143276 480 143304 3318
rect 144460 3256 144512 3262
rect 144460 3198 144512 3204
rect 144472 480 144500 3198
rect 145668 480 145696 7647
rect 146312 6322 146340 31470
rect 147784 17338 147812 31470
rect 148612 30054 148640 31484
rect 149072 31470 149454 31498
rect 148600 30048 148652 30054
rect 148600 29990 148652 29996
rect 148048 19304 148100 19310
rect 148048 19246 148100 19252
rect 147772 17332 147824 17338
rect 147772 17274 147824 17280
rect 147588 14612 147640 14618
rect 147588 14554 147640 14560
rect 146300 6316 146352 6322
rect 146300 6258 146352 6264
rect 145840 3800 145892 3806
rect 145840 3742 145892 3748
rect 145852 3466 145880 3742
rect 145932 3732 145984 3738
rect 145932 3674 145984 3680
rect 145944 3618 145972 3674
rect 145944 3590 146156 3618
rect 146128 3466 146156 3590
rect 145840 3460 145892 3466
rect 145840 3402 145892 3408
rect 146116 3460 146168 3466
rect 146116 3402 146168 3408
rect 147600 3330 147628 14554
rect 148060 11898 148088 19246
rect 148048 11892 148100 11898
rect 148048 11834 148100 11840
rect 149072 6390 149100 31470
rect 149532 26738 149560 31606
rect 149348 26710 149560 26738
rect 150452 31470 151202 31498
rect 151832 31470 152122 31498
rect 152476 31470 152950 31498
rect 153212 31470 153778 31498
rect 149348 13190 149376 26710
rect 149336 13184 149388 13190
rect 149336 13126 149388 13132
rect 150348 13116 150400 13122
rect 150348 13058 150400 13064
rect 149060 6384 149112 6390
rect 149060 6326 149112 6332
rect 150360 3738 150388 13058
rect 149244 3732 149296 3738
rect 149244 3674 149296 3680
rect 150348 3732 150400 3738
rect 150348 3674 150400 3680
rect 148048 3460 148100 3466
rect 148048 3402 148100 3408
rect 146852 3324 146904 3330
rect 146852 3266 146904 3272
rect 147588 3324 147640 3330
rect 147588 3266 147640 3272
rect 146864 480 146892 3266
rect 148060 480 148088 3402
rect 149256 480 149284 3674
rect 150452 3670 150480 31470
rect 151726 14648 151782 14657
rect 151726 14583 151782 14592
rect 151544 9036 151596 9042
rect 151544 8978 151596 8984
rect 150440 3664 150492 3670
rect 150440 3606 150492 3612
rect 150532 3664 150584 3670
rect 150532 3606 150584 3612
rect 150544 3534 150572 3606
rect 150532 3528 150584 3534
rect 150532 3470 150584 3476
rect 150716 3528 150768 3534
rect 150716 3470 150768 3476
rect 150440 3324 150492 3330
rect 150440 3266 150492 3272
rect 150452 480 150480 3266
rect 150728 3262 150756 3470
rect 150716 3256 150768 3262
rect 150716 3198 150768 3204
rect 151556 480 151584 8978
rect 151740 3330 151768 14583
rect 151832 6458 151860 31470
rect 152476 26738 152504 31470
rect 152016 26710 152504 26738
rect 152016 19310 152044 26710
rect 152004 19304 152056 19310
rect 152004 19246 152056 19252
rect 153108 13184 153160 13190
rect 153108 13126 153160 13132
rect 151820 6452 151872 6458
rect 151820 6394 151872 6400
rect 151728 3324 151780 3330
rect 151728 3266 151780 3272
rect 153120 626 153148 13126
rect 153212 3670 153240 31470
rect 154580 26784 154632 26790
rect 154580 26726 154632 26732
rect 154488 14544 154540 14550
rect 154488 14486 154540 14492
rect 154500 3738 154528 14486
rect 154592 6526 154620 26726
rect 154684 20058 154712 31484
rect 155144 31470 155526 31498
rect 155144 26790 155172 31470
rect 156432 28354 156460 31484
rect 156420 28348 156472 28354
rect 156420 28290 156472 28296
rect 155132 26784 155184 26790
rect 156524 26738 156552 31606
rect 155132 26726 155184 26732
rect 156064 26710 156552 26738
rect 157352 31470 158194 31498
rect 158732 31470 159022 31498
rect 156064 21418 156092 26710
rect 156052 21412 156104 21418
rect 156052 21354 156104 21360
rect 154672 20052 154724 20058
rect 154672 19994 154724 20000
rect 156328 8968 156380 8974
rect 156328 8910 156380 8916
rect 154580 6520 154632 6526
rect 154580 6462 154632 6468
rect 153936 3732 153988 3738
rect 153936 3674 153988 3680
rect 154488 3732 154540 3738
rect 154488 3674 154540 3680
rect 153200 3664 153252 3670
rect 153200 3606 153252 3612
rect 152752 598 153148 626
rect 152752 480 152780 598
rect 153948 480 153976 3674
rect 155132 3460 155184 3466
rect 155132 3402 155184 3408
rect 155144 480 155172 3402
rect 156340 480 156368 8910
rect 157352 6662 157380 31470
rect 158732 15978 158760 31470
rect 159100 28914 159128 31606
rect 160112 31470 160770 31498
rect 161492 31470 161598 31498
rect 159364 29844 159416 29850
rect 159364 29786 159416 29792
rect 158824 28886 159128 28914
rect 158824 22778 158852 28886
rect 158812 22772 158864 22778
rect 158812 22714 158864 22720
rect 158720 15972 158772 15978
rect 158720 15914 158772 15920
rect 158626 14784 158682 14793
rect 158626 14719 158682 14728
rect 157340 6656 157392 6662
rect 157340 6598 157392 6604
rect 158640 3194 158668 14719
rect 159376 3806 159404 29786
rect 160008 16720 160060 16726
rect 160008 16662 160060 16668
rect 159916 7608 159968 7614
rect 159916 7550 159968 7556
rect 159364 3800 159416 3806
rect 159364 3742 159416 3748
rect 157524 3188 157576 3194
rect 157524 3130 157576 3136
rect 158628 3188 158680 3194
rect 158628 3130 158680 3136
rect 157536 480 157564 3130
rect 158720 2984 158772 2990
rect 158720 2926 158772 2932
rect 158732 480 158760 2926
rect 159928 480 159956 7550
rect 160020 2990 160048 16662
rect 160112 6594 160140 31470
rect 161492 24138 161520 31470
rect 161676 28914 161704 31606
rect 161584 28886 161704 28914
rect 162872 31470 163346 31498
rect 161584 25566 161612 28886
rect 161572 25560 161624 25566
rect 161572 25502 161624 25508
rect 161480 24132 161532 24138
rect 161480 24074 161532 24080
rect 162872 6730 162900 31470
rect 164252 26994 164280 31484
rect 164240 26988 164292 26994
rect 164240 26930 164292 26936
rect 164344 26874 164372 31606
rect 165632 31470 166014 31498
rect 166276 31470 166842 31498
rect 167012 31470 167670 31498
rect 168392 31470 168590 31498
rect 164884 29912 164936 29918
rect 164884 29854 164936 29860
rect 164252 26846 164372 26874
rect 164252 24206 164280 26846
rect 164240 24200 164292 24206
rect 164240 24142 164292 24148
rect 164148 16788 164200 16794
rect 164148 16730 164200 16736
rect 162860 6724 162912 6730
rect 162860 6666 162912 6672
rect 160100 6588 160152 6594
rect 160100 6530 160152 6536
rect 161112 6316 161164 6322
rect 161112 6258 161164 6264
rect 160008 2984 160060 2990
rect 160008 2926 160060 2932
rect 161124 480 161152 6258
rect 164160 3670 164188 16730
rect 164896 3874 164924 29854
rect 165526 11792 165582 11801
rect 165526 11727 165582 11736
rect 164884 3868 164936 3874
rect 164884 3810 164936 3816
rect 165540 3670 165568 11727
rect 165632 6798 165660 31470
rect 166276 29866 166304 31470
rect 165908 29838 166304 29866
rect 165908 22846 165936 29838
rect 166264 29776 166316 29782
rect 166264 29718 166316 29724
rect 165896 22840 165948 22846
rect 165896 22782 165948 22788
rect 165620 6792 165672 6798
rect 165620 6734 165672 6740
rect 166276 3942 166304 29718
rect 167012 14686 167040 31470
rect 167000 14680 167052 14686
rect 167000 14622 167052 14628
rect 168196 9104 168248 9110
rect 168196 9046 168248 9052
rect 167092 4820 167144 4826
rect 167092 4762 167144 4768
rect 166264 3936 166316 3942
rect 166264 3878 166316 3884
rect 165896 3800 165948 3806
rect 165896 3742 165948 3748
rect 163504 3664 163556 3670
rect 163504 3606 163556 3612
rect 164148 3664 164200 3670
rect 164148 3606 164200 3612
rect 164700 3664 164752 3670
rect 164700 3606 164752 3612
rect 165528 3664 165580 3670
rect 165528 3606 165580 3612
rect 162308 2168 162360 2174
rect 162308 2110 162360 2116
rect 162320 480 162348 2110
rect 163516 480 163544 3606
rect 164712 480 164740 3606
rect 165908 480 165936 3742
rect 167104 480 167132 4762
rect 168208 480 168236 9046
rect 168392 6866 168420 31470
rect 169024 29708 169076 29714
rect 169024 29650 169076 29656
rect 168380 6860 168432 6866
rect 168380 6802 168432 6808
rect 169036 4010 169064 29650
rect 169404 25634 169432 31484
rect 169772 31470 170338 31498
rect 169392 25628 169444 25634
rect 169392 25570 169444 25576
rect 169772 9178 169800 31470
rect 169760 9172 169812 9178
rect 169760 9114 169812 9120
rect 171152 6118 171180 31484
rect 171244 31470 172086 31498
rect 172532 31470 172914 31498
rect 171244 21486 171272 31470
rect 171784 29640 171836 29646
rect 171784 29582 171836 29588
rect 171232 21480 171284 21486
rect 171232 21422 171284 21428
rect 171140 6112 171192 6118
rect 171140 6054 171192 6060
rect 171796 4162 171824 29582
rect 172426 13152 172482 13161
rect 172426 13087 172482 13096
rect 171612 4134 171824 4162
rect 171612 4078 171640 4134
rect 172440 4078 172468 13087
rect 172532 4894 172560 31470
rect 172992 26738 173020 31606
rect 172716 26710 173020 26738
rect 173912 31470 174662 31498
rect 175292 31470 175490 31498
rect 172716 12458 172744 26710
rect 173912 20126 173940 31470
rect 173900 20120 173952 20126
rect 173900 20062 173952 20068
rect 172624 12430 172744 12458
rect 172624 6050 172652 12430
rect 172612 6044 172664 6050
rect 172612 5986 172664 5992
rect 175292 4962 175320 31470
rect 175568 22114 175596 31606
rect 175476 22098 175596 22114
rect 175464 22092 175596 22098
rect 175516 22086 175596 22092
rect 176672 31470 177238 31498
rect 178052 31470 178158 31498
rect 175464 22034 175516 22040
rect 175556 22024 175608 22030
rect 175556 21966 175608 21972
rect 175370 6216 175426 6225
rect 175370 6151 175426 6160
rect 175280 4956 175332 4962
rect 175280 4898 175332 4904
rect 172520 4888 172572 4894
rect 172520 4830 172572 4836
rect 171600 4072 171652 4078
rect 171600 4014 171652 4020
rect 171784 4072 171836 4078
rect 171784 4014 171836 4020
rect 172428 4072 172480 4078
rect 172428 4014 172480 4020
rect 169024 4004 169076 4010
rect 169024 3946 169076 3952
rect 169390 2000 169446 2009
rect 169390 1935 169446 1944
rect 169404 480 169432 1935
rect 170600 598 170812 626
rect 170600 480 170628 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 170784 66 170812 598
rect 171796 480 171824 4014
rect 172980 4004 173032 4010
rect 172980 3946 173032 3952
rect 172992 480 173020 3946
rect 174176 3732 174228 3738
rect 174176 3674 174228 3680
rect 174188 480 174216 3674
rect 175384 480 175412 6151
rect 175568 5982 175596 21966
rect 176672 18698 176700 31470
rect 176660 18692 176712 18698
rect 176660 18634 176712 18640
rect 177762 9072 177818 9081
rect 177762 9007 177818 9016
rect 175556 5976 175608 5982
rect 175556 5918 175608 5924
rect 176566 2136 176622 2145
rect 176566 2071 176622 2080
rect 176580 480 176608 2071
rect 177776 480 177804 9007
rect 178052 5030 178080 31470
rect 178236 26738 178264 31606
rect 179800 29850 179828 31484
rect 179788 29844 179840 29850
rect 179788 29786 179840 29792
rect 179892 26738 179920 31606
rect 178144 26710 178264 26738
rect 179432 26710 179920 26738
rect 178144 21554 178172 26710
rect 179432 21978 179460 26710
rect 181548 25702 181576 31484
rect 182284 31470 182482 31498
rect 182928 31470 183310 31498
rect 181536 25696 181588 25702
rect 181536 25638 181588 25644
rect 182180 23792 182232 23798
rect 182180 23734 182232 23740
rect 179432 21950 179552 21978
rect 178132 21548 178184 21554
rect 178132 21490 178184 21496
rect 179524 5098 179552 21950
rect 180708 16176 180760 16182
rect 180708 16118 180760 16124
rect 179512 5092 179564 5098
rect 179512 5034 179564 5040
rect 178040 5024 178092 5030
rect 178040 4966 178092 4972
rect 178960 4888 179012 4894
rect 178960 4830 179012 4836
rect 178972 480 179000 4830
rect 180720 3670 180748 16118
rect 181352 9240 181404 9246
rect 181352 9182 181404 9188
rect 180156 3664 180208 3670
rect 180156 3606 180208 3612
rect 180708 3664 180760 3670
rect 180708 3606 180760 3612
rect 180168 480 180196 3606
rect 181364 480 181392 9182
rect 182192 5234 182220 23734
rect 182284 10470 182312 31470
rect 182928 23798 182956 31470
rect 182916 23792 182968 23798
rect 182916 23734 182968 23740
rect 184216 22914 184244 31484
rect 185044 29918 185072 31484
rect 185136 31470 185886 31498
rect 186332 31470 186806 31498
rect 187344 31470 187634 31498
rect 187712 31470 188554 31498
rect 189184 31470 189382 31498
rect 185032 29912 185084 29918
rect 185032 29854 185084 29860
rect 185136 26738 185164 31470
rect 185044 26710 185164 26738
rect 184204 22908 184256 22914
rect 184204 22850 184256 22856
rect 185044 21978 185072 26710
rect 185044 21950 185164 21978
rect 184848 16856 184900 16862
rect 184848 16798 184900 16804
rect 182272 10464 182324 10470
rect 182272 10406 182324 10412
rect 182548 9172 182600 9178
rect 182548 9114 182600 9120
rect 182180 5228 182232 5234
rect 182180 5170 182232 5176
rect 182560 480 182588 9114
rect 183744 2916 183796 2922
rect 183744 2858 183796 2864
rect 183756 480 183784 2858
rect 184860 480 184888 16798
rect 185136 5166 185164 21950
rect 186044 9308 186096 9314
rect 186044 9250 186096 9256
rect 185124 5160 185176 5166
rect 185124 5102 185176 5108
rect 186056 480 186084 9250
rect 186332 7818 186360 31470
rect 187344 26314 187372 31470
rect 186504 26308 186556 26314
rect 186504 26250 186556 26256
rect 187332 26308 187384 26314
rect 187332 26250 187384 26256
rect 186516 14754 186544 26250
rect 187608 16244 187660 16250
rect 187608 16186 187660 16192
rect 186504 14748 186556 14754
rect 186504 14690 186556 14696
rect 186320 7812 186372 7818
rect 186320 7754 186372 7760
rect 187620 3482 187648 16186
rect 187712 5302 187740 31470
rect 189184 24274 189212 31470
rect 190288 29782 190316 31484
rect 190472 31470 191130 31498
rect 191852 31470 192050 31498
rect 190276 29776 190328 29782
rect 190276 29718 190328 29724
rect 189172 24268 189224 24274
rect 189172 24210 189224 24216
rect 190368 13320 190420 13326
rect 190368 13262 190420 13268
rect 187700 5296 187752 5302
rect 187700 5238 187752 5244
rect 190380 3670 190408 13262
rect 190472 5370 190500 31470
rect 191852 7886 191880 31470
rect 192128 28914 192156 31606
rect 191944 28886 192156 28914
rect 193232 31470 193706 31498
rect 194626 31470 194732 31498
rect 191944 26194 191972 28886
rect 191944 26166 192156 26194
rect 192128 21622 192156 26166
rect 192116 21616 192168 21622
rect 192116 21558 192168 21564
rect 193128 16924 193180 16930
rect 193128 16866 193180 16872
rect 191840 7880 191892 7886
rect 191840 7822 191892 7828
rect 191746 6352 191802 6361
rect 191746 6287 191802 6296
rect 190460 5364 190512 5370
rect 190460 5306 190512 5312
rect 189632 3664 189684 3670
rect 189632 3606 189684 3612
rect 190368 3664 190420 3670
rect 190368 3606 190420 3612
rect 187252 3454 187648 3482
rect 187252 480 187280 3454
rect 188448 598 188660 626
rect 188448 480 188476 598
rect 170772 60 170824 66
rect 170772 2 170824 8
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 188632 134 188660 598
rect 189644 480 189672 3606
rect 191760 3398 191788 6287
rect 193140 3398 193168 16866
rect 193232 5438 193260 31470
rect 194704 7954 194732 31470
rect 195440 29714 195468 31484
rect 195992 31470 196374 31498
rect 195428 29708 195480 29714
rect 195428 29650 195480 29656
rect 194692 7948 194744 7954
rect 194692 7890 194744 7896
rect 193310 7848 193366 7857
rect 193310 7783 193366 7792
rect 193220 5432 193272 5438
rect 193220 5374 193272 5380
rect 193324 3482 193352 7783
rect 195992 4758 196020 31470
rect 197188 27062 197216 31484
rect 198108 30190 198136 31484
rect 198752 31470 198950 31498
rect 199028 31470 199778 31498
rect 198096 30184 198148 30190
rect 198096 30126 198148 30132
rect 197176 27056 197228 27062
rect 197176 26998 197228 27004
rect 198752 5506 198780 31470
rect 199028 28966 199056 31470
rect 200684 29646 200712 31484
rect 200672 29640 200724 29646
rect 200672 29582 200724 29588
rect 199016 28960 199068 28966
rect 199016 28902 199068 28908
rect 199108 28960 199160 28966
rect 199108 28902 199160 28908
rect 199120 19378 199148 28902
rect 201512 28422 201540 31484
rect 201604 31470 202446 31498
rect 201500 28416 201552 28422
rect 201500 28358 201552 28364
rect 199108 19372 199160 19378
rect 199108 19314 199160 19320
rect 199200 19372 199252 19378
rect 199200 19314 199252 19320
rect 199212 8022 199240 19314
rect 201406 13288 201462 13297
rect 201406 13223 201462 13232
rect 199200 8016 199252 8022
rect 199200 7958 199252 7964
rect 198740 5500 198792 5506
rect 198740 5442 198792 5448
rect 198186 5128 198242 5137
rect 198186 5063 198242 5072
rect 195980 4752 196032 4758
rect 195980 4694 196032 4700
rect 198200 4146 198228 5063
rect 201420 4146 201448 13223
rect 201604 8158 201632 31470
rect 203260 30258 203288 31484
rect 203248 30252 203300 30258
rect 203248 30194 203300 30200
rect 204180 27130 204208 31484
rect 204272 31470 205022 31498
rect 204168 27124 204220 27130
rect 204168 27066 204220 27072
rect 202788 16992 202840 16998
rect 202788 16934 202840 16940
rect 202800 9654 202828 16934
rect 202788 9648 202840 9654
rect 202788 9590 202840 9596
rect 202512 9580 202564 9586
rect 202512 9522 202564 9528
rect 201592 8152 201644 8158
rect 201592 8094 201644 8100
rect 198188 4140 198240 4146
rect 198188 4082 198240 4088
rect 200396 4140 200448 4146
rect 200396 4082 200448 4088
rect 201408 4140 201460 4146
rect 201408 4082 201460 4088
rect 198004 4072 198056 4078
rect 198004 4014 198056 4020
rect 196808 3936 196860 3942
rect 196808 3878 196860 3884
rect 193232 3454 193352 3482
rect 191748 3392 191800 3398
rect 191748 3334 191800 3340
rect 192024 3392 192076 3398
rect 192024 3334 192076 3340
rect 193128 3392 193180 3398
rect 193128 3334 193180 3340
rect 190828 3052 190880 3058
rect 190828 2994 190880 3000
rect 190840 480 190868 2994
rect 192036 480 192064 3334
rect 193232 480 193260 3454
rect 194416 2236 194468 2242
rect 194416 2178 194468 2184
rect 194428 480 194456 2178
rect 195624 598 195836 626
rect 195624 480 195652 598
rect 188620 128 188672 134
rect 188620 70 188672 76
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 195808 202 195836 598
rect 196820 480 196848 3878
rect 198016 480 198044 4014
rect 199212 598 199424 626
rect 199212 480 199240 598
rect 195796 196 195848 202
rect 195796 138 195848 144
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 199396 270 199424 598
rect 200408 480 200436 4082
rect 201500 2304 201552 2310
rect 201500 2246 201552 2252
rect 201512 480 201540 2246
rect 202524 610 202552 9522
rect 203892 9376 203944 9382
rect 203892 9318 203944 9324
rect 202512 604 202564 610
rect 202512 546 202564 552
rect 202696 604 202748 610
rect 202696 546 202748 552
rect 202708 480 202736 546
rect 203904 480 203932 9318
rect 204272 8090 204300 31470
rect 205836 29578 205864 31484
rect 206020 31470 206770 31498
rect 207032 31470 207598 31498
rect 205824 29572 205876 29578
rect 205824 29514 205876 29520
rect 206020 26738 206048 31470
rect 205836 26710 206048 26738
rect 205836 20194 205864 26710
rect 205824 20188 205876 20194
rect 205824 20130 205876 20136
rect 204352 9444 204404 9450
rect 204352 9386 204404 9392
rect 204260 8084 204312 8090
rect 204260 8026 204312 8032
rect 204364 3942 204392 9386
rect 206284 6180 206336 6186
rect 206284 6122 206336 6128
rect 204352 3936 204404 3942
rect 204352 3878 204404 3884
rect 205088 3256 205140 3262
rect 205088 3198 205140 3204
rect 205100 480 205128 3198
rect 206296 480 206324 6122
rect 207032 4690 207060 31470
rect 208504 29510 208532 31484
rect 208492 29504 208544 29510
rect 208492 29446 208544 29452
rect 208780 26738 208808 31606
rect 210252 28286 210280 31484
rect 211080 29442 211108 31484
rect 231964 30326 231992 38542
rect 284588 30326 284616 31484
rect 231952 30320 232004 30326
rect 231952 30262 232004 30268
rect 284576 30320 284628 30326
rect 284576 30262 284628 30268
rect 211068 29436 211120 29442
rect 211068 29378 211120 29384
rect 210240 28280 210292 28286
rect 210240 28222 210292 28228
rect 411916 27577 411944 222838
rect 412008 49881 412036 225558
rect 412100 83570 412128 502930
rect 414032 502846 414184 502874
rect 414032 496126 414060 502846
rect 416148 500274 416176 502982
rect 417424 501628 417476 501634
rect 417424 501570 417476 501576
rect 416136 500268 416188 500274
rect 416136 500210 416188 500216
rect 414020 496120 414072 496126
rect 414020 496062 414072 496068
rect 417436 327078 417464 501570
rect 420840 500954 420868 502982
rect 433444 502982 433596 503010
rect 435560 502982 435712 503010
rect 442000 502982 442152 503010
rect 446324 502982 446476 503010
rect 480824 502982 481312 503010
rect 574008 502998 574060 503004
rect 422832 502846 423168 502874
rect 424948 502846 425008 502874
rect 427064 502846 427124 502874
rect 429272 502846 429332 502874
rect 431388 502846 431448 502874
rect 423140 500954 423168 502846
rect 424980 500954 425008 502846
rect 427096 500954 427124 502846
rect 429304 500954 429332 502846
rect 431420 500954 431448 502846
rect 433444 500954 433472 502982
rect 435560 500954 435588 502982
rect 437584 502846 437920 502874
rect 439700 502846 440036 502874
rect 437584 500954 437612 502846
rect 439700 500954 439728 502846
rect 442000 500954 442028 502982
rect 444360 502846 444420 502874
rect 444392 500954 444420 502846
rect 446324 500954 446352 502982
rect 448532 502846 448684 502874
rect 450464 502846 450800 502874
rect 453008 502846 453344 502874
rect 455124 502846 455368 502874
rect 457332 502846 457392 502874
rect 459448 502846 459508 502874
rect 448532 500954 448560 502846
rect 450464 500954 450492 502846
rect 453316 500954 453344 502846
rect 455340 500954 455368 502846
rect 457364 500954 457392 502846
rect 459480 502722 459508 502846
rect 461228 502846 461900 502874
rect 463772 502846 464108 502874
rect 465888 502846 465948 502874
rect 468096 502846 468156 502874
rect 470212 502846 470272 502874
rect 472420 502846 472756 502874
rect 474536 502846 474688 502874
rect 477756 502846 477816 502874
rect 461228 502722 461256 502846
rect 459468 502716 459520 502722
rect 459468 502658 459520 502664
rect 461216 502716 461268 502722
rect 461216 502658 461268 502664
rect 461872 500954 461900 502846
rect 464080 500954 464108 502846
rect 465920 500954 465948 502846
rect 468128 500954 468156 502846
rect 470244 500954 470272 502846
rect 472728 500954 472756 502846
rect 474660 500954 474688 502846
rect 477788 500954 477816 502846
rect 480824 500954 480852 502982
rect 481284 502926 481312 502982
rect 481272 502920 481324 502926
rect 484308 502920 484360 502926
rect 481272 502862 481324 502868
rect 484196 502868 484308 502874
rect 484196 502862 484360 502868
rect 487160 502920 487212 502926
rect 487212 502868 487508 502874
rect 487160 502862 487508 502868
rect 484196 502846 484348 502862
rect 487172 502846 487508 502862
rect 491740 502846 491892 502874
rect 492844 502846 493180 502874
rect 493948 502846 494008 502874
rect 495052 502846 495388 502874
rect 496064 502846 496768 502874
rect 497168 502846 497504 502874
rect 498272 502846 498608 502874
rect 499284 502846 499436 502874
rect 500388 502846 500908 502874
rect 501492 502846 501828 502874
rect 502596 502846 502932 502874
rect 420828 500948 420880 500954
rect 420828 500890 420880 500896
rect 423128 500948 423180 500954
rect 423128 500890 423180 500896
rect 424968 500948 425020 500954
rect 424968 500890 425020 500896
rect 427084 500948 427136 500954
rect 427084 500890 427136 500896
rect 429292 500948 429344 500954
rect 429292 500890 429344 500896
rect 431408 500948 431460 500954
rect 431408 500890 431460 500896
rect 433432 500948 433484 500954
rect 433432 500890 433484 500896
rect 435548 500948 435600 500954
rect 435548 500890 435600 500896
rect 437572 500948 437624 500954
rect 437572 500890 437624 500896
rect 439688 500948 439740 500954
rect 439688 500890 439740 500896
rect 441988 500948 442040 500954
rect 441988 500890 442040 500896
rect 444380 500948 444432 500954
rect 444380 500890 444432 500896
rect 446312 500948 446364 500954
rect 446312 500890 446364 500896
rect 448520 500948 448572 500954
rect 448520 500890 448572 500896
rect 450452 500948 450504 500954
rect 450452 500890 450504 500896
rect 453304 500948 453356 500954
rect 453304 500890 453356 500896
rect 455328 500948 455380 500954
rect 455328 500890 455380 500896
rect 457352 500948 457404 500954
rect 457352 500890 457404 500896
rect 461860 500948 461912 500954
rect 461860 500890 461912 500896
rect 464068 500948 464120 500954
rect 464068 500890 464120 500896
rect 465908 500948 465960 500954
rect 465908 500890 465960 500896
rect 468116 500948 468168 500954
rect 468116 500890 468168 500896
rect 470232 500948 470284 500954
rect 470232 500890 470284 500896
rect 472716 500948 472768 500954
rect 472716 500890 472768 500896
rect 474648 500948 474700 500954
rect 474648 500890 474700 500896
rect 477776 500948 477828 500954
rect 477776 500890 477828 500896
rect 480812 500948 480864 500954
rect 480812 500890 480864 500896
rect 491864 500857 491892 502846
rect 493152 500857 493180 502846
rect 491850 500848 491906 500857
rect 491850 500783 491906 500792
rect 493138 500848 493194 500857
rect 493138 500783 493194 500792
rect 443644 490612 443696 490618
rect 443644 490554 443696 490560
rect 418158 473784 418214 473793
rect 418080 473742 418158 473770
rect 418080 473657 418108 473742
rect 418158 473719 418214 473728
rect 437386 473784 437442 473793
rect 437570 473784 437626 473793
rect 437442 473742 437570 473770
rect 437386 473719 437442 473728
rect 437570 473719 437626 473728
rect 418066 473648 418122 473657
rect 418066 473583 418122 473592
rect 427726 473376 427782 473385
rect 427910 473376 427966 473385
rect 427782 473334 427910 473362
rect 427726 473311 427782 473320
rect 427910 473311 427966 473320
rect 443656 450673 443684 490554
rect 493980 475561 494008 502846
rect 493966 475552 494022 475561
rect 493966 475487 494022 475496
rect 495360 475425 495388 502846
rect 496740 487801 496768 502846
rect 497476 500410 497504 502846
rect 497464 500404 497516 500410
rect 497464 500346 497516 500352
rect 498108 500404 498160 500410
rect 498108 500346 498160 500352
rect 496726 487792 496782 487801
rect 496726 487727 496782 487736
rect 495346 475416 495402 475425
rect 495346 475351 495402 475360
rect 498120 474026 498148 500346
rect 498580 500274 498608 502846
rect 498568 500268 498620 500274
rect 498568 500210 498620 500216
rect 499408 476785 499436 502846
rect 499488 500268 499540 500274
rect 499488 500210 499540 500216
rect 499394 476776 499450 476785
rect 499394 476711 499450 476720
rect 499500 475386 499528 500210
rect 500880 475697 500908 502846
rect 501800 500002 501828 502846
rect 502904 500954 502932 502846
rect 503594 502602 503622 502860
rect 504712 502846 505048 502874
rect 505816 502846 506428 502874
rect 506828 502846 507164 502874
rect 507932 502846 508268 502874
rect 509036 502846 509188 502874
rect 510140 502846 510568 502874
rect 511152 502846 511488 502874
rect 512256 502846 512592 502874
rect 513360 502846 513696 502874
rect 514372 502846 514616 502874
rect 515476 502846 516088 502874
rect 516580 502846 516916 502874
rect 517684 502846 518020 502874
rect 518696 502846 518848 502874
rect 519800 502846 520228 502874
rect 520904 502846 521608 502874
rect 521916 502846 522252 502874
rect 523020 502846 523356 502874
rect 524124 502846 524276 502874
rect 525228 502846 525748 502874
rect 526240 502846 526576 502874
rect 527344 502846 527680 502874
rect 528448 502846 528508 502874
rect 529460 502846 529888 502874
rect 530564 502846 531268 502874
rect 531668 502846 532004 502874
rect 532772 502846 533108 502874
rect 533784 502846 534028 502874
rect 534888 502846 535224 502874
rect 535992 502846 536328 502874
rect 537004 502846 537340 502874
rect 538108 502846 538168 502874
rect 539212 502846 539548 502874
rect 540316 502846 540928 502874
rect 541328 502846 541664 502874
rect 542432 502846 542676 502874
rect 543536 502846 543688 502874
rect 544548 502846 545068 502874
rect 545652 502846 545988 502874
rect 546756 502846 547092 502874
rect 547860 502846 548196 502874
rect 548872 502846 549208 502874
rect 549976 502846 550128 502874
rect 551080 502846 551416 502874
rect 552092 502846 552428 502874
rect 553196 502846 553348 502874
rect 554300 502846 554728 502874
rect 555404 502846 555556 502874
rect 503548 502574 503622 502602
rect 502892 500948 502944 500954
rect 502892 500890 502944 500896
rect 501788 499996 501840 500002
rect 501788 499938 501840 499944
rect 502248 499996 502300 500002
rect 502248 499938 502300 499944
rect 501604 498840 501656 498846
rect 501604 498782 501656 498788
rect 500866 475688 500922 475697
rect 500866 475623 500922 475632
rect 499488 475380 499540 475386
rect 499488 475322 499540 475328
rect 501616 474774 501644 498782
rect 502260 476921 502288 499938
rect 503548 477057 503576 502574
rect 503628 500948 503680 500954
rect 503628 500890 503680 500896
rect 503534 477048 503590 477057
rect 503534 476983 503590 476992
rect 502246 476912 502302 476921
rect 502246 476847 502302 476856
rect 503640 475833 503668 500890
rect 503626 475824 503682 475833
rect 503626 475759 503682 475768
rect 499304 474768 499356 474774
rect 499304 474710 499356 474716
rect 501604 474768 501656 474774
rect 501604 474710 501656 474716
rect 498108 474020 498160 474026
rect 498108 473962 498160 473968
rect 481638 473784 481694 473793
rect 481638 473719 481640 473728
rect 481692 473719 481694 473728
rect 490656 473748 490708 473754
rect 481640 473690 481692 473696
rect 490656 473690 490708 473696
rect 490668 473657 490696 473690
rect 490654 473648 490710 473657
rect 499316 473620 499344 474710
rect 505020 474065 505048 502846
rect 506400 477193 506428 502846
rect 507136 500410 507164 502846
rect 508240 500857 508268 502846
rect 508226 500848 508282 500857
rect 508226 500783 508282 500792
rect 507124 500404 507176 500410
rect 507124 500346 507176 500352
rect 507768 500404 507820 500410
rect 507768 500346 507820 500352
rect 506386 477184 506442 477193
rect 506386 477119 506442 477128
rect 507780 475969 507808 500346
rect 509160 476105 509188 502846
rect 510540 476814 510568 502846
rect 511460 500954 511488 502846
rect 511448 500948 511500 500954
rect 511448 500890 511500 500896
rect 511908 500948 511960 500954
rect 511908 500890 511960 500896
rect 510528 476808 510580 476814
rect 510528 476750 510580 476756
rect 508502 476096 508558 476105
rect 508502 476031 508558 476040
rect 509146 476096 509202 476105
rect 509146 476031 509202 476040
rect 507766 475960 507822 475969
rect 507766 475895 507822 475904
rect 505006 474056 505062 474065
rect 505006 473991 505062 474000
rect 505006 473648 505062 473657
rect 490654 473583 490710 473592
rect 505006 473583 505008 473592
rect 505060 473583 505062 473592
rect 505008 473554 505060 473560
rect 491850 473512 491906 473521
rect 491850 473447 491852 473456
rect 491904 473447 491906 473456
rect 493138 473512 493194 473521
rect 508516 473482 508544 476031
rect 511920 474094 511948 500890
rect 512564 500682 512592 502846
rect 513668 500682 513696 502846
rect 512552 500676 512604 500682
rect 512552 500618 512604 500624
rect 513288 500676 513340 500682
rect 513288 500618 513340 500624
rect 513656 500676 513708 500682
rect 513656 500618 513708 500624
rect 513300 474201 513328 500618
rect 514588 476882 514616 502846
rect 514668 500676 514720 500682
rect 514668 500618 514720 500624
rect 514576 476876 514628 476882
rect 514576 476818 514628 476824
rect 513286 474192 513342 474201
rect 514680 474162 514708 500618
rect 516060 474230 516088 502846
rect 516888 500954 516916 502846
rect 516876 500948 516928 500954
rect 516876 500890 516928 500896
rect 517428 500948 517480 500954
rect 517428 500890 517480 500896
rect 517440 476950 517468 500890
rect 517992 500857 518020 502846
rect 517978 500848 518034 500857
rect 517978 500783 518034 500792
rect 518820 477018 518848 502846
rect 518808 477012 518860 477018
rect 518808 476954 518860 476960
rect 517428 476944 517480 476950
rect 517428 476886 517480 476892
rect 520200 474337 520228 502846
rect 521580 477086 521608 502846
rect 522224 500274 522252 502846
rect 523328 500954 523356 502846
rect 523316 500948 523368 500954
rect 523316 500890 523368 500896
rect 524248 500342 524276 502846
rect 524328 500948 524380 500954
rect 524328 500890 524380 500896
rect 524236 500336 524288 500342
rect 524236 500278 524288 500284
rect 522212 500268 522264 500274
rect 522212 500210 522264 500216
rect 521568 477080 521620 477086
rect 521568 477022 521620 477028
rect 524340 475454 524368 500890
rect 525720 475522 525748 502846
rect 526548 500410 526576 502846
rect 526536 500404 526588 500410
rect 526536 500346 526588 500352
rect 527652 500206 527680 502846
rect 528480 500478 528508 502846
rect 528468 500472 528520 500478
rect 528468 500414 528520 500420
rect 527640 500200 527692 500206
rect 527640 500142 527692 500148
rect 528468 500200 528520 500206
rect 528468 500142 528520 500148
rect 528480 475590 528508 500142
rect 528468 475584 528520 475590
rect 528468 475526 528520 475532
rect 525708 475516 525760 475522
rect 525708 475458 525760 475464
rect 524328 475448 524380 475454
rect 524328 475390 524380 475396
rect 520186 474328 520242 474337
rect 529860 474298 529888 502846
rect 531240 477154 531268 502846
rect 531976 500546 532004 502846
rect 533080 500546 533108 502846
rect 531964 500540 532016 500546
rect 531964 500482 532016 500488
rect 532608 500540 532660 500546
rect 532608 500482 532660 500488
rect 533068 500540 533120 500546
rect 533068 500482 533120 500488
rect 531228 477148 531280 477154
rect 531228 477090 531280 477096
rect 532620 475658 532648 500482
rect 532608 475652 532660 475658
rect 532608 475594 532660 475600
rect 534000 474366 534028 502846
rect 535196 500614 535224 502846
rect 535184 500608 535236 500614
rect 535184 500550 535236 500556
rect 536300 500206 536328 502846
rect 537312 500682 537340 502846
rect 537300 500676 537352 500682
rect 537300 500618 537352 500624
rect 536288 500200 536340 500206
rect 536288 500142 536340 500148
rect 536748 500200 536800 500206
rect 536748 500142 536800 500148
rect 536760 475726 536788 500142
rect 538140 475794 538168 502846
rect 539520 500750 539548 502846
rect 539508 500744 539560 500750
rect 539508 500686 539560 500692
rect 538128 475788 538180 475794
rect 538128 475730 538180 475736
rect 536748 475720 536800 475726
rect 536748 475662 536800 475668
rect 540900 474434 540928 502846
rect 541636 500818 541664 502846
rect 542648 500857 542676 502846
rect 543660 500886 543688 502846
rect 543648 500880 543700 500886
rect 542634 500848 542690 500857
rect 541624 500812 541676 500818
rect 543648 500822 543700 500828
rect 542634 500783 542690 500792
rect 541624 500754 541676 500760
rect 542910 476232 542966 476241
rect 542910 476167 542966 476176
rect 540888 474428 540940 474434
rect 540888 474370 540940 474376
rect 533988 474360 534040 474366
rect 533988 474302 534040 474308
rect 520186 474263 520242 474272
rect 529848 474292 529900 474298
rect 529848 474234 529900 474240
rect 516048 474224 516100 474230
rect 516048 474166 516100 474172
rect 513286 474127 513342 474136
rect 514668 474156 514720 474162
rect 514668 474098 514720 474104
rect 511908 474088 511960 474094
rect 511908 474030 511960 474036
rect 520738 473920 520794 473929
rect 520738 473855 520794 473864
rect 512642 473784 512698 473793
rect 512642 473719 512698 473728
rect 512656 473618 512684 473719
rect 520556 473680 520608 473686
rect 520556 473622 520608 473628
rect 512644 473612 512696 473618
rect 512644 473554 512696 473560
rect 520464 473612 520516 473618
rect 520464 473554 520516 473560
rect 520476 473482 520504 473554
rect 520568 473482 520596 473622
rect 520752 473482 520780 473855
rect 522672 473680 522724 473686
rect 522672 473622 522724 473628
rect 522684 473482 522712 473622
rect 522856 473612 522908 473618
rect 522856 473554 522908 473560
rect 522868 473482 522896 473554
rect 542924 473482 542952 476167
rect 545040 474502 545068 502846
rect 545960 500954 545988 502846
rect 545948 500948 546000 500954
rect 545948 500890 546000 500896
rect 547064 500206 547092 502846
rect 547972 500336 548024 500342
rect 547972 500278 548024 500284
rect 547052 500200 547104 500206
rect 547052 500142 547104 500148
rect 547984 500138 548012 500278
rect 548168 500274 548196 502846
rect 548156 500268 548208 500274
rect 548156 500210 548208 500216
rect 547972 500132 548024 500138
rect 547972 500074 548024 500080
rect 547328 476944 547380 476950
rect 547328 476886 547380 476892
rect 547340 476610 547368 476886
rect 547328 476604 547380 476610
rect 547328 476546 547380 476552
rect 549180 475590 549208 502846
rect 550100 500857 550128 502846
rect 550086 500848 550142 500857
rect 550086 500783 550142 500792
rect 551388 500546 551416 502846
rect 552400 500954 552428 502846
rect 552112 500948 552164 500954
rect 552112 500890 552164 500896
rect 552388 500948 552440 500954
rect 552388 500890 552440 500896
rect 552124 500750 552152 500890
rect 552020 500744 552072 500750
rect 552020 500686 552072 500692
rect 552112 500744 552164 500750
rect 552112 500686 552164 500692
rect 551192 500540 551244 500546
rect 551192 500482 551244 500488
rect 551376 500540 551428 500546
rect 551376 500482 551428 500488
rect 551928 500540 551980 500546
rect 551928 500482 551980 500488
rect 551204 500070 551232 500482
rect 551284 500404 551336 500410
rect 551284 500346 551336 500352
rect 551376 500404 551428 500410
rect 551376 500346 551428 500352
rect 551192 500064 551244 500070
rect 551192 500006 551244 500012
rect 549168 475584 549220 475590
rect 549168 475526 549220 475532
rect 547420 475448 547472 475454
rect 547420 475390 547472 475396
rect 547432 474570 547460 475390
rect 547420 474564 547472 474570
rect 547420 474506 547472 474512
rect 545028 474496 545080 474502
rect 545028 474438 545080 474444
rect 493138 473447 493140 473456
rect 491852 473418 491904 473424
rect 493192 473447 493194 473456
rect 508504 473476 508556 473482
rect 493140 473418 493192 473424
rect 508504 473418 508556 473424
rect 520464 473476 520516 473482
rect 520464 473418 520516 473424
rect 520556 473476 520608 473482
rect 520556 473418 520608 473424
rect 520740 473476 520792 473482
rect 520740 473418 520792 473424
rect 522672 473476 522724 473482
rect 522672 473418 522724 473424
rect 522856 473476 522908 473482
rect 522856 473418 522908 473424
rect 542912 473476 542964 473482
rect 542912 473418 542964 473424
rect 447784 473408 447836 473414
rect 447784 473350 447836 473356
rect 443642 450664 443698 450673
rect 443642 450599 443698 450608
rect 447796 426426 447824 473350
rect 551296 456362 551324 500346
rect 551388 457042 551416 500346
rect 551940 477018 551968 500482
rect 551928 477012 551980 477018
rect 551928 476954 551980 476960
rect 551928 476876 551980 476882
rect 551928 476818 551980 476824
rect 551744 475788 551796 475794
rect 551744 475730 551796 475736
rect 551652 475652 551704 475658
rect 551652 475594 551704 475600
rect 551560 475584 551612 475590
rect 551560 475526 551612 475532
rect 551468 473340 551520 473346
rect 551468 473282 551520 473288
rect 551480 472258 551508 473282
rect 551572 472326 551600 475526
rect 551560 472320 551612 472326
rect 551560 472262 551612 472268
rect 551468 472252 551520 472258
rect 551468 472194 551520 472200
rect 551560 472184 551612 472190
rect 551560 472126 551612 472132
rect 551572 471594 551600 472126
rect 551664 471850 551692 475594
rect 551756 472190 551784 475730
rect 551836 474360 551888 474366
rect 551836 474302 551888 474308
rect 551744 472184 551796 472190
rect 551744 472126 551796 472132
rect 551744 472048 551796 472054
rect 551744 471990 551796 471996
rect 551652 471844 551704 471850
rect 551652 471786 551704 471792
rect 551480 471566 551600 471594
rect 551480 459320 551508 471566
rect 551756 471458 551784 471990
rect 551572 471430 551784 471458
rect 551572 459898 551600 471430
rect 551744 471232 551796 471238
rect 551664 471180 551744 471186
rect 551664 471174 551796 471180
rect 551664 471158 551784 471174
rect 551664 466290 551692 471158
rect 551848 470694 551876 474302
rect 551836 470688 551888 470694
rect 551836 470630 551888 470636
rect 551940 470506 551968 476818
rect 551756 470478 551968 470506
rect 551756 466410 551784 470478
rect 551744 466404 551796 466410
rect 551744 466346 551796 466352
rect 551664 466262 551876 466290
rect 551744 466200 551796 466206
rect 551744 466142 551796 466148
rect 551756 460766 551784 466142
rect 551848 460902 551876 466262
rect 551836 460896 551888 460902
rect 551836 460838 551888 460844
rect 551744 460760 551796 460766
rect 551744 460702 551796 460708
rect 551572 459882 551784 459898
rect 551572 459876 551796 459882
rect 551572 459870 551744 459876
rect 551744 459818 551796 459824
rect 551928 459876 551980 459882
rect 551928 459818 551980 459824
rect 551744 459332 551796 459338
rect 551480 459292 551744 459320
rect 551744 459274 551796 459280
rect 551388 457014 551784 457042
rect 551756 456822 551784 457014
rect 551744 456816 551796 456822
rect 551744 456758 551796 456764
rect 551296 456346 551784 456362
rect 551296 456340 551796 456346
rect 551296 456334 551744 456340
rect 551744 456282 551796 456288
rect 551744 454912 551796 454918
rect 551480 454872 551744 454900
rect 551480 451058 551508 454872
rect 551744 454854 551796 454860
rect 551744 454776 551796 454782
rect 551572 454724 551744 454730
rect 551572 454718 551796 454724
rect 551572 454702 551784 454718
rect 551572 451194 551600 454702
rect 551940 451738 551968 459818
rect 552032 454170 552060 500686
rect 553320 500342 553348 502846
rect 553492 500948 553544 500954
rect 553492 500890 553544 500896
rect 553308 500336 553360 500342
rect 553308 500278 553360 500284
rect 552664 500200 552716 500206
rect 552664 500142 552716 500148
rect 552112 476944 552164 476950
rect 552112 476886 552164 476892
rect 552124 472666 552152 476886
rect 552676 476338 552704 500142
rect 552756 477148 552808 477154
rect 552756 477090 552808 477096
rect 552664 476332 552716 476338
rect 552664 476274 552716 476280
rect 552478 475552 552534 475561
rect 552478 475487 552534 475496
rect 552294 474600 552350 474609
rect 552294 474535 552350 474544
rect 552204 472864 552256 472870
rect 552204 472806 552256 472812
rect 552112 472660 552164 472666
rect 552112 472602 552164 472608
rect 552110 472560 552166 472569
rect 552110 472495 552166 472504
rect 552124 472462 552152 472495
rect 552112 472456 552164 472462
rect 552216 472433 552244 472806
rect 552112 472398 552164 472404
rect 552202 472424 552258 472433
rect 552202 472359 552258 472368
rect 552112 472320 552164 472326
rect 552112 472262 552164 472268
rect 552020 454164 552072 454170
rect 552020 454106 552072 454112
rect 552018 451752 552074 451761
rect 551940 451710 552018 451738
rect 552018 451687 552074 451696
rect 552018 451208 552074 451217
rect 551572 451166 552018 451194
rect 552018 451143 552074 451152
rect 551480 451030 551600 451058
rect 551572 447658 551600 451030
rect 552018 447672 552074 447681
rect 551572 447630 552018 447658
rect 552018 447607 552074 447616
rect 552124 441697 552152 472262
rect 552204 472252 552256 472258
rect 552204 472194 552256 472200
rect 552216 452062 552244 472194
rect 552308 470801 552336 474535
rect 552388 474020 552440 474026
rect 552388 473962 552440 473968
rect 552294 470792 552350 470801
rect 552294 470727 552350 470736
rect 552296 470688 552348 470694
rect 552296 470630 552348 470636
rect 552308 453234 552336 470630
rect 552400 470121 552428 473962
rect 552492 471889 552520 475487
rect 552572 475380 552624 475386
rect 552572 475322 552624 475328
rect 552478 471880 552534 471889
rect 552478 471815 552534 471824
rect 552480 471776 552532 471782
rect 552480 471718 552532 471724
rect 552386 470112 552442 470121
rect 552386 470047 552442 470056
rect 552388 470008 552440 470014
rect 552388 469950 552440 469956
rect 552400 461650 552428 469950
rect 552492 466410 552520 471718
rect 552584 469577 552612 475322
rect 552664 474224 552716 474230
rect 552664 474166 552716 474172
rect 552570 469568 552626 469577
rect 552570 469503 552626 469512
rect 552676 469418 552704 474166
rect 552768 472054 552796 477090
rect 553216 477080 553268 477086
rect 553216 477022 553268 477028
rect 553124 476808 553176 476814
rect 553124 476750 553176 476756
rect 552848 475516 552900 475522
rect 552848 475458 552900 475464
rect 552756 472048 552808 472054
rect 552756 471990 552808 471996
rect 552756 471912 552808 471918
rect 552756 471854 552808 471860
rect 552584 469390 552704 469418
rect 552480 466404 552532 466410
rect 552480 466346 552532 466352
rect 552584 463162 552612 469390
rect 552768 466478 552796 471854
rect 552860 470014 552888 475458
rect 552940 475448 552992 475454
rect 552940 475390 552992 475396
rect 552952 471782 552980 475390
rect 553032 472932 553084 472938
rect 553032 472874 553084 472880
rect 553044 472705 553072 472874
rect 553030 472696 553086 472705
rect 553030 472631 553086 472640
rect 553032 472592 553084 472598
rect 553032 472534 553084 472540
rect 552940 471776 552992 471782
rect 552940 471718 552992 471724
rect 553044 471578 553072 472534
rect 552940 471572 552992 471578
rect 552940 471514 552992 471520
rect 553032 471572 553084 471578
rect 553032 471514 553084 471520
rect 552848 470008 552900 470014
rect 552848 469950 552900 469956
rect 552952 469826 552980 471514
rect 553136 471458 553164 476750
rect 553228 471918 553256 477022
rect 553308 476604 553360 476610
rect 553308 476546 553360 476552
rect 553216 471912 553268 471918
rect 553216 471854 553268 471860
rect 553320 471730 553348 476546
rect 553400 474496 553452 474502
rect 553400 474438 553452 474444
rect 552860 469798 552980 469826
rect 553044 471430 553164 471458
rect 553228 471702 553348 471730
rect 552664 466472 552716 466478
rect 552664 466414 552716 466420
rect 552756 466472 552808 466478
rect 552756 466414 552808 466420
rect 552676 463758 552704 466414
rect 552664 463752 552716 463758
rect 552664 463694 552716 463700
rect 552756 463752 552808 463758
rect 552756 463694 552808 463700
rect 552584 463134 552704 463162
rect 552388 461644 552440 461650
rect 552388 461586 552440 461592
rect 552572 461644 552624 461650
rect 552572 461586 552624 461592
rect 552388 460760 552440 460766
rect 552386 460728 552388 460737
rect 552440 460728 552442 460737
rect 552386 460663 552442 460672
rect 552388 460624 552440 460630
rect 552388 460566 552440 460572
rect 552400 454753 552428 460566
rect 552480 459332 552532 459338
rect 552480 459274 552532 459280
rect 552492 454918 552520 459274
rect 552480 454912 552532 454918
rect 552480 454854 552532 454860
rect 552386 454744 552442 454753
rect 552386 454679 552442 454688
rect 552480 454164 552532 454170
rect 552480 454106 552532 454112
rect 552308 453206 552428 453234
rect 552204 452056 552256 452062
rect 552204 451998 552256 452004
rect 552204 451920 552256 451926
rect 552204 451862 552256 451868
rect 552216 447001 552244 451862
rect 552400 449993 552428 453206
rect 552492 451926 552520 454106
rect 552584 453529 552612 461586
rect 552676 460057 552704 463134
rect 552662 460048 552718 460057
rect 552662 459983 552718 459992
rect 552664 456816 552716 456822
rect 552664 456758 552716 456764
rect 552768 456770 552796 463694
rect 552860 458017 552888 469798
rect 552940 468444 552992 468450
rect 552940 468386 552992 468392
rect 552952 459241 552980 468386
rect 553044 462777 553072 471430
rect 553228 468450 553256 471702
rect 553216 468444 553268 468450
rect 553216 468386 553268 468392
rect 553124 466404 553176 466410
rect 553124 466346 553176 466352
rect 553030 462768 553086 462777
rect 553030 462703 553086 462712
rect 553032 460896 553084 460902
rect 553032 460838 553084 460844
rect 552938 459232 552994 459241
rect 552938 459167 552994 459176
rect 552846 458008 552902 458017
rect 552846 457943 552902 457952
rect 552846 456784 552902 456793
rect 552570 453520 552626 453529
rect 552570 453455 552626 453464
rect 552676 452985 552704 456758
rect 552768 456742 552846 456770
rect 552846 456719 552902 456728
rect 552756 456340 552808 456346
rect 552756 456282 552808 456288
rect 552768 454209 552796 456282
rect 553044 454782 553072 460838
rect 553136 460630 553164 466346
rect 553124 460624 553176 460630
rect 553124 460566 553176 460572
rect 553032 454776 553084 454782
rect 553032 454718 553084 454724
rect 552754 454200 552810 454209
rect 552754 454135 552810 454144
rect 552662 452976 552718 452985
rect 552662 452911 552718 452920
rect 552572 452056 552624 452062
rect 552572 451998 552624 452004
rect 552480 451920 552532 451926
rect 552480 451862 552532 451868
rect 552386 449984 552442 449993
rect 552386 449919 552442 449928
rect 552202 446992 552258 447001
rect 552202 446927 552258 446936
rect 552584 445233 552612 451998
rect 552570 445224 552626 445233
rect 552570 445159 552626 445168
rect 553412 443737 553440 474438
rect 553398 443728 553454 443737
rect 553398 443663 553454 443672
rect 552110 441688 552166 441697
rect 552110 441623 552166 441632
rect 553504 439657 553532 500890
rect 553768 500880 553820 500886
rect 553768 500822 553820 500828
rect 553676 500744 553728 500750
rect 553676 500686 553728 500692
rect 553584 500268 553636 500274
rect 553584 500210 553636 500216
rect 553596 441969 553624 500210
rect 553688 443193 553716 500686
rect 553780 444417 553808 500822
rect 553860 500812 553912 500818
rect 553860 500754 553912 500760
rect 553872 445505 553900 500754
rect 553952 500676 554004 500682
rect 553952 500618 554004 500624
rect 553964 447953 553992 500618
rect 554044 500608 554096 500614
rect 554044 500550 554096 500556
rect 554056 449041 554084 500550
rect 554228 500336 554280 500342
rect 554228 500278 554280 500284
rect 554136 477012 554188 477018
rect 554136 476954 554188 476960
rect 554042 449032 554098 449041
rect 554042 448967 554098 448976
rect 553950 447944 554006 447953
rect 553950 447879 554006 447888
rect 553858 445496 553914 445505
rect 553858 445431 553914 445440
rect 553766 444408 553822 444417
rect 553766 444343 553822 444352
rect 553674 443184 553730 443193
rect 553674 443119 553730 443128
rect 553582 441960 553638 441969
rect 553582 441895 553638 441904
rect 554148 440201 554176 476954
rect 554134 440192 554190 440201
rect 554134 440127 554190 440136
rect 553490 439648 553546 439657
rect 553490 439583 553546 439592
rect 554240 438977 554268 500278
rect 554320 475720 554372 475726
rect 554320 475662 554372 475668
rect 554332 448497 554360 475662
rect 554700 474094 554728 502846
rect 555056 500404 555108 500410
rect 555056 500346 555108 500352
rect 554964 500132 555016 500138
rect 554964 500074 555016 500080
rect 554688 474088 554740 474094
rect 554688 474030 554740 474036
rect 554872 469192 554924 469198
rect 554872 469134 554924 469140
rect 554884 455569 554912 469134
rect 554870 455560 554926 455569
rect 554870 455495 554926 455504
rect 554976 455025 555004 500074
rect 555068 456249 555096 500346
rect 555424 500064 555476 500070
rect 555424 500006 555476 500012
rect 555240 476332 555292 476338
rect 555240 476274 555292 476280
rect 555148 474088 555200 474094
rect 555148 474030 555200 474036
rect 555054 456240 555110 456249
rect 555054 456175 555110 456184
rect 554962 455016 555018 455025
rect 554962 454951 555018 454960
rect 554318 448488 554374 448497
rect 554318 448423 554374 448432
rect 554226 438968 554282 438977
rect 554226 438903 554282 438912
rect 554872 438932 554924 438938
rect 554872 438874 554924 438880
rect 554780 437300 554832 437306
rect 554780 437242 554832 437248
rect 551744 436960 551796 436966
rect 551480 436908 551744 436914
rect 551480 436902 551796 436908
rect 551480 436886 551784 436902
rect 499316 426426 499344 427516
rect 551480 426426 551508 436886
rect 554792 436665 554820 437242
rect 554884 436966 554912 438874
rect 555160 438433 555188 474030
rect 555252 442513 555280 476274
rect 555332 474564 555384 474570
rect 555332 474506 555384 474512
rect 555344 469198 555372 474506
rect 555332 469192 555384 469198
rect 555332 469134 555384 469140
rect 555332 469056 555384 469062
rect 555332 468998 555384 469004
rect 555344 446185 555372 468998
rect 555436 450265 555464 500006
rect 555422 450256 555478 450265
rect 555422 450191 555478 450200
rect 555330 446176 555386 446185
rect 555330 446111 555386 446120
rect 555238 442504 555294 442513
rect 555238 442439 555294 442448
rect 555146 438424 555202 438433
rect 555146 438359 555202 438368
rect 555528 437889 555556 502846
rect 556172 502846 556416 502874
rect 557520 502846 557672 502874
rect 555608 474428 555660 474434
rect 555608 474370 555660 474376
rect 555620 469062 555648 474370
rect 555792 474292 555844 474298
rect 555792 474234 555844 474240
rect 555700 471980 555752 471986
rect 555700 471922 555752 471928
rect 555608 469056 555660 469062
rect 555608 468998 555660 469004
rect 555608 468920 555660 468926
rect 555608 468862 555660 468868
rect 555620 452033 555648 468862
rect 555712 458561 555740 471922
rect 555804 468926 555832 474234
rect 555884 474156 555936 474162
rect 555884 474098 555936 474104
rect 555792 468920 555844 468926
rect 555792 468862 555844 468868
rect 555896 468738 555924 474098
rect 556068 474020 556120 474026
rect 556068 473962 556120 473968
rect 555804 468710 555924 468738
rect 555804 461009 555832 468710
rect 556080 468602 556108 473962
rect 555896 468574 556108 468602
rect 555896 462097 555924 468574
rect 555882 462088 555938 462097
rect 555882 462023 555938 462032
rect 555790 461000 555846 461009
rect 555790 460935 555846 460944
rect 555698 458552 555754 458561
rect 555698 458487 555754 458496
rect 555606 452024 555662 452033
rect 555606 451959 555662 451968
rect 555514 437880 555570 437889
rect 555514 437815 555570 437824
rect 556066 437200 556122 437209
rect 556172 437186 556200 502846
rect 556804 500268 556856 500274
rect 556804 500210 556856 500216
rect 556122 437158 556200 437186
rect 556066 437135 556122 437144
rect 554872 436960 554924 436966
rect 554872 436902 554924 436908
rect 554778 436656 554834 436665
rect 554778 436591 554834 436600
rect 554780 436552 554832 436558
rect 554780 436494 554832 436500
rect 554792 436121 554820 436494
rect 554778 436112 554834 436121
rect 554778 436047 554834 436056
rect 554872 436076 554924 436082
rect 554872 436018 554924 436024
rect 554780 436008 554832 436014
rect 554780 435950 554832 435956
rect 554792 435441 554820 435950
rect 554778 435432 554834 435441
rect 554778 435367 554834 435376
rect 554884 434897 554912 436018
rect 554870 434888 554926 434897
rect 554870 434823 554926 434832
rect 554872 434716 554924 434722
rect 554872 434658 554924 434664
rect 554780 434648 554832 434654
rect 554780 434590 554832 434596
rect 554792 434217 554820 434590
rect 554778 434208 554834 434217
rect 554778 434143 554834 434152
rect 554884 433673 554912 434658
rect 554870 433664 554926 433673
rect 554870 433599 554926 433608
rect 554872 433288 554924 433294
rect 554872 433230 554924 433236
rect 554780 433220 554832 433226
rect 554780 433162 554832 433168
rect 554792 433129 554820 433162
rect 554778 433120 554834 433129
rect 554778 433055 554834 433064
rect 554884 432449 554912 433230
rect 554870 432440 554926 432449
rect 554870 432375 554926 432384
rect 554964 431928 555016 431934
rect 554778 431896 554834 431905
rect 554964 431870 555016 431876
rect 554778 431831 554780 431840
rect 554832 431831 554834 431840
rect 554780 431802 554832 431808
rect 554872 431792 554924 431798
rect 554872 431734 554924 431740
rect 554884 431361 554912 431734
rect 554870 431352 554926 431361
rect 554870 431287 554926 431296
rect 554976 430681 555004 431870
rect 554962 430672 555018 430681
rect 554962 430607 555018 430616
rect 554872 430568 554924 430574
rect 554872 430510 554924 430516
rect 554780 430500 554832 430506
rect 554780 430442 554832 430448
rect 554792 430137 554820 430442
rect 554778 430128 554834 430137
rect 554778 430063 554834 430072
rect 554884 429593 554912 430510
rect 554870 429584 554926 429593
rect 554870 429519 554926 429528
rect 554780 429140 554832 429146
rect 554780 429082 554832 429088
rect 554792 428369 554820 429082
rect 556816 428942 556844 500210
rect 556896 462392 556948 462398
rect 556896 462334 556948 462340
rect 556908 438938 556936 462334
rect 556896 438932 556948 438938
rect 556896 438874 556948 438880
rect 557644 437306 557672 502846
rect 557736 502846 558624 502874
rect 558932 502846 559636 502874
rect 560312 502846 560740 502874
rect 557632 437300 557684 437306
rect 557632 437242 557684 437248
rect 557736 436558 557764 502846
rect 558552 467832 558604 467838
rect 558552 467774 558604 467780
rect 558564 462398 558592 467774
rect 558552 462392 558604 462398
rect 558552 462334 558604 462340
rect 557724 436552 557776 436558
rect 557724 436494 557776 436500
rect 558932 436014 558960 502846
rect 559564 479528 559616 479534
rect 559564 479470 559616 479476
rect 559576 467838 559604 479470
rect 559564 467832 559616 467838
rect 559564 467774 559616 467780
rect 560312 436082 560340 502846
rect 561830 502602 561858 502860
rect 561784 502574 561858 502602
rect 562612 502846 562948 502874
rect 563072 502846 563960 502874
rect 564452 502846 565064 502874
rect 565832 502846 566168 502874
rect 567180 502846 567240 502874
rect 561680 501220 561732 501226
rect 561680 501162 561732 501168
rect 560944 499588 560996 499594
rect 560944 499530 560996 499536
rect 560392 482860 560444 482866
rect 560392 482802 560444 482808
rect 560404 479534 560432 482802
rect 560392 479528 560444 479534
rect 560392 479470 560444 479476
rect 560300 436076 560352 436082
rect 560300 436018 560352 436024
rect 558920 436008 558972 436014
rect 558920 435950 558972 435956
rect 560956 431798 560984 499530
rect 561692 434722 561720 501162
rect 561680 434716 561732 434722
rect 561680 434658 561732 434664
rect 561784 434654 561812 502574
rect 562612 501226 562640 502846
rect 562600 501220 562652 501226
rect 562600 501162 562652 501168
rect 561772 434648 561824 434654
rect 561772 434590 561824 434596
rect 563072 433226 563100 502846
rect 563704 493332 563756 493338
rect 563704 493274 563756 493280
rect 563716 482866 563744 493274
rect 563704 482860 563756 482866
rect 563704 482802 563756 482808
rect 563704 462392 563756 462398
rect 563704 462334 563756 462340
rect 563060 433220 563112 433226
rect 563060 433162 563112 433168
rect 560944 431792 560996 431798
rect 560944 431734 560996 431740
rect 554872 428936 554924 428942
rect 554870 428904 554872 428913
rect 556804 428936 556856 428942
rect 554924 428904 554926 428913
rect 556804 428878 556856 428884
rect 554870 428839 554926 428848
rect 554778 428360 554834 428369
rect 554778 428295 554834 428304
rect 554778 427816 554834 427825
rect 554778 427751 554780 427760
rect 554832 427751 554834 427760
rect 554780 427722 554832 427728
rect 447784 426420 447836 426426
rect 447784 426362 447836 426368
rect 499304 426420 499356 426426
rect 499304 426362 499356 426368
rect 551468 426420 551520 426426
rect 551468 426362 551520 426368
rect 417424 327072 417476 327078
rect 417424 327014 417476 327020
rect 563716 325650 563744 462334
rect 564452 433294 564480 502846
rect 564440 433288 564492 433294
rect 564440 433230 564492 433236
rect 565832 431866 565860 502846
rect 567212 499594 567240 502846
rect 567304 502846 568284 502874
rect 568592 502846 569388 502874
rect 569972 502846 570492 502874
rect 571352 502846 571504 502874
rect 571628 502846 572608 502874
rect 572732 502846 573712 502874
rect 567200 499588 567252 499594
rect 567200 499530 567252 499536
rect 567304 431934 567332 502846
rect 567292 431928 567344 431934
rect 567292 431870 567344 431876
rect 565820 431860 565872 431866
rect 565820 431802 565872 431808
rect 568592 430506 568620 502846
rect 569972 430574 570000 502846
rect 571352 500274 571380 502846
rect 571340 500268 571392 500274
rect 571340 500210 571392 500216
rect 571340 495508 571392 495514
rect 571340 495450 571392 495456
rect 571352 493338 571380 495450
rect 571340 493332 571392 493338
rect 571340 493274 571392 493280
rect 569960 430568 570012 430574
rect 569960 430510 570012 430516
rect 568580 430500 568632 430506
rect 568580 430442 568632 430448
rect 571628 429146 571656 502846
rect 571616 429140 571668 429146
rect 571616 429082 571668 429088
rect 572732 427786 572760 502846
rect 573454 502752 573510 502761
rect 573454 502687 573510 502696
rect 573364 502376 573416 502382
rect 573364 502318 573416 502324
rect 572720 427780 572772 427786
rect 572720 427722 572772 427728
rect 563704 325644 563756 325650
rect 563704 325586 563756 325592
rect 560944 306400 560996 306406
rect 560944 306342 560996 306348
rect 412088 83564 412140 83570
rect 412088 83506 412140 83512
rect 487620 62824 487672 62830
rect 487620 62766 487672 62772
rect 487632 60860 487660 62766
rect 411994 49872 412050 49881
rect 411994 49807 412050 49816
rect 560956 41410 560984 306342
rect 573376 62830 573404 502318
rect 573468 495514 573496 502687
rect 574020 502382 574048 502998
rect 574112 502846 574724 502874
rect 574008 502376 574060 502382
rect 574008 502318 574060 502324
rect 574112 498846 574140 502846
rect 574100 498840 574152 498846
rect 574100 498782 574152 498788
rect 573456 495508 573508 495514
rect 573456 495450 573508 495456
rect 576136 95198 576164 696934
rect 580354 686352 580410 686361
rect 580354 686287 580410 686296
rect 579618 651128 579674 651137
rect 579618 651063 579674 651072
rect 579632 650078 579660 651063
rect 577504 650072 577556 650078
rect 577504 650014 577556 650020
rect 579620 650072 579672 650078
rect 579620 650014 579672 650020
rect 576124 95192 576176 95198
rect 576124 95134 576176 95140
rect 577516 93770 577544 650014
rect 580262 639432 580318 639441
rect 580262 639367 580318 639376
rect 578882 604208 578938 604217
rect 578882 604143 578938 604152
rect 578896 93838 578924 604143
rect 579802 557288 579858 557297
rect 579802 557223 579858 557232
rect 579816 556238 579844 557223
rect 579804 556232 579856 556238
rect 579804 556174 579856 556180
rect 580170 463448 580226 463457
rect 580170 463383 580226 463392
rect 580184 462398 580212 463383
rect 580172 462392 580224 462398
rect 580172 462334 580224 462340
rect 580170 416528 580226 416537
rect 580170 416463 580226 416472
rect 580184 415478 580212 416463
rect 580172 415472 580224 415478
rect 580172 415414 580224 415420
rect 580170 369608 580226 369617
rect 580170 369543 580226 369552
rect 580184 368558 580212 369543
rect 580172 368552 580224 368558
rect 580172 368494 580224 368500
rect 580170 322688 580226 322697
rect 580170 322623 580226 322632
rect 580184 321638 580212 322623
rect 580172 321632 580224 321638
rect 580172 321574 580224 321580
rect 580172 276004 580224 276010
rect 580172 275946 580224 275952
rect 580184 275777 580212 275946
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 579988 229084 580040 229090
rect 579988 229026 580040 229032
rect 580000 228857 580028 229026
rect 579986 228848 580042 228857
rect 579986 228783 580042 228792
rect 579988 182164 580040 182170
rect 579988 182106 580040 182112
rect 580000 181937 580028 182106
rect 579986 181928 580042 181937
rect 579986 181863 580042 181872
rect 580172 135244 580224 135250
rect 580172 135186 580224 135192
rect 580184 134881 580212 135186
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 578884 93832 578936 93838
rect 578884 93774 578936 93780
rect 577504 93764 577556 93770
rect 577504 93706 577556 93712
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 87961 580212 88266
rect 580170 87952 580226 87961
rect 580170 87887 580226 87896
rect 580276 83502 580304 639367
rect 580368 502994 580396 686287
rect 580538 592512 580594 592521
rect 580538 592447 580594 592456
rect 580446 580816 580502 580825
rect 580446 580751 580502 580760
rect 580460 503062 580488 580751
rect 580552 569226 580580 592447
rect 580540 569220 580592 569226
rect 580540 569162 580592 569168
rect 580906 545592 580962 545601
rect 580906 545527 580962 545536
rect 580538 510368 580594 510377
rect 580538 510303 580594 510312
rect 580448 503056 580500 503062
rect 580448 502998 580500 503004
rect 580356 502988 580408 502994
rect 580356 502930 580408 502936
rect 580552 501634 580580 510303
rect 580540 501628 580592 501634
rect 580540 501570 580592 501576
rect 580920 498681 580948 545527
rect 580906 498672 580962 498681
rect 580906 498607 580962 498616
rect 580920 451761 580948 498607
rect 580906 451752 580962 451761
rect 580906 451687 580962 451696
rect 580920 404841 580948 451687
rect 580906 404832 580962 404841
rect 580906 404767 580962 404776
rect 580920 357921 580948 404767
rect 580906 357912 580962 357921
rect 580906 357847 580962 357856
rect 580920 310865 580948 357847
rect 580354 310856 580410 310865
rect 580354 310791 580410 310800
rect 580906 310856 580962 310865
rect 580906 310791 580962 310800
rect 580368 303618 580396 310791
rect 580356 303612 580408 303618
rect 580356 303554 580408 303560
rect 580368 263945 580396 303554
rect 580354 263936 580410 263945
rect 580354 263871 580410 263880
rect 580906 263936 580962 263945
rect 580906 263871 580962 263880
rect 580920 217025 580948 263871
rect 580906 217016 580962 217025
rect 580906 216951 580962 216960
rect 580920 170105 580948 216951
rect 580906 170096 580962 170105
rect 580906 170031 580962 170040
rect 580920 123185 580948 170031
rect 580906 123176 580962 123185
rect 580906 123111 580962 123120
rect 580264 83496 580316 83502
rect 580264 83438 580316 83444
rect 580920 76265 580948 123111
rect 580906 76256 580962 76265
rect 580906 76191 580962 76200
rect 573364 62824 573416 62830
rect 573364 62766 573416 62772
rect 560944 41404 560996 41410
rect 560944 41346 560996 41352
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 563702 38720 563758 38729
rect 563702 38655 563758 38664
rect 411902 27568 411958 27577
rect 411902 27503 411958 27512
rect 208688 26710 208808 26738
rect 208688 19310 208716 26710
rect 208492 19304 208544 19310
rect 208492 19246 208544 19252
rect 208676 19304 208728 19310
rect 208676 19246 208728 19252
rect 208504 9722 208532 19246
rect 406476 18012 406528 18018
rect 406476 17954 406528 17960
rect 287060 17400 287112 17406
rect 270512 17338 270632 17354
rect 287060 17342 287112 17348
rect 296536 17400 296588 17406
rect 296536 17342 296588 17348
rect 393964 17400 394016 17406
rect 393964 17342 394016 17348
rect 246948 17332 247000 17338
rect 246948 17274 247000 17280
rect 270500 17332 270632 17338
rect 270552 17326 270632 17332
rect 270500 17274 270552 17280
rect 217968 17060 218020 17066
rect 217968 17002 218020 17008
rect 215206 13424 215262 13433
rect 215206 13359 215262 13368
rect 208492 9716 208544 9722
rect 208492 9658 208544 9664
rect 208768 9716 208820 9722
rect 208768 9658 208820 9664
rect 207020 4684 207072 4690
rect 207020 4626 207072 4632
rect 208780 4622 208808 9658
rect 211066 7984 211122 7993
rect 211066 7919 211122 7928
rect 208768 4616 208820 4622
rect 208768 4558 208820 4564
rect 208676 3936 208728 3942
rect 208676 3878 208728 3884
rect 207480 3664 207532 3670
rect 207480 3606 207532 3612
rect 207492 480 207520 3606
rect 208688 480 208716 3878
rect 209872 3868 209924 3874
rect 209872 3810 209924 3816
rect 209884 480 209912 3810
rect 211080 480 211108 7919
rect 212262 4856 212318 4865
rect 212262 4791 212318 4800
rect 212276 480 212304 4791
rect 215220 4146 215248 13359
rect 215852 4956 215904 4962
rect 215852 4898 215904 4904
rect 214656 4140 214708 4146
rect 214656 4082 214708 4088
rect 215208 4140 215260 4146
rect 215208 4082 215260 4088
rect 213472 598 213684 626
rect 213472 480 213500 598
rect 199384 264 199436 270
rect 199384 206 199436 212
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 213656 338 213684 598
rect 214668 480 214696 4082
rect 215864 480 215892 4898
rect 217980 3398 218008 17002
rect 246302 15464 246358 15473
rect 246302 15399 246358 15408
rect 234528 15360 234580 15366
rect 234528 15302 234580 15308
rect 226248 13388 226300 13394
rect 226248 13330 226300 13336
rect 220728 10396 220780 10402
rect 220728 10338 220780 10344
rect 218152 9512 218204 9518
rect 218152 9454 218204 9460
rect 217048 3392 217100 3398
rect 217048 3334 217100 3340
rect 217968 3392 218020 3398
rect 217968 3334 218020 3340
rect 217060 480 217088 3334
rect 218164 480 218192 9454
rect 219348 5024 219400 5030
rect 219348 4966 219400 4972
rect 219360 480 219388 4966
rect 220740 610 220768 10338
rect 224866 10296 224922 10305
rect 224866 10231 224922 10240
rect 221740 6248 221792 6254
rect 221740 6190 221792 6196
rect 220544 604 220596 610
rect 220544 546 220596 552
rect 220728 604 220780 610
rect 220728 546 220780 552
rect 220556 480 220584 546
rect 221752 480 221780 6190
rect 222934 4992 222990 5001
rect 222934 4927 222990 4936
rect 222948 480 222976 4927
rect 224880 3398 224908 10231
rect 226260 3398 226288 13330
rect 231768 10532 231820 10538
rect 231768 10474 231820 10480
rect 229008 10464 229060 10470
rect 229008 10406 229060 10412
rect 228916 9580 228968 9586
rect 228916 9522 228968 9528
rect 226524 5092 226576 5098
rect 226524 5034 226576 5040
rect 224132 3392 224184 3398
rect 224132 3334 224184 3340
rect 224868 3392 224920 3398
rect 224868 3334 224920 3340
rect 225328 3392 225380 3398
rect 225328 3334 225380 3340
rect 226248 3392 226300 3398
rect 226248 3334 226300 3340
rect 224144 480 224172 3334
rect 225340 480 225368 3334
rect 226536 480 226564 5034
rect 227720 3392 227772 3398
rect 227720 3334 227772 3340
rect 227732 480 227760 3334
rect 228928 480 228956 9522
rect 229020 3398 229048 10406
rect 230112 5160 230164 5166
rect 230112 5102 230164 5108
rect 229008 3392 229060 3398
rect 229008 3334 229060 3340
rect 230124 480 230152 5102
rect 231780 3398 231808 10474
rect 232502 8120 232558 8129
rect 232502 8055 232558 8064
rect 231308 3392 231360 3398
rect 231308 3334 231360 3340
rect 231768 3392 231820 3398
rect 231768 3334 231820 3340
rect 231320 480 231348 3334
rect 232516 480 232544 8055
rect 234540 3398 234568 15302
rect 244186 11928 244242 11937
rect 244186 11863 244242 11872
rect 240048 10668 240100 10674
rect 240048 10610 240100 10616
rect 235908 10600 235960 10606
rect 235908 10542 235960 10548
rect 235920 3398 235948 10542
rect 238666 10432 238722 10441
rect 238666 10367 238722 10376
rect 236000 5228 236052 5234
rect 236000 5170 236052 5176
rect 233700 3392 233752 3398
rect 233700 3334 233752 3340
rect 234528 3392 234580 3398
rect 234528 3334 234580 3340
rect 234804 3392 234856 3398
rect 234804 3334 234856 3340
rect 235908 3392 235960 3398
rect 235908 3334 235960 3340
rect 233712 480 233740 3334
rect 234816 480 234844 3334
rect 236012 480 236040 5170
rect 238680 3482 238708 10367
rect 238404 3454 238708 3482
rect 237196 2372 237248 2378
rect 237196 2314 237248 2320
rect 237208 480 237236 2314
rect 238404 480 238432 3454
rect 240060 3398 240088 10610
rect 242806 10568 242862 10577
rect 242806 10503 242862 10512
rect 242820 3398 242848 10503
rect 244200 3398 244228 11863
rect 245568 10736 245620 10742
rect 245568 10678 245620 10684
rect 239588 3392 239640 3398
rect 239588 3334 239640 3340
rect 240048 3392 240100 3398
rect 240048 3334 240100 3340
rect 241980 3392 242032 3398
rect 241980 3334 242032 3340
rect 242808 3392 242860 3398
rect 242808 3334 242860 3340
rect 243176 3392 243228 3398
rect 243176 3334 243228 3340
rect 244188 3392 244240 3398
rect 244188 3334 244240 3340
rect 239600 480 239628 3334
rect 240784 3188 240836 3194
rect 240784 3130 240836 3136
rect 240796 480 240824 3130
rect 241992 480 242020 3334
rect 243188 480 243216 3334
rect 244372 2440 244424 2446
rect 244372 2382 244424 2388
rect 244384 480 244412 2382
rect 245580 480 245608 10678
rect 246316 3806 246344 15399
rect 246304 3800 246356 3806
rect 246304 3742 246356 3748
rect 246960 3482 246988 17274
rect 267648 17196 267700 17202
rect 267648 17138 267700 17144
rect 250442 15600 250498 15609
rect 250442 15535 250498 15544
rect 248328 15428 248380 15434
rect 248328 15370 248380 15376
rect 248340 3482 248368 15370
rect 249708 10804 249760 10810
rect 249708 10746 249760 10752
rect 246776 3454 246988 3482
rect 247972 3454 248368 3482
rect 246776 480 246804 3454
rect 247972 480 248000 3454
rect 249720 3398 249748 10746
rect 250456 4010 250484 15535
rect 259368 15496 259420 15502
rect 259368 15438 259420 15444
rect 250536 14680 250588 14686
rect 250536 14622 250588 14628
rect 250548 6322 250576 14622
rect 253848 10872 253900 10878
rect 253848 10814 253900 10820
rect 253756 9648 253808 9654
rect 253756 9590 253808 9596
rect 250536 6316 250588 6322
rect 250536 6258 250588 6264
rect 250444 4004 250496 4010
rect 250444 3946 250496 3952
rect 250536 4004 250588 4010
rect 250536 3946 250588 3952
rect 249156 3392 249208 3398
rect 249156 3334 249208 3340
rect 249708 3392 249760 3398
rect 249708 3334 249760 3340
rect 249168 480 249196 3334
rect 250548 1986 250576 3946
rect 252652 3800 252704 3806
rect 252652 3742 252704 3748
rect 251456 2984 251508 2990
rect 251456 2926 251508 2932
rect 250364 1958 250576 1986
rect 250364 480 250392 1958
rect 251468 480 251496 2926
rect 252664 480 252692 3742
rect 253768 3482 253796 9590
rect 253860 3806 253888 10814
rect 256240 5364 256292 5370
rect 256240 5306 256292 5312
rect 255044 5296 255096 5302
rect 255044 5238 255096 5244
rect 253848 3800 253900 3806
rect 253848 3742 253900 3748
rect 253768 3454 253888 3482
rect 253860 480 253888 3454
rect 255056 480 255084 5238
rect 256252 480 256280 5306
rect 258448 4004 258500 4010
rect 258448 3946 258500 3952
rect 258540 4004 258592 4010
rect 258540 3946 258592 3952
rect 258460 3806 258488 3946
rect 258448 3800 258500 3806
rect 258448 3742 258500 3748
rect 258552 3602 258580 3946
rect 259380 3602 259408 15438
rect 263508 10940 263560 10946
rect 263508 10882 263560 10888
rect 261024 6316 261076 6322
rect 261024 6258 261076 6264
rect 258540 3596 258592 3602
rect 258540 3538 258592 3544
rect 258632 3596 258684 3602
rect 258632 3538 258684 3544
rect 259368 3596 259420 3602
rect 259368 3538 259420 3544
rect 257436 3324 257488 3330
rect 257436 3266 257488 3272
rect 256700 2916 256752 2922
rect 256700 2858 256752 2864
rect 256712 2689 256740 2858
rect 256698 2680 256754 2689
rect 256698 2615 256754 2624
rect 257448 480 257476 3266
rect 258644 480 258672 3538
rect 259828 604 259880 610
rect 259828 546 259880 552
rect 259840 480 259868 546
rect 261036 480 261064 6258
rect 263520 3482 263548 10882
rect 263600 5500 263652 5506
rect 263600 5442 263652 5448
rect 263612 4010 263640 5442
rect 263600 4004 263652 4010
rect 263600 3946 263652 3952
rect 267660 3602 267688 17138
rect 270604 17134 270632 17326
rect 278688 17264 278740 17270
rect 278688 17206 278740 17212
rect 270592 17128 270644 17134
rect 270592 17070 270644 17076
rect 275284 15632 275336 15638
rect 275284 15574 275336 15580
rect 269028 13456 269080 13462
rect 269028 13398 269080 13404
rect 267740 4004 267792 4010
rect 267740 3946 267792 3952
rect 267752 3806 267780 3946
rect 267740 3800 267792 3806
rect 267740 3742 267792 3748
rect 269040 3602 269068 13398
rect 273166 9208 273222 9217
rect 273166 9143 273222 9152
rect 272890 6488 272946 6497
rect 272890 6423 272946 6432
rect 269304 6384 269356 6390
rect 269304 6326 269356 6332
rect 267004 3596 267056 3602
rect 267004 3538 267056 3544
rect 267648 3596 267700 3602
rect 267648 3538 267700 3544
rect 268108 3596 268160 3602
rect 268108 3538 268160 3544
rect 269028 3596 269080 3602
rect 269028 3538 269080 3544
rect 263428 3454 263548 3482
rect 262220 2848 262272 2854
rect 262220 2790 262272 2796
rect 262232 480 262260 2790
rect 263428 480 263456 3454
rect 264612 3392 264664 3398
rect 264612 3334 264664 3340
rect 263600 3052 263652 3058
rect 263600 2994 263652 3000
rect 263612 1698 263640 2994
rect 263600 1692 263652 1698
rect 263600 1634 263652 1640
rect 264624 480 264652 3334
rect 265808 604 265860 610
rect 265808 546 265860 552
rect 265820 480 265848 546
rect 267016 480 267044 3538
rect 268120 480 268148 3538
rect 269316 480 269344 6326
rect 271696 4140 271748 4146
rect 271696 4082 271748 4088
rect 270500 604 270552 610
rect 270500 546 270552 552
rect 270512 480 270540 546
rect 271708 480 271736 4082
rect 272904 480 272932 6423
rect 273180 3738 273208 9143
rect 275296 4078 275324 15574
rect 276480 6452 276532 6458
rect 276480 6394 276532 6400
rect 275284 4072 275336 4078
rect 275284 4014 275336 4020
rect 273168 3732 273220 3738
rect 273168 3674 273220 3680
rect 275282 3496 275338 3505
rect 275282 3431 275338 3440
rect 274088 2508 274140 2514
rect 274088 2450 274140 2456
rect 274100 480 274128 2450
rect 275296 480 275324 3431
rect 276492 480 276520 6394
rect 278700 4078 278728 17206
rect 287072 17134 287100 17342
rect 296548 17134 296576 17342
rect 300768 17332 300820 17338
rect 300768 17274 300820 17280
rect 287060 17128 287112 17134
rect 287060 17070 287112 17076
rect 296536 17128 296588 17134
rect 296536 17070 296588 17076
rect 282184 15700 282236 15706
rect 282184 15642 282236 15648
rect 280068 15564 280120 15570
rect 280068 15506 280120 15512
rect 279976 6520 280028 6526
rect 279976 6462 280028 6468
rect 277676 4072 277728 4078
rect 277676 4014 277728 4020
rect 278688 4072 278740 4078
rect 278688 4014 278740 4020
rect 278872 4072 278924 4078
rect 278872 4014 278924 4020
rect 277688 480 277716 4014
rect 278884 480 278912 4014
rect 279988 3890 280016 6462
rect 280080 4078 280108 15506
rect 281264 11008 281316 11014
rect 281264 10950 281316 10956
rect 280068 4072 280120 4078
rect 280068 4014 280120 4020
rect 279988 3862 280108 3890
rect 280080 480 280108 3862
rect 281276 480 281304 10950
rect 282196 3262 282224 15642
rect 293868 13728 293920 13734
rect 293868 13670 293920 13676
rect 291936 11960 291988 11966
rect 291936 11902 291988 11908
rect 288348 11892 288400 11898
rect 288348 11834 288400 11840
rect 284760 11824 284812 11830
rect 284760 11766 284812 11772
rect 283656 6588 283708 6594
rect 283656 6530 283708 6536
rect 282736 4004 282788 4010
rect 282736 3946 282788 3952
rect 282748 3602 282776 3946
rect 282828 3936 282880 3942
rect 282920 3936 282972 3942
rect 282880 3896 282920 3924
rect 282828 3878 282880 3884
rect 282920 3878 282972 3884
rect 282736 3596 282788 3602
rect 282736 3538 282788 3544
rect 282458 3360 282514 3369
rect 282458 3295 282514 3304
rect 282184 3256 282236 3262
rect 282184 3198 282236 3204
rect 282472 480 282500 3295
rect 283668 480 283696 6530
rect 284772 480 284800 11766
rect 285956 7676 286008 7682
rect 285956 7618 286008 7624
rect 285968 480 285996 7618
rect 287152 6656 287204 6662
rect 287152 6598 287204 6604
rect 287164 480 287192 6598
rect 288360 480 288388 11834
rect 290740 6724 290792 6730
rect 290740 6666 290792 6672
rect 289818 5264 289874 5273
rect 289818 5199 289874 5208
rect 289832 3942 289860 5199
rect 289820 3936 289872 3942
rect 289820 3878 289872 3884
rect 289728 3664 289780 3670
rect 289542 3632 289598 3641
rect 289912 3664 289964 3670
rect 289780 3612 289912 3618
rect 289728 3606 289964 3612
rect 289542 3567 289598 3576
rect 289636 3596 289688 3602
rect 289556 480 289584 3567
rect 289740 3590 289952 3606
rect 289636 3538 289688 3544
rect 289648 3262 289676 3538
rect 289636 3256 289688 3262
rect 289636 3198 289688 3204
rect 290752 480 290780 6666
rect 291948 480 291976 11902
rect 293880 4078 293908 13670
rect 299112 12164 299164 12170
rect 299112 12106 299164 12112
rect 295524 12028 295576 12034
rect 295524 11970 295576 11976
rect 294328 6792 294380 6798
rect 294328 6734 294380 6740
rect 293132 4072 293184 4078
rect 293132 4014 293184 4020
rect 293868 4072 293920 4078
rect 293868 4014 293920 4020
rect 293144 480 293172 4014
rect 294340 480 294368 6734
rect 295536 480 295564 11970
rect 297916 6860 297968 6866
rect 297916 6802 297968 6808
rect 296718 3768 296774 3777
rect 296718 3703 296774 3712
rect 296732 480 296760 3703
rect 297928 480 297956 6802
rect 298020 3602 298140 3618
rect 298020 3596 298152 3602
rect 298020 3590 298100 3596
rect 298020 3262 298048 3590
rect 298100 3538 298152 3544
rect 298008 3256 298060 3262
rect 298008 3198 298060 3204
rect 299124 480 299152 12106
rect 300780 4078 300808 17274
rect 393976 17202 394004 17342
rect 393964 17196 394016 17202
rect 393964 17138 394016 17144
rect 406488 16969 406516 17954
rect 414388 17672 414440 17678
rect 414388 17614 414440 17620
rect 414296 17468 414348 17474
rect 414296 17410 414348 17416
rect 410524 17400 410576 17406
rect 410616 17400 410668 17406
rect 410576 17348 410616 17354
rect 410524 17342 410668 17348
rect 410536 17326 410656 17342
rect 414308 17270 414336 17410
rect 414400 17338 414428 17614
rect 414388 17332 414440 17338
rect 414388 17274 414440 17280
rect 414296 17264 414348 17270
rect 414296 17206 414348 17212
rect 459112 17066 459402 17082
rect 462608 17066 462898 17082
rect 470060 17066 470166 17082
rect 424600 17060 424652 17066
rect 424600 17002 424652 17008
rect 439412 17060 439464 17066
rect 439412 17002 439464 17008
rect 459100 17060 459402 17066
rect 459152 17054 459402 17060
rect 462596 17060 462898 17066
rect 459100 17002 459152 17008
rect 462648 17054 462898 17060
rect 470048 17060 470166 17066
rect 462596 17002 462648 17008
rect 470100 17054 470166 17060
rect 470048 17002 470100 17008
rect 418712 16992 418764 16998
rect 406474 16960 406530 16969
rect 406474 16895 406530 16904
rect 414662 16960 414718 16969
rect 414718 16918 414966 16946
rect 424612 16969 424640 17002
rect 425612 16992 425664 16998
rect 418712 16934 418764 16940
rect 424598 16960 424654 16969
rect 414662 16895 414718 16904
rect 415412 16658 415702 16674
rect 418724 16658 418752 16934
rect 439424 16969 439452 17002
rect 425612 16934 425664 16940
rect 435362 16960 435418 16969
rect 424598 16895 424654 16904
rect 424232 16720 424284 16726
rect 424284 16668 424534 16674
rect 424232 16662 424534 16668
rect 415400 16652 415702 16658
rect 415452 16646 415702 16652
rect 418712 16652 418764 16658
rect 415400 16594 415452 16600
rect 424244 16646 424534 16662
rect 425624 16658 425652 16934
rect 430028 16924 430080 16930
rect 435362 16895 435418 16904
rect 439410 16960 439466 16969
rect 439410 16895 439466 16904
rect 452566 16960 452622 16969
rect 452622 16918 452870 16946
rect 452566 16895 452622 16904
rect 430028 16866 430080 16872
rect 429936 16856 429988 16862
rect 425808 16794 426098 16810
rect 429936 16798 429988 16804
rect 425796 16788 426098 16794
rect 425848 16782 426098 16788
rect 425796 16730 425848 16736
rect 429948 16658 429976 16798
rect 425612 16652 425664 16658
rect 418712 16594 418764 16600
rect 425612 16594 425664 16600
rect 429936 16652 429988 16658
rect 429936 16594 429988 16600
rect 430040 16590 430068 16866
rect 435376 16794 435404 16895
rect 435364 16788 435416 16794
rect 435364 16730 435416 16736
rect 443000 16788 443052 16794
rect 443000 16730 443052 16736
rect 438400 16720 438452 16726
rect 432708 16658 432998 16674
rect 443012 16674 443040 16730
rect 438452 16668 438702 16674
rect 438400 16662 438702 16668
rect 432696 16652 432998 16658
rect 432748 16646 432998 16652
rect 438412 16646 438702 16662
rect 443012 16646 443302 16674
rect 432696 16594 432748 16600
rect 430028 16584 430080 16590
rect 430028 16526 430080 16532
rect 434996 16584 435048 16590
rect 435048 16532 435298 16538
rect 434996 16526 435298 16532
rect 435008 16510 435298 16526
rect 479812 16510 480102 16538
rect 535012 16510 535302 16538
rect 479812 16454 479840 16510
rect 535012 16454 535040 16510
rect 479064 16448 479116 16454
rect 387708 16108 387760 16114
rect 387708 16050 387760 16056
rect 376208 16040 376260 16046
rect 376208 15982 376260 15988
rect 311164 15972 311216 15978
rect 311164 15914 311216 15920
rect 307206 14920 307262 14929
rect 307206 14855 307262 14864
rect 306196 12232 306248 12238
rect 306196 12174 306248 12180
rect 302608 12164 302660 12170
rect 302608 12106 302660 12112
rect 301412 6112 301464 6118
rect 301412 6054 301464 6060
rect 300308 4072 300360 4078
rect 300308 4014 300360 4020
rect 300768 4072 300820 4078
rect 300768 4014 300820 4020
rect 300320 480 300348 4014
rect 300768 2984 300820 2990
rect 300768 2926 300820 2932
rect 300780 2718 300808 2926
rect 300768 2712 300820 2718
rect 300768 2654 300820 2660
rect 301424 480 301452 6054
rect 302620 480 302648 12106
rect 303804 5432 303856 5438
rect 303804 5374 303856 5380
rect 303816 480 303844 5374
rect 305000 4004 305052 4010
rect 305000 3946 305052 3952
rect 305012 480 305040 3946
rect 306208 480 306236 12174
rect 307220 8362 307248 14855
rect 307758 9344 307814 9353
rect 307758 9279 307814 9288
rect 307208 8356 307260 8362
rect 307208 8298 307260 8304
rect 307392 8356 307444 8362
rect 307392 8298 307444 8304
rect 307404 8242 307432 8298
rect 307312 8214 307432 8242
rect 307312 610 307340 8214
rect 307772 3874 307800 9279
rect 309784 3936 309836 3942
rect 309784 3878 309836 3884
rect 307760 3868 307812 3874
rect 307760 3810 307812 3816
rect 307668 3800 307720 3806
rect 307668 3742 307720 3748
rect 307680 3602 307708 3742
rect 307668 3596 307720 3602
rect 307668 3538 307720 3544
rect 308588 2576 308640 2582
rect 308588 2518 308640 2524
rect 307300 604 307352 610
rect 307300 546 307352 552
rect 307392 604 307444 610
rect 307392 546 307444 552
rect 307404 480 307432 546
rect 308600 480 308628 2518
rect 309796 480 309824 3878
rect 310980 3256 311032 3262
rect 310980 3198 311032 3204
rect 310992 480 311020 3198
rect 311176 3194 311204 15914
rect 339408 15904 339460 15910
rect 339408 15846 339460 15852
rect 326344 15836 326396 15842
rect 326344 15778 326396 15784
rect 314568 14748 314620 14754
rect 314568 14690 314620 14696
rect 313372 12368 313424 12374
rect 313372 12310 313424 12316
rect 311164 3188 311216 3194
rect 311164 3130 311216 3136
rect 312176 604 312228 610
rect 312176 546 312228 552
rect 312188 480 312216 546
rect 313384 480 313412 12310
rect 313924 4072 313976 4078
rect 313924 4014 313976 4020
rect 313936 3806 313964 4014
rect 313924 3800 313976 3806
rect 313924 3742 313976 3748
rect 314580 480 314608 14690
rect 320088 13660 320140 13666
rect 320088 13602 320140 13608
rect 316960 12368 317012 12374
rect 316960 12310 317012 12316
rect 316684 12300 316736 12306
rect 316684 12242 316736 12248
rect 316696 11626 316724 12242
rect 316684 11620 316736 11626
rect 316684 11562 316736 11568
rect 316592 3596 316644 3602
rect 316592 3538 316644 3544
rect 316604 3262 316632 3538
rect 316592 3256 316644 3262
rect 316592 3198 316644 3204
rect 315764 672 315816 678
rect 315764 614 315816 620
rect 315776 480 315804 614
rect 316972 480 317000 12310
rect 318064 3868 318116 3874
rect 318064 3810 318116 3816
rect 318076 480 318104 3810
rect 320100 2990 320128 13602
rect 320456 12436 320508 12442
rect 320456 12378 320508 12384
rect 319260 2984 319312 2990
rect 319260 2926 319312 2932
rect 320088 2984 320140 2990
rect 320088 2926 320140 2932
rect 318708 2848 318760 2854
rect 318708 2790 318760 2796
rect 318720 1970 318748 2790
rect 318708 1964 318760 1970
rect 318708 1906 318760 1912
rect 319272 480 319300 2926
rect 320468 480 320496 12378
rect 325608 12096 325660 12102
rect 325608 12038 325660 12044
rect 324228 11688 324280 11694
rect 324228 11630 324280 11636
rect 322848 10260 322900 10266
rect 322848 10202 322900 10208
rect 322860 3738 322888 10202
rect 323032 4072 323084 4078
rect 323032 4014 323084 4020
rect 323044 3874 323072 4014
rect 323032 3868 323084 3874
rect 323032 3810 323084 3816
rect 321652 3732 321704 3738
rect 321652 3674 321704 3680
rect 322848 3732 322900 3738
rect 322848 3674 322900 3680
rect 321664 480 321692 3674
rect 324240 3482 324268 11630
rect 325620 11626 325648 12038
rect 325608 11620 325660 11626
rect 325608 11562 325660 11568
rect 325240 4072 325292 4078
rect 325240 4014 325292 4020
rect 324056 3454 324268 3482
rect 322848 740 322900 746
rect 322848 682 322900 688
rect 322860 480 322888 682
rect 324056 480 324084 3454
rect 325252 480 325280 4014
rect 326356 4010 326384 15778
rect 333244 15768 333296 15774
rect 333244 15710 333296 15716
rect 329748 14816 329800 14822
rect 329748 14758 329800 14764
rect 327632 6044 327684 6050
rect 327632 5986 327684 5992
rect 326344 4004 326396 4010
rect 326344 3946 326396 3952
rect 326436 808 326488 814
rect 326436 750 326488 756
rect 326448 480 326476 750
rect 327644 480 327672 5986
rect 329760 3262 329788 14758
rect 331220 4752 331272 4758
rect 331220 4694 331272 4700
rect 328828 3256 328880 3262
rect 328828 3198 328880 3204
rect 329748 3256 329800 3262
rect 329748 3198 329800 3204
rect 330024 3256 330076 3262
rect 330024 3198 330076 3204
rect 328840 480 328868 3198
rect 330036 480 330064 3198
rect 331232 480 331260 4694
rect 332416 3868 332468 3874
rect 332416 3810 332468 3816
rect 332428 480 332456 3810
rect 333256 3262 333284 15710
rect 335360 12096 335412 12102
rect 335360 12038 335412 12044
rect 335372 11626 335400 12038
rect 335360 11620 335412 11626
rect 335360 11562 335412 11568
rect 336004 11552 336056 11558
rect 336004 11494 336056 11500
rect 334716 8900 334768 8906
rect 334716 8842 334768 8848
rect 333244 3256 333296 3262
rect 333244 3198 333296 3204
rect 333612 2644 333664 2650
rect 333612 2586 333664 2592
rect 333624 480 333652 2586
rect 334728 480 334756 8842
rect 336016 4010 336044 11494
rect 338028 9988 338080 9994
rect 338028 9930 338080 9936
rect 336004 4004 336056 4010
rect 336004 3946 336056 3952
rect 335268 3936 335320 3942
rect 335268 3878 335320 3884
rect 337752 3936 337804 3942
rect 337752 3878 337804 3884
rect 335280 3806 335308 3878
rect 335268 3800 335320 3806
rect 335268 3742 335320 3748
rect 337764 3670 337792 3878
rect 337752 3664 337804 3670
rect 337752 3606 337804 3612
rect 335912 3256 335964 3262
rect 335912 3198 335964 3204
rect 335924 480 335952 3198
rect 338040 3058 338068 9930
rect 339420 3670 339448 15846
rect 368664 15156 368716 15162
rect 368664 15098 368716 15104
rect 368388 15020 368440 15026
rect 368388 14962 368440 14968
rect 357348 14952 357400 14958
rect 357348 14894 357400 14900
rect 350172 14884 350224 14890
rect 350172 14826 350224 14832
rect 342996 12096 343048 12102
rect 340142 12064 340198 12073
rect 342996 12038 343048 12044
rect 340142 11999 340198 12008
rect 339500 4004 339552 4010
rect 339500 3946 339552 3952
rect 338304 3664 338356 3670
rect 338304 3606 338356 3612
rect 339408 3664 339460 3670
rect 339408 3606 339460 3612
rect 337108 3052 337160 3058
rect 337108 2994 337160 3000
rect 338028 3052 338080 3058
rect 338028 2994 338080 3000
rect 337120 480 337148 2994
rect 338316 480 338344 3606
rect 339512 480 339540 3946
rect 340156 3942 340184 11999
rect 343008 11626 343036 12038
rect 342996 11620 343048 11626
rect 342996 11562 343048 11568
rect 349068 11620 349120 11626
rect 349068 11562 349120 11568
rect 345664 8832 345716 8838
rect 345664 8774 345716 8780
rect 344284 7744 344336 7750
rect 344284 7686 344336 7692
rect 340696 7336 340748 7342
rect 340696 7278 340748 7284
rect 340328 4004 340380 4010
rect 340328 3946 340380 3952
rect 340144 3936 340196 3942
rect 340144 3878 340196 3884
rect 340340 3262 340368 3946
rect 340328 3256 340380 3262
rect 340328 3198 340380 3204
rect 340708 480 340736 7278
rect 343088 2916 343140 2922
rect 343088 2858 343140 2864
rect 341892 876 341944 882
rect 341892 818 341944 824
rect 341904 480 341932 818
rect 343100 480 343128 2858
rect 344296 480 344324 7686
rect 345676 4010 345704 8774
rect 347872 7812 347924 7818
rect 347872 7754 347924 7760
rect 345664 4004 345716 4010
rect 345664 3946 345716 3952
rect 346676 4004 346728 4010
rect 346676 3946 346728 3952
rect 345480 2032 345532 2038
rect 345480 1974 345532 1980
rect 345492 480 345520 1974
rect 346688 480 346716 3946
rect 347884 480 347912 7754
rect 349080 480 349108 11562
rect 350184 4842 350212 14826
rect 355324 12096 355376 12102
rect 355324 12038 355376 12044
rect 355336 11490 355364 12038
rect 355324 11484 355376 11490
rect 355324 11426 355376 11432
rect 352564 10192 352616 10198
rect 352564 10134 352616 10140
rect 351368 7880 351420 7886
rect 351368 7822 351420 7828
rect 350184 4814 350304 4842
rect 350276 480 350304 4814
rect 351380 480 351408 7822
rect 352576 480 352604 10134
rect 354956 7948 355008 7954
rect 354956 7890 355008 7896
rect 353760 5976 353812 5982
rect 353760 5918 353812 5924
rect 353772 480 353800 5918
rect 354968 480 354996 7890
rect 356152 5908 356204 5914
rect 356152 5850 356204 5856
rect 356058 2952 356114 2961
rect 356058 2887 356060 2896
rect 356112 2887 356114 2896
rect 356060 2858 356112 2864
rect 356164 480 356192 5850
rect 357360 480 357388 14894
rect 364248 13592 364300 13598
rect 364248 13534 364300 13540
rect 360108 13524 360160 13530
rect 360108 13466 360160 13472
rect 358544 8016 358596 8022
rect 358544 7958 358596 7964
rect 358556 480 358584 7958
rect 360120 626 360148 13466
rect 364156 12096 364208 12102
rect 364156 12038 364208 12044
rect 364168 11490 364196 12038
rect 364156 11484 364208 11490
rect 364156 11426 364208 11432
rect 362132 8084 362184 8090
rect 362132 8026 362184 8032
rect 360936 3188 360988 3194
rect 360936 3130 360988 3136
rect 359752 598 360148 626
rect 359752 480 359780 598
rect 360948 480 360976 3130
rect 362144 480 362172 8026
rect 364260 3670 364288 13534
rect 364984 10124 365036 10130
rect 364984 10066 365036 10072
rect 364340 4004 364392 4010
rect 364340 3946 364392 3952
rect 363328 3664 363380 3670
rect 363328 3606 363380 3612
rect 364248 3664 364300 3670
rect 364248 3606 364300 3612
rect 363340 480 363368 3606
rect 364352 3126 364380 3946
rect 364996 3330 365024 10066
rect 365720 8152 365772 8158
rect 365720 8094 365772 8100
rect 364984 3324 365036 3330
rect 364984 3266 365036 3272
rect 364524 3256 364576 3262
rect 364524 3198 364576 3204
rect 364340 3120 364392 3126
rect 364340 3062 364392 3068
rect 364536 480 364564 3198
rect 365732 480 365760 8094
rect 368400 3346 368428 14962
rect 368676 13666 368704 15098
rect 375196 13796 375248 13802
rect 375196 13738 375248 13744
rect 368664 13660 368716 13666
rect 368664 13602 368716 13608
rect 371148 13660 371200 13666
rect 371148 13602 371200 13608
rect 369216 8220 369268 8226
rect 369216 8162 369268 8168
rect 368032 3318 368428 3346
rect 366916 944 366968 950
rect 366916 886 366968 892
rect 366928 480 366956 886
rect 368032 480 368060 3318
rect 369122 2952 369178 2961
rect 369122 2887 369124 2896
rect 369176 2887 369178 2896
rect 369124 2858 369176 2864
rect 369228 480 369256 8162
rect 371160 4010 371188 13602
rect 374644 12096 374696 12102
rect 374644 12038 374696 12044
rect 374656 11490 374684 12038
rect 374644 11484 374696 11490
rect 374644 11426 374696 11432
rect 371424 8628 371476 8634
rect 371424 8570 371476 8576
rect 370412 4004 370464 4010
rect 370412 3946 370464 3952
rect 371148 4004 371200 4010
rect 371148 3946 371200 3952
rect 370424 480 370452 3946
rect 371436 3806 371464 8570
rect 372804 8288 372856 8294
rect 372804 8230 372856 8236
rect 371424 3800 371476 3806
rect 371424 3742 371476 3748
rect 371608 3324 371660 3330
rect 371608 3266 371660 3272
rect 371620 480 371648 3266
rect 372816 480 372844 8230
rect 375208 4010 375236 13738
rect 376220 9722 376248 15982
rect 378048 14272 378100 14278
rect 378048 14214 378100 14220
rect 378060 13734 378088 14214
rect 384120 14204 384172 14210
rect 384120 14146 384172 14152
rect 378048 13728 378100 13734
rect 378048 13670 378100 13676
rect 378140 13728 378192 13734
rect 378140 13670 378192 13676
rect 378152 13546 378180 13670
rect 378060 13518 378180 13546
rect 376208 9716 376260 9722
rect 376208 9658 376260 9664
rect 376392 9716 376444 9722
rect 376392 9658 376444 9664
rect 375288 4684 375340 4690
rect 375288 4626 375340 4632
rect 374000 4004 374052 4010
rect 374000 3946 374052 3952
rect 375196 4004 375248 4010
rect 375196 3946 375248 3952
rect 374012 480 374040 3946
rect 374090 2952 374146 2961
rect 374090 2887 374092 2896
rect 374144 2887 374146 2896
rect 374092 2858 374144 2864
rect 375300 2394 375328 4626
rect 375208 2366 375328 2394
rect 375208 480 375236 2366
rect 376404 480 376432 9658
rect 378060 4010 378088 13518
rect 384132 13258 384160 14146
rect 384120 13252 384172 13258
rect 384120 13194 384172 13200
rect 384488 13252 384540 13258
rect 384488 13194 384540 13200
rect 382188 13048 382240 13054
rect 382188 12990 382240 12996
rect 378140 4548 378192 4554
rect 378140 4490 378192 4496
rect 377588 4004 377640 4010
rect 377588 3946 377640 3952
rect 378048 4004 378100 4010
rect 378048 3946 378100 3952
rect 377600 480 377628 3946
rect 378152 3398 378180 4490
rect 382200 4146 382228 12990
rect 384304 12096 384356 12102
rect 384304 12038 384356 12044
rect 384316 11490 384344 12038
rect 384304 11484 384356 11490
rect 384304 11426 384356 11432
rect 384500 8362 384528 13194
rect 384488 8356 384540 8362
rect 384488 8298 384540 8304
rect 384672 8356 384724 8362
rect 384672 8298 384724 8304
rect 383568 7540 383620 7546
rect 383568 7482 383620 7488
rect 381176 4140 381228 4146
rect 381176 4082 381228 4088
rect 382188 4140 382240 4146
rect 382188 4082 382240 4088
rect 378232 4004 378284 4010
rect 378232 3946 378284 3952
rect 378140 3392 378192 3398
rect 378140 3334 378192 3340
rect 378244 3126 378272 3946
rect 378876 3664 378928 3670
rect 378876 3606 378928 3612
rect 378232 3120 378284 3126
rect 378232 3062 378284 3068
rect 378888 1850 378916 3606
rect 378966 2952 379022 2961
rect 378966 2887 379022 2896
rect 378980 2854 379008 2887
rect 378968 2848 379020 2854
rect 378968 2790 379020 2796
rect 378796 1822 378916 1850
rect 379980 1896 380032 1902
rect 379980 1838 380032 1844
rect 378796 480 378824 1822
rect 379992 480 380020 1838
rect 381188 480 381216 4082
rect 382372 3052 382424 3058
rect 382372 2994 382424 3000
rect 382384 480 382412 2994
rect 383580 480 383608 7482
rect 384304 4004 384356 4010
rect 384304 3946 384356 3952
rect 384316 3398 384344 3946
rect 384304 3392 384356 3398
rect 384304 3334 384356 3340
rect 383672 2922 383884 2938
rect 383660 2916 383896 2922
rect 383712 2910 383844 2916
rect 383660 2858 383712 2864
rect 383844 2858 383896 2864
rect 384684 480 384712 8298
rect 385040 7268 385092 7274
rect 385040 7210 385092 7216
rect 384856 4412 384908 4418
rect 384856 4354 384908 4360
rect 384868 3534 384896 4354
rect 385052 4146 385080 7210
rect 387720 4146 387748 16050
rect 405648 15292 405700 15298
rect 405648 15234 405700 15240
rect 398748 15224 398800 15230
rect 398748 15166 398800 15172
rect 390468 15088 390520 15094
rect 390468 15030 390520 15036
rect 389088 12980 389140 12986
rect 389088 12922 389140 12928
rect 385040 4140 385092 4146
rect 385040 4082 385092 4088
rect 387064 4140 387116 4146
rect 387064 4082 387116 4088
rect 387708 4140 387760 4146
rect 387708 4082 387760 4088
rect 385868 3800 385920 3806
rect 385868 3742 385920 3748
rect 384856 3528 384908 3534
rect 384856 3470 384908 3476
rect 385880 480 385908 3742
rect 387076 480 387104 4082
rect 389100 3126 389128 12922
rect 389272 4276 389324 4282
rect 389272 4218 389324 4224
rect 389284 4078 389312 4218
rect 390480 4146 390508 15030
rect 397368 14408 397420 14414
rect 397368 14350 397420 14356
rect 391848 12912 391900 12918
rect 391848 12854 391900 12860
rect 389456 4140 389508 4146
rect 389456 4082 389508 4088
rect 390468 4140 390520 4146
rect 390468 4082 390520 4088
rect 389272 4072 389324 4078
rect 389272 4014 389324 4020
rect 388260 3120 388312 3126
rect 388260 3062 388312 3068
rect 389088 3120 389140 3126
rect 389088 3062 389140 3068
rect 388272 480 388300 3062
rect 389468 480 389496 4082
rect 390652 1828 390704 1834
rect 390652 1770 390704 1776
rect 390664 480 390692 1770
rect 391860 480 391888 12854
rect 395988 12708 396040 12714
rect 395988 12650 396040 12656
rect 393964 12096 394016 12102
rect 393964 12038 394016 12044
rect 393976 11422 394004 12038
rect 393964 11416 394016 11422
rect 393964 11358 394016 11364
rect 393226 10704 393282 10713
rect 393226 10639 393282 10648
rect 393240 4418 393268 10639
rect 394240 5840 394292 5846
rect 394240 5782 394292 5788
rect 393228 4412 393280 4418
rect 393228 4354 393280 4360
rect 393964 4004 394016 4010
rect 393964 3946 394016 3952
rect 393044 3528 393096 3534
rect 393044 3470 393096 3476
rect 393056 480 393084 3470
rect 393976 3398 394004 3946
rect 393964 3392 394016 3398
rect 393964 3334 394016 3340
rect 394252 480 394280 5782
rect 396000 4146 396028 12650
rect 397380 4146 397408 14350
rect 395436 4140 395488 4146
rect 395436 4082 395488 4088
rect 395988 4140 396040 4146
rect 395988 4082 396040 4088
rect 396632 4140 396684 4146
rect 396632 4082 396684 4088
rect 397368 4140 397420 4146
rect 397368 4082 397420 4088
rect 397460 4140 397512 4146
rect 397460 4082 397512 4088
rect 395448 480 395476 4082
rect 396644 480 396672 4082
rect 397472 3534 397500 4082
rect 398760 3534 398788 15166
rect 403624 12096 403676 12102
rect 403624 12038 403676 12044
rect 400220 11484 400272 11490
rect 400220 11426 400272 11432
rect 399024 8764 399076 8770
rect 399024 8706 399076 8712
rect 397460 3528 397512 3534
rect 397460 3470 397512 3476
rect 397828 3528 397880 3534
rect 397828 3470 397880 3476
rect 398748 3528 398800 3534
rect 398748 3470 398800 3476
rect 397840 480 397868 3470
rect 398840 2984 398892 2990
rect 398760 2932 398840 2938
rect 398760 2926 398892 2932
rect 398760 2922 398880 2926
rect 398748 2916 398880 2922
rect 398800 2910 398880 2916
rect 398748 2858 398800 2864
rect 399036 480 399064 8706
rect 400232 480 400260 11426
rect 403636 11422 403664 12038
rect 403624 11416 403676 11422
rect 403624 11358 403676 11364
rect 403716 4616 403768 4622
rect 403716 4558 403768 4564
rect 403624 4004 403676 4010
rect 403624 3946 403676 3952
rect 402520 3392 402572 3398
rect 402520 3334 402572 3340
rect 401324 1760 401376 1766
rect 401324 1702 401376 1708
rect 401336 480 401364 1702
rect 402532 480 402560 3334
rect 403636 3126 403664 3946
rect 403624 3120 403676 3126
rect 403624 3062 403676 3068
rect 403728 480 403756 4558
rect 405660 4010 405688 15234
rect 414216 14521 414244 16388
rect 414202 14512 414258 14521
rect 414202 14447 414258 14456
rect 408408 14340 408460 14346
rect 408408 14282 408460 14288
rect 407028 12844 407080 12850
rect 407028 12786 407080 12792
rect 407040 4010 407068 12786
rect 408420 4010 408448 14282
rect 411260 14068 411312 14074
rect 411260 14010 411312 14016
rect 409144 13184 409196 13190
rect 409144 13126 409196 13132
rect 409156 12646 409184 13126
rect 409144 12640 409196 12646
rect 409144 12582 409196 12588
rect 409696 11416 409748 11422
rect 409696 11358 409748 11364
rect 408500 7472 408552 7478
rect 408500 7414 408552 7420
rect 404912 4004 404964 4010
rect 404912 3946 404964 3952
rect 405648 4004 405700 4010
rect 405648 3946 405700 3952
rect 406108 4004 406160 4010
rect 406108 3946 406160 3952
rect 407028 4004 407080 4010
rect 407028 3946 407080 3952
rect 407304 4004 407356 4010
rect 407304 3946 407356 3952
rect 408408 4004 408460 4010
rect 408408 3946 408460 3952
rect 404924 480 404952 3946
rect 406120 480 406148 3946
rect 407316 480 407344 3946
rect 408512 480 408540 7414
rect 409708 480 409736 11358
rect 411272 9042 411300 14010
rect 413284 12096 413336 12102
rect 413284 12038 413336 12044
rect 413296 11354 413324 12038
rect 413284 11348 413336 11354
rect 413284 11290 413336 11296
rect 411260 9036 411312 9042
rect 411260 8978 411312 8984
rect 414480 9036 414532 9042
rect 414480 8978 414532 8984
rect 412088 8696 412140 8702
rect 412088 8638 412140 8644
rect 411168 4480 411220 4486
rect 411168 4422 411220 4428
rect 410892 3528 410944 3534
rect 410892 3470 410944 3476
rect 410904 480 410932 3470
rect 411180 3466 411208 4422
rect 411168 3460 411220 3466
rect 411168 3402 411220 3408
rect 412100 480 412128 8638
rect 413192 7404 413244 7410
rect 413192 7346 413244 7352
rect 412638 3088 412694 3097
rect 412638 3023 412694 3032
rect 412652 2990 412680 3023
rect 412640 2984 412692 2990
rect 412640 2926 412692 2932
rect 413204 2802 413232 7346
rect 413284 4004 413336 4010
rect 413284 3946 413336 3952
rect 413296 3126 413324 3946
rect 413284 3120 413336 3126
rect 413284 3062 413336 3068
rect 414202 3088 414258 3097
rect 414202 3023 414258 3032
rect 414216 2854 414244 3023
rect 414204 2848 414256 2854
rect 413204 2774 413324 2802
rect 414204 2790 414256 2796
rect 413296 480 413324 2774
rect 414492 480 414520 8978
rect 414584 7585 414612 16388
rect 415320 15337 415348 16388
rect 415306 15328 415362 15337
rect 415306 15263 415362 15272
rect 415308 12776 415360 12782
rect 415308 12718 415360 12724
rect 415320 12646 415348 12718
rect 415308 12640 415360 12646
rect 415308 12582 415360 12588
rect 416056 11762 416084 16388
rect 416332 16374 416530 16402
rect 416044 11756 416096 11762
rect 416044 11698 416096 11704
rect 414570 7576 414626 7585
rect 414570 7511 414626 7520
rect 416332 7426 416360 16374
rect 416688 11756 416740 11762
rect 416688 11698 416740 11704
rect 415596 7398 416360 7426
rect 415596 2106 415624 7398
rect 416700 3466 416728 11698
rect 416884 10334 416912 16388
rect 417252 13025 417280 16388
rect 417528 16374 417634 16402
rect 417238 13016 417294 13025
rect 417238 12951 417294 12960
rect 416872 10328 416924 10334
rect 416872 10270 416924 10276
rect 417056 10328 417108 10334
rect 417056 10270 417108 10276
rect 415676 3460 415728 3466
rect 415676 3402 415728 3408
rect 416688 3460 416740 3466
rect 416688 3402 416740 3408
rect 415584 2100 415636 2106
rect 415584 2042 415636 2048
rect 415688 480 415716 3402
rect 417068 2802 417096 10270
rect 417528 5137 417556 16374
rect 417988 8945 418016 16388
rect 418356 14210 418384 16388
rect 418632 16374 418830 16402
rect 418344 14204 418396 14210
rect 418344 14146 418396 14152
rect 418528 14204 418580 14210
rect 418528 14146 418580 14152
rect 418540 9042 418568 14146
rect 418528 9036 418580 9042
rect 418528 8978 418580 8984
rect 417974 8936 418030 8945
rect 418632 8922 418660 16374
rect 419184 11665 419212 16388
rect 419448 14680 419500 14686
rect 419448 14622 419500 14628
rect 419460 14074 419488 14622
rect 419552 14482 419580 16388
rect 419632 14612 419684 14618
rect 419632 14554 419684 14560
rect 419540 14476 419592 14482
rect 419540 14418 419592 14424
rect 419540 14136 419592 14142
rect 419540 14078 419592 14084
rect 419448 14068 419500 14074
rect 419448 14010 419500 14016
rect 419170 11656 419226 11665
rect 419170 11591 419226 11600
rect 418804 10056 418856 10062
rect 418804 9998 418856 10004
rect 417974 8871 418030 8880
rect 418264 8894 418660 8922
rect 418264 6361 418292 8894
rect 418250 6352 418306 6361
rect 418250 6287 418306 6296
rect 417514 5128 417570 5137
rect 417514 5063 417570 5072
rect 418816 3398 418844 9998
rect 419552 9994 419580 14078
rect 419540 9988 419592 9994
rect 419540 9930 419592 9936
rect 419172 9036 419224 9042
rect 419172 8978 419224 8984
rect 418804 3392 418856 3398
rect 418804 3334 418856 3340
rect 416884 2774 417096 2802
rect 416884 480 416912 2774
rect 417976 2100 418028 2106
rect 417976 2042 418028 2048
rect 417988 480 418016 2042
rect 419184 480 419212 8978
rect 419644 7342 419672 14554
rect 419920 10713 419948 16388
rect 419906 10704 419962 10713
rect 419906 10639 419962 10648
rect 420288 7721 420316 16388
rect 420656 14686 420684 16388
rect 420644 14680 420696 14686
rect 420644 14622 420696 14628
rect 420920 14544 420972 14550
rect 420920 14486 420972 14492
rect 420932 8702 420960 14486
rect 420920 8696 420972 8702
rect 420920 8638 420972 8644
rect 420274 7712 420330 7721
rect 420274 7647 420330 7656
rect 419632 7336 419684 7342
rect 419632 7278 419684 7284
rect 420368 7336 420420 7342
rect 420368 7278 420420 7284
rect 420380 480 420408 7278
rect 421116 5506 421144 16388
rect 421484 13122 421512 16388
rect 421852 14657 421880 16388
rect 421838 14648 421894 14657
rect 421838 14583 421894 14592
rect 422220 14006 422248 16388
rect 422208 14000 422260 14006
rect 422208 13942 422260 13948
rect 421472 13116 421524 13122
rect 421472 13058 421524 13064
rect 422588 12782 422616 16388
rect 422956 14482 422984 16388
rect 423048 16374 423430 16402
rect 422944 14476 422996 14482
rect 422944 14418 422996 14424
rect 422576 12776 422628 12782
rect 422576 12718 422628 12724
rect 422760 12776 422812 12782
rect 422760 12718 422812 12724
rect 421564 12708 421616 12714
rect 421564 12650 421616 12656
rect 421104 5500 421156 5506
rect 421104 5442 421156 5448
rect 421576 3210 421604 12650
rect 422772 12617 422800 12718
rect 422298 12608 422354 12617
rect 422298 12543 422300 12552
rect 422352 12543 422354 12552
rect 422758 12608 422814 12617
rect 422758 12543 422814 12552
rect 422300 12514 422352 12520
rect 422208 12096 422260 12102
rect 422208 12038 422260 12044
rect 422220 11354 422248 12038
rect 423048 11642 423076 16374
rect 423128 14476 423180 14482
rect 423128 14418 423180 14424
rect 423140 11801 423168 14418
rect 423126 11792 423182 11801
rect 423126 11727 423182 11736
rect 422312 11614 423076 11642
rect 422208 11348 422260 11354
rect 422208 11290 422260 11296
rect 422312 4486 422340 11614
rect 423784 8974 423812 16388
rect 424152 14793 424180 16388
rect 424138 14784 424194 14793
rect 424138 14719 424194 14728
rect 423772 8968 423824 8974
rect 423772 8910 423824 8916
rect 422760 8696 422812 8702
rect 422760 8638 422812 8644
rect 422300 4480 422352 4486
rect 422300 4422 422352 4428
rect 422300 4004 422352 4010
rect 422300 3946 422352 3952
rect 421484 3194 421604 3210
rect 422312 3194 422340 3946
rect 421472 3188 421604 3194
rect 421524 3182 421604 3188
rect 422300 3188 422352 3194
rect 421472 3130 421524 3136
rect 422300 3130 422352 3136
rect 421564 3120 421616 3126
rect 421564 3062 421616 3068
rect 421576 480 421604 3062
rect 422772 480 422800 8638
rect 424888 7614 424916 16388
rect 425256 14074 425284 16388
rect 425532 16374 425730 16402
rect 425244 14068 425296 14074
rect 425244 14010 425296 14016
rect 425060 13932 425112 13938
rect 425060 13874 425112 13880
rect 425072 13161 425100 13874
rect 425058 13152 425114 13161
rect 424968 13116 425020 13122
rect 425058 13087 425114 13096
rect 424968 13058 425020 13064
rect 424876 7608 424928 7614
rect 424876 7550 424928 7556
rect 424980 3466 425008 13058
rect 425532 11354 425560 16374
rect 426452 14482 426480 16388
rect 426820 15473 426848 16388
rect 426912 16374 427202 16402
rect 427280 16374 427570 16402
rect 427924 16374 428030 16402
rect 428108 16374 428398 16402
rect 426806 15464 426862 15473
rect 426806 15399 426862 15408
rect 426440 14476 426492 14482
rect 426440 14418 426492 14424
rect 426912 12866 426940 16374
rect 426992 14680 427044 14686
rect 426992 14622 427044 14628
rect 426544 12838 426940 12866
rect 425060 11348 425112 11354
rect 425060 11290 425112 11296
rect 425520 11348 425572 11354
rect 425520 11290 425572 11296
rect 423956 3460 424008 3466
rect 423956 3402 424008 3408
rect 424968 3460 425020 3466
rect 424968 3402 425020 3408
rect 423968 480 423996 3402
rect 425072 2174 425100 11290
rect 426348 8968 426400 8974
rect 426348 8910 426400 8916
rect 426256 7608 426308 7614
rect 426256 7550 426308 7556
rect 425152 3392 425204 3398
rect 425152 3334 425204 3340
rect 425060 2168 425112 2174
rect 425060 2110 425112 2116
rect 425164 480 425192 3334
rect 426268 3058 426296 7550
rect 426256 3052 426308 3058
rect 426256 2994 426308 3000
rect 426360 480 426388 8910
rect 426544 4826 426572 12838
rect 427004 12730 427032 14622
rect 426728 12702 427032 12730
rect 427084 12708 427136 12714
rect 426728 7857 426756 12702
rect 427084 12650 427136 12656
rect 427096 12510 427124 12650
rect 427084 12504 427136 12510
rect 427084 12446 427136 12452
rect 427280 9110 427308 16374
rect 427268 9104 427320 9110
rect 427268 9046 427320 9052
rect 427544 9104 427596 9110
rect 427544 9046 427596 9052
rect 426714 7848 426770 7857
rect 426714 7783 426770 7792
rect 426532 4820 426584 4826
rect 426532 4762 426584 4768
rect 427084 4480 427136 4486
rect 427084 4422 427136 4428
rect 427096 3505 427124 4422
rect 427082 3496 427138 3505
rect 427082 3431 427138 3440
rect 427556 480 427584 9046
rect 427924 2009 427952 16374
rect 428004 12708 428056 12714
rect 428004 12650 428056 12656
rect 428016 12510 428044 12650
rect 428004 12504 428056 12510
rect 428004 12446 428056 12452
rect 427910 2000 427966 2009
rect 427910 1935 427966 1944
rect 213644 332 213696 338
rect 213644 274 213696 280
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428108 66 428136 16374
rect 428464 14544 428516 14550
rect 428464 14486 428516 14492
rect 428476 4894 428504 14486
rect 428752 13938 428780 16388
rect 429120 15609 429148 16388
rect 429212 16374 429502 16402
rect 429580 16374 429870 16402
rect 430132 16374 430330 16402
rect 429106 15600 429162 15609
rect 429106 15535 429162 15544
rect 428740 13932 428792 13938
rect 428740 13874 428792 13880
rect 429212 9217 429240 16374
rect 429580 11642 429608 16374
rect 429304 11614 429608 11642
rect 429198 9208 429254 9217
rect 429198 9143 429254 9152
rect 429304 6225 429332 11614
rect 430132 6934 430160 16374
rect 430684 9081 430712 16388
rect 431052 14550 431080 16388
rect 431420 16182 431448 16388
rect 431512 16374 431802 16402
rect 431408 16176 431460 16182
rect 431408 16118 431460 16124
rect 431040 14544 431092 14550
rect 431040 14486 431092 14492
rect 431512 9330 431540 16374
rect 431960 12096 432012 12102
rect 431960 12038 432012 12044
rect 431972 11286 432000 12038
rect 431960 11280 432012 11286
rect 431960 11222 432012 11228
rect 431052 9302 431540 9330
rect 431052 9246 431080 9302
rect 431040 9240 431092 9246
rect 431040 9182 431092 9188
rect 431132 9240 431184 9246
rect 431132 9182 431184 9188
rect 430670 9072 430726 9081
rect 430670 9007 430726 9016
rect 429476 6928 429528 6934
rect 429476 6870 429528 6876
rect 430120 6928 430172 6934
rect 430120 6870 430172 6876
rect 429290 6216 429346 6225
rect 429290 6151 429346 6160
rect 428464 4888 428516 4894
rect 428464 4830 428516 4836
rect 428740 3460 428792 3466
rect 428740 3402 428792 3408
rect 428752 480 428780 3402
rect 429488 2145 429516 6870
rect 429936 4820 429988 4826
rect 429936 4762 429988 4768
rect 429474 2136 429530 2145
rect 429474 2071 429530 2080
rect 429948 480 429976 4762
rect 431144 480 431172 9182
rect 432156 9178 432184 16388
rect 432340 16374 432630 16402
rect 432144 9172 432196 9178
rect 432144 9114 432196 9120
rect 432340 9058 432368 16374
rect 433248 14544 433300 14550
rect 433248 14486 433300 14492
rect 432064 9030 432368 9058
rect 431868 4004 431920 4010
rect 431868 3946 431920 3952
rect 431960 4004 432012 4010
rect 431960 3946 432012 3952
rect 431880 3194 431908 3946
rect 431868 3188 431920 3194
rect 431868 3130 431920 3136
rect 431972 3058 432000 3946
rect 431960 3052 432012 3058
rect 431960 2994 432012 3000
rect 431960 2780 432012 2786
rect 431960 2722 432012 2728
rect 431972 2174 432000 2722
rect 432064 2689 432092 9030
rect 433260 3262 433288 14486
rect 433352 9314 433380 16388
rect 433720 16250 433748 16388
rect 433812 16374 434102 16402
rect 433708 16244 433760 16250
rect 433708 16186 433760 16192
rect 433340 9308 433392 9314
rect 433340 9250 433392 9256
rect 433340 8560 433392 8566
rect 433340 8502 433392 8508
rect 433352 3369 433380 8502
rect 433524 4888 433576 4894
rect 433524 4830 433576 4836
rect 433338 3360 433394 3369
rect 433338 3295 433394 3304
rect 432328 3256 432380 3262
rect 432328 3198 432380 3204
rect 433248 3256 433300 3262
rect 433248 3198 433300 3204
rect 432050 2680 432106 2689
rect 432050 2615 432106 2624
rect 431960 2168 432012 2174
rect 431960 2110 432012 2116
rect 432340 480 432368 3198
rect 433536 480 433564 4830
rect 428096 60 428148 66
rect 428096 2 428148 8
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 433812 134 433840 16374
rect 434456 13326 434484 16388
rect 434930 16374 435036 16402
rect 434444 13320 434496 13326
rect 434444 13262 434496 13268
rect 434812 11348 434864 11354
rect 434812 11290 434864 11296
rect 434628 9172 434680 9178
rect 434628 9114 434680 9120
rect 434640 480 434668 9114
rect 434720 3664 434772 3670
rect 434720 3606 434772 3612
rect 434732 3505 434760 3606
rect 434718 3496 434774 3505
rect 434718 3431 434774 3440
rect 434824 2242 434852 11290
rect 434812 2236 434864 2242
rect 434812 2178 434864 2184
rect 435008 1698 435036 16374
rect 435652 14686 435680 16388
rect 435744 16374 436034 16402
rect 436112 16374 436402 16402
rect 436480 16374 436770 16402
rect 435640 14680 435692 14686
rect 435640 14622 435692 14628
rect 435744 11354 435772 16374
rect 435732 11348 435784 11354
rect 435732 11290 435784 11296
rect 435824 3188 435876 3194
rect 435824 3130 435876 3136
rect 434996 1692 435048 1698
rect 434996 1634 435048 1640
rect 435836 480 435864 3130
rect 433800 128 433852 134
rect 433800 70 433852 76
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436112 202 436140 16374
rect 436480 9450 436508 16374
rect 437216 15638 437244 16388
rect 437598 16374 437704 16402
rect 437204 15632 437256 15638
rect 437204 15574 437256 15580
rect 436744 13184 436796 13190
rect 436744 13126 436796 13132
rect 436468 9444 436520 9450
rect 436468 9386 436520 9392
rect 436756 3641 436784 13126
rect 437572 7200 437624 7206
rect 437572 7142 437624 7148
rect 437020 5500 437072 5506
rect 437020 5442 437072 5448
rect 436742 3632 436798 3641
rect 436742 3567 436798 3576
rect 437032 480 437060 5442
rect 437584 2310 437612 7142
rect 437572 2304 437624 2310
rect 437572 2246 437624 2252
rect 436100 196 436152 202
rect 436100 138 436152 144
rect 436990 -960 437102 480
rect 437676 270 437704 16374
rect 437952 13297 437980 16388
rect 438044 16374 438334 16402
rect 437938 13288 437994 13297
rect 437938 13223 437994 13232
rect 438044 7206 438072 16374
rect 439056 9382 439084 16388
rect 439516 15706 439544 16388
rect 439608 16374 439898 16402
rect 439504 15700 439556 15706
rect 439504 15642 439556 15648
rect 439044 9376 439096 9382
rect 439044 9318 439096 9324
rect 438216 9308 438268 9314
rect 438216 9250 438268 9256
rect 438032 7200 438084 7206
rect 438032 7142 438084 7148
rect 438228 480 438256 9250
rect 439608 6186 439636 16374
rect 440252 12073 440280 16388
rect 440528 16374 440634 16402
rect 440424 14680 440476 14686
rect 440424 14622 440476 14628
rect 440238 12064 440294 12073
rect 440238 11999 440294 12008
rect 440436 10402 440464 14622
rect 440424 10396 440476 10402
rect 440424 10338 440476 10344
rect 439780 9444 439832 9450
rect 439780 9386 439832 9392
rect 439596 6180 439648 6186
rect 439596 6122 439648 6128
rect 439044 5772 439096 5778
rect 439044 5714 439096 5720
rect 439056 4078 439084 5714
rect 439044 4072 439096 4078
rect 439044 4014 439096 4020
rect 439320 4004 439372 4010
rect 439320 3946 439372 3952
rect 439332 3058 439360 3946
rect 439596 3732 439648 3738
rect 439596 3674 439648 3680
rect 439502 3496 439558 3505
rect 439502 3431 439504 3440
rect 439556 3431 439558 3440
rect 439504 3402 439556 3408
rect 439320 3052 439372 3058
rect 439320 2994 439372 3000
rect 439412 3052 439464 3058
rect 439412 2994 439464 3000
rect 439424 480 439452 2994
rect 439608 2990 439636 3674
rect 439688 3460 439740 3466
rect 439688 3402 439740 3408
rect 439700 3330 439728 3402
rect 439688 3324 439740 3330
rect 439688 3266 439740 3272
rect 439792 3262 439820 9386
rect 440528 5273 440556 16374
rect 440608 10396 440660 10402
rect 440608 10338 440660 10344
rect 440514 5264 440570 5273
rect 440514 5199 440570 5208
rect 439780 3256 439832 3262
rect 439780 3198 439832 3204
rect 439596 2984 439648 2990
rect 439596 2926 439648 2932
rect 440620 480 440648 10338
rect 440988 9353 441016 16388
rect 440974 9344 441030 9353
rect 440974 9279 441030 9288
rect 441356 7993 441384 16388
rect 441724 16374 441830 16402
rect 441908 16374 442198 16402
rect 441724 11082 441752 16374
rect 441712 11076 441764 11082
rect 441712 11018 441764 11024
rect 441908 10146 441936 16374
rect 442552 13433 442580 16388
rect 442736 16374 442934 16402
rect 442538 13424 442594 13433
rect 442538 13359 442594 13368
rect 442264 12096 442316 12102
rect 442264 12038 442316 12044
rect 442276 11286 442304 12038
rect 442264 11280 442316 11286
rect 442264 11222 442316 11228
rect 441988 11076 442040 11082
rect 441988 11018 442040 11024
rect 441724 10118 441936 10146
rect 441342 7984 441398 7993
rect 441342 7919 441398 7928
rect 441528 2780 441580 2786
rect 441528 2722 441580 2728
rect 441540 2174 441568 2722
rect 441528 2168 441580 2174
rect 441528 2110 441580 2116
rect 441724 626 441752 10118
rect 442000 4865 442028 11018
rect 442356 9988 442408 9994
rect 442356 9930 442408 9936
rect 441986 4856 442042 4865
rect 441986 4791 442042 4800
rect 442368 4078 442396 9930
rect 442736 4962 442764 16374
rect 443656 9518 443684 16388
rect 443840 16374 444130 16402
rect 443644 9512 443696 9518
rect 443644 9454 443696 9460
rect 443840 5030 443868 16374
rect 444484 14686 444512 16388
rect 444668 16374 444866 16402
rect 445036 16374 445234 16402
rect 444472 14680 444524 14686
rect 444472 14622 444524 14628
rect 444380 12708 444432 12714
rect 444380 12650 444432 12656
rect 444392 12578 444420 12650
rect 444380 12572 444432 12578
rect 444380 12514 444432 12520
rect 444668 6254 444696 16374
rect 444656 6248 444708 6254
rect 444656 6190 444708 6196
rect 443828 5024 443880 5030
rect 445036 5001 445064 16374
rect 445588 10305 445616 16388
rect 445956 13394 445984 16388
rect 446140 16374 446430 16402
rect 445944 13388 445996 13394
rect 445944 13330 445996 13336
rect 445574 10296 445630 10305
rect 445574 10231 445630 10240
rect 445760 9920 445812 9926
rect 445760 9862 445812 9868
rect 445392 9376 445444 9382
rect 445392 9318 445444 9324
rect 443828 4966 443880 4972
rect 445022 4992 445078 5001
rect 442724 4956 442776 4962
rect 442724 4898 442776 4904
rect 443920 4956 443972 4962
rect 445022 4927 445078 4936
rect 443920 4898 443972 4904
rect 443000 4412 443052 4418
rect 443000 4354 443052 4360
rect 441804 4072 441856 4078
rect 441804 4014 441856 4020
rect 442356 4072 442408 4078
rect 442356 4014 442408 4020
rect 441632 598 441752 626
rect 437664 264 437716 270
rect 437664 206 437716 212
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441632 338 441660 598
rect 441816 480 441844 4014
rect 443012 3777 443040 4354
rect 442998 3768 443054 3777
rect 442998 3703 443054 3712
rect 443000 2848 443052 2854
rect 443000 2790 443052 2796
rect 443012 480 443040 2790
rect 443932 2530 443960 4898
rect 444286 3496 444342 3505
rect 444024 3454 444236 3482
rect 444024 3398 444052 3454
rect 444208 3398 444236 3454
rect 444286 3431 444288 3440
rect 444340 3431 444342 3440
rect 444288 3402 444340 3408
rect 444012 3392 444064 3398
rect 444012 3334 444064 3340
rect 444196 3392 444248 3398
rect 444196 3334 444248 3340
rect 444196 3256 444248 3262
rect 444196 3198 444248 3204
rect 444208 2854 444236 3198
rect 444196 2848 444248 2854
rect 444196 2790 444248 2796
rect 443932 2502 444236 2530
rect 444208 480 444236 2502
rect 445404 480 445432 9318
rect 445772 3602 445800 9862
rect 446140 5098 446168 16374
rect 446784 10470 446812 16388
rect 447048 12776 447100 12782
rect 447048 12718 447100 12724
rect 447060 12510 447088 12718
rect 447048 12504 447100 12510
rect 447048 12446 447100 12452
rect 446772 10464 446824 10470
rect 446772 10406 446824 10412
rect 447152 9586 447180 16388
rect 447428 16374 447534 16402
rect 447612 16374 447902 16402
rect 447140 9580 447192 9586
rect 447140 9522 447192 9528
rect 447428 5166 447456 16374
rect 447612 10538 447640 16374
rect 447600 10532 447652 10538
rect 447600 10474 447652 10480
rect 448152 10532 448204 10538
rect 448152 10474 448204 10480
rect 447416 5160 447468 5166
rect 447416 5102 447468 5108
rect 446128 5092 446180 5098
rect 446128 5034 446180 5040
rect 447784 5024 447836 5030
rect 447784 4966 447836 4972
rect 446588 4072 446640 4078
rect 446588 4014 446640 4020
rect 446404 3664 446456 3670
rect 446402 3632 446404 3641
rect 446456 3632 446458 3641
rect 445760 3596 445812 3602
rect 446402 3567 446458 3576
rect 445760 3538 445812 3544
rect 446600 480 446628 4014
rect 447796 480 447824 4966
rect 448164 3058 448192 10474
rect 448256 8129 448284 16388
rect 448716 15366 448744 16388
rect 448808 16374 449098 16402
rect 449176 16374 449466 16402
rect 449636 16374 449834 16402
rect 448704 15360 448756 15366
rect 448704 15302 448756 15308
rect 448808 10606 448836 16374
rect 448796 10600 448848 10606
rect 448796 10542 448848 10548
rect 448980 10464 449032 10470
rect 448980 10406 449032 10412
rect 448242 8120 448298 8129
rect 448242 8055 448298 8064
rect 448704 7200 448756 7206
rect 448704 7142 448756 7148
rect 448152 3052 448204 3058
rect 448152 2994 448204 3000
rect 448716 2378 448744 7142
rect 448704 2372 448756 2378
rect 448704 2314 448756 2320
rect 448992 480 449020 10406
rect 449176 5234 449204 16374
rect 449636 7206 449664 16374
rect 450188 10441 450216 16388
rect 450556 10674 450584 16388
rect 451016 15978 451044 16388
rect 451004 15972 451056 15978
rect 451004 15914 451056 15920
rect 450544 10668 450596 10674
rect 450544 10610 450596 10616
rect 451384 10577 451412 16388
rect 451752 11937 451780 16388
rect 451738 11928 451794 11937
rect 451738 11863 451794 11872
rect 451370 10568 451426 10577
rect 451370 10503 451426 10512
rect 450174 10432 450230 10441
rect 450174 10367 450230 10376
rect 450084 9852 450136 9858
rect 450084 9794 450136 9800
rect 449624 7200 449676 7206
rect 449624 7142 449676 7148
rect 449164 5228 449216 5234
rect 449164 5170 449216 5176
rect 450096 2990 450124 9794
rect 452120 9722 452148 16388
rect 452488 10742 452516 16388
rect 453316 15434 453344 16388
rect 453304 15428 453356 15434
rect 453304 15370 453356 15376
rect 453684 10810 453712 16388
rect 453672 10804 453724 10810
rect 453672 10746 453724 10752
rect 452476 10736 452528 10742
rect 452476 10678 452528 10684
rect 452660 10736 452712 10742
rect 452660 10678 452712 10684
rect 452476 10600 452528 10606
rect 452476 10542 452528 10548
rect 451832 9716 451884 9722
rect 451832 9658 451884 9664
rect 452108 9716 452160 9722
rect 452108 9658 452160 9664
rect 451280 5092 451332 5098
rect 451280 5034 451332 5040
rect 450176 3052 450228 3058
rect 450176 2994 450228 3000
rect 450084 2984 450136 2990
rect 450084 2926 450136 2932
rect 450188 480 450216 2994
rect 451292 480 451320 5034
rect 451844 2802 451872 9658
rect 451568 2774 451872 2802
rect 451568 2446 451596 2774
rect 451556 2440 451608 2446
rect 451556 2382 451608 2388
rect 452488 480 452516 10542
rect 452672 3874 452700 10678
rect 454052 8634 454080 16388
rect 454328 16374 454434 16402
rect 454132 9512 454184 9518
rect 454132 9454 454184 9460
rect 454040 8628 454092 8634
rect 454040 8570 454092 8576
rect 452660 3868 452712 3874
rect 452660 3810 452712 3816
rect 454144 3330 454172 9454
rect 454132 3324 454184 3330
rect 454132 3266 454184 3272
rect 453672 2984 453724 2990
rect 453672 2926 453724 2932
rect 453684 480 453712 2926
rect 454328 2718 454356 16374
rect 454788 10878 454816 16388
rect 454776 10872 454828 10878
rect 454776 10814 454828 10820
rect 455156 9654 455184 16388
rect 455524 16374 455630 16402
rect 455800 16374 455998 16402
rect 455144 9648 455196 9654
rect 455144 9590 455196 9596
rect 455524 5302 455552 16374
rect 455800 5370 455828 16374
rect 456064 10668 456116 10674
rect 456064 10610 456116 10616
rect 455972 5636 456024 5642
rect 455972 5578 456024 5584
rect 455788 5364 455840 5370
rect 455788 5306 455840 5312
rect 455512 5296 455564 5302
rect 455512 5238 455564 5244
rect 454868 5160 454920 5166
rect 454868 5102 454920 5108
rect 454316 2712 454368 2718
rect 454316 2654 454368 2660
rect 454880 480 454908 5102
rect 455984 3942 456012 5578
rect 455972 3936 456024 3942
rect 455972 3878 456024 3884
rect 455972 3664 456024 3670
rect 455970 3632 455972 3641
rect 456024 3632 456026 3641
rect 455970 3567 456026 3576
rect 456076 480 456104 10610
rect 456352 10130 456380 16388
rect 456720 15502 456748 16388
rect 456708 15496 456760 15502
rect 456708 15438 456760 15444
rect 456984 13320 457036 13326
rect 456984 13262 457036 13268
rect 456340 10124 456392 10130
rect 456340 10066 456392 10072
rect 456800 7676 456852 7682
rect 456800 7618 456852 7624
rect 456892 7676 456944 7682
rect 456892 7618 456944 7624
rect 456812 7206 456840 7618
rect 456800 7200 456852 7206
rect 456800 7142 456852 7148
rect 456904 1970 456932 7618
rect 456996 6322 457024 13262
rect 456984 6316 457036 6322
rect 456984 6258 457036 6264
rect 456892 1964 456944 1970
rect 456892 1906 456944 1912
rect 441620 332 441672 338
rect 441620 274 441672 280
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457088 406 457116 16388
rect 457456 13326 457484 16388
rect 457640 16374 457930 16402
rect 457444 13320 457496 13326
rect 457444 13262 457496 13268
rect 457640 7682 457668 16374
rect 458284 10946 458312 16388
rect 458468 16374 458666 16402
rect 458272 10940 458324 10946
rect 458272 10882 458324 10888
rect 457628 7676 457680 7682
rect 457628 7618 457680 7624
rect 457260 5704 457312 5710
rect 457260 5646 457312 5652
rect 457272 480 457300 5646
rect 458468 5386 458496 16374
rect 459020 9722 459048 16388
rect 459756 13462 459784 16388
rect 459848 16374 460230 16402
rect 459744 13456 459796 13462
rect 459744 13398 459796 13404
rect 458640 9716 458692 9722
rect 458640 9658 458692 9664
rect 459008 9716 459060 9722
rect 459008 9658 459060 9664
rect 458376 5358 458496 5386
rect 458376 4554 458404 5358
rect 458456 5228 458508 5234
rect 458456 5170 458508 5176
rect 458364 4548 458416 4554
rect 458364 4490 458416 4496
rect 458468 480 458496 5170
rect 457076 400 457128 406
rect 457076 342 457128 348
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 458652 474 458680 9658
rect 459848 6390 459876 16374
rect 460584 9722 460612 16388
rect 460966 16374 461256 16402
rect 459928 9716 459980 9722
rect 459928 9658 459980 9664
rect 460572 9716 460624 9722
rect 460572 9658 460624 9664
rect 459836 6384 459888 6390
rect 459836 6326 459888 6332
rect 459652 6180 459704 6186
rect 459652 6122 459704 6128
rect 459664 480 459692 6122
rect 459940 2802 459968 9658
rect 461228 7274 461256 16374
rect 461216 7268 461268 7274
rect 461216 7210 461268 7216
rect 461320 6497 461348 16388
rect 461412 16374 461702 16402
rect 461780 16374 462070 16402
rect 462424 16374 462530 16402
rect 461306 6488 461362 6497
rect 461306 6423 461362 6432
rect 461412 6338 461440 16374
rect 461492 12096 461544 12102
rect 461492 12038 461544 12044
rect 461504 11286 461532 12038
rect 461492 11280 461544 11286
rect 461492 11222 461544 11228
rect 461320 6310 461440 6338
rect 460848 3868 460900 3874
rect 460848 3810 460900 3816
rect 459848 2774 459968 2802
rect 459848 542 459876 2774
rect 459836 536 459888 542
rect 458640 468 458692 474
rect 458640 410 458692 416
rect 459622 -960 459734 480
rect 459836 478 459888 484
rect 460860 480 460888 3810
rect 461320 2514 461348 6310
rect 461780 4486 461808 16374
rect 462320 6452 462372 6458
rect 462320 6394 462372 6400
rect 462044 5296 462096 5302
rect 462044 5238 462096 5244
rect 461768 4480 461820 4486
rect 461768 4422 461820 4428
rect 461584 3596 461636 3602
rect 461584 3538 461636 3544
rect 461596 2990 461624 3538
rect 461584 2984 461636 2990
rect 461584 2926 461636 2932
rect 461308 2508 461360 2514
rect 461308 2450 461360 2456
rect 462056 480 462084 5238
rect 462332 4010 462360 6394
rect 462424 6390 462452 16374
rect 463252 15570 463280 16388
rect 463344 16374 463634 16402
rect 463240 15564 463292 15570
rect 463240 15506 463292 15512
rect 463344 6526 463372 16374
rect 463988 11014 464016 16388
rect 463976 11008 464028 11014
rect 463976 10950 464028 10956
rect 464356 8566 464384 16388
rect 464448 16374 464830 16402
rect 464344 8560 464396 8566
rect 464344 8502 464396 8508
rect 464448 6594 464476 16374
rect 464988 14680 465040 14686
rect 464988 14622 465040 14628
rect 464436 6588 464488 6594
rect 464436 6530 464488 6536
rect 463332 6520 463384 6526
rect 463332 6462 463384 6468
rect 462412 6384 462464 6390
rect 462412 6326 462464 6332
rect 463240 6248 463292 6254
rect 463240 6190 463292 6196
rect 462320 4004 462372 4010
rect 462320 3946 462372 3952
rect 463252 480 463280 6190
rect 465000 4010 465028 14622
rect 465184 11830 465212 16388
rect 465172 11824 465224 11830
rect 465172 11766 465224 11772
rect 465552 7206 465580 16388
rect 465644 16374 465934 16402
rect 465540 7200 465592 7206
rect 465540 7142 465592 7148
rect 465644 6662 465672 16374
rect 466184 12640 466236 12646
rect 466182 12608 466184 12617
rect 466236 12608 466238 12617
rect 466182 12543 466238 12552
rect 466288 11898 466316 16388
rect 466656 13190 466684 16388
rect 466932 16374 467130 16402
rect 466644 13184 466696 13190
rect 466644 13126 466696 13132
rect 466276 11892 466328 11898
rect 466276 11834 466328 11840
rect 466828 11824 466880 11830
rect 466828 11766 466880 11772
rect 465632 6656 465684 6662
rect 465632 6598 465684 6604
rect 465632 5364 465684 5370
rect 465632 5306 465684 5312
rect 464436 4004 464488 4010
rect 464436 3946 464488 3952
rect 464988 4004 465040 4010
rect 464988 3946 465040 3952
rect 464448 480 464476 3946
rect 465644 480 465672 5306
rect 466840 480 466868 11766
rect 466932 6730 466960 16374
rect 467484 12034 467512 16388
rect 467852 14278 467880 16388
rect 467944 16374 468234 16402
rect 467840 14272 467892 14278
rect 467840 14214 467892 14220
rect 467472 12028 467524 12034
rect 467472 11970 467524 11976
rect 467944 6798 467972 16374
rect 468588 12102 468616 16388
rect 468680 16374 468970 16402
rect 468576 12096 468628 12102
rect 468576 12038 468628 12044
rect 468300 11348 468352 11354
rect 468300 11290 468352 11296
rect 467932 6792 467984 6798
rect 467932 6734 467984 6740
rect 466920 6724 466972 6730
rect 466920 6666 466972 6672
rect 467932 3324 467984 3330
rect 467932 3266 467984 3272
rect 467944 480 467972 3266
rect 468312 3058 468340 11290
rect 468680 4418 468708 16374
rect 469416 6866 469444 16388
rect 469784 11286 469812 16388
rect 470244 16374 470534 16402
rect 469772 11280 469824 11286
rect 469772 11222 469824 11228
rect 469404 6860 469456 6866
rect 469404 6802 469456 6808
rect 470244 6118 470272 16374
rect 470888 12170 470916 16388
rect 470876 12164 470928 12170
rect 470876 12106 470928 12112
rect 470508 11892 470560 11898
rect 470508 11834 470560 11840
rect 470232 6112 470284 6118
rect 470232 6054 470284 6060
rect 469128 4548 469180 4554
rect 469128 4490 469180 4496
rect 468668 4412 468720 4418
rect 468668 4354 468720 4360
rect 469036 3732 469088 3738
rect 469036 3674 469088 3680
rect 469048 3641 469076 3674
rect 469034 3632 469090 3641
rect 469034 3567 469090 3576
rect 468300 3052 468352 3058
rect 468300 2994 468352 3000
rect 469140 480 469168 4490
rect 470520 626 470548 11834
rect 471256 9722 471284 16388
rect 471716 15842 471744 16388
rect 471704 15836 471756 15842
rect 471704 15778 471756 15784
rect 471980 14272 472032 14278
rect 471980 14214 472032 14220
rect 471888 12640 471940 12646
rect 471886 12608 471888 12617
rect 471940 12608 471942 12617
rect 471886 12543 471942 12552
rect 471992 9722 472020 14214
rect 472084 12238 472112 16388
rect 472452 14929 472480 16388
rect 472438 14920 472494 14929
rect 472438 14855 472494 14864
rect 472072 12232 472124 12238
rect 472072 12174 472124 12180
rect 472716 11960 472768 11966
rect 472716 11902 472768 11908
rect 470600 9716 470652 9722
rect 470600 9658 470652 9664
rect 471244 9716 471296 9722
rect 471244 9658 471296 9664
rect 471520 9716 471572 9722
rect 471520 9658 471572 9664
rect 471980 9716 472032 9722
rect 471980 9658 472032 9664
rect 472164 9716 472216 9722
rect 472164 9658 472216 9664
rect 470612 5438 470640 9658
rect 470600 5432 470652 5438
rect 470600 5374 470652 5380
rect 470336 598 470548 626
rect 470336 480 470364 598
rect 471532 480 471560 9658
rect 471888 3664 471940 3670
rect 472072 3664 472124 3670
rect 471940 3624 472072 3652
rect 471888 3606 471940 3612
rect 472072 3606 472124 3612
rect 472176 2582 472204 9658
rect 472164 2576 472216 2582
rect 472164 2518 472216 2524
rect 472728 480 472756 11902
rect 472820 9722 472848 16388
rect 473188 11558 473216 16388
rect 473452 12232 473504 12238
rect 473452 12174 473504 12180
rect 473176 11552 473228 11558
rect 473176 11494 473228 11500
rect 472808 9716 472860 9722
rect 472808 9658 472860 9664
rect 473464 610 473492 12174
rect 473556 9926 473584 16388
rect 474016 12238 474044 16388
rect 474384 12306 474412 16388
rect 474752 14754 474780 16388
rect 474936 16374 475134 16402
rect 474740 14748 474792 14754
rect 474740 14690 474792 14696
rect 474372 12300 474424 12306
rect 474372 12242 474424 12248
rect 474004 12232 474056 12238
rect 474004 12174 474056 12180
rect 473912 12028 473964 12034
rect 473912 11970 473964 11976
rect 473544 9920 473596 9926
rect 473544 9862 473596 9868
rect 473452 604 473504 610
rect 473452 546 473504 552
rect 473924 480 473952 11970
rect 474740 10872 474792 10878
rect 474740 10814 474792 10820
rect 474752 3126 474780 10814
rect 474740 3120 474792 3126
rect 474740 3062 474792 3068
rect 474936 678 474964 16374
rect 475488 12374 475516 16388
rect 475476 12368 475528 12374
rect 475476 12310 475528 12316
rect 475856 9858 475884 16388
rect 476316 15162 476344 16388
rect 476304 15156 476356 15162
rect 476304 15098 476356 15104
rect 476028 12776 476080 12782
rect 476028 12718 476080 12724
rect 476040 12646 476068 12718
rect 476028 12640 476080 12646
rect 476028 12582 476080 12588
rect 476684 12442 476712 16388
rect 476672 12436 476724 12442
rect 476672 12378 476724 12384
rect 477052 10266 477080 16388
rect 477236 16374 477434 16402
rect 477512 16374 477802 16402
rect 477880 16374 478170 16402
rect 478340 16374 478630 16402
rect 479064 16390 479116 16396
rect 479800 16448 479852 16454
rect 534356 16448 534408 16454
rect 479800 16390 479852 16396
rect 477040 10260 477092 10266
rect 477040 10202 477092 10208
rect 475844 9852 475896 9858
rect 475844 9794 475896 9800
rect 477236 6934 477264 16374
rect 477512 11694 477540 16374
rect 477500 11688 477552 11694
rect 477880 11642 477908 16374
rect 477500 11630 477552 11636
rect 477604 11614 477908 11642
rect 476212 6928 476264 6934
rect 476212 6870 476264 6876
rect 477224 6928 477276 6934
rect 477224 6870 477276 6876
rect 475108 3936 475160 3942
rect 475108 3878 475160 3884
rect 474924 672 474976 678
rect 474924 614 474976 620
rect 475120 480 475148 3878
rect 476224 746 476252 6870
rect 476304 6316 476356 6322
rect 476304 6258 476356 6264
rect 476212 740 476264 746
rect 476212 682 476264 688
rect 476316 480 476344 6258
rect 477604 5778 477632 11614
rect 478340 11370 478368 16374
rect 478788 14748 478840 14754
rect 478788 14690 478840 14696
rect 478696 12096 478748 12102
rect 478696 12038 478748 12044
rect 477696 11342 478368 11370
rect 477592 5772 477644 5778
rect 477592 5714 477644 5720
rect 477500 3732 477552 3738
rect 477500 3674 477552 3680
rect 477512 480 477540 3674
rect 477696 814 477724 11342
rect 478708 3738 478736 12038
rect 478696 3732 478748 3738
rect 478696 3674 478748 3680
rect 478800 3482 478828 14690
rect 478984 6050 479012 16388
rect 478972 6044 479024 6050
rect 478972 5986 479024 5992
rect 479076 4758 479104 16390
rect 479352 14822 479380 16388
rect 479720 15774 479748 16388
rect 479708 15768 479760 15774
rect 479708 15710 479760 15716
rect 479340 14816 479392 14822
rect 479340 14758 479392 14764
rect 480456 10742 480484 16388
rect 480640 16374 480930 16402
rect 480444 10736 480496 10742
rect 480444 10678 480496 10684
rect 480640 10554 480668 16374
rect 480364 10526 480668 10554
rect 479892 6384 479944 6390
rect 479892 6326 479944 6332
rect 479064 4752 479116 4758
rect 479064 4694 479116 4700
rect 478708 3454 478828 3482
rect 477684 808 477736 814
rect 477684 750 477736 756
rect 478708 480 478736 3454
rect 479904 480 479932 6326
rect 480364 2650 480392 10526
rect 481284 8906 481312 16388
rect 481548 10736 481600 10742
rect 481548 10678 481600 10684
rect 481272 8900 481324 8906
rect 481272 8842 481324 8848
rect 481560 3738 481588 10678
rect 481652 8838 481680 16388
rect 482020 14142 482048 16388
rect 482388 15910 482416 16388
rect 482572 16374 482770 16402
rect 482376 15904 482428 15910
rect 482376 15846 482428 15852
rect 482008 14136 482060 14142
rect 482008 14078 482060 14084
rect 482572 11642 482600 16374
rect 482928 14816 482980 14822
rect 482928 14758 482980 14764
rect 481744 11614 482600 11642
rect 481640 8832 481692 8838
rect 481640 8774 481692 8780
rect 481744 5642 481772 11614
rect 481732 5636 481784 5642
rect 481732 5578 481784 5584
rect 482940 4758 482968 14758
rect 483216 14618 483244 16388
rect 483308 16374 483598 16402
rect 483676 16374 483966 16402
rect 484044 16374 484334 16402
rect 483204 14612 483256 14618
rect 483204 14554 483256 14560
rect 483112 11688 483164 11694
rect 483112 11630 483164 11636
rect 482284 4752 482336 4758
rect 482284 4694 482336 4700
rect 482928 4752 482980 4758
rect 482928 4694 482980 4700
rect 481088 3732 481140 3738
rect 481088 3674 481140 3680
rect 481548 3732 481600 3738
rect 481548 3674 481600 3680
rect 480352 2644 480404 2650
rect 480352 2586 480404 2592
rect 481100 480 481128 3674
rect 482296 480 482324 4694
rect 483018 3768 483074 3777
rect 483018 3703 483020 3712
rect 483072 3703 483074 3712
rect 483020 3674 483072 3680
rect 483020 3460 483072 3466
rect 483020 3402 483072 3408
rect 483032 3369 483060 3402
rect 483018 3360 483074 3369
rect 483018 3295 483074 3304
rect 483124 2718 483152 11630
rect 483204 3528 483256 3534
rect 483202 3496 483204 3505
rect 483256 3496 483258 3505
rect 483202 3431 483258 3440
rect 483112 2712 483164 2718
rect 483112 2654 483164 2660
rect 483308 882 483336 16374
rect 483676 11694 483704 16374
rect 483664 11688 483716 11694
rect 483664 11630 483716 11636
rect 484044 7750 484072 16374
rect 484492 12300 484544 12306
rect 484492 12242 484544 12248
rect 484308 12164 484360 12170
rect 484308 12106 484360 12112
rect 484032 7744 484084 7750
rect 484032 7686 484084 7692
rect 484320 3738 484348 12106
rect 484504 6458 484532 12242
rect 484492 6452 484544 6458
rect 484492 6394 484544 6400
rect 484584 6452 484636 6458
rect 484584 6394 484636 6400
rect 484398 3768 484454 3777
rect 483480 3732 483532 3738
rect 483480 3674 483532 3680
rect 484308 3732 484360 3738
rect 484398 3703 484400 3712
rect 484308 3674 484360 3680
rect 484452 3703 484454 3712
rect 484400 3674 484452 3680
rect 483388 3528 483440 3534
rect 483386 3496 483388 3505
rect 483440 3496 483442 3505
rect 483386 3431 483442 3440
rect 483296 876 483348 882
rect 483296 818 483348 824
rect 483492 480 483520 3674
rect 483572 3460 483624 3466
rect 483572 3402 483624 3408
rect 483584 3369 483612 3402
rect 483570 3360 483626 3369
rect 483570 3295 483626 3304
rect 484596 480 484624 6394
rect 484688 2038 484716 16388
rect 485056 12306 485084 16388
rect 485044 12300 485096 12306
rect 485044 12242 485096 12248
rect 485516 7818 485544 16388
rect 485884 11626 485912 16388
rect 486252 14890 486280 16388
rect 486240 14884 486292 14890
rect 486240 14826 486292 14832
rect 485872 11620 485924 11626
rect 485872 11562 485924 11568
rect 486620 7886 486648 16388
rect 486988 10198 487016 16388
rect 487172 16374 487370 16402
rect 487068 10804 487120 10810
rect 487068 10746 487120 10752
rect 486976 10192 487028 10198
rect 486976 10134 487028 10140
rect 486608 7880 486660 7886
rect 486608 7822 486660 7828
rect 485504 7812 485556 7818
rect 485504 7754 485556 7760
rect 485780 7676 485832 7682
rect 485780 7618 485832 7624
rect 484676 2032 484728 2038
rect 484676 1974 484728 1980
rect 485792 480 485820 7618
rect 487080 626 487108 10746
rect 487172 5982 487200 16374
rect 487816 7954 487844 16388
rect 488000 16374 488198 16402
rect 487804 7948 487856 7954
rect 487804 7890 487856 7896
rect 488000 7834 488028 16374
rect 488552 14958 488580 16388
rect 488540 14952 488592 14958
rect 488540 14894 488592 14900
rect 488920 8022 488948 16388
rect 489288 13530 489316 16388
rect 489276 13524 489328 13530
rect 489276 13466 489328 13472
rect 489656 12714 489684 16388
rect 489644 12708 489696 12714
rect 489644 12650 489696 12656
rect 489920 11008 489972 11014
rect 489920 10950 489972 10956
rect 489932 10810 489960 10950
rect 489920 10804 489972 10810
rect 489920 10746 489972 10752
rect 490116 8090 490144 16388
rect 490484 13598 490512 16388
rect 490472 13592 490524 13598
rect 490472 13534 490524 13540
rect 490576 12850 490788 12866
rect 490564 12844 490800 12850
rect 490616 12838 490748 12844
rect 490564 12786 490616 12792
rect 490748 12786 490800 12792
rect 490852 9450 490880 16388
rect 490840 9444 490892 9450
rect 490840 9386 490892 9392
rect 491220 8158 491248 16388
rect 491496 16374 491602 16402
rect 491208 8152 491260 8158
rect 491208 8094 491260 8100
rect 490104 8084 490156 8090
rect 490104 8026 490156 8032
rect 488908 8016 488960 8022
rect 488908 7958 488960 7964
rect 487264 7806 488028 7834
rect 490564 7812 490616 7818
rect 487160 5976 487212 5982
rect 487160 5918 487212 5924
rect 487264 5914 487292 7806
rect 490564 7754 490616 7760
rect 489368 7744 489420 7750
rect 489368 7686 489420 7692
rect 488172 6520 488224 6526
rect 488172 6462 488224 6468
rect 487252 5908 487304 5914
rect 487252 5850 487304 5856
rect 486988 598 487108 626
rect 486988 480 487016 598
rect 488184 480 488212 6462
rect 489380 480 489408 7686
rect 490576 480 490604 7754
rect 491496 950 491524 16374
rect 491956 15026 491984 16388
rect 491944 15020 491996 15026
rect 491944 14962 491996 14968
rect 491944 14884 491996 14890
rect 491944 14826 491996 14832
rect 491760 6588 491812 6594
rect 491760 6530 491812 6536
rect 491484 944 491536 950
rect 491484 886 491536 892
rect 491772 480 491800 6530
rect 491956 5710 491984 14826
rect 492416 8226 492444 16388
rect 492784 13666 492812 16388
rect 492772 13660 492824 13666
rect 492772 13602 492824 13608
rect 493152 9518 493180 16388
rect 493140 9512 493192 9518
rect 493140 9454 493192 9460
rect 493520 8294 493548 16388
rect 493888 13802 493916 16388
rect 494164 16374 494270 16402
rect 493876 13796 493928 13802
rect 493876 13738 493928 13744
rect 493508 8288 493560 8294
rect 493508 8230 493560 8236
rect 492404 8220 492456 8226
rect 492404 8162 492456 8168
rect 493876 7880 493928 7886
rect 493876 7822 493928 7828
rect 493692 6860 493744 6866
rect 493692 6802 493744 6808
rect 491944 5704 491996 5710
rect 491944 5646 491996 5652
rect 492956 4004 493008 4010
rect 492956 3946 493008 3952
rect 492968 480 492996 3946
rect 493704 1834 493732 6802
rect 493888 3398 493916 7822
rect 494164 4690 494192 16374
rect 494716 16046 494744 16388
rect 494704 16040 494756 16046
rect 494704 15982 494756 15988
rect 495084 13734 495112 16388
rect 495466 16374 495572 16402
rect 495072 13728 495124 13734
rect 495072 13670 495124 13676
rect 495348 13184 495400 13190
rect 495348 13126 495400 13132
rect 495256 6656 495308 6662
rect 495256 6598 495308 6604
rect 494152 4684 494204 4690
rect 494152 4626 494204 4632
rect 494152 3460 494204 3466
rect 494152 3402 494204 3408
rect 493876 3392 493928 3398
rect 493876 3334 493928 3340
rect 493692 1828 493744 1834
rect 493692 1770 493744 1776
rect 494164 480 494192 3402
rect 495268 3346 495296 6598
rect 495360 3466 495388 13126
rect 495544 3670 495572 16374
rect 495728 16374 495834 16402
rect 495532 3664 495584 3670
rect 495532 3606 495584 3612
rect 495348 3460 495400 3466
rect 495348 3402 495400 3408
rect 495268 3318 495388 3346
rect 495360 480 495388 3318
rect 495728 1902 495756 16374
rect 496188 13054 496216 16388
rect 496176 13048 496228 13054
rect 496176 12990 496228 12996
rect 496556 7614 496584 16388
rect 496728 13320 496780 13326
rect 496728 13262 496780 13268
rect 496544 7608 496596 7614
rect 496544 7550 496596 7556
rect 495716 1896 495768 1902
rect 495716 1838 495768 1844
rect 496740 610 496768 13262
rect 497016 7546 497044 16388
rect 497384 13258 497412 16388
rect 497372 13252 497424 13258
rect 497372 13194 497424 13200
rect 497752 9722 497780 16388
rect 498120 16114 498148 16388
rect 498108 16108 498160 16114
rect 498108 16050 498160 16056
rect 498108 13252 498160 13258
rect 498108 13194 498160 13200
rect 497096 9716 497148 9722
rect 497096 9658 497148 9664
rect 497740 9716 497792 9722
rect 497740 9658 497792 9664
rect 497004 7540 497056 7546
rect 497004 7482 497056 7488
rect 497108 3806 497136 9658
rect 497096 3800 497148 3806
rect 497096 3742 497148 3748
rect 498120 626 498148 13194
rect 498488 12986 498516 16388
rect 498856 15094 498884 16388
rect 498948 16374 499330 16402
rect 498844 15088 498896 15094
rect 498844 15030 498896 15036
rect 498476 12980 498528 12986
rect 498476 12922 498528 12928
rect 498948 6866 498976 16374
rect 499120 13456 499172 13462
rect 499120 13398 499172 13404
rect 498936 6860 498988 6866
rect 498936 6802 498988 6808
rect 498936 6724 498988 6730
rect 498936 6666 498988 6672
rect 496544 604 496596 610
rect 496544 546 496596 552
rect 496728 604 496780 610
rect 496728 546 496780 552
rect 497752 598 498148 626
rect 496556 480 496584 546
rect 497752 480 497780 598
rect 498948 480 498976 6666
rect 499132 3398 499160 13398
rect 499684 12782 499712 16388
rect 499776 16374 500066 16402
rect 500144 16374 500434 16402
rect 499672 12776 499724 12782
rect 499672 12718 499724 12724
rect 499776 4146 499804 16374
rect 500144 5846 500172 16374
rect 500224 13388 500276 13394
rect 500224 13330 500276 13336
rect 500132 5840 500184 5846
rect 500132 5782 500184 5788
rect 499764 4140 499816 4146
rect 499764 4082 499816 4088
rect 500132 3460 500184 3466
rect 500132 3402 500184 3408
rect 499120 3392 499172 3398
rect 499120 3334 499172 3340
rect 500144 480 500172 3402
rect 500236 3194 500264 13330
rect 500788 12714 500816 16388
rect 501156 14414 501184 16388
rect 501616 15230 501644 16388
rect 501604 15224 501656 15230
rect 501604 15166 501656 15172
rect 501144 14408 501196 14414
rect 501144 14350 501196 14356
rect 500776 12708 500828 12714
rect 500776 12650 500828 12656
rect 501236 12232 501288 12238
rect 501236 12174 501288 12180
rect 500316 3596 500368 3602
rect 500316 3538 500368 3544
rect 500328 3398 500356 3538
rect 500316 3392 500368 3398
rect 500316 3334 500368 3340
rect 500224 3188 500276 3194
rect 500224 3130 500276 3136
rect 501248 480 501276 12174
rect 501984 8770 502012 16388
rect 502352 11490 502380 16388
rect 502628 16374 502734 16402
rect 502340 11484 502392 11490
rect 502340 11426 502392 11432
rect 501972 8764 502024 8770
rect 501972 8706 502024 8712
rect 502432 6792 502484 6798
rect 502432 6734 502484 6740
rect 502444 480 502472 6734
rect 502628 1766 502656 16374
rect 503088 10062 503116 16388
rect 503180 16374 503470 16402
rect 503076 10056 503128 10062
rect 503076 9998 503128 10004
rect 503180 4622 503208 16374
rect 503916 15298 503944 16388
rect 503904 15292 503956 15298
rect 503904 15234 503956 15240
rect 503628 14612 503680 14618
rect 503628 14554 503680 14560
rect 503168 4616 503220 4622
rect 503168 4558 503220 4564
rect 502616 1760 502668 1766
rect 502616 1702 502668 1708
rect 503640 480 503668 14554
rect 504284 12850 504312 16388
rect 504652 14346 504680 16388
rect 504744 16374 505034 16402
rect 504640 14340 504692 14346
rect 504640 14282 504692 14288
rect 504364 13524 504416 13530
rect 504364 13466 504416 13472
rect 504272 12844 504324 12850
rect 504272 12786 504324 12792
rect 504376 3262 504404 13466
rect 504744 7478 504772 16374
rect 505388 11422 505416 16388
rect 505572 16374 505770 16402
rect 505376 11416 505428 11422
rect 505376 11358 505428 11364
rect 505572 11234 505600 16374
rect 506216 14482 506244 16388
rect 506204 14476 506256 14482
rect 506204 14418 506256 14424
rect 505296 11206 505600 11234
rect 504824 7608 504876 7614
rect 504824 7550 504876 7556
rect 504732 7472 504784 7478
rect 504732 7414 504784 7420
rect 504364 3256 504416 3262
rect 504364 3198 504416 3204
rect 504836 480 504864 7550
rect 505296 3602 505324 11206
rect 506388 10940 506440 10946
rect 506388 10882 506440 10888
rect 505284 3596 505336 3602
rect 505284 3538 505336 3544
rect 506400 626 506428 10882
rect 506584 7410 506612 16388
rect 506952 14210 506980 16388
rect 506940 14204 506992 14210
rect 506940 14146 506992 14152
rect 507320 11762 507348 16388
rect 507308 11756 507360 11762
rect 507308 11698 507360 11704
rect 507688 10334 507716 16388
rect 507768 14476 507820 14482
rect 507768 14418 507820 14424
rect 507676 10328 507728 10334
rect 507676 10270 507728 10276
rect 506572 7404 506624 7410
rect 506572 7346 506624 7352
rect 507780 3534 507808 14418
rect 507216 3528 507268 3534
rect 507216 3470 507268 3476
rect 507768 3528 507820 3534
rect 507768 3470 507820 3476
rect 506032 598 506428 626
rect 506032 480 506060 598
rect 507228 480 507256 3470
rect 508056 2106 508084 16388
rect 508516 9042 508544 16388
rect 508504 9036 508556 9042
rect 508504 8978 508556 8984
rect 508884 7342 508912 16388
rect 509148 11008 509200 11014
rect 509148 10950 509200 10956
rect 509160 10810 509188 10950
rect 509252 10878 509280 16388
rect 509240 10872 509292 10878
rect 509240 10814 509292 10820
rect 509148 10804 509200 10810
rect 509148 10746 509200 10752
rect 509240 9648 509292 9654
rect 509240 9590 509292 9596
rect 508872 7336 508924 7342
rect 508872 7278 508924 7284
rect 508412 5432 508464 5438
rect 508412 5374 508464 5380
rect 508044 2100 508096 2106
rect 508044 2042 508096 2048
rect 508424 480 508452 5374
rect 509252 4078 509280 9590
rect 509620 8702 509648 16388
rect 509988 13122 510016 16388
rect 509976 13116 510028 13122
rect 509976 13058 510028 13064
rect 509608 8696 509660 8702
rect 509608 8638 509660 8644
rect 510356 8022 510384 16388
rect 510620 9444 510672 9450
rect 510620 9386 510672 9392
rect 510344 8016 510396 8022
rect 510344 7958 510396 7964
rect 509608 7880 509660 7886
rect 509608 7822 509660 7828
rect 509240 4072 509292 4078
rect 509240 4014 509292 4020
rect 509620 480 509648 7822
rect 510632 3874 510660 9386
rect 510816 8974 510844 16388
rect 511184 9110 511212 16388
rect 511552 13462 511580 16388
rect 511828 16374 511934 16402
rect 511540 13456 511592 13462
rect 511540 13398 511592 13404
rect 511172 9104 511224 9110
rect 511172 9046 511224 9052
rect 510804 8968 510856 8974
rect 510804 8910 510856 8916
rect 511828 8838 511856 16374
rect 511908 14952 511960 14958
rect 511908 14894 511960 14900
rect 510804 8832 510856 8838
rect 510804 8774 510856 8780
rect 511816 8832 511868 8838
rect 511816 8774 511868 8780
rect 510816 4826 510844 8774
rect 510804 4820 510856 4826
rect 510804 4762 510856 4768
rect 510620 3868 510672 3874
rect 510620 3810 510672 3816
rect 511920 3534 511948 14894
rect 512092 11688 512144 11694
rect 512092 11630 512144 11636
rect 512104 4894 512132 11630
rect 512288 9246 512316 16388
rect 512656 14550 512684 16388
rect 512932 16374 513130 16402
rect 512644 14544 512696 14550
rect 512644 14486 512696 14492
rect 512932 11694 512960 16374
rect 512920 11688 512972 11694
rect 512920 11630 512972 11636
rect 512276 9240 512328 9246
rect 512276 9182 512328 9188
rect 513484 9178 513512 16388
rect 513852 13394 513880 16388
rect 514036 16374 514234 16402
rect 513840 13388 513892 13394
rect 513840 13330 513892 13336
rect 514036 11642 514064 16374
rect 513576 11614 514064 11642
rect 513472 9172 513524 9178
rect 513472 9114 513524 9120
rect 513196 8968 513248 8974
rect 513196 8910 513248 8916
rect 512092 4888 512144 4894
rect 512092 4830 512144 4836
rect 512000 4820 512052 4826
rect 512000 4762 512052 4768
rect 510804 3528 510856 3534
rect 510804 3470 510856 3476
rect 511908 3528 511960 3534
rect 511908 3470 511960 3476
rect 510816 480 510844 3470
rect 512012 480 512040 4762
rect 513208 480 513236 8910
rect 513576 5506 513604 11614
rect 514588 9314 514616 16388
rect 514956 10538 514984 16388
rect 514944 10532 514996 10538
rect 514944 10474 514996 10480
rect 515416 10402 515444 16388
rect 515404 10396 515456 10402
rect 515404 10338 515456 10344
rect 515784 9994 515812 16388
rect 516152 13530 516180 16388
rect 516336 16374 516534 16402
rect 516140 13524 516192 13530
rect 516140 13466 516192 13472
rect 515772 9988 515824 9994
rect 515772 9930 515824 9936
rect 514576 9308 514628 9314
rect 514576 9250 514628 9256
rect 514668 9308 514720 9314
rect 514668 9250 514720 9256
rect 513564 5500 513616 5506
rect 513564 5442 513616 5448
rect 514392 3596 514444 3602
rect 514392 3538 514444 3544
rect 514404 480 514432 3538
rect 514680 3534 514708 9250
rect 516336 4962 516364 16374
rect 516888 9382 516916 16388
rect 517256 9654 517284 16388
rect 517624 16374 517730 16402
rect 517428 13116 517480 13122
rect 517428 13058 517480 13064
rect 517244 9648 517296 9654
rect 517244 9590 517296 9596
rect 516876 9376 516928 9382
rect 516876 9318 516928 9324
rect 516324 4956 516376 4962
rect 516324 4898 516376 4904
rect 515588 4888 515640 4894
rect 515588 4830 515640 4836
rect 514668 3528 514720 3534
rect 514668 3470 514720 3476
rect 515600 480 515628 4830
rect 517440 4146 517468 13058
rect 517624 5030 517652 16374
rect 518084 10470 518112 16388
rect 518452 11354 518480 16388
rect 518636 16374 518834 16402
rect 518912 16374 519202 16402
rect 518440 11348 518492 11354
rect 518440 11290 518492 11296
rect 518072 10464 518124 10470
rect 518072 10406 518124 10412
rect 518636 5098 518664 16374
rect 518912 10606 518940 16374
rect 518900 10600 518952 10606
rect 518900 10542 518952 10548
rect 519556 9314 519584 16388
rect 519648 16374 520030 16402
rect 520292 16374 520398 16402
rect 519544 9308 519596 9314
rect 519544 9250 519596 9256
rect 519084 9036 519136 9042
rect 519084 8978 519136 8984
rect 518624 5092 518676 5098
rect 518624 5034 518676 5040
rect 517612 5024 517664 5030
rect 517612 4966 517664 4972
rect 516784 4140 516836 4146
rect 516784 4082 516836 4088
rect 517428 4140 517480 4146
rect 517428 4082 517480 4088
rect 516796 480 516824 4082
rect 517888 3868 517940 3874
rect 517888 3810 517940 3816
rect 517900 480 517928 3810
rect 519096 480 519124 8978
rect 519648 5166 519676 16374
rect 520292 10674 520320 16374
rect 520752 14890 520780 16388
rect 520936 16374 521134 16402
rect 521212 16374 521502 16402
rect 520740 14884 520792 14890
rect 520740 14826 520792 14832
rect 520280 10668 520332 10674
rect 520280 10610 520332 10616
rect 520280 9172 520332 9178
rect 520280 9114 520332 9120
rect 519636 5160 519688 5166
rect 519636 5102 519688 5108
rect 520292 480 520320 9114
rect 520936 5234 520964 16374
rect 521212 6186 521240 16374
rect 521856 9450 521884 16388
rect 522040 16374 522330 16402
rect 522408 16374 522698 16402
rect 521844 9444 521896 9450
rect 521844 9386 521896 9392
rect 521200 6180 521252 6186
rect 521200 6122 521252 6128
rect 522040 5302 522068 16374
rect 522408 6254 522436 16374
rect 523052 14686 523080 16388
rect 523144 16374 523434 16402
rect 523040 14680 523092 14686
rect 523040 14622 523092 14628
rect 522672 10328 522724 10334
rect 522672 10270 522724 10276
rect 522396 6248 522448 6254
rect 522396 6190 522448 6196
rect 522028 5296 522080 5302
rect 522028 5238 522080 5244
rect 520924 5228 520976 5234
rect 520924 5170 520976 5176
rect 521476 3664 521528 3670
rect 521476 3606 521528 3612
rect 521488 480 521516 3606
rect 522684 480 522712 10270
rect 523144 5370 523172 16374
rect 523788 11830 523816 16388
rect 523880 16374 524170 16402
rect 523776 11824 523828 11830
rect 523776 11766 523828 11772
rect 523132 5364 523184 5370
rect 523132 5306 523184 5312
rect 523880 3754 523908 16374
rect 523960 14408 524012 14414
rect 523960 14350 524012 14356
rect 523972 4010 524000 14350
rect 524616 4554 524644 16388
rect 524984 11898 525012 16388
rect 525064 15156 525116 15162
rect 525064 15098 525116 15104
rect 524972 11892 525024 11898
rect 524972 11834 525024 11840
rect 524604 4548 524656 4554
rect 524604 4490 524656 4496
rect 525076 4298 525104 15098
rect 525352 14278 525380 16388
rect 525444 16374 525734 16402
rect 525340 14272 525392 14278
rect 525340 14214 525392 14220
rect 525444 11966 525472 16374
rect 525708 14544 525760 14550
rect 525708 14486 525760 14492
rect 525432 11960 525484 11966
rect 525432 11902 525484 11908
rect 524984 4270 525104 4298
rect 523960 4004 524012 4010
rect 523960 3946 524012 3952
rect 523788 3726 523908 3754
rect 523788 3330 523816 3726
rect 523868 3596 523920 3602
rect 523868 3538 523920 3544
rect 523776 3324 523828 3330
rect 523776 3266 523828 3272
rect 523880 480 523908 3538
rect 524984 3466 525012 4270
rect 525720 4146 525748 14486
rect 526088 12034 526116 16388
rect 526272 16374 526470 16402
rect 526640 16374 526930 16402
rect 526076 12028 526128 12034
rect 526076 11970 526128 11976
rect 525064 4140 525116 4146
rect 525064 4082 525116 4088
rect 525708 4140 525760 4146
rect 525708 4082 525760 4088
rect 524972 3460 525024 3466
rect 524972 3402 525024 3408
rect 525076 480 525104 4082
rect 526272 3942 526300 16374
rect 526444 11756 526496 11762
rect 526444 11698 526496 11704
rect 526260 3936 526312 3942
rect 526260 3878 526312 3884
rect 526456 3602 526484 11698
rect 526640 6322 526668 16374
rect 527284 12102 527312 16388
rect 527652 14754 527680 16388
rect 527744 16374 528034 16402
rect 527640 14748 527692 14754
rect 527640 14690 527692 14696
rect 527272 12096 527324 12102
rect 527272 12038 527324 12044
rect 527744 6390 527772 16374
rect 527916 15088 527968 15094
rect 527916 15030 527968 15036
rect 527824 14884 527876 14890
rect 527824 14826 527876 14832
rect 527732 6384 527784 6390
rect 527732 6326 527784 6332
rect 526628 6316 526680 6322
rect 526628 6258 526680 6264
rect 527456 4140 527508 4146
rect 527456 4082 527508 4088
rect 526444 3596 526496 3602
rect 526444 3538 526496 3544
rect 526260 3460 526312 3466
rect 526260 3402 526312 3408
rect 526272 480 526300 3402
rect 527468 480 527496 4082
rect 527836 3874 527864 14826
rect 527824 3868 527876 3874
rect 527824 3810 527876 3816
rect 527928 3738 527956 15030
rect 528388 10742 528416 16388
rect 528756 14822 528784 16388
rect 528744 14816 528796 14822
rect 528744 14758 528796 14764
rect 528468 14680 528520 14686
rect 528468 14622 528520 14628
rect 528376 10736 528428 10742
rect 528376 10678 528428 10684
rect 528480 4146 528508 14622
rect 528652 14408 528704 14414
rect 528652 14350 528704 14356
rect 528664 6458 528692 14350
rect 529216 12170 529244 16388
rect 529308 16374 529598 16402
rect 529308 14414 529336 16374
rect 529296 14408 529348 14414
rect 529296 14350 529348 14356
rect 529204 12164 529256 12170
rect 529204 12106 529256 12112
rect 529848 11824 529900 11830
rect 529848 11766 529900 11772
rect 528652 6452 528704 6458
rect 528652 6394 528704 6400
rect 528468 4140 528520 4146
rect 528468 4082 528520 4088
rect 527916 3732 527968 3738
rect 527916 3674 527968 3680
rect 528652 3188 528704 3194
rect 528652 3130 528704 3136
rect 528664 480 528692 3130
rect 529860 480 529888 11766
rect 529952 7682 529980 16388
rect 530320 10878 530348 16388
rect 530584 15020 530636 15026
rect 530584 14962 530636 14968
rect 530308 10872 530360 10878
rect 530308 10814 530360 10820
rect 530124 9716 530176 9722
rect 530124 9658 530176 9664
rect 529940 7676 529992 7682
rect 529940 7618 529992 7624
rect 530136 6526 530164 9658
rect 530124 6520 530176 6526
rect 530124 6462 530176 6468
rect 530596 3670 530624 14962
rect 530688 9722 530716 16388
rect 530676 9716 530728 9722
rect 530676 9658 530728 9664
rect 531056 7750 531084 16388
rect 531228 14748 531280 14754
rect 531228 14690 531280 14696
rect 531044 7744 531096 7750
rect 531044 7686 531096 7692
rect 530584 3664 530636 3670
rect 530584 3606 530636 3612
rect 531240 626 531268 14690
rect 531320 9308 531372 9314
rect 531320 9250 531372 9256
rect 531332 9178 531360 9250
rect 531320 9172 531372 9178
rect 531320 9114 531372 9120
rect 531516 7818 531544 16388
rect 531700 16374 531898 16402
rect 531504 7812 531556 7818
rect 531504 7754 531556 7760
rect 531700 6594 531728 16374
rect 531964 14816 532016 14822
rect 531964 14758 532016 14764
rect 531688 6588 531740 6594
rect 531688 6530 531740 6536
rect 531976 3194 532004 14758
rect 532252 14346 532280 16388
rect 532240 14340 532292 14346
rect 532240 14282 532292 14288
rect 532620 13190 532648 16388
rect 532896 16374 533002 16402
rect 534356 16390 534408 16396
rect 535000 16448 535052 16454
rect 535000 16390 535052 16396
rect 532608 13184 532660 13190
rect 532608 13126 532660 13132
rect 532896 6662 532924 16374
rect 533356 13326 533384 16388
rect 533344 13320 533396 13326
rect 533344 13262 533396 13268
rect 533816 13258 533844 16388
rect 533804 13252 533856 13258
rect 533804 13194 533856 13200
rect 533988 13184 534040 13190
rect 533988 13126 534040 13132
rect 532884 6656 532936 6662
rect 532884 6598 532936 6604
rect 534000 4146 534028 13126
rect 534184 6730 534212 16388
rect 534368 6798 534396 16390
rect 534552 15162 534580 16388
rect 534540 15156 534592 15162
rect 534540 15098 534592 15104
rect 534920 12238 534948 16388
rect 535368 15156 535420 15162
rect 535368 15098 535420 15104
rect 534908 12232 534960 12238
rect 534908 12174 534960 12180
rect 534356 6792 534408 6798
rect 534356 6734 534408 6740
rect 534172 6724 534224 6730
rect 534172 6666 534224 6672
rect 535276 5636 535328 5642
rect 535276 5578 535328 5584
rect 533436 4140 533488 4146
rect 533436 4082 533488 4088
rect 533988 4140 534040 4146
rect 533988 4082 534040 4088
rect 532240 3324 532292 3330
rect 532240 3266 532292 3272
rect 531964 3188 532016 3194
rect 531964 3130 532016 3136
rect 531056 598 531268 626
rect 531056 480 531084 598
rect 532252 480 532280 3266
rect 533448 480 533476 4082
rect 534540 3528 534592 3534
rect 534540 3470 534592 3476
rect 534552 480 534580 3470
rect 535288 3466 535316 5578
rect 535380 3534 535408 15098
rect 535656 14618 535684 16388
rect 535840 16374 536130 16402
rect 535644 14612 535696 14618
rect 535644 14554 535696 14560
rect 535840 7614 535868 16374
rect 536104 14408 536156 14414
rect 536104 14350 536156 14356
rect 535828 7608 535880 7614
rect 535828 7550 535880 7556
rect 535736 4004 535788 4010
rect 535736 3946 535788 3952
rect 535368 3528 535420 3534
rect 535368 3470 535420 3476
rect 535276 3460 535328 3466
rect 535276 3402 535328 3408
rect 535748 480 535776 3946
rect 536116 3330 536144 14350
rect 536484 10946 536512 16388
rect 536748 14612 536800 14618
rect 536748 14554 536800 14560
rect 536472 10940 536524 10946
rect 536472 10882 536524 10888
rect 536760 4010 536788 14554
rect 536852 14482 536880 16388
rect 537036 16374 537234 16402
rect 536840 14476 536892 14482
rect 536840 14418 536892 14424
rect 537036 5438 537064 16374
rect 537588 7886 537616 16388
rect 537956 14958 537984 16388
rect 537944 14952 537996 14958
rect 537944 14894 537996 14900
rect 538128 14476 538180 14482
rect 538128 14418 538180 14424
rect 537576 7880 537628 7886
rect 537576 7822 537628 7828
rect 537024 5432 537076 5438
rect 537024 5374 537076 5380
rect 536748 4004 536800 4010
rect 536748 3946 536800 3952
rect 536932 3596 536984 3602
rect 536932 3538 536984 3544
rect 536104 3324 536156 3330
rect 536104 3266 536156 3272
rect 536944 480 536972 3538
rect 538140 480 538168 14418
rect 538416 4826 538444 16388
rect 538784 8974 538812 16388
rect 539152 15094 539180 16388
rect 539244 16374 539534 16402
rect 539140 15088 539192 15094
rect 539140 15030 539192 15036
rect 538772 8968 538824 8974
rect 538772 8910 538824 8916
rect 539244 4894 539272 16374
rect 539888 13122 539916 16388
rect 540256 14890 540284 16388
rect 540244 14884 540296 14890
rect 540244 14826 540296 14832
rect 539876 13116 539928 13122
rect 539876 13058 539928 13064
rect 540716 9042 540744 16388
rect 541084 9314 541112 16388
rect 541452 15026 541480 16388
rect 541440 15020 541492 15026
rect 541440 14962 541492 14968
rect 541820 10334 541848 16388
rect 542188 11762 542216 16388
rect 542556 14550 542584 16388
rect 542740 16374 543030 16402
rect 542544 14544 542596 14550
rect 542544 14486 542596 14492
rect 542176 11756 542228 11762
rect 542176 11698 542228 11704
rect 541808 10328 541860 10334
rect 541808 10270 541860 10276
rect 540888 9308 540940 9314
rect 540888 9250 540940 9256
rect 541072 9308 541124 9314
rect 541072 9250 541124 9256
rect 540900 9110 540928 9250
rect 540888 9104 540940 9110
rect 540888 9046 540940 9052
rect 540704 9036 540756 9042
rect 540704 8978 540756 8984
rect 542740 5642 542768 16374
rect 543384 14686 543412 16388
rect 543752 14822 543780 16388
rect 543740 14816 543792 14822
rect 543740 14758 543792 14764
rect 543372 14680 543424 14686
rect 543372 14622 543424 14628
rect 543648 14204 543700 14210
rect 543648 14146 543700 14152
rect 542728 5636 542780 5642
rect 542728 5578 542780 5584
rect 539232 4888 539284 4894
rect 539232 4830 539284 4836
rect 538404 4820 538456 4826
rect 538404 4762 538456 4768
rect 543660 4146 543688 14146
rect 544120 11830 544148 16388
rect 544488 14754 544516 16388
rect 544476 14748 544528 14754
rect 544476 14690 544528 14696
rect 544856 14414 544884 16388
rect 544844 14408 544896 14414
rect 544844 14350 544896 14356
rect 545028 14136 545080 14142
rect 545028 14078 545080 14084
rect 544384 13932 544436 13938
rect 544384 13874 544436 13880
rect 544108 11824 544160 11830
rect 544108 11766 544160 11772
rect 542912 4140 542964 4146
rect 542912 4082 542964 4088
rect 543648 4140 543700 4146
rect 543648 4082 543700 4088
rect 539324 3460 539376 3466
rect 539324 3402 539376 3408
rect 539336 480 539364 3402
rect 540520 3256 540572 3262
rect 540520 3198 540572 3204
rect 540532 480 540560 3198
rect 541716 2916 541768 2922
rect 541716 2858 541768 2864
rect 541728 480 541756 2858
rect 542924 480 542952 4082
rect 544396 3602 544424 13874
rect 544384 3596 544436 3602
rect 544384 3538 544436 3544
rect 545040 3534 545068 14078
rect 545316 13190 545344 16388
rect 545684 15162 545712 16388
rect 545672 15156 545724 15162
rect 545672 15098 545724 15104
rect 546052 14618 546080 16388
rect 546040 14612 546092 14618
rect 546040 14554 546092 14560
rect 546316 14068 546368 14074
rect 546316 14010 546368 14016
rect 545764 13864 545816 13870
rect 545764 13806 545816 13812
rect 545304 13184 545356 13190
rect 545304 13126 545356 13132
rect 544108 3528 544160 3534
rect 544108 3470 544160 3476
rect 545028 3528 545080 3534
rect 545028 3470 545080 3476
rect 545304 3528 545356 3534
rect 545304 3470 545356 3476
rect 544120 480 544148 3470
rect 545316 480 545344 3470
rect 545776 3466 545804 13806
rect 546328 3534 546356 14010
rect 546420 13938 546448 16388
rect 546788 14482 546816 16388
rect 546776 14476 546828 14482
rect 546776 14418 546828 14424
rect 546408 13932 546460 13938
rect 546408 13874 546460 13880
rect 547156 13870 547184 16388
rect 547340 16374 547630 16402
rect 547998 16374 548104 16402
rect 547144 13864 547196 13870
rect 547144 13806 547196 13812
rect 547340 11642 547368 16374
rect 547696 14000 547748 14006
rect 547696 13942 547748 13948
rect 546604 11614 547368 11642
rect 546316 3528 546368 3534
rect 546316 3470 546368 3476
rect 545764 3460 545816 3466
rect 545764 3402 545816 3408
rect 546500 3392 546552 3398
rect 546500 3334 546552 3340
rect 546512 480 546540 3334
rect 546604 3262 546632 11614
rect 546592 3256 546644 3262
rect 546592 3198 546644 3204
rect 547708 480 547736 13942
rect 547788 13932 547840 13938
rect 547788 13874 547840 13880
rect 547800 3398 547828 13874
rect 547788 3392 547840 3398
rect 547788 3334 547840 3340
rect 548076 2922 548104 16374
rect 548352 14210 548380 16388
rect 548340 14204 548392 14210
rect 548340 14146 548392 14152
rect 548720 14142 548748 16388
rect 548708 14136 548760 14142
rect 548708 14078 548760 14084
rect 549088 14074 549116 16388
rect 549076 14068 549128 14074
rect 549076 14010 549128 14016
rect 549456 13938 549484 16388
rect 549916 14006 549944 16388
rect 549904 14000 549956 14006
rect 549904 13942 549956 13948
rect 549444 13932 549496 13938
rect 549444 13874 549496 13880
rect 550284 13870 550312 16388
rect 549168 13864 549220 13870
rect 549168 13806 549220 13812
rect 550272 13864 550324 13870
rect 550652 13818 550680 16388
rect 550272 13806 550324 13812
rect 548064 2916 548116 2922
rect 548064 2858 548116 2864
rect 549180 626 549208 13806
rect 550560 13790 550680 13818
rect 550836 16374 551034 16402
rect 550560 3534 550588 13790
rect 550088 3528 550140 3534
rect 550088 3470 550140 3476
rect 550548 3528 550600 3534
rect 550548 3470 550600 3476
rect 548904 598 549208 626
rect 548904 480 548932 598
rect 550100 480 550128 3470
rect 550836 626 550864 16374
rect 551388 13938 551416 16388
rect 551376 13932 551428 13938
rect 551376 13874 551428 13880
rect 551756 13870 551784 16388
rect 552216 14142 552244 16388
rect 552204 14136 552256 14142
rect 552204 14078 552256 14084
rect 552584 13938 552612 16388
rect 552952 14074 552980 16388
rect 552940 14068 552992 14074
rect 552940 14010 552992 14016
rect 553320 14006 553348 16388
rect 553688 14346 553716 16388
rect 553676 14340 553728 14346
rect 553676 14282 553728 14288
rect 554056 14278 554084 16388
rect 554044 14272 554096 14278
rect 554044 14214 554096 14220
rect 554516 14210 554544 16388
rect 554884 14618 554912 16388
rect 554872 14612 554924 14618
rect 554872 14554 554924 14560
rect 555252 14550 555280 16388
rect 555620 14686 555648 16388
rect 556002 16374 556108 16402
rect 555608 14680 555660 14686
rect 555608 14622 555660 14628
rect 555240 14544 555292 14550
rect 555240 14486 555292 14492
rect 554504 14204 554556 14210
rect 554504 14146 554556 14152
rect 555240 14136 555292 14142
rect 555240 14078 555292 14084
rect 553308 14000 553360 14006
rect 553308 13942 553360 13948
rect 551836 13932 551888 13938
rect 551836 13874 551888 13880
rect 552572 13932 552624 13938
rect 552572 13874 552624 13880
rect 554872 13932 554924 13938
rect 554872 13874 554924 13880
rect 551744 13864 551796 13870
rect 551744 13806 551796 13812
rect 551848 3534 551876 13874
rect 553400 13864 553452 13870
rect 553400 13806 553452 13812
rect 551836 3528 551888 3534
rect 551836 3470 551888 3476
rect 552388 3528 552440 3534
rect 552388 3470 552440 3476
rect 550836 598 551232 626
rect 551204 480 551232 598
rect 552400 480 552428 3470
rect 553412 626 553440 13806
rect 554884 3602 554912 13874
rect 554872 3596 554924 3602
rect 554872 3538 554924 3544
rect 555252 3380 555280 14078
rect 555516 14068 555568 14074
rect 555516 14010 555568 14016
rect 555424 14000 555476 14006
rect 555424 13942 555476 13948
rect 554792 3352 555280 3380
rect 553412 598 553624 626
rect 553596 480 553624 598
rect 554792 480 554820 3352
rect 555436 2922 555464 13942
rect 555528 3534 555556 14010
rect 555976 3596 556028 3602
rect 555976 3538 556028 3544
rect 555516 3528 555568 3534
rect 555516 3470 555568 3476
rect 555424 2916 555476 2922
rect 555424 2858 555476 2864
rect 555988 480 556016 3538
rect 556080 3398 556108 16374
rect 556356 13870 556384 16388
rect 556620 14272 556672 14278
rect 556620 14214 556672 14220
rect 556344 13864 556396 13870
rect 556344 13806 556396 13812
rect 556632 11642 556660 14214
rect 556816 11762 556844 16388
rect 557198 16374 557396 16402
rect 556988 14340 557040 14346
rect 556988 14282 557040 14288
rect 556896 14204 556948 14210
rect 556896 14146 556948 14152
rect 556804 11756 556856 11762
rect 556804 11698 556856 11704
rect 556632 11614 556844 11642
rect 556816 3466 556844 11614
rect 556908 3602 556936 14146
rect 557000 3874 557028 14282
rect 557264 13864 557316 13870
rect 557264 13806 557316 13812
rect 556988 3868 557040 3874
rect 556988 3810 557040 3816
rect 556896 3596 556948 3602
rect 556896 3538 556948 3544
rect 557172 3528 557224 3534
rect 557172 3470 557224 3476
rect 556804 3460 556856 3466
rect 556804 3402 556856 3408
rect 556068 3392 556120 3398
rect 556068 3334 556120 3340
rect 557184 480 557212 3470
rect 557276 3330 557304 13806
rect 557368 4078 557396 16374
rect 557552 13938 557580 16388
rect 557920 14482 557948 16388
rect 557908 14476 557960 14482
rect 557908 14418 557960 14424
rect 557540 13932 557592 13938
rect 557540 13874 557592 13880
rect 558288 13870 558316 16388
rect 558276 13864 558328 13870
rect 558276 13806 558328 13812
rect 557356 4072 557408 4078
rect 557356 4014 557408 4020
rect 558656 3942 558684 16388
rect 559116 13938 559144 16388
rect 558736 13932 558788 13938
rect 558736 13874 558788 13880
rect 559104 13932 559156 13938
rect 559104 13874 559156 13880
rect 558748 4146 558776 13874
rect 559484 13870 559512 16388
rect 559852 14006 559880 16388
rect 559944 16374 560234 16402
rect 559840 14000 559892 14006
rect 559840 13942 559892 13948
rect 558828 13864 558880 13870
rect 558828 13806 558880 13812
rect 559472 13864 559524 13870
rect 559472 13806 559524 13812
rect 558736 4140 558788 4146
rect 558736 4082 558788 4088
rect 558840 4010 558868 13806
rect 558828 4004 558880 4010
rect 558828 3946 558880 3952
rect 558644 3936 558696 3942
rect 558644 3878 558696 3884
rect 559564 3868 559616 3874
rect 559564 3810 559616 3816
rect 557264 3324 557316 3330
rect 557264 3266 557316 3272
rect 558368 2916 558420 2922
rect 558368 2858 558420 2864
rect 558380 480 558408 2858
rect 559576 480 559604 3810
rect 559944 3194 559972 16374
rect 560208 14000 560260 14006
rect 560208 13942 560260 13948
rect 560024 13932 560076 13938
rect 560024 13874 560076 13880
rect 560036 3874 560064 13874
rect 560116 13864 560168 13870
rect 560116 13806 560168 13812
rect 560024 3868 560076 3874
rect 560024 3810 560076 3816
rect 560128 3806 560156 13806
rect 560116 3800 560168 3806
rect 560116 3742 560168 3748
rect 560220 3738 560248 13942
rect 560588 13870 560616 16388
rect 560970 16374 561536 16402
rect 560576 13864 560628 13870
rect 560576 13806 560628 13812
rect 560208 3732 560260 3738
rect 560208 3674 560260 3680
rect 560760 3528 560812 3534
rect 560760 3470 560812 3476
rect 559932 3188 559984 3194
rect 559932 3130 559984 3136
rect 560772 480 560800 3470
rect 561508 3466 561536 16374
rect 561680 14680 561732 14686
rect 561680 14622 561732 14628
rect 561588 13864 561640 13870
rect 561588 13806 561640 13812
rect 561600 3670 561628 13806
rect 561692 12850 561720 14622
rect 563152 14612 563204 14618
rect 563152 14554 563204 14560
rect 563060 14544 563112 14550
rect 563060 14486 563112 14492
rect 561680 12844 561732 12850
rect 561680 12786 561732 12792
rect 561588 3664 561640 3670
rect 561588 3606 561640 3612
rect 561956 3596 562008 3602
rect 561956 3538 562008 3544
rect 561496 3460 561548 3466
rect 561496 3402 561548 3408
rect 561968 480 561996 3538
rect 563072 3534 563100 14486
rect 563060 3528 563112 3534
rect 563060 3470 563112 3476
rect 563164 480 563192 14554
rect 563716 3602 563744 38655
rect 580920 29345 580948 76191
rect 580906 29336 580962 29345
rect 580906 29271 580962 29280
rect 570604 14476 570656 14482
rect 570604 14418 570656 14424
rect 564440 12844 564492 12850
rect 564440 12786 564492 12792
rect 563704 3596 563756 3602
rect 563704 3538 563756 3544
rect 564348 3528 564400 3534
rect 564348 3470 564400 3476
rect 564360 480 564388 3470
rect 564452 610 564480 12786
rect 568580 11756 568632 11762
rect 568580 11698 568632 11704
rect 568592 3482 568620 11698
rect 570616 5574 570644 14418
rect 570604 5568 570656 5574
rect 570604 5510 570656 5516
rect 572628 5568 572680 5574
rect 572628 5510 572680 5516
rect 571432 4140 571484 4146
rect 571432 4082 571484 4088
rect 570236 4072 570288 4078
rect 570236 4014 570288 4020
rect 564532 3460 564584 3466
rect 568592 3454 569080 3482
rect 564532 3402 564584 3408
rect 564544 3194 564572 3402
rect 566740 3392 566792 3398
rect 566740 3334 566792 3340
rect 564532 3188 564584 3194
rect 564532 3130 564584 3136
rect 564440 604 564492 610
rect 564440 546 564492 552
rect 565544 604 565596 610
rect 565544 546 565596 552
rect 565556 480 565584 546
rect 566752 480 566780 3334
rect 567844 3324 567896 3330
rect 567844 3266 567896 3272
rect 567856 480 567884 3266
rect 569052 480 569080 3454
rect 570248 480 570276 4014
rect 571444 480 571472 4082
rect 572640 480 572668 5510
rect 573824 4004 573876 4010
rect 573824 3946 573876 3952
rect 573836 480 573864 3946
rect 575020 3936 575072 3942
rect 575020 3878 575072 3884
rect 575032 480 575060 3878
rect 576216 3868 576268 3874
rect 576216 3810 576268 3816
rect 576228 480 576256 3810
rect 577412 3800 577464 3806
rect 577412 3742 577464 3748
rect 577424 480 577452 3742
rect 578608 3732 578660 3738
rect 578608 3674 578660 3680
rect 578620 480 578648 3674
rect 581000 3664 581052 3670
rect 581000 3606 581052 3612
rect 579804 3460 579856 3466
rect 579804 3402 579856 3408
rect 579816 480 579844 3402
rect 581012 480 581040 3606
rect 583392 3596 583444 3602
rect 583392 3538 583444 3544
rect 582196 3528 582248 3534
rect 582196 3470 582248 3476
rect 582208 480 582236 3470
rect 583404 480 583432 3538
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3514 682216 3570 682272
rect 3054 653520 3110 653576
rect 3422 624824 3478 624880
rect 3330 610408 3386 610464
rect 3146 553016 3202 553072
rect 2870 509904 2926 509960
rect 3514 595992 3570 596048
rect 3514 567296 3570 567352
rect 3514 538600 3570 538656
rect 3514 495508 3570 495544
rect 3514 495488 3516 495508
rect 3516 495488 3568 495508
rect 3568 495488 3570 495508
rect 3146 481072 3202 481128
rect 3422 452376 3478 452432
rect 3514 437960 3570 438016
rect 3422 423700 3478 423736
rect 3422 423680 3424 423700
rect 3424 423680 3476 423700
rect 3476 423680 3478 423700
rect 4802 394984 4858 395040
rect 2778 380568 2834 380624
rect 2778 366152 2834 366208
rect 3146 337456 3202 337512
rect 2778 323040 2834 323096
rect 2778 309032 2834 309088
rect 3422 309032 3478 309088
rect 2778 308760 2834 308816
rect 3422 294344 3478 294400
rect 2778 280064 2834 280120
rect 2778 265648 2834 265704
rect 2778 236952 2834 237008
rect 2778 222536 2834 222592
rect 2778 193840 2834 193896
rect 2778 179424 2834 179480
rect 4802 173712 4858 173768
rect 2778 150728 2834 150784
rect 2778 136312 2834 136368
rect 2778 107616 2834 107672
rect 2778 93200 2834 93256
rect 6182 65456 6238 65512
rect 2778 64504 2834 64560
rect 2778 50088 2834 50144
rect 72974 700304 73030 700360
rect 30194 617752 30250 617808
rect 28630 616936 28686 616992
rect 28630 616564 28632 616584
rect 28632 616564 28684 616584
rect 28684 616564 28686 616584
rect 28630 616528 28686 616564
rect 30286 617616 30342 617672
rect 91098 619520 91154 619576
rect 95882 619520 95938 619576
rect 31482 617500 31538 617536
rect 31482 617480 31484 617500
rect 31484 617480 31536 617500
rect 31536 617480 31538 617500
rect 28630 615848 28686 615904
rect 27526 608912 27582 608968
rect 27434 607688 27490 607744
rect 25226 606600 25282 606656
rect 27342 602384 27398 602440
rect 24766 601704 24822 601760
rect 24674 583752 24730 583808
rect 24582 572872 24638 572928
rect 24490 572328 24546 572384
rect 24122 571920 24178 571976
rect 27250 599936 27306 599992
rect 25778 598712 25834 598768
rect 25226 596400 25282 596456
rect 25134 582528 25190 582584
rect 25042 577088 25098 577144
rect 24950 575320 25006 575376
rect 25318 587696 25374 587752
rect 25686 580760 25742 580816
rect 25410 578312 25466 578368
rect 25318 570560 25374 570616
rect 25502 574096 25558 574152
rect 25594 571784 25650 571840
rect 27158 597488 27214 597544
rect 27066 595176 27122 595232
rect 26054 591504 26110 591560
rect 25962 586744 26018 586800
rect 25870 583072 25926 583128
rect 26974 590280 27030 590336
rect 26882 585520 26938 585576
rect 26146 584976 26202 585032
rect 26606 580080 26662 580136
rect 26146 578856 26202 578912
rect 26330 573552 26386 573608
rect 26698 577768 26754 577824
rect 26790 576544 26846 576600
rect 27986 603744 28042 603800
rect 27618 603608 27674 603664
rect 27710 596944 27766 597000
rect 27802 593272 27858 593328
rect 27894 590688 27950 590744
rect 28354 604832 28410 604888
rect 28538 600072 28594 600128
rect 28446 598984 28502 599040
rect 28354 596672 28410 596728
rect 28262 595312 28318 595368
rect 28170 593408 28226 593464
rect 28078 591640 28134 591696
rect 28078 581440 28134 581496
rect 28354 594632 28410 594688
rect 28354 591912 28410 591968
rect 28354 588648 28410 588704
rect 28262 578992 28318 579048
rect 28262 575612 28318 575648
rect 28262 575592 28264 575612
rect 28264 575592 28316 575612
rect 28316 575592 28318 575612
rect 28262 574232 28318 574288
rect 28630 598304 28686 598360
rect 28630 594088 28686 594144
rect 28538 593408 28594 593464
rect 28630 592320 28686 592376
rect 28538 591232 28594 591288
rect 28630 589328 28686 589384
rect 28538 588104 28594 588160
rect 28630 587696 28686 587752
rect 28630 587424 28686 587480
rect 28630 585656 28686 585712
rect 28630 583888 28686 583944
rect 28538 580896 28594 580952
rect 29090 567432 29146 567488
rect 29090 558320 29146 558376
rect 29182 547576 29238 547632
rect 29182 531528 29238 531584
rect 30010 557368 30066 557424
rect 30010 557096 30066 557152
rect 30470 540912 30526 540968
rect 30470 533568 30526 533624
rect 76010 570560 76066 570616
rect 70582 530848 70638 530904
rect 74906 531664 74962 531720
rect 219070 679088 219126 679144
rect 218978 676232 219034 676288
rect 279146 619520 279202 619576
rect 139582 594768 139638 594824
rect 78678 547032 78734 547088
rect 91006 534928 91062 534984
rect 88890 534792 88946 534848
rect 84566 533840 84622 533896
rect 83462 531800 83518 531856
rect 82450 530712 82506 530768
rect 86682 533704 86738 533760
rect 93214 534656 93270 534712
rect 92110 532616 92166 532672
rect 101770 533568 101826 533624
rect 94226 532480 94282 532536
rect 96434 532344 96490 532400
rect 95330 531256 95386 531312
rect 98550 532208 98606 532264
rect 97538 530576 97594 530632
rect 99654 532072 99710 532128
rect 100758 531936 100814 531992
rect 102874 533432 102930 533488
rect 103978 533296 104034 533352
rect 105082 531256 105138 531312
rect 106094 529896 106150 529952
rect 111522 531392 111578 531448
rect 114742 534112 114798 534168
rect 131946 534248 132002 534304
rect 129830 532752 129886 532808
rect 135258 531528 135314 531584
rect 138478 531664 138534 531720
rect 141698 534384 141754 534440
rect 157890 532888 157946 532944
rect 161110 533024 161166 533080
rect 182178 528400 182234 528456
rect 183926 528400 183982 528456
rect 175922 528264 175978 528320
rect 177946 528264 178002 528320
rect 181902 528264 181958 528320
rect 185950 528300 185952 528320
rect 185952 528300 186004 528320
rect 186004 528300 186006 528320
rect 185950 528264 186006 528300
rect 207570 528264 207626 528320
rect 251822 528420 251878 528456
rect 251822 528400 251824 528420
rect 251824 528400 251876 528420
rect 251876 528400 251878 528420
rect 251822 528264 251878 528320
rect 253846 528420 253902 528456
rect 253846 528400 253848 528420
rect 253848 528400 253900 528420
rect 253900 528400 253902 528420
rect 254306 528264 254362 528320
rect 207018 528216 207074 528218
rect 207018 528164 207020 528216
rect 207020 528164 207072 528216
rect 207072 528164 207074 528216
rect 207018 528162 207074 528164
rect 281538 515888 281594 515944
rect 3422 35844 3424 35864
rect 3424 35844 3476 35864
rect 3476 35844 3478 35864
rect 3422 35808 3478 35844
rect 2778 21392 2834 21448
rect 2778 7112 2834 7168
rect 12622 443536 12678 443592
rect 107198 500384 107254 500440
rect 107658 497528 107714 497584
rect 109038 497392 109094 497448
rect 110602 497800 110658 497856
rect 110418 497664 110474 497720
rect 114742 500656 114798 500712
rect 113638 500248 113694 500304
rect 112626 500112 112682 500168
rect 116858 500520 116914 500576
rect 114558 497936 114614 497992
rect 117962 500384 118018 500440
rect 124218 498072 124274 498128
rect 125598 497256 125654 497312
rect 130934 500792 130990 500848
rect 141698 500792 141754 500848
rect 142710 500656 142766 500712
rect 142710 499840 142766 499896
rect 143814 499704 143870 499760
rect 128358 497120 128414 497176
rect 154302 502288 154358 502344
rect 154394 502152 154450 502208
rect 153566 500792 153622 500848
rect 147034 499568 147090 499624
rect 148138 499568 148194 499624
rect 149242 499568 149298 499624
rect 150346 499568 150402 499624
rect 151358 499568 151414 499624
rect 152462 499568 152518 499624
rect 153198 497664 153254 497720
rect 146850 492632 146906 492688
rect 131026 401376 131082 401432
rect 129646 401240 129702 401296
rect 126886 401104 126942 401160
rect 125506 400968 125562 401024
rect 118606 400832 118662 400888
rect 78586 377304 78642 377360
rect 21362 357312 21418 357368
rect 114006 351736 114062 351792
rect 111706 351600 111762 351656
rect 110694 351464 110750 351520
rect 108670 351328 108726 351384
rect 107566 351056 107622 351112
rect 109590 351192 109646 351248
rect 117134 350920 117190 350976
rect 115110 350784 115166 350840
rect 122654 351736 122710 351792
rect 122654 350648 122710 350704
rect 142618 351192 142674 351248
rect 142802 351192 142858 351248
rect 142802 350920 142858 350976
rect 142618 350648 142674 350704
rect 147126 389408 147182 389464
rect 147126 386416 147182 386472
rect 147586 351872 147642 351928
rect 146942 351736 146998 351792
rect 147218 351736 147274 351792
rect 146298 350920 146354 350976
rect 147218 351464 147274 351520
rect 147678 351736 147734 351792
rect 148046 351736 148102 351792
rect 149426 351736 149482 351792
rect 150070 351736 150126 351792
rect 151174 351736 151230 351792
rect 152370 351736 152426 351792
rect 147678 351464 147734 351520
rect 147586 350512 147642 350568
rect 149058 350784 149114 350840
rect 153198 351328 153254 351384
rect 154210 492632 154266 492688
rect 155406 499704 155462 499760
rect 155866 482976 155922 483032
rect 155774 463664 155830 463720
rect 155682 405728 155738 405784
rect 155682 376624 155738 376680
rect 155774 369688 155830 369744
rect 156142 482976 156198 483032
rect 156050 465296 156106 465352
rect 156142 463664 156198 463720
rect 156142 405864 156198 405920
rect 185582 450880 185638 450936
rect 190182 500792 190238 500848
rect 191286 500792 191342 500848
rect 189078 500656 189134 500712
rect 280158 471280 280214 471336
rect 281538 430480 281594 430536
rect 282182 430480 282238 430536
rect 281630 421232 281686 421288
rect 189446 351736 189502 351792
rect 191194 351736 191250 351792
rect 189906 351600 189962 351656
rect 282182 335960 282238 336016
rect 17130 274896 17186 274952
rect 113178 295296 113234 295352
rect 113914 254496 113970 254552
rect 116398 221176 116454 221232
rect 116122 219952 116178 220008
rect 104806 219272 104862 219328
rect 116398 218864 116454 218920
rect 104806 217948 104808 217968
rect 104808 217948 104860 217968
rect 104860 217948 104862 217968
rect 104806 217912 104862 217948
rect 116398 217640 116454 217696
rect 104806 216588 104808 216608
rect 104808 216588 104860 216608
rect 104860 216588 104862 216608
rect 104806 216552 104862 216588
rect 115938 216552 115994 216608
rect 104806 215600 104862 215656
rect 116398 215348 116454 215384
rect 116398 215328 116400 215348
rect 116400 215328 116452 215348
rect 116452 215328 116454 215348
rect 104806 214648 104862 214704
rect 116398 214104 116454 214160
rect 104806 213424 104862 213480
rect 115938 213016 115994 213072
rect 104438 212064 104494 212120
rect 116306 211792 116362 211848
rect 104806 210840 104862 210896
rect 116306 210704 116362 210760
rect 104806 209480 104862 209536
rect 116030 209480 116086 209536
rect 115938 208256 115994 208312
rect 104806 208120 104862 208176
rect 104806 206916 104862 206952
rect 104806 206896 104808 206916
rect 104808 206896 104860 206916
rect 104860 206896 104862 206916
rect 116030 207168 116086 207224
rect 104714 206216 104770 206272
rect 115938 205944 115994 206000
rect 104806 204992 104862 205048
rect 116398 204856 116454 204912
rect 104806 203632 104862 203688
rect 116306 203632 116362 203688
rect 104806 202408 104862 202464
rect 116122 202408 116178 202464
rect 116122 201320 116178 201376
rect 104806 201048 104862 201104
rect 115938 200132 115940 200152
rect 115940 200132 115992 200152
rect 115992 200132 115994 200152
rect 104806 199824 104862 199880
rect 104806 198464 104862 198520
rect 115938 200096 115994 200132
rect 116398 199008 116454 199064
rect 116398 197784 116454 197840
rect 104806 197276 104808 197296
rect 104808 197276 104860 197296
rect 104860 197276 104862 197296
rect 104806 197240 104862 197276
rect 116398 196696 116454 196752
rect 104530 196560 104586 196616
rect 115938 195472 115994 195528
rect 104806 195336 104862 195392
rect 116122 194248 116178 194304
rect 104806 193976 104862 194032
rect 116398 193160 116454 193216
rect 104438 192752 104494 192808
rect 116030 191956 116086 191992
rect 116030 191936 116032 191956
rect 116032 191936 116084 191956
rect 116084 191936 116086 191956
rect 104806 191392 104862 191448
rect 116490 190848 116546 190904
rect 104714 190168 104770 190224
rect 116398 189624 116454 189680
rect 104806 188808 104862 188864
rect 104806 187448 104862 187504
rect 116214 188400 116270 188456
rect 116306 187312 116362 187368
rect 104806 186260 104808 186280
rect 104808 186260 104860 186280
rect 104860 186260 104862 186280
rect 104806 186224 104862 186260
rect 116030 186088 116086 186144
rect 104530 185544 104586 185600
rect 104806 184320 104862 184376
rect 104806 182960 104862 183016
rect 104806 181736 104862 181792
rect 116398 185020 116454 185056
rect 116398 185000 116400 185020
rect 116400 185000 116452 185020
rect 116452 185000 116454 185020
rect 116398 183776 116454 183832
rect 115938 182552 115994 182608
rect 115938 181464 115994 181520
rect 104806 180376 104862 180432
rect 116398 180240 116454 180296
rect 104806 179016 104862 179072
rect 115938 179152 115994 179208
rect 104162 177792 104218 177848
rect 104162 176432 104218 176488
rect 115938 177928 115994 177984
rect 116398 176840 116454 176896
rect 104806 175108 104808 175128
rect 104808 175108 104860 175128
rect 104860 175108 104862 175128
rect 104806 175072 104862 175108
rect 104438 174664 104494 174720
rect 116398 175616 116454 175672
rect 115938 174392 115994 174448
rect 104806 173304 104862 173360
rect 104438 172080 104494 172136
rect 116398 173304 116454 173360
rect 116122 172080 116178 172136
rect 104806 170720 104862 170776
rect 104162 168136 104218 168192
rect 116306 170992 116362 171048
rect 104806 169360 104862 169416
rect 104254 166912 104310 166968
rect 116398 169788 116454 169824
rect 116398 169768 116400 169788
rect 116400 169768 116452 169788
rect 116452 169768 116454 169788
rect 116398 168544 116454 168600
rect 115938 167456 115994 167512
rect 104806 165552 104862 165608
rect 104622 164872 104678 164928
rect 115938 166232 115994 166288
rect 116122 165144 116178 165200
rect 104806 163648 104862 163704
rect 104806 162288 104862 162344
rect 116398 163920 116454 163976
rect 116214 162696 116270 162752
rect 104806 160928 104862 160984
rect 103702 158616 103758 158672
rect 116398 161608 116454 161664
rect 116398 160384 116454 160440
rect 104806 159704 104862 159760
rect 116398 159296 116454 159352
rect 104254 157256 104310 157312
rect 116398 158072 116454 158128
rect 116030 156984 116086 157040
rect 104806 155896 104862 155952
rect 104346 154400 104402 154456
rect 104622 153856 104678 153912
rect 116030 155760 116086 155816
rect 116398 154572 116400 154592
rect 116400 154572 116452 154592
rect 116452 154572 116454 154592
rect 116398 154536 116454 154572
rect 115938 153448 115994 153504
rect 104806 152632 104862 152688
rect 116398 152224 116454 152280
rect 104162 151544 104218 151600
rect 116398 151136 116454 151192
rect 103794 150320 103850 150376
rect 103702 148960 103758 149016
rect 116398 149912 116454 149968
rect 104346 147600 104402 147656
rect 116398 148688 116454 148744
rect 104438 146240 104494 146296
rect 104162 142976 104218 143032
rect 103518 140528 103574 140584
rect 115938 147600 115994 147656
rect 116398 146376 116454 146432
rect 116030 145288 116086 145344
rect 104806 144744 104862 144800
rect 104622 144200 104678 144256
rect 116398 144064 116454 144120
rect 116398 142840 116454 142896
rect 104530 141752 104586 141808
rect 116398 141752 116454 141808
rect 103702 139304 103758 139360
rect 116398 140528 116454 140584
rect 116306 139476 116308 139496
rect 116308 139476 116360 139496
rect 116360 139476 116362 139496
rect 104346 137944 104402 138000
rect 104806 136584 104862 136640
rect 116306 139440 116362 139476
rect 115846 138216 115902 138272
rect 104806 135088 104862 135144
rect 104806 133728 104862 133784
rect 104714 133184 104770 133240
rect 104346 131960 104402 132016
rect 116398 137128 116454 137184
rect 115938 135904 115994 135960
rect 116398 134680 116454 134736
rect 103978 130600 104034 130656
rect 104806 129240 104862 129296
rect 116122 132368 116178 132424
rect 116398 131280 116454 131336
rect 116398 128832 116454 128888
rect 104806 128016 104862 128072
rect 116398 127744 116454 127800
rect 116398 126520 116454 126576
rect 116398 125432 116454 125488
rect 32218 125024 32274 125080
rect 185582 274896 185638 274952
rect 189078 320320 189134 320376
rect 193402 320320 193458 320376
rect 190182 320184 190238 320240
rect 191286 320184 191342 320240
rect 192390 320184 192446 320240
rect 194506 320184 194562 320240
rect 348790 700576 348846 700632
rect 283010 684392 283066 684448
rect 283102 678816 283158 678872
rect 283010 585928 283066 585984
rect 283194 568520 283250 568576
rect 283378 568520 283434 568576
rect 282918 511944 282974 512000
rect 283102 511980 283104 512000
rect 283104 511980 283156 512000
rect 283156 511980 283158 512000
rect 283102 511944 283158 511980
rect 282918 454008 282974 454064
rect 283194 454008 283250 454064
rect 282734 434696 282790 434752
rect 282918 434696 282974 434752
rect 283194 403552 283250 403608
rect 284390 608776 284446 608832
rect 284390 392672 284446 392728
rect 284298 369552 284354 369608
rect 282274 322088 282330 322144
rect 280158 295840 280214 295896
rect 281538 253952 281594 254008
rect 282182 253952 282238 254008
rect 235262 235184 235318 235240
rect 207754 224848 207810 224904
rect 206650 224576 206706 224632
rect 204534 224440 204590 224496
rect 205638 224304 205694 224360
rect 208858 224712 208914 224768
rect 209870 224168 209926 224224
rect 214378 212608 214434 212664
rect 214194 210296 214250 210352
rect 214194 208800 214250 208856
rect 214286 207168 214342 207224
rect 214378 205672 214434 205728
rect 214286 201728 214342 201784
rect 214378 200912 214434 200968
rect 214102 199280 214158 199336
rect 214102 197784 214158 197840
rect 214378 196152 214434 196208
rect 214286 190712 214342 190768
rect 214378 189216 214434 189272
rect 214010 188400 214066 188456
rect 213918 185272 213974 185328
rect 214470 184456 214526 184512
rect 214194 183640 214250 183696
rect 214194 181328 214250 181384
rect 214102 180512 214158 180568
rect 214010 179696 214066 179752
rect 213918 179016 213974 179072
rect 214102 178200 214158 178256
rect 214102 174256 214158 174312
rect 214286 172760 214342 172816
rect 214286 171944 214342 172000
rect 213918 168036 213920 168056
rect 213920 168036 213972 168056
rect 213972 168036 213974 168056
rect 213918 168000 213974 168036
rect 214286 167184 214342 167240
rect 214378 165688 214434 165744
rect 214102 164872 214158 164928
rect 214378 163240 214434 163296
rect 214286 161744 214342 161800
rect 214378 155488 214434 155544
rect 214010 152360 214066 152416
rect 214378 151544 214434 151600
rect 214378 149912 214434 149968
rect 214470 144472 214526 144528
rect 214378 139848 214434 139904
rect 214470 139032 214526 139088
rect 214286 137400 214342 137456
rect 214194 135904 214250 135960
rect 117134 133592 117190 133648
rect 214010 132776 214066 132832
rect 214378 131960 214434 132016
rect 214194 130328 214250 130384
rect 116674 130056 116730 130112
rect 214194 129648 214250 129704
rect 214010 128832 214066 128888
rect 116582 122984 116638 123040
rect 116398 121896 116454 121952
rect 116398 120672 116454 120728
rect 94778 97960 94834 98016
rect 94686 97144 94742 97200
rect 94870 96192 94926 96248
rect 94594 95376 94650 95432
rect 94502 94424 94558 94480
rect 94410 92656 94466 92712
rect 94410 87216 94466 87272
rect 94502 86400 94558 86456
rect 94042 83680 94098 83736
rect 94226 82864 94282 82920
rect 94410 80960 94466 81016
rect 94870 93472 94926 93528
rect 95146 98948 95148 98968
rect 95148 98948 95200 98968
rect 95200 98948 95202 98968
rect 95146 98912 95202 98948
rect 95146 91704 95202 91760
rect 94962 90888 95018 90944
rect 95054 89936 95110 89992
rect 95146 89120 95202 89176
rect 95146 88204 95148 88224
rect 95148 88204 95200 88224
rect 95200 88204 95202 88224
rect 95146 88168 95202 88204
rect 94870 85484 94872 85504
rect 94872 85484 94924 85504
rect 94924 85484 94926 85504
rect 94870 85448 94926 85484
rect 95146 84632 95202 84688
rect 95146 81912 95202 81968
rect 94686 80144 94742 80200
rect 94594 78376 94650 78432
rect 94410 77424 94466 77480
rect 94226 76472 94282 76528
rect 94594 75692 94596 75712
rect 94596 75692 94648 75712
rect 94648 75692 94650 75712
rect 94594 75656 94650 75692
rect 95146 79192 95202 79248
rect 94962 74704 95018 74760
rect 94042 72936 94098 72992
rect 94410 72120 94466 72176
rect 94226 71168 94282 71224
rect 94042 68448 94098 68504
rect 94134 65900 94136 65920
rect 94136 65900 94188 65920
rect 94188 65900 94190 65920
rect 94134 65864 94190 65900
rect 94410 64912 94466 64968
rect 94318 61376 94374 61432
rect 95146 73888 95202 73944
rect 94594 63960 94650 64016
rect 94502 60424 94558 60480
rect 94318 59472 94374 59528
rect 94410 57704 94466 57760
rect 94042 49680 94098 49736
rect 94870 70252 94872 70272
rect 94872 70252 94924 70272
rect 94924 70252 94926 70272
rect 94870 70216 94926 70252
rect 95054 69400 95110 69456
rect 95146 67632 95202 67688
rect 95146 66680 95202 66736
rect 94778 62192 94834 62248
rect 94686 58656 94742 58712
rect 94594 55120 94650 55176
rect 94594 54168 94650 54224
rect 95146 63180 95148 63200
rect 95148 63180 95200 63200
rect 95200 63180 95202 63200
rect 95146 63144 95202 63180
rect 94870 56888 94926 56944
rect 94778 53216 94834 53272
rect 94134 48864 94190 48920
rect 116398 119584 116454 119640
rect 214194 119448 214250 119504
rect 116398 118360 116454 118416
rect 214286 117816 214342 117872
rect 116306 117136 116362 117192
rect 116398 116048 116454 116104
rect 116398 114824 116454 114880
rect 214010 113872 214066 113928
rect 116398 113736 116454 113792
rect 116398 112512 116454 112568
rect 214378 112376 214434 112432
rect 116398 111424 116454 111480
rect 95146 55936 95202 55992
rect 95146 52420 95202 52456
rect 95146 52400 95148 52420
rect 95148 52400 95200 52420
rect 95200 52400 95202 52420
rect 94962 51448 95018 51504
rect 94870 47912 94926 47968
rect 94778 46960 94834 47016
rect 94410 44376 94466 44432
rect 95146 50632 95202 50688
rect 116398 110200 116454 110256
rect 214470 109248 214526 109304
rect 116306 108976 116362 109032
rect 116398 107888 116454 107944
rect 214194 106936 214250 106992
rect 116398 106664 116454 106720
rect 116398 105576 116454 105632
rect 214378 105304 214434 105360
rect 116398 104352 116454 104408
rect 214378 103808 214434 103864
rect 116306 103128 116362 103184
rect 116674 102040 116730 102096
rect 116398 100816 116454 100872
rect 116398 99728 116454 99784
rect 116398 98504 116454 98560
rect 116398 97280 116454 97336
rect 116306 96192 116362 96248
rect 116582 94968 116638 95024
rect 116398 93900 116454 93936
rect 116398 93880 116400 93900
rect 116400 93880 116452 93900
rect 116452 93880 116454 93900
rect 116398 92656 116454 92712
rect 116398 91568 116454 91624
rect 116398 90344 116454 90400
rect 115938 89120 115994 89176
rect 116398 88032 116454 88088
rect 116122 86808 116178 86864
rect 116398 85720 116454 85776
rect 116398 83272 116454 83328
rect 115938 82184 115994 82240
rect 116398 80960 116454 81016
rect 214470 99864 214526 99920
rect 214102 97416 214158 97472
rect 214838 170312 214894 170368
rect 215114 221312 215170 221368
rect 227626 221312 227682 221368
rect 226338 220804 226340 220824
rect 226340 220804 226392 220824
rect 226392 220804 226394 220824
rect 226338 220768 226394 220804
rect 215206 220496 215262 220552
rect 226338 220108 226394 220144
rect 226338 220088 226340 220108
rect 226340 220088 226392 220108
rect 226392 220088 226394 220108
rect 215114 219680 215170 219736
rect 226430 219544 226486 219600
rect 226338 219000 226394 219056
rect 215114 218864 215170 218920
rect 226430 218320 226486 218376
rect 215206 218184 215262 218240
rect 226338 217776 226394 217832
rect 215114 217368 215170 217424
rect 226430 217232 226486 217288
rect 215114 216588 215116 216608
rect 215116 216588 215168 216608
rect 215168 216588 215170 216608
rect 215114 216552 215170 216588
rect 226338 216552 226394 216608
rect 226430 216008 226486 216064
rect 215114 215736 215170 215792
rect 226338 215464 226394 215520
rect 215114 215056 215170 215112
rect 226430 214784 226486 214840
rect 215206 214240 215262 214296
rect 226338 214240 226394 214296
rect 226430 213560 226486 213616
rect 215114 213424 215170 213480
rect 226338 213016 226394 213072
rect 226522 212472 226578 212528
rect 215114 211928 215170 211984
rect 226154 211792 226210 211848
rect 215206 211112 215262 211168
rect 226062 210704 226118 210760
rect 225970 210024 226026 210080
rect 215114 209480 215170 209536
rect 226246 211248 226302 211304
rect 226154 209480 226210 209536
rect 226246 208936 226302 208992
rect 215114 207984 215170 208040
rect 225878 207712 225934 207768
rect 225786 206488 225842 206544
rect 215114 206352 215170 206408
rect 225602 205264 225658 205320
rect 215114 204856 215170 204912
rect 215114 204040 215170 204096
rect 215206 203224 215262 203280
rect 215114 202408 215170 202464
rect 225694 202952 225750 203008
rect 215114 200096 215170 200152
rect 215114 198636 215116 198656
rect 215116 198636 215168 198656
rect 215168 198636 215170 198656
rect 215114 198600 215170 198636
rect 215114 196968 215170 197024
rect 215114 195472 215170 195528
rect 215206 194656 215262 194712
rect 215114 193840 215170 193896
rect 215114 193024 215170 193080
rect 215206 192344 215262 192400
rect 215114 191528 215170 191584
rect 215114 189896 215170 189952
rect 215206 187584 215262 187640
rect 215206 186768 215262 186824
rect 215114 185952 215170 186008
rect 215114 182824 215170 182880
rect 215206 182144 215262 182200
rect 215022 177384 215078 177440
rect 215114 176604 215116 176624
rect 215116 176604 215168 176624
rect 215168 176604 215170 176624
rect 215114 176568 215170 176604
rect 215114 175888 215170 175944
rect 215114 175108 215116 175128
rect 215116 175108 215168 175128
rect 215168 175108 215170 175128
rect 215114 175072 215170 175108
rect 215206 173440 215262 173496
rect 215022 171128 215078 171184
rect 215114 169496 215170 169552
rect 215114 168816 215170 168872
rect 215206 166368 215262 166424
rect 214930 164092 214932 164112
rect 214932 164092 214984 164112
rect 214984 164092 214986 164112
rect 214930 164056 214986 164092
rect 225970 207168 226026 207224
rect 226154 207984 226210 208040
rect 226062 205944 226118 206000
rect 225970 203496 226026 203552
rect 225878 202408 225934 202464
rect 225786 199960 225842 200016
rect 226154 204720 226210 204776
rect 226246 204176 226302 204232
rect 226154 201728 226210 201784
rect 226062 200640 226118 200696
rect 226338 201184 226394 201240
rect 226430 199416 226486 199472
rect 226338 198872 226394 198928
rect 226430 198192 226486 198248
rect 226338 197648 226394 197704
rect 226614 196968 226670 197024
rect 226706 196424 226762 196480
rect 226338 195880 226394 195936
rect 226614 195200 226670 195256
rect 226430 194112 226486 194168
rect 226338 193432 226394 193488
rect 226430 192888 226486 192944
rect 226338 192344 226394 192400
rect 226338 191664 226394 191720
rect 226522 191120 226578 191176
rect 226982 194656 227038 194712
rect 226338 190476 226340 190496
rect 226340 190476 226392 190496
rect 226392 190476 226394 190496
rect 226338 190440 226394 190476
rect 226338 189896 226394 189952
rect 225786 189352 225842 189408
rect 225602 186904 225658 186960
rect 226338 188672 226394 188728
rect 226430 188128 226486 188184
rect 226338 187584 226394 187640
rect 226338 186380 226394 186416
rect 226338 186360 226340 186380
rect 226340 186360 226392 186380
rect 226392 186360 226394 186380
rect 226338 185816 226394 185872
rect 226982 185136 227038 185192
rect 226338 184592 226394 184648
rect 226522 184048 226578 184104
rect 226522 183368 226578 183424
rect 226430 182824 226486 182880
rect 226338 182180 226340 182200
rect 226340 182180 226392 182200
rect 226392 182180 226394 182200
rect 226338 182144 226394 182180
rect 226338 181056 226394 181112
rect 226338 180376 226394 180432
rect 226430 179832 226486 179888
rect 226430 178608 226486 178664
rect 226706 178064 226762 178120
rect 226338 177520 226394 177576
rect 227074 179288 227130 179344
rect 226982 175752 227038 175808
rect 227626 181600 227682 181656
rect 227350 176840 227406 176896
rect 227442 176296 227498 176352
rect 215114 162560 215170 162616
rect 288898 317056 288954 317112
rect 304262 328208 304318 328264
rect 303618 326304 303674 326360
rect 289726 325216 289782 325272
rect 303618 324400 303674 324456
rect 304354 322496 304410 322552
rect 304446 320592 304502 320648
rect 303618 318688 303674 318744
rect 304354 316920 304410 316976
rect 304262 315016 304318 315072
rect 303618 313112 303674 313168
rect 303618 311208 303674 311264
rect 303618 309304 303674 309360
rect 289634 308896 289690 308952
rect 303618 307400 303674 307456
rect 300858 305496 300914 305552
rect 292578 302776 292634 302832
rect 309046 473864 309102 473920
rect 309046 473320 309102 473376
rect 312542 613400 312598 613456
rect 312542 462712 312598 462768
rect 313278 439592 313334 439648
rect 478510 700440 478566 700496
rect 543462 700304 543518 700360
rect 580170 697992 580226 698048
rect 506018 663856 506074 663912
rect 553398 649576 553454 649632
rect 551742 638152 551798 638208
rect 456062 635160 456118 635216
rect 455418 591640 455474 591696
rect 385406 528808 385462 528864
rect 387338 528808 387394 528864
rect 398838 528944 398894 529000
rect 315302 528400 315358 528456
rect 315210 528284 315266 528320
rect 315210 528264 315212 528284
rect 315212 528264 315264 528284
rect 315264 528264 315266 528284
rect 320086 528400 320142 528456
rect 324226 528284 324282 528320
rect 324226 528264 324228 528284
rect 324228 528264 324280 528284
rect 324280 528264 324282 528284
rect 385682 528672 385738 528728
rect 386234 528672 386290 528728
rect 385958 528536 386014 528592
rect 385866 528400 385922 528456
rect 385774 528300 385776 528320
rect 385776 528300 385828 528320
rect 385828 528300 385830 528320
rect 385774 528264 385830 528300
rect 386510 528536 386566 528592
rect 386418 528400 386474 528456
rect 386326 528300 386328 528320
rect 386328 528300 386380 528320
rect 386380 528300 386382 528320
rect 386326 528264 386382 528300
rect 399206 528944 399262 529000
rect 435362 533024 435418 533080
rect 438950 532888 439006 532944
rect 454774 534384 454830 534440
rect 456798 616256 456854 616312
rect 458178 531664 458234 531720
rect 464526 534248 464582 534304
rect 461214 531528 461270 531584
rect 466642 532752 466698 532808
rect 481730 534112 481786 534168
rect 501786 533432 501842 533488
rect 499394 533296 499450 533352
rect 498566 532344 498622 532400
rect 496358 532072 496414 532128
rect 484950 531392 485006 531448
rect 493046 531256 493102 531312
rect 492034 531120 492090 531176
rect 490378 529896 490434 529952
rect 495346 530576 495402 530632
rect 493782 529896 493838 529952
rect 497462 531936 497518 531992
rect 500682 532208 500738 532264
rect 502890 532480 502946 532536
rect 520186 547032 520242 547088
rect 506110 533568 506166 533624
rect 507122 532616 507178 532672
rect 398838 528556 398894 528592
rect 398838 528536 398840 528556
rect 398840 528536 398892 528556
rect 398892 528536 398894 528556
rect 403714 528536 403770 528592
rect 422298 528420 422354 528456
rect 422298 528400 422300 528420
rect 422300 528400 422352 528420
rect 422352 528400 422354 528420
rect 431774 528400 431830 528456
rect 408222 528264 408278 528320
rect 422206 528300 422208 528320
rect 422208 528300 422260 528320
rect 422260 528300 422262 528320
rect 422206 528264 422262 528300
rect 509054 530712 509110 530768
rect 511446 531800 511502 531856
rect 515770 531664 515826 531720
rect 524234 530848 524290 530904
rect 551006 567704 551062 567760
rect 551006 559136 551062 559192
rect 550730 539552 550786 539608
rect 550914 539552 550970 539608
rect 551374 636928 551430 636984
rect 551374 633528 551430 633584
rect 551466 630808 551522 630864
rect 551374 628360 551430 628416
rect 551466 627952 551522 628008
rect 551558 623736 551614 623792
rect 551466 616256 551522 616312
rect 551650 618568 551706 618624
rect 552018 621288 552074 621344
rect 551834 616256 551890 616312
rect 551834 612856 551890 612912
rect 551742 603064 551798 603120
rect 551926 604288 551982 604344
rect 551834 588512 551890 588568
rect 552110 614352 552166 614408
rect 552202 611904 552258 611960
rect 552294 609456 552350 609512
rect 552386 607008 552442 607064
rect 552478 604560 552534 604616
rect 552570 602112 552626 602168
rect 552938 600888 552994 600944
rect 552754 599664 552810 599720
rect 552662 594768 552718 594824
rect 552846 597216 552902 597272
rect 553030 598440 553086 598496
rect 554410 648352 554466 648408
rect 553490 644680 553546 644736
rect 554042 643456 554098 643512
rect 553582 642232 553638 642288
rect 553674 639920 553730 639976
rect 553766 635024 553822 635080
rect 553858 632576 553914 632632
rect 553950 630128 554006 630184
rect 554870 627680 554926 627736
rect 554226 625232 554282 625288
rect 554134 610680 554190 610736
rect 554042 593952 554098 594008
rect 554042 593680 554098 593736
rect 554134 592456 554190 592512
rect 554778 617888 554834 617944
rect 554410 605784 554466 605840
rect 554318 588784 554374 588840
rect 554318 587560 554374 587616
rect 554318 585148 554320 585168
rect 554320 585148 554372 585168
rect 554372 585148 554374 585168
rect 554318 585112 554374 585148
rect 554318 583888 554374 583944
rect 554318 581440 554374 581496
rect 554318 580216 554374 580272
rect 554318 578992 554374 579048
rect 554318 577768 554374 577824
rect 554594 595992 554650 596048
rect 554502 591232 554558 591288
rect 554502 590008 554558 590064
rect 554502 586336 554558 586392
rect 554410 576544 554466 576600
rect 554318 575320 554374 575376
rect 554410 574116 554466 574152
rect 554410 574096 554412 574116
rect 554412 574096 554464 574116
rect 554464 574096 554466 574116
rect 554410 572872 554466 572928
rect 554226 571648 554282 571704
rect 554410 570560 554466 570616
rect 555146 622784 555202 622840
rect 555054 620336 555110 620392
rect 554962 613128 555018 613184
rect 555330 615576 555386 615632
rect 555238 608232 555294 608288
rect 555422 582664 555478 582720
rect 508502 528264 508558 528320
rect 315946 515752 316002 515808
rect 389822 473864 389878 473920
rect 408590 473728 408646 473784
rect 389822 473592 389878 473648
rect 408406 473592 408462 473648
rect 314658 439592 314714 439648
rect 338118 428712 338174 428768
rect 338394 428576 338450 428632
rect 338118 198600 338174 198656
rect 283378 173848 283434 173904
rect 232226 173168 232282 173224
rect 283378 173168 283434 173224
rect 215114 160928 215170 160984
rect 214930 160112 214986 160168
rect 214838 158616 214894 158672
rect 214746 157800 214802 157856
rect 215114 156984 215170 157040
rect 214746 156304 214802 156360
rect 215114 154672 215170 154728
rect 215206 153856 215262 153912
rect 215114 153212 215116 153232
rect 215116 153212 215168 153232
rect 215168 153212 215170 153232
rect 215114 153176 215170 153212
rect 215114 150728 215170 150784
rect 215114 149232 215170 149288
rect 215114 148416 215170 148472
rect 214838 147600 214894 147656
rect 215206 146784 215262 146840
rect 215022 146104 215078 146160
rect 215206 145288 215262 145344
rect 215206 143676 215262 143712
rect 215206 143656 215208 143676
rect 215208 143656 215260 143676
rect 215260 143656 215262 143676
rect 215114 142976 215170 143032
rect 215206 142196 215208 142216
rect 215208 142196 215260 142216
rect 215260 142196 215262 142216
rect 215206 142160 215262 142196
rect 215114 141344 215170 141400
rect 215114 140528 215170 140584
rect 215114 138216 215170 138272
rect 215114 136740 215170 136776
rect 215114 136720 215116 136740
rect 215116 136720 215168 136740
rect 215168 136720 215170 136740
rect 215206 135088 215262 135144
rect 215114 134272 215170 134328
rect 215114 133456 215170 133512
rect 215114 131180 215116 131200
rect 215116 131180 215168 131200
rect 215168 131180 215170 131200
rect 215114 131144 215170 131180
rect 215114 128016 215170 128072
rect 215114 127200 215170 127256
rect 215114 126520 215170 126576
rect 215114 125704 215170 125760
rect 215114 124908 215170 124944
rect 215114 124888 215116 124908
rect 215116 124888 215168 124908
rect 215168 124888 215170 124908
rect 215114 124108 215116 124128
rect 215116 124108 215168 124128
rect 215168 124108 215170 124128
rect 215114 124072 215170 124108
rect 215114 123428 215116 123448
rect 215116 123428 215168 123448
rect 215168 123428 215170 123448
rect 215114 123392 215170 123428
rect 215114 122576 215170 122632
rect 215114 121760 215170 121816
rect 215114 120944 215170 121000
rect 215114 120264 215170 120320
rect 215114 118632 215170 118688
rect 215114 117000 215170 117056
rect 215206 116320 215262 116376
rect 215114 115504 215170 115560
rect 215206 114688 215262 114744
rect 215114 113192 215170 113248
rect 215114 111560 215170 111616
rect 215206 110744 215262 110800
rect 215114 110064 215170 110120
rect 215114 108432 215170 108488
rect 215206 107616 215262 107672
rect 215114 106120 215170 106176
rect 215114 104488 215170 104544
rect 215206 102992 215262 103048
rect 215114 102176 215170 102232
rect 215114 101360 215170 101416
rect 215114 100580 215116 100600
rect 215116 100580 215168 100600
rect 215168 100580 215170 100600
rect 215114 100544 215170 100580
rect 214654 98232 214710 98288
rect 214562 96736 214618 96792
rect 214286 95920 214342 95976
rect 215114 99048 215170 99104
rect 232318 154536 232374 154592
rect 232502 154536 232558 154592
rect 227442 149368 227498 149424
rect 227442 148824 227498 148880
rect 227534 148144 227590 148200
rect 225602 147600 225658 147656
rect 226706 146920 226762 146976
rect 226522 146376 226578 146432
rect 227442 145832 227498 145888
rect 226706 145152 226762 145208
rect 226522 143928 226578 143984
rect 226890 142840 226946 142896
rect 226706 141616 226762 141672
rect 227442 144608 227498 144664
rect 227442 143420 227444 143440
rect 227444 143420 227496 143440
rect 227496 143420 227498 143440
rect 227442 143384 227498 143420
rect 227258 140936 227314 140992
rect 226522 136720 226578 136776
rect 227074 140392 227130 140448
rect 227626 142160 227682 142216
rect 227534 139712 227590 139768
rect 227442 139168 227498 139224
rect 227350 138624 227406 138680
rect 226706 137400 226762 137456
rect 226614 136176 226670 136232
rect 226430 135632 226486 135688
rect 227442 137964 227498 138000
rect 227442 137944 227444 137964
rect 227444 137944 227496 137964
rect 227496 137944 227498 137964
rect 226798 134952 226854 135008
rect 226522 133184 226578 133240
rect 227442 134408 227498 134464
rect 227258 133728 227314 133784
rect 226706 131960 226762 132016
rect 227534 132504 227590 132560
rect 227442 131416 227498 131472
rect 227350 130736 227406 130792
rect 227074 130192 227130 130248
rect 226522 129512 226578 129568
rect 227534 128968 227590 129024
rect 227442 128424 227498 128480
rect 226338 127744 226394 127800
rect 227442 127200 227498 127256
rect 227442 126520 227498 126576
rect 227442 125976 227498 126032
rect 227442 125296 227498 125352
rect 227258 124752 227314 124808
rect 227258 124208 227314 124264
rect 227258 123528 227314 123584
rect 227442 122984 227498 123040
rect 227442 122304 227498 122360
rect 227442 121760 227498 121816
rect 227442 121216 227498 121272
rect 227442 120536 227498 120592
rect 226430 119992 226486 120048
rect 226338 119312 226394 119368
rect 226246 118768 226302 118824
rect 226154 117544 226210 117600
rect 227442 118088 227498 118144
rect 227442 117000 227498 117056
rect 226246 116320 226302 116376
rect 226154 115096 226210 115152
rect 226062 114552 226118 114608
rect 225970 113328 226026 113384
rect 225786 112104 225842 112160
rect 225694 110336 225750 110392
rect 225602 109112 225658 109168
rect 227074 115776 227130 115832
rect 226246 114008 226302 114064
rect 226154 112784 226210 112840
rect 226062 110880 226118 110936
rect 225786 107888 225842 107944
rect 226246 111560 226302 111616
rect 226154 109792 226210 109848
rect 226062 107344 226118 107400
rect 225878 106800 225934 106856
rect 225970 106120 226026 106176
rect 226246 108568 226302 108624
rect 226154 105576 226210 105632
rect 227442 104916 227498 104952
rect 227442 104896 227444 104916
rect 227444 104896 227496 104916
rect 227496 104896 227498 104916
rect 226246 104352 226302 104408
rect 227442 103808 227498 103864
rect 343638 428440 343694 428496
rect 214746 95104 214802 95160
rect 215114 94288 215170 94344
rect 215114 93608 215170 93664
rect 215206 92792 215262 92848
rect 214562 91976 214618 92032
rect 214470 90480 214526 90536
rect 214102 88848 214158 88904
rect 117042 84496 117098 84552
rect 116398 79872 116454 79928
rect 214194 82592 214250 82648
rect 214746 91160 214802 91216
rect 214654 84904 214710 84960
rect 214010 80960 214066 81016
rect 116582 78648 116638 78704
rect 214562 78648 214618 78704
rect 116398 77424 116454 77480
rect 116398 76336 116454 76392
rect 116398 75112 116454 75168
rect 116398 74024 116454 74080
rect 214470 77152 214526 77208
rect 214286 74024 214342 74080
rect 116398 72800 116454 72856
rect 116306 71712 116362 71768
rect 214102 71576 214158 71632
rect 116398 70488 116454 70544
rect 116398 69264 116454 69320
rect 116398 68176 116454 68232
rect 116398 66952 116454 67008
rect 215114 89664 215170 89720
rect 215022 88032 215078 88088
rect 215114 87352 215170 87408
rect 215206 86536 215262 86592
rect 215114 85720 215170 85776
rect 214838 83408 214894 83464
rect 214746 77832 214802 77888
rect 214930 81776 214986 81832
rect 214654 72392 214710 72448
rect 213918 66136 213974 66192
rect 116398 65864 116454 65920
rect 214010 65320 214066 65376
rect 215206 84244 215262 84280
rect 215206 84224 215208 84244
rect 215208 84224 215260 84244
rect 215260 84224 215262 84244
rect 215022 80280 215078 80336
rect 215114 79464 215170 79520
rect 215206 76336 215262 76392
rect 215114 75520 215170 75576
rect 215206 74704 215262 74760
rect 215114 73208 215170 73264
rect 215114 70896 215170 70952
rect 214930 70080 214986 70136
rect 215114 69264 215170 69320
rect 215206 68448 215262 68504
rect 215114 67768 215170 67824
rect 215114 66952 215170 67008
rect 115938 64640 115994 64696
rect 214102 64504 214158 64560
rect 215114 63824 215170 63880
rect 116398 63416 116454 63472
rect 214378 63008 214434 63064
rect 116490 62328 116546 62384
rect 116398 61104 116454 61160
rect 116398 60016 116454 60072
rect 215114 62192 215170 62248
rect 214746 61376 214802 61432
rect 215114 60732 215116 60752
rect 215116 60732 215168 60752
rect 215168 60732 215170 60752
rect 215114 60696 215170 60732
rect 214378 59880 214434 59936
rect 214286 59064 214342 59120
rect 116398 58792 116454 58848
rect 214378 58248 214434 58304
rect 116306 57568 116362 57624
rect 213918 57568 213974 57624
rect 214010 56752 214066 56808
rect 116306 56480 116362 56536
rect 215114 55936 215170 55992
rect 116398 55276 116454 55312
rect 116398 55256 116400 55276
rect 116400 55256 116452 55276
rect 116452 55256 116454 55276
rect 214746 55120 214802 55176
rect 116398 54168 116454 54224
rect 215114 54440 215170 54496
rect 214746 53624 214802 53680
rect 116398 52944 116454 53000
rect 215114 52808 215170 52864
rect 214562 51992 214618 52048
rect 115938 51856 115994 51912
rect 215114 51312 215170 51368
rect 116398 50632 116454 50688
rect 214378 50496 214434 50552
rect 215114 49716 215116 49736
rect 215116 49716 215168 49736
rect 215168 49716 215170 49736
rect 95054 46144 95110 46200
rect 215114 49680 215170 49716
rect 116398 49408 116454 49464
rect 116122 48356 116124 48376
rect 116124 48356 116176 48376
rect 116176 48356 116178 48376
rect 116122 48320 116178 48356
rect 215114 48864 215170 48920
rect 214746 48048 214802 48104
rect 214010 47368 214066 47424
rect 116398 47096 116454 47152
rect 215206 46552 215262 46608
rect 116398 46008 116454 46064
rect 215114 45736 215170 45792
rect 95146 45192 95202 45248
rect 214470 44920 214526 44976
rect 116398 44784 116454 44840
rect 215114 44260 215170 44296
rect 215114 44240 215116 44260
rect 215116 44240 215168 44260
rect 215168 44240 215170 44260
rect 94962 43424 95018 43480
rect 94134 42472 94190 42528
rect 93950 41656 94006 41712
rect 115938 43560 115994 43616
rect 214378 43424 214434 43480
rect 214102 42608 214158 42664
rect 116398 42472 116454 42528
rect 215114 41792 215170 41848
rect 95054 40704 95110 40760
rect 94594 39888 94650 39944
rect 94502 38120 94558 38176
rect 116306 41248 116362 41304
rect 214654 41112 214710 41168
rect 116398 40160 116454 40216
rect 215114 40296 215170 40352
rect 214470 39480 214526 39536
rect 95146 38936 95202 38992
rect 116398 38936 116454 38992
rect 215114 38684 215170 38720
rect 215114 38664 215116 38684
rect 215116 38664 215168 38684
rect 215168 38664 215170 38684
rect 215114 37984 215170 38040
rect 116398 37712 116454 37768
rect 95054 37168 95110 37224
rect 215114 37168 215170 37224
rect 116398 36624 116454 36680
rect 94594 36216 94650 36272
rect 214562 36352 214618 36408
rect 93858 35400 93914 35456
rect 214654 35536 214710 35592
rect 116398 35400 116454 35456
rect 215114 34856 215170 34912
rect 93950 34448 94006 34504
rect 116306 34312 116362 34368
rect 95146 33632 95202 33688
rect 214562 34040 214618 34096
rect 215114 33244 215170 33280
rect 215114 33224 215116 33244
rect 215116 33224 215168 33244
rect 215168 33224 215170 33244
rect 116398 33088 116454 33144
rect 95146 32680 95202 32736
rect 225602 75792 225658 75848
rect 227074 74568 227130 74624
rect 343638 126656 343694 126712
rect 227442 81096 227498 81152
rect 227534 80416 227590 80472
rect 227350 79736 227406 79792
rect 227442 79056 227498 79112
rect 227442 78548 227444 78568
rect 227444 78548 227496 78568
rect 227496 78548 227498 78568
rect 227442 78512 227498 78548
rect 227534 77832 227590 77888
rect 227442 77172 227498 77208
rect 227442 77152 227444 77172
rect 227444 77152 227496 77172
rect 227496 77152 227498 77172
rect 227534 76472 227590 76528
rect 227442 75248 227498 75304
rect 227442 73888 227498 73944
rect 227166 73208 227222 73264
rect 227442 72664 227498 72720
rect 227534 71984 227590 72040
rect 227442 71304 227498 71360
rect 227534 70624 227590 70680
rect 227442 69944 227498 70000
rect 226522 69400 226578 69456
rect 227442 68720 227498 68776
rect 227534 68040 227590 68096
rect 227442 67360 227498 67416
rect 227534 66816 227590 66872
rect 227442 66172 227444 66192
rect 227444 66172 227496 66192
rect 227496 66172 227498 66192
rect 227442 66136 227498 66172
rect 227534 65456 227590 65512
rect 227258 64776 227314 64832
rect 227442 64096 227498 64152
rect 227534 63552 227590 63608
rect 227442 62872 227498 62928
rect 227074 62192 227130 62248
rect 227442 61512 227498 61568
rect 226706 60968 226762 61024
rect 227442 60288 227498 60344
rect 227534 59608 227590 59664
rect 227442 58928 227498 58984
rect 227534 58248 227590 58304
rect 227258 57704 227314 57760
rect 227442 57024 227498 57080
rect 227258 56344 227314 56400
rect 227442 55664 227498 55720
rect 227442 55156 227444 55176
rect 227444 55156 227496 55176
rect 227496 55156 227498 55176
rect 227442 55120 227498 55156
rect 226522 54440 226578 54496
rect 226522 50496 226578 50552
rect 226338 47912 226394 47968
rect 226706 49272 226762 49328
rect 227258 53760 227314 53816
rect 227442 53080 227498 53136
rect 227258 52400 227314 52456
rect 227442 51856 227498 51912
rect 227534 51176 227590 51232
rect 226982 49816 227038 49872
rect 226798 48592 226854 48648
rect 226614 47232 226670 47288
rect 227350 46552 227406 46608
rect 227074 46008 227130 46064
rect 227534 45328 227590 45384
rect 227442 44648 227498 44704
rect 227074 43424 227130 43480
rect 226706 42744 226762 42800
rect 226430 40704 226486 40760
rect 226338 40160 226394 40216
rect 227626 43968 227682 44024
rect 227442 42064 227498 42120
rect 227350 41384 227406 41440
rect 226614 39480 226670 39536
rect 227074 38800 227130 38856
rect 226890 38120 226946 38176
rect 227442 37576 227498 37632
rect 227534 36896 227590 36952
rect 227442 36216 227498 36272
rect 227442 35536 227498 35592
rect 227534 34856 227590 34912
rect 227442 34312 227498 34368
rect 227350 33632 227406 33688
rect 227442 32952 227498 33008
rect 116398 32000 116454 32056
rect 95146 31864 95202 31920
rect 215114 32428 215170 32464
rect 215114 32408 215116 32428
rect 215116 32408 215168 32428
rect 215168 32408 215170 32428
rect 227534 32272 227590 32328
rect 213918 31728 213974 31784
rect 227442 31728 227498 31784
rect 32310 30268 32312 30288
rect 32312 30268 32364 30288
rect 32364 30268 32366 30288
rect 32310 30232 32366 30268
rect 126886 14456 126942 14512
rect 127806 7520 127862 7576
rect 131026 15272 131082 15328
rect 136546 12960 136602 13016
rect 138478 8880 138534 8936
rect 142066 11600 142122 11656
rect 145654 7656 145710 7712
rect 151726 14592 151782 14648
rect 158626 14728 158682 14784
rect 165526 11736 165582 11792
rect 172426 13096 172482 13152
rect 175370 6160 175426 6216
rect 169390 1944 169446 2000
rect 177762 9016 177818 9072
rect 176566 2080 176622 2136
rect 191746 6296 191802 6352
rect 193310 7792 193366 7848
rect 201406 13232 201462 13288
rect 198186 5072 198242 5128
rect 491850 500792 491906 500848
rect 493138 500792 493194 500848
rect 418158 473728 418214 473784
rect 437386 473728 437442 473784
rect 437570 473728 437626 473784
rect 418066 473592 418122 473648
rect 427726 473320 427782 473376
rect 427910 473320 427966 473376
rect 493966 475496 494022 475552
rect 496726 487736 496782 487792
rect 495346 475360 495402 475416
rect 499394 476720 499450 476776
rect 500866 475632 500922 475688
rect 503534 476992 503590 477048
rect 502246 476856 502302 476912
rect 503626 475768 503682 475824
rect 481638 473748 481694 473784
rect 481638 473728 481640 473748
rect 481640 473728 481692 473748
rect 481692 473728 481694 473748
rect 490654 473592 490710 473648
rect 508226 500792 508282 500848
rect 506386 477128 506442 477184
rect 508502 476040 508558 476096
rect 509146 476040 509202 476096
rect 507766 475904 507822 475960
rect 505006 474000 505062 474056
rect 505006 473612 505062 473648
rect 505006 473592 505008 473612
rect 505008 473592 505060 473612
rect 505060 473592 505062 473612
rect 491850 473476 491906 473512
rect 491850 473456 491852 473476
rect 491852 473456 491904 473476
rect 491904 473456 491906 473476
rect 493138 473476 493194 473512
rect 513286 474136 513342 474192
rect 517978 500792 518034 500848
rect 520186 474272 520242 474328
rect 542634 500792 542690 500848
rect 542910 476176 542966 476232
rect 520738 473864 520794 473920
rect 512642 473728 512698 473784
rect 550086 500792 550142 500848
rect 493138 473456 493140 473476
rect 493140 473456 493192 473476
rect 493192 473456 493194 473476
rect 443642 450608 443698 450664
rect 552478 475496 552534 475552
rect 552294 474544 552350 474600
rect 552110 472504 552166 472560
rect 552202 472368 552258 472424
rect 552018 451696 552074 451752
rect 552018 451152 552074 451208
rect 552018 447616 552074 447672
rect 552294 470736 552350 470792
rect 552478 471824 552534 471880
rect 552386 470056 552442 470112
rect 552570 469512 552626 469568
rect 553030 472640 553086 472696
rect 552386 460708 552388 460728
rect 552388 460708 552440 460728
rect 552440 460708 552442 460728
rect 552386 460672 552442 460708
rect 552386 454688 552442 454744
rect 552662 459992 552718 460048
rect 553030 462712 553086 462768
rect 552938 459176 552994 459232
rect 552846 457952 552902 458008
rect 552570 453464 552626 453520
rect 552846 456728 552902 456784
rect 552754 454144 552810 454200
rect 552662 452920 552718 452976
rect 552386 449928 552442 449984
rect 552202 446936 552258 446992
rect 552570 445168 552626 445224
rect 553398 443672 553454 443728
rect 552110 441632 552166 441688
rect 554042 448976 554098 449032
rect 553950 447888 554006 447944
rect 553858 445440 553914 445496
rect 553766 444352 553822 444408
rect 553674 443128 553730 443184
rect 553582 441904 553638 441960
rect 554134 440136 554190 440192
rect 553490 439592 553546 439648
rect 554870 455504 554926 455560
rect 555054 456184 555110 456240
rect 554962 454960 555018 455016
rect 554318 448432 554374 448488
rect 554226 438912 554282 438968
rect 555422 450200 555478 450256
rect 555330 446120 555386 446176
rect 555238 442448 555294 442504
rect 555146 438368 555202 438424
rect 555882 462032 555938 462088
rect 555790 460944 555846 461000
rect 555698 458496 555754 458552
rect 555606 451968 555662 452024
rect 555514 437824 555570 437880
rect 556066 437144 556122 437200
rect 554778 436600 554834 436656
rect 554778 436056 554834 436112
rect 554778 435376 554834 435432
rect 554870 434832 554926 434888
rect 554778 434152 554834 434208
rect 554870 433608 554926 433664
rect 554778 433064 554834 433120
rect 554870 432384 554926 432440
rect 554778 431860 554834 431896
rect 554778 431840 554780 431860
rect 554780 431840 554832 431860
rect 554832 431840 554834 431860
rect 554870 431296 554926 431352
rect 554962 430616 555018 430672
rect 554778 430072 554834 430128
rect 554870 429528 554926 429584
rect 554870 428884 554872 428904
rect 554872 428884 554924 428904
rect 554924 428884 554926 428904
rect 554870 428848 554926 428884
rect 554778 428304 554834 428360
rect 554778 427780 554834 427816
rect 554778 427760 554780 427780
rect 554780 427760 554832 427780
rect 554832 427760 554834 427780
rect 573454 502696 573510 502752
rect 411994 49816 412050 49872
rect 580354 686296 580410 686352
rect 579618 651072 579674 651128
rect 580262 639376 580318 639432
rect 578882 604152 578938 604208
rect 579802 557232 579858 557288
rect 580170 463392 580226 463448
rect 580170 416472 580226 416528
rect 580170 369552 580226 369608
rect 580170 322632 580226 322688
rect 580170 275712 580226 275768
rect 579986 228792 580042 228848
rect 579986 181872 580042 181928
rect 580170 134816 580226 134872
rect 580170 87896 580226 87952
rect 580538 592456 580594 592512
rect 580446 580760 580502 580816
rect 580906 545536 580962 545592
rect 580538 510312 580594 510368
rect 580906 498616 580962 498672
rect 580906 451696 580962 451752
rect 580906 404776 580962 404832
rect 580906 357856 580962 357912
rect 580354 310800 580410 310856
rect 580906 310800 580962 310856
rect 580354 263880 580410 263936
rect 580906 263880 580962 263936
rect 580906 216960 580962 217016
rect 580906 170040 580962 170096
rect 580906 123120 580962 123176
rect 580906 76200 580962 76256
rect 580170 40976 580226 41032
rect 563702 38664 563758 38720
rect 411902 27512 411958 27568
rect 215206 13368 215262 13424
rect 211066 7928 211122 7984
rect 212262 4800 212318 4856
rect 246302 15408 246358 15464
rect 224866 10240 224922 10296
rect 222934 4936 222990 4992
rect 232502 8064 232558 8120
rect 244186 11872 244242 11928
rect 238666 10376 238722 10432
rect 242806 10512 242862 10568
rect 250442 15544 250498 15600
rect 256698 2624 256754 2680
rect 273166 9152 273222 9208
rect 272890 6432 272946 6488
rect 275282 3440 275338 3496
rect 282458 3304 282514 3360
rect 289818 5208 289874 5264
rect 289542 3576 289598 3632
rect 296718 3712 296774 3768
rect 406474 16904 406530 16960
rect 414662 16904 414718 16960
rect 424598 16904 424654 16960
rect 435362 16904 435418 16960
rect 439410 16904 439466 16960
rect 452566 16904 452622 16960
rect 307206 14864 307262 14920
rect 307758 9288 307814 9344
rect 340142 12008 340198 12064
rect 356058 2916 356114 2952
rect 356058 2896 356060 2916
rect 356060 2896 356112 2916
rect 356112 2896 356114 2916
rect 369122 2916 369178 2952
rect 369122 2896 369124 2916
rect 369124 2896 369176 2916
rect 369176 2896 369178 2916
rect 374090 2916 374146 2952
rect 374090 2896 374092 2916
rect 374092 2896 374144 2916
rect 374144 2896 374146 2916
rect 378966 2896 379022 2952
rect 393226 10648 393282 10704
rect 414202 14456 414258 14512
rect 412638 3032 412694 3088
rect 414202 3032 414258 3088
rect 415306 15272 415362 15328
rect 414570 7520 414626 7576
rect 417238 12960 417294 13016
rect 417974 8880 418030 8936
rect 419170 11600 419226 11656
rect 418250 6296 418306 6352
rect 417514 5072 417570 5128
rect 419906 10648 419962 10704
rect 420274 7656 420330 7712
rect 421838 14592 421894 14648
rect 422298 12572 422354 12608
rect 422298 12552 422300 12572
rect 422300 12552 422352 12572
rect 422352 12552 422354 12572
rect 422758 12552 422814 12608
rect 423126 11736 423182 11792
rect 424138 14728 424194 14784
rect 425058 13096 425114 13152
rect 426806 15408 426862 15464
rect 426714 7792 426770 7848
rect 427082 3440 427138 3496
rect 427910 1944 427966 2000
rect 429106 15544 429162 15600
rect 429198 9152 429254 9208
rect 430670 9016 430726 9072
rect 429290 6160 429346 6216
rect 429474 2080 429530 2136
rect 433338 3304 433394 3360
rect 432050 2624 432106 2680
rect 434718 3440 434774 3496
rect 436742 3576 436798 3632
rect 437938 13232 437994 13288
rect 440238 12008 440294 12064
rect 439502 3460 439558 3496
rect 439502 3440 439504 3460
rect 439504 3440 439556 3460
rect 439556 3440 439558 3460
rect 440514 5208 440570 5264
rect 440974 9288 441030 9344
rect 442538 13368 442594 13424
rect 441342 7928 441398 7984
rect 441986 4800 442042 4856
rect 445574 10240 445630 10296
rect 445022 4936 445078 4992
rect 442998 3712 443054 3768
rect 444286 3460 444342 3496
rect 444286 3440 444288 3460
rect 444288 3440 444340 3460
rect 444340 3440 444342 3460
rect 446402 3612 446404 3632
rect 446404 3612 446456 3632
rect 446456 3612 446458 3632
rect 446402 3576 446458 3612
rect 448242 8064 448298 8120
rect 451738 11872 451794 11928
rect 451370 10512 451426 10568
rect 450174 10376 450230 10432
rect 455970 3612 455972 3632
rect 455972 3612 456024 3632
rect 456024 3612 456026 3632
rect 455970 3576 456026 3612
rect 461306 6432 461362 6488
rect 466182 12588 466184 12608
rect 466184 12588 466236 12608
rect 466236 12588 466238 12608
rect 466182 12552 466238 12588
rect 469034 3576 469090 3632
rect 471886 12588 471888 12608
rect 471888 12588 471940 12608
rect 471940 12588 471942 12608
rect 471886 12552 471942 12588
rect 472438 14864 472494 14920
rect 483018 3732 483074 3768
rect 483018 3712 483020 3732
rect 483020 3712 483072 3732
rect 483072 3712 483074 3732
rect 483018 3304 483074 3360
rect 483202 3476 483204 3496
rect 483204 3476 483256 3496
rect 483256 3476 483258 3496
rect 483202 3440 483258 3476
rect 484398 3732 484454 3768
rect 484398 3712 484400 3732
rect 484400 3712 484452 3732
rect 484452 3712 484454 3732
rect 483386 3476 483388 3496
rect 483388 3476 483440 3496
rect 483440 3476 483442 3496
rect 483386 3440 483442 3476
rect 483570 3304 483626 3360
rect 580906 29280 580962 29336
<< metal3 >>
rect 317086 700572 317092 700636
rect 317156 700634 317162 700636
rect 348785 700634 348851 700637
rect 317156 700632 348851 700634
rect 317156 700576 348790 700632
rect 348846 700576 348851 700632
rect 317156 700574 348851 700576
rect 317156 700572 317162 700574
rect 348785 700571 348851 700574
rect 317270 700436 317276 700500
rect 317340 700498 317346 700500
rect 478505 700498 478571 700501
rect 317340 700496 478571 700498
rect 317340 700440 478510 700496
rect 478566 700440 478571 700496
rect 317340 700438 478571 700440
rect 317340 700436 317346 700438
rect 478505 700435 478571 700438
rect 18638 700300 18644 700364
rect 18708 700362 18714 700364
rect 72969 700362 73035 700365
rect 18708 700360 73035 700362
rect 18708 700304 72974 700360
rect 73030 700304 73035 700360
rect 18708 700302 73035 700304
rect 18708 700300 18714 700302
rect 72969 700299 73035 700302
rect 316902 700300 316908 700364
rect 316972 700362 316978 700364
rect 543457 700362 543523 700365
rect 316972 700360 543523 700362
rect 316972 700304 543462 700360
rect 543518 700304 543523 700360
rect 316972 700302 543523 700304
rect 316972 700300 316978 700302
rect 543457 700299 543523 700302
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 580349 686354 580415 686357
rect 583520 686354 584960 686444
rect 580349 686352 584960 686354
rect 580349 686296 580354 686352
rect 580410 686296 584960 686352
rect 580349 686294 584960 686296
rect 580349 686291 580415 686294
rect 583520 686204 584960 686294
rect 283005 684452 283071 684453
rect 283005 684448 283052 684452
rect 283116 684450 283122 684452
rect 283005 684392 283010 684448
rect 283005 684388 283052 684392
rect 283116 684390 283162 684450
rect 283116 684388 283122 684390
rect 283005 684387 283071 684388
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 219065 679148 219131 679149
rect 219014 679146 219020 679148
rect 218974 679086 219020 679146
rect 219084 679144 219131 679148
rect 219126 679088 219131 679144
rect 219014 679084 219020 679086
rect 219084 679084 219131 679088
rect 219065 679083 219131 679084
rect 283097 678876 283163 678877
rect 283046 678874 283052 678876
rect 283006 678814 283052 678874
rect 283116 678872 283163 678876
rect 283158 678816 283163 678872
rect 283046 678812 283052 678814
rect 283116 678812 283163 678816
rect 283097 678811 283163 678812
rect 218973 676292 219039 676293
rect 218973 676288 219020 676292
rect 219084 676290 219090 676292
rect 218973 676232 218978 676288
rect 218973 676228 219020 676232
rect 219084 676230 219130 676290
rect 219084 676228 219090 676230
rect 218973 676227 219039 676228
rect 583520 674508 584960 674748
rect -960 667994 480 668084
rect 280654 667994 280660 667996
rect -960 667934 280660 667994
rect -960 667844 480 667934
rect 280654 667932 280660 667934
rect 280724 667932 280730 667996
rect 492438 663852 492444 663916
rect 492508 663914 492514 663916
rect 506013 663914 506079 663917
rect 492508 663912 506079 663914
rect 492508 663856 506018 663912
rect 506074 663856 506079 663912
rect 492508 663854 506079 663856
rect 492508 663852 492514 663854
rect 506013 663851 506079 663854
rect 583520 662676 584960 662916
rect 493910 662084 493916 662148
rect 493980 662146 493986 662148
rect 493980 662086 551386 662146
rect 493980 662084 493986 662086
rect 551326 661844 551386 662086
rect 551326 660108 551386 660620
rect 551318 660044 551324 660108
rect 551388 660044 551394 660108
rect 553342 659426 553348 659428
rect 551908 659366 553348 659426
rect 553342 659364 553348 659366
rect 553412 659364 553418 659428
rect 551326 657932 551386 658172
rect 551318 657868 551324 657932
rect 551388 657868 551394 657932
rect 553526 656978 553532 656980
rect 551908 656918 553532 656978
rect 553526 656916 553532 656918
rect 553596 656916 553602 656980
rect 551878 655618 551938 655724
rect 552054 655618 552060 655620
rect 551878 655558 552060 655618
rect 552054 655556 552060 655558
rect 552124 655556 552130 655620
rect 553894 654530 553900 654532
rect 551908 654470 553900 654530
rect 553894 654468 553900 654470
rect 553964 654468 553970 654532
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 553710 653306 553716 653308
rect 551908 653246 553716 653306
rect 553710 653244 553716 653246
rect 553780 653244 553786 653308
rect 554078 652082 554084 652084
rect 551908 652022 554084 652082
rect 554078 652020 554084 652022
rect 554148 652020 554154 652084
rect 579613 651130 579679 651133
rect 583520 651130 584960 651220
rect 579613 651128 584960 651130
rect 579613 651072 579618 651128
rect 579674 651072 584960 651128
rect 579613 651070 584960 651072
rect 579613 651067 579679 651070
rect 583520 650980 584960 651070
rect 551326 650588 551386 650828
rect 551318 650524 551324 650588
rect 551388 650524 551394 650588
rect 553393 649634 553459 649637
rect 551908 649632 553459 649634
rect 551908 649576 553398 649632
rect 553454 649576 553459 649632
rect 551908 649574 553459 649576
rect 553393 649571 553459 649574
rect 554405 648410 554471 648413
rect 551908 648408 554471 648410
rect 551908 648352 554410 648408
rect 554466 648352 554471 648408
rect 551908 648350 554471 648352
rect 554405 648347 554471 648350
rect 551510 646644 551570 647156
rect 551502 646580 551508 646644
rect 551572 646580 551578 646644
rect 551326 645828 551386 645932
rect 551318 645764 551324 645828
rect 551388 645764 551394 645828
rect 553485 644738 553551 644741
rect 551908 644736 553551 644738
rect 551908 644680 553490 644736
rect 553546 644680 553551 644736
rect 551908 644678 553551 644680
rect 553485 644675 553551 644678
rect 554037 643514 554103 643517
rect 551908 643512 554103 643514
rect 551908 643456 554042 643512
rect 554098 643456 554103 643512
rect 551908 643454 554103 643456
rect 554037 643451 554103 643454
rect 553577 642290 553643 642293
rect 551908 642288 553643 642290
rect 551908 642232 553582 642288
rect 553638 642232 553643 642288
rect 551908 642230 553643 642232
rect 553577 642227 553643 642230
rect 552238 641066 552244 641068
rect 551908 641006 552244 641066
rect 552238 641004 552244 641006
rect 552308 641004 552314 641068
rect 553669 639978 553735 639981
rect 551908 639976 553735 639978
rect 551908 639920 553674 639976
rect 553730 639920 553735 639976
rect 551908 639918 553735 639920
rect 553669 639915 553735 639918
rect 580257 639434 580323 639437
rect 583520 639434 584960 639524
rect 580257 639432 584960 639434
rect 580257 639376 580262 639432
rect 580318 639376 584960 639432
rect 580257 639374 584960 639376
rect 580257 639371 580323 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 551694 638213 551754 638724
rect 551694 638208 551803 638213
rect 551694 638152 551742 638208
rect 551798 638152 551803 638208
rect 551694 638150 551803 638152
rect 551737 638147 551803 638150
rect 551326 636989 551386 637500
rect 551326 636984 551435 636989
rect 551326 636928 551374 636984
rect 551430 636928 551435 636984
rect 551326 636926 551435 636928
rect 551369 636923 551435 636926
rect 552422 636306 552428 636308
rect 551908 636246 552428 636306
rect 552422 636244 552428 636246
rect 552492 636244 552498 636308
rect 456057 635218 456123 635221
rect 454020 635216 456123 635218
rect 454020 635160 456062 635216
rect 456118 635160 456123 635216
rect 454020 635158 456123 635160
rect 456057 635155 456123 635158
rect 553761 635082 553827 635085
rect 551908 635080 553827 635082
rect 551908 635024 553766 635080
rect 553822 635024 553827 635080
rect 551908 635022 553827 635024
rect 553761 635019 553827 635022
rect 551326 633589 551386 633828
rect 551326 633584 551435 633589
rect 551326 633528 551374 633584
rect 551430 633528 551435 633584
rect 551326 633526 551435 633528
rect 551369 633523 551435 633526
rect 553853 632634 553919 632637
rect 551908 632632 553919 632634
rect 551908 632576 553858 632632
rect 553914 632576 553919 632632
rect 551908 632574 553919 632576
rect 553853 632571 553919 632574
rect 552790 631410 552796 631412
rect 551908 631350 552796 631410
rect 552790 631348 552796 631350
rect 552860 631348 552866 631412
rect 551461 630866 551527 630869
rect 551686 630866 551692 630868
rect 551461 630864 551692 630866
rect 551461 630808 551466 630864
rect 551522 630808 551692 630864
rect 551461 630806 551692 630808
rect 551461 630803 551527 630806
rect 551686 630804 551692 630806
rect 551756 630804 551762 630868
rect 551502 630668 551508 630732
rect 551572 630668 551578 630732
rect 551510 630594 551570 630668
rect 551686 630594 551692 630596
rect 551510 630534 551692 630594
rect 551686 630532 551692 630534
rect 551756 630532 551762 630596
rect 553945 630186 554011 630189
rect 551908 630184 554011 630186
rect 551908 630128 553950 630184
rect 554006 630128 554011 630184
rect 551908 630126 554011 630128
rect 553945 630123 554011 630126
rect 551326 628421 551386 628932
rect 551326 628416 551435 628421
rect 551326 628360 551374 628416
rect 551430 628360 551435 628416
rect 551326 628358 551435 628360
rect 551369 628355 551435 628358
rect 551318 627948 551324 628012
rect 551388 628010 551394 628012
rect 551461 628010 551527 628013
rect 551388 628008 551527 628010
rect 551388 627952 551466 628008
rect 551522 627952 551527 628008
rect 551388 627950 551527 627952
rect 551388 627948 551394 627950
rect 551461 627947 551527 627950
rect 554865 627738 554931 627741
rect 551908 627736 554931 627738
rect 551908 627680 554870 627736
rect 554926 627680 554931 627736
rect 551908 627678 554931 627680
rect 554865 627675 554931 627678
rect 583520 627588 584960 627828
rect 552606 626514 552612 626516
rect 551908 626454 552612 626514
rect 552606 626452 552612 626454
rect 552676 626452 552682 626516
rect 554221 625290 554287 625293
rect 551908 625288 554287 625290
rect 551908 625232 554226 625288
rect 554282 625232 554287 625288
rect 551908 625230 554287 625232
rect 554221 625227 554287 625230
rect -960 624882 480 624972
rect 3417 624882 3483 624885
rect -960 624880 3483 624882
rect -960 624824 3422 624880
rect 3478 624824 3483 624880
rect -960 624822 3483 624824
rect -960 624732 480 624822
rect 3417 624819 3483 624822
rect 551510 623797 551570 624036
rect 551510 623792 551619 623797
rect 551510 623736 551558 623792
rect 551614 623736 551619 623792
rect 551510 623734 551619 623736
rect 551553 623731 551619 623734
rect 555141 622842 555207 622845
rect 551908 622840 555207 622842
rect 551908 622784 555146 622840
rect 555202 622784 555207 622840
rect 551908 622782 555207 622784
rect 555141 622779 555207 622782
rect 551878 621346 551938 621588
rect 552013 621346 552079 621349
rect 551878 621344 552079 621346
rect 551878 621288 552018 621344
rect 552074 621288 552079 621344
rect 551878 621286 552079 621288
rect 552013 621283 552079 621286
rect 555049 620394 555115 620397
rect 551908 620392 555115 620394
rect 551908 620336 555054 620392
rect 555110 620336 555115 620392
rect 551908 620334 555115 620336
rect 555049 620331 555115 620334
rect 91093 619578 91159 619581
rect 95877 619578 95943 619581
rect 91093 619576 95943 619578
rect 91093 619520 91098 619576
rect 91154 619520 95882 619576
rect 95938 619520 95943 619576
rect 91093 619518 95943 619520
rect 91093 619515 91159 619518
rect 95877 619515 95943 619518
rect 279141 619578 279207 619581
rect 280102 619578 280108 619580
rect 279141 619576 280108 619578
rect 279141 619520 279146 619576
rect 279202 619520 280108 619576
rect 279141 619518 280108 619520
rect 279141 619515 279207 619518
rect 280102 619516 280108 619518
rect 280172 619516 280178 619580
rect 551694 618629 551754 619140
rect 551645 618624 551754 618629
rect 551645 618568 551650 618624
rect 551706 618568 551754 618624
rect 551645 618566 551754 618568
rect 551645 618563 551711 618566
rect 554773 617946 554839 617949
rect 551908 617944 554839 617946
rect 551908 617888 554778 617944
rect 554834 617888 554839 617944
rect 551908 617886 554839 617888
rect 554773 617883 554839 617886
rect 30189 617810 30255 617813
rect 31150 617810 31156 617812
rect 30189 617808 31156 617810
rect 30189 617752 30194 617808
rect 30250 617752 31156 617808
rect 30189 617750 31156 617752
rect 30189 617747 30255 617750
rect 31150 617748 31156 617750
rect 31220 617748 31226 617812
rect 30281 617674 30347 617677
rect 31334 617674 31340 617676
rect 30281 617672 31340 617674
rect 30281 617616 30286 617672
rect 30342 617616 31340 617672
rect 30281 617614 31340 617616
rect 30281 617611 30347 617614
rect 31334 617612 31340 617614
rect 31404 617612 31410 617676
rect 31477 617540 31543 617541
rect 30782 617538 30788 617540
rect 28582 617478 30788 617538
rect 28582 617372 28642 617478
rect 30782 617476 30788 617478
rect 30852 617476 30858 617540
rect 31477 617536 31524 617540
rect 31588 617538 31594 617540
rect 31477 617480 31482 617536
rect 31477 617476 31524 617480
rect 31588 617478 31634 617538
rect 31588 617476 31594 617478
rect 31477 617475 31543 617476
rect 28625 616994 28691 616997
rect 28582 616992 28691 616994
rect 28582 616936 28630 616992
rect 28686 616936 28691 616992
rect 28582 616931 28691 616936
rect 28582 616828 28642 616931
rect 28625 616586 28691 616589
rect 28582 616584 28691 616586
rect 28582 616528 28630 616584
rect 28686 616528 28691 616584
rect 28582 616523 28691 616528
rect 28582 616148 28642 616523
rect 551510 616317 551570 616828
rect 456793 616314 456859 616317
rect 456793 616312 460092 616314
rect 456793 616256 456798 616312
rect 456854 616256 460092 616312
rect 456793 616254 460092 616256
rect 551461 616312 551570 616317
rect 551461 616256 551466 616312
rect 551522 616256 551570 616312
rect 551461 616254 551570 616256
rect 456793 616251 456859 616254
rect 551461 616251 551527 616254
rect 551686 616252 551692 616316
rect 551756 616314 551762 616316
rect 551829 616314 551895 616317
rect 551756 616312 551895 616314
rect 551756 616256 551834 616312
rect 551890 616256 551895 616312
rect 551756 616254 551895 616256
rect 551756 616252 551762 616254
rect 551829 616251 551895 616254
rect 28625 615906 28691 615909
rect 28582 615904 28691 615906
rect 28582 615848 28630 615904
rect 28686 615848 28691 615904
rect 28582 615843 28691 615848
rect 28582 615604 28642 615843
rect 583520 615756 584960 615996
rect 555325 615634 555391 615637
rect 551908 615632 555391 615634
rect 551908 615576 555330 615632
rect 555386 615576 555391 615632
rect 551908 615574 555391 615576
rect 555325 615571 555391 615574
rect 27470 614892 27476 614956
rect 27540 614954 27546 614956
rect 27540 614894 28060 614954
rect 27540 614892 27546 614894
rect 27286 614348 27292 614412
rect 27356 614410 27362 614412
rect 552105 614410 552171 614413
rect 27356 614350 28060 614410
rect 551908 614408 552171 614410
rect 551908 614352 552110 614408
rect 552166 614352 552171 614408
rect 551908 614350 552171 614352
rect 27356 614348 27362 614350
rect 552105 614347 552171 614350
rect 28582 613324 28642 613836
rect 312537 613458 312603 613461
rect 312537 613456 316204 613458
rect 312537 613400 312542 613456
rect 312598 613400 316204 613456
rect 312537 613398 316204 613400
rect 312537 613395 312603 613398
rect 28574 613260 28580 613324
rect 28644 613260 28650 613324
rect 27654 613124 27660 613188
rect 27724 613186 27730 613188
rect 554957 613186 555023 613189
rect 27724 613126 28060 613186
rect 551908 613184 555023 613186
rect 551908 613128 554962 613184
rect 555018 613128 555023 613184
rect 551908 613126 555023 613128
rect 27724 613124 27730 613126
rect 554957 613123 555023 613126
rect 551829 612914 551895 612917
rect 551510 612912 551895 612914
rect 551510 612856 551834 612912
rect 551890 612856 551895 612912
rect 551510 612854 551895 612856
rect 551510 612780 551570 612854
rect 551829 612851 551895 612854
rect 551502 612716 551508 612780
rect 551572 612716 551578 612780
rect 26918 612580 26924 612644
rect 26988 612642 26994 612644
rect 26988 612582 28060 612642
rect 26988 612580 26994 612582
rect 24894 611900 24900 611964
rect 24964 611962 24970 611964
rect 552197 611962 552263 611965
rect 24964 611902 28060 611962
rect 551908 611960 552263 611962
rect 551908 611904 552202 611960
rect 552258 611904 552263 611960
rect 551908 611902 552263 611904
rect 24964 611900 24970 611902
rect 552197 611899 552263 611902
rect 27102 611356 27108 611420
rect 27172 611418 27178 611420
rect 27172 611358 28060 611418
rect 27172 611356 27178 611358
rect 27838 610812 27844 610876
rect 27908 610874 27914 610876
rect 27908 610814 28060 610874
rect 27908 610812 27914 610814
rect 554129 610738 554195 610741
rect 551908 610736 554195 610738
rect 551908 610680 554134 610736
rect 554190 610680 554195 610736
rect 551908 610678 554195 610680
rect 554129 610675 554195 610678
rect -960 610466 480 610556
rect 3325 610466 3391 610469
rect -960 610464 3391 610466
rect -960 610408 3330 610464
rect 3386 610408 3391 610464
rect -960 610406 3391 610408
rect -960 610316 480 610406
rect 3325 610403 3391 610406
rect 26734 610132 26740 610196
rect 26804 610194 26810 610196
rect 26804 610134 28060 610194
rect 26804 610132 26810 610134
rect 28030 609108 28090 609620
rect 552289 609514 552355 609517
rect 551908 609512 552355 609514
rect 551908 609456 552294 609512
rect 552350 609456 552355 609512
rect 551908 609454 552355 609456
rect 552289 609451 552355 609454
rect 28022 609044 28028 609108
rect 28092 609044 28098 609108
rect 27521 608970 27587 608973
rect 27521 608968 28060 608970
rect 27521 608912 27526 608968
rect 27582 608912 28060 608968
rect 27521 608910 28060 608912
rect 27521 608907 27587 608910
rect 284385 608834 284451 608837
rect 282686 608832 284451 608834
rect 282686 608776 284390 608832
rect 284446 608776 284451 608832
rect 282686 608774 284451 608776
rect 282686 608668 282746 608774
rect 284385 608771 284451 608774
rect 25998 608364 26004 608428
rect 26068 608426 26074 608428
rect 26068 608366 28060 608426
rect 26068 608364 26074 608366
rect 555233 608290 555299 608293
rect 551908 608288 555299 608290
rect 551908 608232 555238 608288
rect 555294 608232 555299 608288
rect 551908 608230 555299 608232
rect 555233 608227 555299 608230
rect 27429 607746 27495 607749
rect 27429 607744 28060 607746
rect 27429 607688 27434 607744
rect 27490 607688 28060 607744
rect 27429 607686 28060 607688
rect 27429 607683 27495 607686
rect 28214 606796 28274 607172
rect 552381 607066 552447 607069
rect 551908 607064 552447 607066
rect 551908 607008 552386 607064
rect 552442 607008 552447 607064
rect 551908 607006 552447 607008
rect 552381 607003 552447 607006
rect 28206 606732 28212 606796
rect 28276 606732 28282 606796
rect 25221 606658 25287 606661
rect 25221 606656 28060 606658
rect 25221 606600 25226 606656
rect 25282 606600 28060 606656
rect 25221 606598 28060 606600
rect 25221 606595 25287 606598
rect 28398 605708 28458 605948
rect 554405 605842 554471 605845
rect 551908 605840 554471 605842
rect 551908 605784 554410 605840
rect 554466 605784 554471 605840
rect 551908 605782 554471 605784
rect 554405 605779 554471 605782
rect 28390 605644 28396 605708
rect 28460 605644 28466 605708
rect 28398 604893 28458 605404
rect 28349 604888 28458 604893
rect 28349 604832 28354 604888
rect 28410 604832 28458 604888
rect 28349 604830 28458 604832
rect 28349 604827 28415 604830
rect 25630 604692 25636 604756
rect 25700 604754 25706 604756
rect 25700 604694 28060 604754
rect 25700 604692 25706 604694
rect 552473 604618 552539 604621
rect 551908 604616 552539 604618
rect 551908 604560 552478 604616
rect 552534 604560 552539 604616
rect 551908 604558 552539 604560
rect 552473 604555 552539 604558
rect 551732 604284 551738 604348
rect 551802 604346 551808 604348
rect 551921 604346 551987 604349
rect 551802 604344 551987 604346
rect 551802 604288 551926 604344
rect 551982 604288 551987 604344
rect 551802 604286 551987 604288
rect 551802 604284 551808 604286
rect 551921 604283 551987 604286
rect 578877 604210 578943 604213
rect 583520 604210 584960 604300
rect 578877 604208 584960 604210
rect 28030 603805 28090 604180
rect 578877 604152 578882 604208
rect 578938 604152 584960 604208
rect 578877 604150 584960 604152
rect 578877 604147 578943 604150
rect 583520 604060 584960 604150
rect 27981 603800 28090 603805
rect 27981 603744 27986 603800
rect 28042 603744 28090 603800
rect 27981 603742 28090 603744
rect 27981 603739 28047 603742
rect 27613 603666 27679 603669
rect 27613 603664 28060 603666
rect 27613 603608 27618 603664
rect 27674 603608 28060 603664
rect 27613 603606 28060 603608
rect 27613 603603 27679 603606
rect 551694 603125 551754 603364
rect 551694 603120 551803 603125
rect 551694 603064 551742 603120
rect 551798 603064 551803 603120
rect 551694 603062 551803 603064
rect 551737 603059 551803 603062
rect 25814 602924 25820 602988
rect 25884 602986 25890 602988
rect 25884 602926 28060 602986
rect 25884 602924 25890 602926
rect 551318 602788 551324 602852
rect 551388 602850 551394 602852
rect 551686 602850 551692 602852
rect 551388 602790 551692 602850
rect 551388 602788 551394 602790
rect 551686 602788 551692 602790
rect 551756 602788 551762 602852
rect 27337 602442 27403 602445
rect 27337 602440 28060 602442
rect 27337 602384 27342 602440
rect 27398 602384 28060 602440
rect 27337 602382 28060 602384
rect 27337 602379 27403 602382
rect 552565 602170 552631 602173
rect 551908 602168 552631 602170
rect 551908 602112 552570 602168
rect 552626 602112 552631 602168
rect 551908 602110 552631 602112
rect 552565 602107 552631 602110
rect 24761 601762 24827 601765
rect 24761 601760 28060 601762
rect 24761 601704 24766 601760
rect 24822 601704 28060 601760
rect 24761 601702 28060 601704
rect 24761 601699 24827 601702
rect 25262 601156 25268 601220
rect 25332 601218 25338 601220
rect 25332 601158 28060 601218
rect 25332 601156 25338 601158
rect 552933 600946 552999 600949
rect 551908 600944 552999 600946
rect 551908 600888 552938 600944
rect 552994 600888 552999 600944
rect 551908 600886 552999 600888
rect 552933 600883 552999 600886
rect 28582 600133 28642 600508
rect 28533 600128 28642 600133
rect 28533 600072 28538 600128
rect 28594 600072 28642 600128
rect 28533 600070 28642 600072
rect 28533 600067 28599 600070
rect 27245 599994 27311 599997
rect 27245 599992 28060 599994
rect 27245 599936 27250 599992
rect 27306 599936 28060 599992
rect 27245 599934 28060 599936
rect 27245 599931 27311 599934
rect 552749 599722 552815 599725
rect 551908 599720 552815 599722
rect 551908 599664 552754 599720
rect 552810 599664 552815 599720
rect 551908 599662 552815 599664
rect 552749 599659 552815 599662
rect 28398 599045 28458 599420
rect 28398 599040 28507 599045
rect 28398 598984 28446 599040
rect 28502 598984 28507 599040
rect 28398 598982 28507 598984
rect 28441 598979 28507 598982
rect 25773 598770 25839 598773
rect 25773 598768 28060 598770
rect 25773 598712 25778 598768
rect 25834 598712 28060 598768
rect 25773 598710 28060 598712
rect 25773 598707 25839 598710
rect 553025 598498 553091 598501
rect 551908 598496 553091 598498
rect 551908 598440 553030 598496
rect 553086 598440 553091 598496
rect 551908 598438 553091 598440
rect 553025 598435 553091 598438
rect 28625 598364 28691 598365
rect 28620 598362 28626 598364
rect 28534 598302 28626 598362
rect 28620 598300 28626 598302
rect 28690 598300 28696 598364
rect 28625 598299 28691 598300
rect 28582 597684 28642 598196
rect 28574 597620 28580 597684
rect 28644 597620 28650 597684
rect 27153 597546 27219 597549
rect 27153 597544 28060 597546
rect 27153 597488 27158 597544
rect 27214 597488 28060 597544
rect 27153 597486 28060 597488
rect 27153 597483 27219 597486
rect 552841 597274 552907 597277
rect 551908 597272 552907 597274
rect 551908 597216 552846 597272
rect 552902 597216 552907 597272
rect 551908 597214 552907 597216
rect 552841 597211 552907 597214
rect 27705 597002 27771 597005
rect 27705 597000 28060 597002
rect 27705 596944 27710 597000
rect 27766 596944 28060 597000
rect 27705 596942 28060 596944
rect 27705 596939 27771 596942
rect 28349 596730 28415 596733
rect 28574 596730 28580 596732
rect 28349 596728 28580 596730
rect 28349 596672 28354 596728
rect 28410 596672 28580 596728
rect 28349 596670 28580 596672
rect 28349 596667 28415 596670
rect 28574 596668 28580 596670
rect 28644 596668 28650 596732
rect 25221 596458 25287 596461
rect 25221 596456 28060 596458
rect 25221 596400 25226 596456
rect 25282 596400 28060 596456
rect 25221 596398 28060 596400
rect 25221 596395 25287 596398
rect -960 596050 480 596140
rect 3509 596050 3575 596053
rect 554589 596050 554655 596053
rect -960 596048 3575 596050
rect -960 595992 3514 596048
rect 3570 595992 3575 596048
rect -960 595990 3575 595992
rect 551908 596048 554655 596050
rect 551908 595992 554594 596048
rect 554650 595992 554655 596048
rect 551908 595990 554655 595992
rect -960 595900 480 595990
rect 3509 595987 3575 595990
rect 554589 595987 554655 595990
rect 28214 595373 28274 595748
rect 28214 595368 28323 595373
rect 28214 595312 28262 595368
rect 28318 595312 28323 595368
rect 28214 595310 28323 595312
rect 28257 595307 28323 595310
rect 27061 595234 27127 595237
rect 27061 595232 28060 595234
rect 27061 595176 27066 595232
rect 27122 595176 28060 595232
rect 27061 595174 28060 595176
rect 27061 595171 27127 595174
rect 139577 594826 139643 594829
rect 552657 594826 552723 594829
rect 139534 594824 139643 594826
rect 139534 594768 139582 594824
rect 139638 594768 139643 594824
rect 139534 594763 139643 594768
rect 551908 594824 552723 594826
rect 551908 594768 552662 594824
rect 552718 594768 552723 594824
rect 551908 594766 552723 594768
rect 552657 594763 552723 594766
rect 28349 594690 28415 594693
rect 28574 594690 28580 594692
rect 28349 594688 28580 594690
rect 28349 594632 28354 594688
rect 28410 594632 28580 594688
rect 28349 594630 28580 594632
rect 28349 594627 28415 594630
rect 28574 594628 28580 594630
rect 28644 594628 28650 594692
rect 139534 594660 139594 594763
rect 28582 594149 28642 594524
rect 28582 594144 28691 594149
rect 28582 594088 28630 594144
rect 28686 594088 28691 594144
rect 28582 594086 28691 594088
rect 28625 594083 28691 594086
rect 28214 593469 28274 593980
rect 551870 593948 551876 594012
rect 551940 594010 551946 594012
rect 554037 594010 554103 594013
rect 551940 594008 554103 594010
rect 551940 593952 554042 594008
rect 554098 593952 554103 594008
rect 551940 593950 554103 593952
rect 551940 593948 551946 593950
rect 554037 593947 554103 593950
rect 554037 593738 554103 593741
rect 551908 593736 554103 593738
rect 551908 593680 554042 593736
rect 554098 593680 554103 593736
rect 551908 593678 554103 593680
rect 554037 593675 554103 593678
rect 28165 593464 28274 593469
rect 28533 593468 28599 593469
rect 28533 593466 28580 593468
rect 28165 593408 28170 593464
rect 28226 593408 28274 593464
rect 28165 593406 28274 593408
rect 28488 593464 28580 593466
rect 28488 593408 28538 593464
rect 28488 593406 28580 593408
rect 28165 593403 28231 593406
rect 28533 593404 28580 593406
rect 28644 593404 28650 593468
rect 551318 593404 551324 593468
rect 551388 593466 551394 593468
rect 551686 593466 551692 593468
rect 551388 593406 551692 593466
rect 551388 593404 551394 593406
rect 551686 593404 551692 593406
rect 551756 593404 551762 593468
rect 28533 593403 28599 593404
rect 27797 593330 27863 593333
rect 27797 593328 28060 593330
rect 27797 593272 27802 593328
rect 27858 593272 28060 593328
rect 27797 593270 28060 593272
rect 27797 593267 27863 593270
rect 28582 592381 28642 592756
rect 554129 592514 554195 592517
rect 551908 592512 554195 592514
rect 551908 592456 554134 592512
rect 554190 592456 554195 592512
rect 551908 592454 554195 592456
rect 554129 592451 554195 592454
rect 580533 592514 580599 592517
rect 583520 592514 584960 592604
rect 580533 592512 584960 592514
rect 580533 592456 580538 592512
rect 580594 592456 584960 592512
rect 580533 592454 584960 592456
rect 580533 592451 580599 592454
rect 28582 592376 28691 592381
rect 28582 592320 28630 592376
rect 28686 592320 28691 592376
rect 583520 592364 584960 592454
rect 28582 592318 28691 592320
rect 28625 592315 28691 592318
rect 25262 592242 25268 592244
rect 25086 592182 25268 592242
rect 25086 591972 25146 592182
rect 25262 592180 25268 592182
rect 25332 592180 25338 592244
rect 25078 591908 25084 591972
rect 25148 591908 25154 591972
rect 28030 591701 28090 592212
rect 28349 591970 28415 591973
rect 28574 591970 28580 591972
rect 28349 591968 28580 591970
rect 28349 591912 28354 591968
rect 28410 591912 28580 591968
rect 28349 591910 28580 591912
rect 28349 591907 28415 591910
rect 28574 591908 28580 591910
rect 28644 591908 28650 591972
rect 28030 591696 28139 591701
rect 455413 591698 455479 591701
rect 28030 591640 28078 591696
rect 28134 591640 28139 591696
rect 28030 591638 28139 591640
rect 454020 591696 455479 591698
rect 454020 591640 455418 591696
rect 455474 591640 455479 591696
rect 454020 591638 455479 591640
rect 28073 591635 28139 591638
rect 455413 591635 455479 591638
rect 26049 591562 26115 591565
rect 26049 591560 28060 591562
rect 26049 591504 26054 591560
rect 26110 591504 28060 591560
rect 26049 591502 28060 591504
rect 26049 591499 26115 591502
rect 28533 591292 28599 591293
rect 28533 591288 28580 591292
rect 28644 591290 28650 591292
rect 554497 591290 554563 591293
rect 28533 591232 28538 591288
rect 28533 591228 28580 591232
rect 28644 591230 28690 591290
rect 551908 591288 554563 591290
rect 551908 591232 554502 591288
rect 554558 591232 554563 591288
rect 551908 591230 554563 591232
rect 28644 591228 28650 591230
rect 28533 591227 28599 591228
rect 554497 591227 554563 591230
rect 27889 590746 27955 590749
rect 28030 590746 28090 590988
rect 27889 590744 28090 590746
rect 27889 590688 27894 590744
rect 27950 590688 28090 590744
rect 27889 590686 28090 590688
rect 27889 590683 27955 590686
rect 26969 590338 27035 590341
rect 26969 590336 28060 590338
rect 26969 590280 26974 590336
rect 27030 590280 28060 590336
rect 26969 590278 28060 590280
rect 26969 590275 27035 590278
rect 554497 590066 554563 590069
rect 551908 590064 554563 590066
rect 551908 590008 554502 590064
rect 554558 590008 554563 590064
rect 551908 590006 554563 590008
rect 554497 590003 554563 590006
rect 28582 589389 28642 589764
rect 28582 589384 28691 589389
rect 28582 589328 28630 589384
rect 28686 589328 28691 589384
rect 28582 589326 28691 589328
rect 28625 589323 28691 589326
rect 28398 588709 28458 589220
rect 554313 588842 554379 588845
rect 551908 588840 554379 588842
rect 551908 588784 554318 588840
rect 554374 588784 554379 588840
rect 551908 588782 554379 588784
rect 554313 588779 554379 588782
rect 28349 588704 28458 588709
rect 28349 588648 28354 588704
rect 28410 588648 28458 588704
rect 28349 588646 28458 588648
rect 28349 588643 28415 588646
rect 28582 588165 28642 588540
rect 551318 588508 551324 588572
rect 551388 588570 551394 588572
rect 551829 588570 551895 588573
rect 551388 588568 551895 588570
rect 551388 588512 551834 588568
rect 551890 588512 551895 588568
rect 551388 588510 551895 588512
rect 551388 588508 551394 588510
rect 551829 588507 551895 588510
rect 28533 588160 28642 588165
rect 28533 588104 28538 588160
rect 28594 588104 28642 588160
rect 28533 588102 28642 588104
rect 28533 588099 28599 588102
rect 25078 587828 25084 587892
rect 25148 587828 25154 587892
rect 25086 587754 25146 587828
rect 28582 587757 28642 587996
rect 25313 587754 25379 587757
rect 25086 587752 25379 587754
rect 25086 587696 25318 587752
rect 25374 587696 25379 587752
rect 25086 587694 25379 587696
rect 28582 587752 28691 587757
rect 28582 587696 28630 587752
rect 28686 587696 28691 587752
rect 28582 587694 28691 587696
rect 25313 587691 25379 587694
rect 28625 587691 28691 587694
rect 554313 587618 554379 587621
rect 551908 587616 554379 587618
rect 551908 587560 554318 587616
rect 554374 587560 554379 587616
rect 551908 587558 554379 587560
rect 554313 587555 554379 587558
rect 28625 587482 28691 587485
rect 28582 587480 28691 587482
rect 28582 587424 28630 587480
rect 28686 587424 28691 587480
rect 28582 587419 28691 587424
rect 28582 587316 28642 587419
rect 25957 586802 26023 586805
rect 25957 586800 28060 586802
rect 25957 586744 25962 586800
rect 26018 586744 28060 586800
rect 25957 586742 28060 586744
rect 25957 586739 26023 586742
rect 554497 586394 554563 586397
rect 551908 586392 554563 586394
rect 551908 586336 554502 586392
rect 554558 586336 554563 586392
rect 551908 586334 554563 586336
rect 554497 586331 554563 586334
rect 28582 585717 28642 586092
rect 283005 585986 283071 585989
rect 282686 585984 283071 585986
rect 282686 585928 283010 585984
rect 283066 585928 283071 585984
rect 282686 585926 283071 585928
rect 28582 585712 28691 585717
rect 28582 585656 28630 585712
rect 28686 585656 28691 585712
rect 28582 585654 28691 585656
rect 28625 585651 28691 585654
rect 26877 585578 26943 585581
rect 26877 585576 28060 585578
rect 26877 585520 26882 585576
rect 26938 585520 28060 585576
rect 282686 585548 282746 585926
rect 283005 585923 283071 585926
rect 26877 585518 28060 585520
rect 26877 585515 26943 585518
rect 554313 585170 554379 585173
rect 551908 585168 554379 585170
rect 551908 585112 554318 585168
rect 554374 585112 554379 585168
rect 551908 585110 554379 585112
rect 554313 585107 554379 585110
rect 26141 585034 26207 585037
rect 26141 585032 28060 585034
rect 26141 584976 26146 585032
rect 26202 584976 28060 585032
rect 26141 584974 28060 584976
rect 26141 584971 26207 584974
rect 28582 583949 28642 584324
rect 28582 583944 28691 583949
rect 554313 583946 554379 583949
rect 28582 583888 28630 583944
rect 28686 583888 28691 583944
rect 28582 583886 28691 583888
rect 551908 583944 554379 583946
rect 551908 583888 554318 583944
rect 554374 583888 554379 583944
rect 551908 583886 554379 583888
rect 28625 583883 28691 583886
rect 554313 583883 554379 583886
rect 24669 583810 24735 583813
rect 24669 583808 28060 583810
rect 24669 583752 24674 583808
rect 24730 583752 28060 583808
rect 24669 583750 28060 583752
rect 24669 583747 24735 583750
rect 25865 583130 25931 583133
rect 25865 583128 28060 583130
rect 25865 583072 25870 583128
rect 25926 583072 28060 583128
rect 25865 583070 28060 583072
rect 25865 583067 25931 583070
rect 555417 582722 555483 582725
rect 551908 582720 555483 582722
rect 551908 582664 555422 582720
rect 555478 582664 555483 582720
rect 551908 582662 555483 582664
rect 555417 582659 555483 582662
rect 25129 582586 25195 582589
rect 25129 582584 28060 582586
rect 25129 582528 25134 582584
rect 25190 582528 28060 582584
rect 25129 582526 28060 582528
rect 25129 582523 25195 582526
rect 551686 582524 551692 582588
rect 551756 582524 551762 582588
rect 551694 582314 551754 582524
rect 551870 582314 551876 582316
rect 551694 582254 551876 582314
rect 551870 582252 551876 582254
rect 551940 582252 551946 582316
rect -960 581620 480 581860
rect 28030 581501 28090 582012
rect 28030 581496 28139 581501
rect 554313 581498 554379 581501
rect 28030 581440 28078 581496
rect 28134 581440 28139 581496
rect 28030 581438 28139 581440
rect 551908 581496 554379 581498
rect 551908 581440 554318 581496
rect 554374 581440 554379 581496
rect 551908 581438 554379 581440
rect 28073 581435 28139 581438
rect 554313 581435 554379 581438
rect 28582 580957 28642 581332
rect 28533 580952 28642 580957
rect 28533 580896 28538 580952
rect 28594 580896 28642 580952
rect 28533 580894 28642 580896
rect 28533 580891 28599 580894
rect 25681 580818 25747 580821
rect 580441 580818 580507 580821
rect 583520 580818 584960 580908
rect 25681 580816 28060 580818
rect 25681 580760 25686 580816
rect 25742 580760 28060 580816
rect 25681 580758 28060 580760
rect 580441 580816 584960 580818
rect 580441 580760 580446 580816
rect 580502 580760 584960 580816
rect 580441 580758 584960 580760
rect 25681 580755 25747 580758
rect 580441 580755 580507 580758
rect 583520 580668 584960 580758
rect 554313 580274 554379 580277
rect 551908 580272 554379 580274
rect 551908 580216 554318 580272
rect 554374 580216 554379 580272
rect 551908 580214 554379 580216
rect 554313 580211 554379 580214
rect 26601 580138 26667 580141
rect 26601 580136 28060 580138
rect 26601 580080 26606 580136
rect 26662 580080 28060 580136
rect 26601 580078 28060 580080
rect 26601 580075 26667 580078
rect 28214 579053 28274 579564
rect 28214 579048 28323 579053
rect 554313 579050 554379 579053
rect 28214 578992 28262 579048
rect 28318 578992 28323 579048
rect 28214 578990 28323 578992
rect 551908 579048 554379 579050
rect 551908 578992 554318 579048
rect 554374 578992 554379 579048
rect 551908 578990 554379 578992
rect 28257 578987 28323 578990
rect 554313 578987 554379 578990
rect 26141 578914 26207 578917
rect 26141 578912 28060 578914
rect 26141 578856 26146 578912
rect 26202 578856 28060 578912
rect 26141 578854 28060 578856
rect 26141 578851 26207 578854
rect 25405 578370 25471 578373
rect 25405 578368 28060 578370
rect 25405 578312 25410 578368
rect 25466 578312 28060 578368
rect 25405 578310 28060 578312
rect 25405 578307 25471 578310
rect 26693 577826 26759 577829
rect 554313 577826 554379 577829
rect 26693 577824 28060 577826
rect 26693 577768 26698 577824
rect 26754 577768 28060 577824
rect 26693 577766 28060 577768
rect 551908 577824 554379 577826
rect 551908 577768 554318 577824
rect 554374 577768 554379 577824
rect 551908 577766 554379 577768
rect 26693 577763 26759 577766
rect 554313 577763 554379 577766
rect 25037 577146 25103 577149
rect 25037 577144 28060 577146
rect 25037 577088 25042 577144
rect 25098 577088 28060 577144
rect 25037 577086 28060 577088
rect 25037 577083 25103 577086
rect 551318 576948 551324 577012
rect 551388 577010 551394 577012
rect 551686 577010 551692 577012
rect 551388 576950 551692 577010
rect 551388 576948 551394 576950
rect 551686 576948 551692 576950
rect 551756 576948 551762 577012
rect 25630 576540 25636 576604
rect 25700 576602 25706 576604
rect 26366 576602 26372 576604
rect 25700 576542 26372 576602
rect 25700 576540 25706 576542
rect 26366 576540 26372 576542
rect 26436 576540 26442 576604
rect 26785 576602 26851 576605
rect 554405 576602 554471 576605
rect 26785 576600 28060 576602
rect 26785 576544 26790 576600
rect 26846 576544 28060 576600
rect 26785 576542 28060 576544
rect 551908 576600 554471 576602
rect 551908 576544 554410 576600
rect 554466 576544 554471 576600
rect 551908 576542 554471 576544
rect 26785 576539 26851 576542
rect 554405 576539 554471 576542
rect 28214 575653 28274 575892
rect 28214 575648 28323 575653
rect 28214 575592 28262 575648
rect 28318 575592 28323 575648
rect 28214 575590 28323 575592
rect 28257 575587 28323 575590
rect 24945 575378 25011 575381
rect 554313 575378 554379 575381
rect 24945 575376 28060 575378
rect 24945 575320 24950 575376
rect 25006 575320 28060 575376
rect 24945 575318 28060 575320
rect 551908 575376 554379 575378
rect 551908 575320 554318 575376
rect 554374 575320 554379 575376
rect 551908 575318 554379 575320
rect 24945 575315 25011 575318
rect 554313 575315 554379 575318
rect 28214 574293 28274 574804
rect 28214 574288 28323 574293
rect 28214 574232 28262 574288
rect 28318 574232 28323 574288
rect 28214 574230 28323 574232
rect 28257 574227 28323 574230
rect 25497 574154 25563 574157
rect 554405 574154 554471 574157
rect 25497 574152 28060 574154
rect 25497 574096 25502 574152
rect 25558 574096 28060 574152
rect 25497 574094 28060 574096
rect 551908 574152 554471 574154
rect 551908 574096 554410 574152
rect 554466 574096 554471 574152
rect 551908 574094 554471 574096
rect 25497 574091 25563 574094
rect 554405 574091 554471 574094
rect 26325 573610 26391 573613
rect 26325 573608 28060 573610
rect 26325 573552 26330 573608
rect 26386 573552 28060 573608
rect 26325 573550 28060 573552
rect 26325 573547 26391 573550
rect 551502 573412 551508 573476
rect 551572 573474 551578 573476
rect 551870 573474 551876 573476
rect 551572 573414 551876 573474
rect 551572 573412 551578 573414
rect 551870 573412 551876 573414
rect 551940 573412 551946 573476
rect 24577 572930 24643 572933
rect 554405 572930 554471 572933
rect 24577 572928 28060 572930
rect 24577 572872 24582 572928
rect 24638 572872 28060 572928
rect 24577 572870 28060 572872
rect 551908 572928 554471 572930
rect 551908 572872 554410 572928
rect 554466 572872 554471 572928
rect 551908 572870 554471 572872
rect 24577 572867 24643 572870
rect 554405 572867 554471 572870
rect 24485 572386 24551 572389
rect 24485 572384 28060 572386
rect 24485 572328 24490 572384
rect 24546 572328 28060 572384
rect 24485 572326 28060 572328
rect 24485 572323 24551 572326
rect 20478 571916 20484 571980
rect 20548 571978 20554 571980
rect 24117 571978 24183 571981
rect 20548 571976 24183 571978
rect 20548 571920 24122 571976
rect 24178 571920 24183 571976
rect 20548 571918 24183 571920
rect 20548 571916 20554 571918
rect 24117 571915 24183 571918
rect 25589 571842 25655 571845
rect 25589 571840 28060 571842
rect 25589 571784 25594 571840
rect 25650 571784 28060 571840
rect 25589 571782 28060 571784
rect 25589 571779 25655 571782
rect 554221 571706 554287 571709
rect 551908 571704 554287 571706
rect 551908 571648 554226 571704
rect 554282 571648 554287 571704
rect 551908 571646 554287 571648
rect 554221 571643 554287 571646
rect 29494 571372 29500 571436
rect 29564 571434 29570 571436
rect 30414 571434 30420 571436
rect 29564 571374 30420 571434
rect 29564 571372 29570 571374
rect 30414 571372 30420 571374
rect 30484 571372 30490 571436
rect 25313 570618 25379 570621
rect 76005 570618 76071 570621
rect 554405 570618 554471 570621
rect 25313 570616 76071 570618
rect 25313 570560 25318 570616
rect 25374 570560 76010 570616
rect 76066 570560 76071 570616
rect 25313 570558 76071 570560
rect 551908 570616 554471 570618
rect 551908 570560 554410 570616
rect 554466 570560 554471 570616
rect 551908 570558 554471 570560
rect 25313 570555 25379 570558
rect 76005 570555 76071 570558
rect 554405 570555 554471 570558
rect 550766 570420 550772 570484
rect 550836 570482 550842 570484
rect 551686 570482 551692 570484
rect 550836 570422 551692 570482
rect 550836 570420 550842 570422
rect 551686 570420 551692 570422
rect 551756 570420 551762 570484
rect 551502 570012 551508 570076
rect 551572 570074 551578 570076
rect 551870 570074 551876 570076
rect 551572 570014 551876 570074
rect 551572 570012 551578 570014
rect 551870 570012 551876 570014
rect 551940 570012 551946 570076
rect 583520 568836 584960 569076
rect 283189 568578 283255 568581
rect 283373 568578 283439 568581
rect 283189 568576 283439 568578
rect 283189 568520 283194 568576
rect 283250 568520 283378 568576
rect 283434 568520 283439 568576
rect 283189 568518 283439 568520
rect 283189 568515 283255 568518
rect 283373 568515 283439 568518
rect 29310 567836 29316 567900
rect 29380 567898 29386 567900
rect 29862 567898 29868 567900
rect 29380 567838 29868 567898
rect 29380 567836 29386 567838
rect 29862 567836 29868 567838
rect 29932 567836 29938 567900
rect 551001 567762 551067 567765
rect 551870 567762 551876 567764
rect 551001 567760 551876 567762
rect 551001 567704 551006 567760
rect 551062 567704 551876 567760
rect 551001 567702 551876 567704
rect 551001 567699 551067 567702
rect 551870 567700 551876 567702
rect 551940 567700 551946 567764
rect 550582 567564 550588 567628
rect 550652 567626 550658 567628
rect 551870 567626 551876 567628
rect 550652 567566 551876 567626
rect 550652 567564 550658 567566
rect 551870 567564 551876 567566
rect 551940 567564 551946 567628
rect 29085 567492 29151 567493
rect 29085 567490 29132 567492
rect 29040 567488 29132 567490
rect -960 567354 480 567444
rect 29040 567432 29090 567488
rect 29040 567430 29132 567432
rect 29085 567428 29132 567430
rect 29196 567428 29202 567492
rect 29085 567427 29151 567428
rect 3509 567354 3575 567357
rect -960 567352 3575 567354
rect -960 567296 3514 567352
rect 3570 567296 3575 567352
rect -960 567294 3575 567296
rect -960 567204 480 567294
rect 3509 567291 3575 567294
rect 29678 565660 29684 565724
rect 29748 565660 29754 565724
rect 29126 565388 29132 565452
rect 29196 565450 29202 565452
rect 29686 565450 29746 565660
rect 29196 565390 29746 565450
rect 29196 565388 29202 565390
rect 551318 563212 551324 563276
rect 551388 563212 551394 563276
rect 551326 563004 551386 563212
rect 551318 562940 551324 563004
rect 551388 562940 551394 563004
rect 29310 560764 29316 560828
rect 29380 560826 29386 560828
rect 29862 560826 29868 560828
rect 29380 560766 29868 560826
rect 29380 560764 29386 560766
rect 29862 560764 29868 560766
rect 29932 560764 29938 560828
rect 551001 559194 551067 559197
rect 551001 559192 551570 559194
rect 551001 559136 551006 559192
rect 551062 559136 551570 559192
rect 551001 559134 551570 559136
rect 551001 559131 551067 559134
rect 551510 559060 551570 559134
rect 551502 558996 551508 559060
rect 551572 558996 551578 559060
rect 28942 558452 28948 558516
rect 29012 558514 29018 558516
rect 29494 558514 29500 558516
rect 29012 558454 29500 558514
rect 29012 558452 29018 558454
rect 29494 558452 29500 558454
rect 29564 558452 29570 558516
rect 29085 558378 29151 558381
rect 29494 558378 29500 558380
rect 29085 558376 29500 558378
rect 29085 558320 29090 558376
rect 29146 558320 29500 558376
rect 29085 558318 29500 558320
rect 29085 558315 29151 558318
rect 29494 558316 29500 558318
rect 29564 558316 29570 558380
rect 550582 558180 550588 558244
rect 550652 558242 550658 558244
rect 551686 558242 551692 558244
rect 550652 558182 551692 558242
rect 550652 558180 550658 558182
rect 551686 558180 551692 558182
rect 551756 558180 551762 558244
rect 30005 557428 30071 557429
rect 30005 557424 30052 557428
rect 30116 557426 30122 557428
rect 30005 557368 30010 557424
rect 30005 557364 30052 557368
rect 30116 557366 30162 557426
rect 30116 557364 30122 557366
rect 30005 557363 30071 557364
rect 579797 557290 579863 557293
rect 583520 557290 584960 557380
rect 579797 557288 584960 557290
rect 579797 557232 579802 557288
rect 579858 557232 584960 557288
rect 579797 557230 584960 557232
rect 579797 557227 579863 557230
rect 30005 557154 30071 557157
rect 30230 557154 30236 557156
rect 30005 557152 30236 557154
rect 30005 557096 30010 557152
rect 30066 557096 30236 557152
rect 30005 557094 30236 557096
rect 30005 557091 30071 557094
rect 30230 557092 30236 557094
rect 30300 557092 30306 557156
rect 583520 557140 584960 557230
rect 550766 553964 550772 554028
rect 550836 554026 550842 554028
rect 551502 554026 551508 554028
rect 550836 553966 551508 554026
rect 550836 553964 550842 553966
rect 551502 553964 551508 553966
rect 551572 553964 551578 554028
rect -960 553074 480 553164
rect 3141 553074 3207 553077
rect -960 553072 3207 553074
rect -960 553016 3146 553072
rect 3202 553016 3207 553072
rect -960 553014 3207 553016
rect -960 552924 480 553014
rect 3141 553011 3207 553014
rect 28942 547708 28948 547772
rect 29012 547708 29018 547772
rect 28950 547634 29010 547708
rect 29177 547634 29243 547637
rect 28950 547632 29243 547634
rect 28950 547576 29182 547632
rect 29238 547576 29243 547632
rect 28950 547574 29243 547576
rect 29177 547571 29243 547574
rect 25814 547028 25820 547092
rect 25884 547090 25890 547092
rect 78673 547090 78739 547093
rect 25884 547088 78739 547090
rect 25884 547032 78678 547088
rect 78734 547032 78739 547088
rect 25884 547030 78739 547032
rect 25884 547028 25890 547030
rect 78673 547027 78739 547030
rect 520181 547090 520247 547093
rect 552790 547090 552796 547092
rect 520181 547088 552796 547090
rect 520181 547032 520186 547088
rect 520242 547032 552796 547088
rect 520181 547030 552796 547032
rect 520181 547027 520247 547030
rect 552790 547028 552796 547030
rect 552860 547028 552866 547092
rect 29126 545804 29132 545868
rect 29196 545866 29202 545868
rect 29678 545866 29684 545868
rect 29196 545806 29684 545866
rect 29196 545804 29202 545806
rect 29678 545804 29684 545806
rect 29748 545804 29754 545868
rect 580901 545594 580967 545597
rect 583520 545594 584960 545684
rect 580901 545592 584960 545594
rect 580901 545536 580906 545592
rect 580962 545536 584960 545592
rect 580901 545534 584960 545536
rect 580901 545531 580967 545534
rect 583520 545444 584960 545534
rect 551134 543764 551140 543828
rect 551204 543826 551210 543828
rect 551870 543826 551876 543828
rect 551204 543766 551876 543826
rect 551204 543764 551210 543766
rect 551870 543764 551876 543766
rect 551940 543764 551946 543828
rect 551134 543628 551140 543692
rect 551204 543690 551210 543692
rect 551502 543690 551508 543692
rect 551204 543630 551508 543690
rect 551204 543628 551210 543630
rect 551502 543628 551508 543630
rect 551572 543628 551578 543692
rect 30046 540908 30052 540972
rect 30116 540970 30122 540972
rect 30465 540970 30531 540973
rect 30116 540968 30531 540970
rect 30116 540912 30470 540968
rect 30526 540912 30531 540968
rect 30116 540910 30531 540912
rect 30116 540908 30122 540910
rect 30465 540907 30531 540910
rect 550725 539610 550791 539613
rect 550909 539610 550975 539613
rect 550725 539608 550975 539610
rect 550725 539552 550730 539608
rect 550786 539552 550914 539608
rect 550970 539552 550975 539608
rect 550725 539550 550975 539552
rect 550725 539547 550791 539550
rect 550909 539547 550975 539550
rect -960 538658 480 538748
rect 3509 538658 3575 538661
rect -960 538656 3575 538658
rect -960 538600 3514 538656
rect 3570 538600 3575 538656
rect -960 538598 3575 538600
rect -960 538508 480 538598
rect 3509 538595 3575 538598
rect 29310 538324 29316 538388
rect 29380 538386 29386 538388
rect 29380 538326 29562 538386
rect 29380 538324 29386 538326
rect 29502 538252 29562 538326
rect 29494 538188 29500 538252
rect 29564 538188 29570 538252
rect 28022 534924 28028 534988
rect 28092 534986 28098 534988
rect 91001 534986 91067 534989
rect 28092 534984 91067 534986
rect 28092 534928 91006 534984
rect 91062 534928 91067 534984
rect 28092 534926 91067 534928
rect 28092 534924 28098 534926
rect 91001 534923 91067 534926
rect 25998 534788 26004 534852
rect 26068 534850 26074 534852
rect 88885 534850 88951 534853
rect 26068 534848 88951 534850
rect 26068 534792 88890 534848
rect 88946 534792 88951 534848
rect 26068 534790 88951 534792
rect 26068 534788 26074 534790
rect 88885 534787 88951 534790
rect 27838 534652 27844 534716
rect 27908 534714 27914 534716
rect 93209 534714 93275 534717
rect 27908 534712 93275 534714
rect 27908 534656 93214 534712
rect 93270 534656 93275 534712
rect 27908 534654 93275 534656
rect 27908 534652 27914 534654
rect 93209 534651 93275 534654
rect 141693 534442 141759 534445
rect 454769 534442 454835 534445
rect 141693 534440 454835 534442
rect 141693 534384 141698 534440
rect 141754 534384 454774 534440
rect 454830 534384 454835 534440
rect 141693 534382 454835 534384
rect 141693 534379 141759 534382
rect 454769 534379 454835 534382
rect 131941 534306 132007 534309
rect 464521 534306 464587 534309
rect 131941 534304 464587 534306
rect 131941 534248 131946 534304
rect 132002 534248 464526 534304
rect 464582 534248 464587 534304
rect 131941 534246 464587 534248
rect 131941 534243 132007 534246
rect 464521 534243 464587 534246
rect 114737 534170 114803 534173
rect 481725 534170 481791 534173
rect 114737 534168 481791 534170
rect 114737 534112 114742 534168
rect 114798 534112 481730 534168
rect 481786 534112 481791 534168
rect 114737 534110 481791 534112
rect 114737 534107 114803 534110
rect 481725 534107 481791 534110
rect 28390 533836 28396 533900
rect 28460 533898 28466 533900
rect 84561 533898 84627 533901
rect 28460 533896 84627 533898
rect 28460 533840 84566 533896
rect 84622 533840 84627 533896
rect 28460 533838 84627 533840
rect 28460 533836 28466 533838
rect 84561 533835 84627 533838
rect 28206 533700 28212 533764
rect 28276 533762 28282 533764
rect 86677 533762 86743 533765
rect 28276 533760 86743 533762
rect 28276 533704 86682 533760
rect 86738 533704 86743 533760
rect 583520 533748 584960 533988
rect 28276 533702 86743 533704
rect 28276 533700 28282 533702
rect 86677 533699 86743 533702
rect 30230 533564 30236 533628
rect 30300 533626 30306 533628
rect 30465 533626 30531 533629
rect 30300 533624 30531 533626
rect 30300 533568 30470 533624
rect 30526 533568 30531 533624
rect 30300 533566 30531 533568
rect 30300 533564 30306 533566
rect 30465 533563 30531 533566
rect 31150 533564 31156 533628
rect 31220 533626 31226 533628
rect 101765 533626 101831 533629
rect 31220 533624 101831 533626
rect 31220 533568 101770 533624
rect 101826 533568 101831 533624
rect 31220 533566 101831 533568
rect 31220 533564 31226 533566
rect 101765 533563 101831 533566
rect 506105 533626 506171 533629
rect 551502 533626 551508 533628
rect 506105 533624 551508 533626
rect 506105 533568 506110 533624
rect 506166 533568 551508 533624
rect 506105 533566 551508 533568
rect 506105 533563 506171 533566
rect 551502 533564 551508 533566
rect 551572 533564 551578 533628
rect 31334 533428 31340 533492
rect 31404 533490 31410 533492
rect 102869 533490 102935 533493
rect 31404 533488 102935 533490
rect 31404 533432 102874 533488
rect 102930 533432 102935 533488
rect 31404 533430 102935 533432
rect 31404 533428 31410 533430
rect 102869 533427 102935 533430
rect 501781 533490 501847 533493
rect 554078 533490 554084 533492
rect 501781 533488 554084 533490
rect 501781 533432 501786 533488
rect 501842 533432 554084 533488
rect 501781 533430 554084 533432
rect 501781 533427 501847 533430
rect 554078 533428 554084 533430
rect 554148 533428 554154 533492
rect 31518 533292 31524 533356
rect 31588 533354 31594 533356
rect 103973 533354 104039 533357
rect 31588 533352 104039 533354
rect 31588 533296 103978 533352
rect 104034 533296 104039 533352
rect 31588 533294 104039 533296
rect 31588 533292 31594 533294
rect 103973 533291 104039 533294
rect 499389 533354 499455 533357
rect 553894 533354 553900 533356
rect 499389 533352 553900 533354
rect 499389 533296 499394 533352
rect 499450 533296 553900 533352
rect 499389 533294 553900 533296
rect 499389 533291 499455 533294
rect 553894 533292 553900 533294
rect 553964 533292 553970 533356
rect 161105 533082 161171 533085
rect 435357 533082 435423 533085
rect 161105 533080 435423 533082
rect 161105 533024 161110 533080
rect 161166 533024 435362 533080
rect 435418 533024 435423 533080
rect 161105 533022 435423 533024
rect 161105 533019 161171 533022
rect 435357 533019 435423 533022
rect 157885 532946 157951 532949
rect 438945 532946 439011 532949
rect 157885 532944 439011 532946
rect 157885 532888 157890 532944
rect 157946 532888 438950 532944
rect 439006 532888 439011 532944
rect 157885 532886 439011 532888
rect 157885 532883 157951 532886
rect 438945 532883 439011 532886
rect 129825 532810 129891 532813
rect 466637 532810 466703 532813
rect 129825 532808 466703 532810
rect 129825 532752 129830 532808
rect 129886 532752 466642 532808
rect 466698 532752 466703 532808
rect 129825 532750 466703 532752
rect 129825 532747 129891 532750
rect 466637 532747 466703 532750
rect 26734 532612 26740 532676
rect 26804 532674 26810 532676
rect 92105 532674 92171 532677
rect 26804 532672 92171 532674
rect 26804 532616 92110 532672
rect 92166 532616 92171 532672
rect 26804 532614 92171 532616
rect 26804 532612 26810 532614
rect 92105 532611 92171 532614
rect 507117 532674 507183 532677
rect 550950 532674 550956 532676
rect 507117 532672 550956 532674
rect 507117 532616 507122 532672
rect 507178 532616 550956 532672
rect 507117 532614 550956 532616
rect 507117 532611 507183 532614
rect 550950 532612 550956 532614
rect 551020 532612 551026 532676
rect 27102 532476 27108 532540
rect 27172 532538 27178 532540
rect 94221 532538 94287 532541
rect 27172 532536 94287 532538
rect 27172 532480 94226 532536
rect 94282 532480 94287 532536
rect 27172 532478 94287 532480
rect 27172 532476 27178 532478
rect 94221 532475 94287 532478
rect 502885 532538 502951 532541
rect 550766 532538 550772 532540
rect 502885 532536 550772 532538
rect 502885 532480 502890 532536
rect 502946 532480 550772 532536
rect 502885 532478 550772 532480
rect 502885 532475 502951 532478
rect 550766 532476 550772 532478
rect 550836 532476 550842 532540
rect 26918 532340 26924 532404
rect 26988 532402 26994 532404
rect 96429 532402 96495 532405
rect 26988 532400 96495 532402
rect 26988 532344 96434 532400
rect 96490 532344 96495 532400
rect 26988 532342 96495 532344
rect 26988 532340 26994 532342
rect 96429 532339 96495 532342
rect 498561 532402 498627 532405
rect 552054 532402 552060 532404
rect 498561 532400 552060 532402
rect 498561 532344 498566 532400
rect 498622 532344 552060 532400
rect 498561 532342 552060 532344
rect 498561 532339 498627 532342
rect 552054 532340 552060 532342
rect 552124 532340 552130 532404
rect 29494 532204 29500 532268
rect 29564 532266 29570 532268
rect 98545 532266 98611 532269
rect 29564 532264 98611 532266
rect 29564 532208 98550 532264
rect 98606 532208 98611 532264
rect 29564 532206 98611 532208
rect 29564 532204 29570 532206
rect 98545 532203 98611 532206
rect 500677 532266 500743 532269
rect 553710 532266 553716 532268
rect 500677 532264 553716 532266
rect 500677 532208 500682 532264
rect 500738 532208 553716 532264
rect 500677 532206 553716 532208
rect 500677 532203 500743 532206
rect 553710 532204 553716 532206
rect 553780 532204 553786 532268
rect 27286 532068 27292 532132
rect 27356 532130 27362 532132
rect 99649 532130 99715 532133
rect 27356 532128 99715 532130
rect 27356 532072 99654 532128
rect 99710 532072 99715 532128
rect 27356 532070 99715 532072
rect 27356 532068 27362 532070
rect 99649 532067 99715 532070
rect 496353 532130 496419 532133
rect 550582 532130 550588 532132
rect 496353 532128 550588 532130
rect 496353 532072 496358 532128
rect 496414 532072 550588 532128
rect 496353 532070 550588 532072
rect 496353 532067 496419 532070
rect 550582 532068 550588 532070
rect 550652 532068 550658 532132
rect 27470 531932 27476 531996
rect 27540 531994 27546 531996
rect 100753 531994 100819 531997
rect 27540 531992 100819 531994
rect 27540 531936 100758 531992
rect 100814 531936 100819 531992
rect 27540 531934 100819 531936
rect 27540 531932 27546 531934
rect 100753 531931 100819 531934
rect 497457 531994 497523 531997
rect 553526 531994 553532 531996
rect 497457 531992 553532 531994
rect 497457 531936 497462 531992
rect 497518 531936 553532 531992
rect 497457 531934 553532 531936
rect 497457 531931 497523 531934
rect 553526 531932 553532 531934
rect 553596 531932 553602 531996
rect 29678 531796 29684 531860
rect 29748 531858 29754 531860
rect 83457 531858 83523 531861
rect 29748 531856 83523 531858
rect 29748 531800 83462 531856
rect 83518 531800 83523 531856
rect 29748 531798 83523 531800
rect 29748 531796 29754 531798
rect 83457 531795 83523 531798
rect 511441 531858 511507 531861
rect 552238 531858 552244 531860
rect 511441 531856 552244 531858
rect 511441 531800 511446 531856
rect 511502 531800 552244 531856
rect 511441 531798 552244 531800
rect 511441 531795 511507 531798
rect 552238 531796 552244 531798
rect 552308 531796 552314 531860
rect 29862 531660 29868 531724
rect 29932 531722 29938 531724
rect 74901 531722 74967 531725
rect 29932 531720 74967 531722
rect 29932 531664 74906 531720
rect 74962 531664 74967 531720
rect 29932 531662 74967 531664
rect 29932 531660 29938 531662
rect 74901 531659 74967 531662
rect 138473 531722 138539 531725
rect 458173 531722 458239 531725
rect 138473 531720 458239 531722
rect 138473 531664 138478 531720
rect 138534 531664 458178 531720
rect 458234 531664 458239 531720
rect 138473 531662 458239 531664
rect 138473 531659 138539 531662
rect 458173 531659 458239 531662
rect 515765 531722 515831 531725
rect 552422 531722 552428 531724
rect 515765 531720 552428 531722
rect 515765 531664 515770 531720
rect 515826 531664 552428 531720
rect 515765 531662 552428 531664
rect 515765 531659 515831 531662
rect 552422 531660 552428 531662
rect 552492 531660 552498 531724
rect 29177 531586 29243 531589
rect 29134 531584 29243 531586
rect 29134 531528 29182 531584
rect 29238 531528 29243 531584
rect 29134 531523 29243 531528
rect 135253 531586 135319 531589
rect 461209 531586 461275 531589
rect 135253 531584 461275 531586
rect 135253 531528 135258 531584
rect 135314 531528 461214 531584
rect 461270 531528 461275 531584
rect 135253 531526 461275 531528
rect 135253 531523 135319 531526
rect 461209 531523 461275 531526
rect 29134 531452 29194 531523
rect 29126 531388 29132 531452
rect 29196 531388 29202 531452
rect 111517 531450 111583 531453
rect 484945 531450 485011 531453
rect 111517 531448 485011 531450
rect 111517 531392 111522 531448
rect 111578 531392 484950 531448
rect 485006 531392 485011 531448
rect 111517 531390 485011 531392
rect 111517 531387 111583 531390
rect 484945 531387 485011 531390
rect 95182 531252 95188 531316
rect 95252 531314 95258 531316
rect 95325 531314 95391 531317
rect 95252 531312 95391 531314
rect 95252 531256 95330 531312
rect 95386 531256 95391 531312
rect 95252 531254 95391 531256
rect 95252 531252 95258 531254
rect 95325 531251 95391 531254
rect 104934 531252 104940 531316
rect 105004 531314 105010 531316
rect 105077 531314 105143 531317
rect 105004 531312 105143 531314
rect 105004 531256 105082 531312
rect 105138 531256 105143 531312
rect 105004 531254 105143 531256
rect 105004 531252 105010 531254
rect 105077 531251 105143 531254
rect 493041 531314 493107 531317
rect 493910 531314 493916 531316
rect 493041 531312 493916 531314
rect 493041 531256 493046 531312
rect 493102 531256 493916 531312
rect 493041 531254 493916 531256
rect 493041 531251 493107 531254
rect 493910 531252 493916 531254
rect 493980 531252 493986 531316
rect 492029 531178 492095 531181
rect 492438 531178 492444 531180
rect 492029 531176 492444 531178
rect 492029 531120 492034 531176
rect 492090 531120 492444 531176
rect 492029 531118 492444 531120
rect 492029 531115 492095 531118
rect 492438 531116 492444 531118
rect 492508 531116 492514 531180
rect 30230 530844 30236 530908
rect 30300 530906 30306 530908
rect 70577 530906 70643 530909
rect 30300 530904 70643 530906
rect 30300 530848 70582 530904
rect 70638 530848 70643 530904
rect 30300 530846 70643 530848
rect 30300 530844 30306 530846
rect 70577 530843 70643 530846
rect 524229 530906 524295 530909
rect 552606 530906 552612 530908
rect 524229 530904 552612 530906
rect 524229 530848 524234 530904
rect 524290 530848 552612 530904
rect 524229 530846 552612 530848
rect 524229 530843 524295 530846
rect 552606 530844 552612 530846
rect 552676 530844 552682 530908
rect 29126 530708 29132 530772
rect 29196 530770 29202 530772
rect 82445 530770 82511 530773
rect 29196 530768 82511 530770
rect 29196 530712 82450 530768
rect 82506 530712 82511 530768
rect 29196 530710 82511 530712
rect 29196 530708 29202 530710
rect 82445 530707 82511 530710
rect 509049 530770 509115 530773
rect 551318 530770 551324 530772
rect 509049 530768 551324 530770
rect 509049 530712 509054 530768
rect 509110 530712 551324 530768
rect 509049 530710 551324 530712
rect 509049 530707 509115 530710
rect 551318 530708 551324 530710
rect 551388 530708 551394 530772
rect 27654 530572 27660 530636
rect 27724 530634 27730 530636
rect 97533 530634 97599 530637
rect 27724 530632 97599 530634
rect 27724 530576 97538 530632
rect 97594 530576 97599 530632
rect 27724 530574 97599 530576
rect 27724 530572 27730 530574
rect 97533 530571 97599 530574
rect 495341 530634 495407 530637
rect 553342 530634 553348 530636
rect 495341 530632 553348 530634
rect 495341 530576 495346 530632
rect 495402 530576 553348 530632
rect 495341 530574 553348 530576
rect 495341 530571 495407 530574
rect 553342 530572 553348 530574
rect 553412 530572 553418 530636
rect 106089 529954 106155 529957
rect 490373 529954 490439 529957
rect 106089 529952 490439 529954
rect 106089 529896 106094 529952
rect 106150 529896 490378 529952
rect 490434 529896 490439 529952
rect 106089 529894 490439 529896
rect 106089 529891 106155 529894
rect 490373 529891 490439 529894
rect 493542 529892 493548 529956
rect 493612 529954 493618 529956
rect 493777 529954 493843 529957
rect 493612 529952 493843 529954
rect 493612 529896 493782 529952
rect 493838 529896 493843 529952
rect 493612 529894 493843 529896
rect 493612 529892 493618 529894
rect 493777 529891 493843 529894
rect 398833 529002 398899 529005
rect 399201 529002 399267 529005
rect 398833 529000 399267 529002
rect 398833 528944 398838 529000
rect 398894 528944 399206 529000
rect 399262 528944 399267 529000
rect 398833 528942 399267 528944
rect 398833 528939 398899 528942
rect 399201 528939 399267 528942
rect 385401 528866 385467 528869
rect 387333 528866 387399 528869
rect 385401 528864 387399 528866
rect 385401 528808 385406 528864
rect 385462 528808 387338 528864
rect 387394 528808 387399 528864
rect 385401 528806 387399 528808
rect 385401 528803 385467 528806
rect 387333 528803 387399 528806
rect 385677 528730 385743 528733
rect 386229 528730 386295 528733
rect 385677 528728 386295 528730
rect 385677 528672 385682 528728
rect 385738 528672 386234 528728
rect 386290 528672 386295 528728
rect 385677 528670 386295 528672
rect 385677 528667 385743 528670
rect 386229 528667 386295 528670
rect 385953 528594 386019 528597
rect 386505 528594 386571 528597
rect 385953 528592 386571 528594
rect 385953 528536 385958 528592
rect 386014 528536 386510 528592
rect 386566 528536 386571 528592
rect 385953 528534 386571 528536
rect 385953 528531 386019 528534
rect 386505 528531 386571 528534
rect 398833 528594 398899 528597
rect 403709 528594 403775 528597
rect 398833 528592 403775 528594
rect 398833 528536 398838 528592
rect 398894 528536 403714 528592
rect 403770 528536 403775 528592
rect 398833 528534 403775 528536
rect 398833 528531 398899 528534
rect 403709 528531 403775 528534
rect 182173 528458 182239 528461
rect 183921 528458 183987 528461
rect 182173 528456 183987 528458
rect 182173 528400 182178 528456
rect 182234 528400 183926 528456
rect 183982 528400 183987 528456
rect 182173 528398 183987 528400
rect 182173 528395 182239 528398
rect 183921 528395 183987 528398
rect 251817 528458 251883 528461
rect 253841 528458 253907 528461
rect 251817 528456 253907 528458
rect 251817 528400 251822 528456
rect 251878 528400 253846 528456
rect 253902 528400 253907 528456
rect 251817 528398 253907 528400
rect 251817 528395 251883 528398
rect 253841 528395 253907 528398
rect 315297 528458 315363 528461
rect 320081 528458 320147 528461
rect 315297 528456 320147 528458
rect 315297 528400 315302 528456
rect 315358 528400 320086 528456
rect 320142 528400 320147 528456
rect 315297 528398 320147 528400
rect 315297 528395 315363 528398
rect 320081 528395 320147 528398
rect 385861 528458 385927 528461
rect 386413 528458 386479 528461
rect 385861 528456 386479 528458
rect 385861 528400 385866 528456
rect 385922 528400 386418 528456
rect 386474 528400 386479 528456
rect 385861 528398 386479 528400
rect 385861 528395 385927 528398
rect 386413 528395 386479 528398
rect 422293 528458 422359 528461
rect 431769 528458 431835 528461
rect 422293 528456 431835 528458
rect 422293 528400 422298 528456
rect 422354 528400 431774 528456
rect 431830 528400 431835 528456
rect 422293 528398 431835 528400
rect 422293 528395 422359 528398
rect 431769 528395 431835 528398
rect 175917 528322 175983 528325
rect 177941 528322 178007 528325
rect 175917 528320 176026 528322
rect 175917 528264 175922 528320
rect 175978 528264 176026 528320
rect 175917 528259 176026 528264
rect 175966 528186 176026 528259
rect 177806 528320 178007 528322
rect 177806 528264 177946 528320
rect 178002 528264 178007 528320
rect 177806 528262 178007 528264
rect 177806 528186 177866 528262
rect 177941 528259 178007 528262
rect 181897 528322 181963 528325
rect 185945 528322 186011 528325
rect 207565 528322 207631 528325
rect 181897 528320 186011 528322
rect 181897 528264 181902 528320
rect 181958 528264 185950 528320
rect 186006 528264 186011 528320
rect 181897 528262 186011 528264
rect 181897 528259 181963 528262
rect 185945 528259 186011 528262
rect 207062 528320 207631 528322
rect 207062 528264 207570 528320
rect 207626 528264 207631 528320
rect 207062 528262 207631 528264
rect 207062 528223 207122 528262
rect 207565 528259 207631 528262
rect 251817 528322 251883 528325
rect 254301 528322 254367 528325
rect 251817 528320 254367 528322
rect 251817 528264 251822 528320
rect 251878 528264 254306 528320
rect 254362 528264 254367 528320
rect 251817 528262 254367 528264
rect 251817 528259 251883 528262
rect 254301 528259 254367 528262
rect 315205 528322 315271 528325
rect 324221 528322 324287 528325
rect 315205 528320 324287 528322
rect 315205 528264 315210 528320
rect 315266 528264 324226 528320
rect 324282 528264 324287 528320
rect 315205 528262 324287 528264
rect 315205 528259 315271 528262
rect 324221 528259 324287 528262
rect 385769 528322 385835 528325
rect 386321 528322 386387 528325
rect 385769 528320 386387 528322
rect 385769 528264 385774 528320
rect 385830 528264 386326 528320
rect 386382 528264 386387 528320
rect 385769 528262 386387 528264
rect 385769 528259 385835 528262
rect 386321 528259 386387 528262
rect 408217 528322 408283 528325
rect 422201 528322 422267 528325
rect 508497 528322 508563 528325
rect 408217 528320 422267 528322
rect 408217 528264 408222 528320
rect 408278 528264 422206 528320
rect 422262 528264 422267 528320
rect 408217 528262 422267 528264
rect 408217 528259 408283 528262
rect 422201 528259 422267 528262
rect 508454 528320 508563 528322
rect 508454 528264 508502 528320
rect 508558 528264 508563 528320
rect 508454 528259 508563 528264
rect 175966 528126 177866 528186
rect 207013 528218 207122 528223
rect 207013 528162 207018 528218
rect 207074 528162 207122 528218
rect 207013 528160 207122 528162
rect 207013 528157 207079 528160
rect 508454 527778 508514 528259
rect 574870 527778 574876 527780
rect 508454 527718 574876 527778
rect 574870 527716 574876 527718
rect 574940 527716 574946 527780
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 281533 515946 281599 515949
rect 279036 515944 281599 515946
rect 279036 515888 281538 515944
rect 281594 515888 281599 515944
rect 279036 515886 281599 515888
rect 281533 515883 281599 515886
rect 315941 515810 316007 515813
rect 315941 515808 317676 515810
rect 315941 515752 315946 515808
rect 316002 515752 317676 515808
rect 315941 515750 317676 515752
rect 315941 515747 316007 515750
rect 282913 512002 282979 512005
rect 283097 512002 283163 512005
rect 282913 512000 283163 512002
rect 282913 511944 282918 512000
rect 282974 511944 283102 512000
rect 283158 511944 283163 512000
rect 282913 511942 283163 511944
rect 282913 511939 282979 511942
rect 283097 511939 283163 511942
rect 580533 510370 580599 510373
rect 583520 510370 584960 510460
rect 580533 510368 584960 510370
rect 580533 510312 580538 510368
rect 580594 510312 584960 510368
rect 580533 510310 584960 510312
rect 580533 510307 580599 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 2865 509962 2931 509965
rect -960 509960 2931 509962
rect -960 509904 2870 509960
rect 2926 509904 2931 509960
rect -960 509902 2931 509904
rect -960 509812 480 509902
rect 2865 509899 2931 509902
rect 573449 502754 573515 502757
rect 574870 502754 574876 502756
rect 573449 502752 574876 502754
rect 573449 502696 573454 502752
rect 573510 502696 574876 502752
rect 573449 502694 574876 502696
rect 573449 502691 573515 502694
rect 574870 502692 574876 502694
rect 574940 502692 574946 502756
rect 154297 502346 154363 502349
rect 154254 502344 154363 502346
rect 154254 502288 154302 502344
rect 154358 502288 154363 502344
rect 154254 502283 154363 502288
rect 154254 502210 154314 502283
rect 154389 502210 154455 502213
rect 154254 502208 154455 502210
rect 154254 502152 154394 502208
rect 154450 502152 154455 502208
rect 154254 502150 154455 502152
rect 154389 502147 154455 502150
rect 130694 500788 130700 500852
rect 130764 500850 130770 500852
rect 130929 500850 130995 500853
rect 130764 500848 130995 500850
rect 130764 500792 130934 500848
rect 130990 500792 130995 500848
rect 130764 500790 130995 500792
rect 130764 500788 130770 500790
rect 130929 500787 130995 500790
rect 141693 500850 141759 500853
rect 153561 500850 153627 500853
rect 141693 500848 153627 500850
rect 141693 500792 141698 500848
rect 141754 500792 153566 500848
rect 153622 500792 153627 500848
rect 141693 500790 153627 500792
rect 141693 500787 141759 500790
rect 153561 500787 153627 500790
rect 189574 500788 189580 500852
rect 189644 500850 189650 500852
rect 190177 500850 190243 500853
rect 189644 500848 190243 500850
rect 189644 500792 190182 500848
rect 190238 500792 190243 500848
rect 189644 500790 190243 500792
rect 189644 500788 189650 500790
rect 190177 500787 190243 500790
rect 191046 500788 191052 500852
rect 191116 500850 191122 500852
rect 191281 500850 191347 500853
rect 191116 500848 191347 500850
rect 191116 500792 191286 500848
rect 191342 500792 191347 500848
rect 191116 500790 191347 500792
rect 191116 500788 191122 500790
rect 191281 500787 191347 500790
rect 491845 500852 491911 500853
rect 493133 500852 493199 500853
rect 491845 500848 491892 500852
rect 491956 500850 491962 500852
rect 491845 500792 491850 500848
rect 491845 500788 491892 500792
rect 491956 500790 492002 500850
rect 493133 500848 493180 500852
rect 493244 500850 493250 500852
rect 508221 500850 508287 500853
rect 517973 500852 518039 500853
rect 508446 500850 508452 500852
rect 493133 500792 493138 500848
rect 491956 500788 491962 500790
rect 493133 500788 493180 500792
rect 493244 500790 493290 500850
rect 508221 500848 508452 500850
rect 508221 500792 508226 500848
rect 508282 500792 508452 500848
rect 508221 500790 508452 500792
rect 493244 500788 493250 500790
rect 491845 500787 491911 500788
rect 493133 500787 493199 500788
rect 508221 500787 508287 500790
rect 508446 500788 508452 500790
rect 508516 500788 508522 500852
rect 517973 500848 518020 500852
rect 518084 500850 518090 500852
rect 542629 500850 542695 500853
rect 542854 500850 542860 500852
rect 517973 500792 517978 500848
rect 517973 500788 518020 500792
rect 518084 500790 518130 500850
rect 542629 500848 542860 500850
rect 542629 500792 542634 500848
rect 542690 500792 542860 500848
rect 542629 500790 542860 500792
rect 518084 500788 518090 500790
rect 517973 500787 518039 500788
rect 542629 500787 542695 500790
rect 542854 500788 542860 500790
rect 542924 500788 542930 500852
rect 550081 500850 550147 500853
rect 550214 500850 550220 500852
rect 550081 500848 550220 500850
rect 550081 500792 550086 500848
rect 550142 500792 550220 500848
rect 550081 500790 550220 500792
rect 550081 500787 550147 500790
rect 550214 500788 550220 500790
rect 550284 500788 550290 500852
rect 114737 500714 114803 500717
rect 142705 500714 142771 500717
rect 114737 500712 142771 500714
rect 114737 500656 114742 500712
rect 114798 500656 142710 500712
rect 142766 500656 142771 500712
rect 114737 500654 142771 500656
rect 114737 500651 114803 500654
rect 142705 500651 142771 500654
rect 189073 500714 189139 500717
rect 189758 500714 189764 500716
rect 189073 500712 189764 500714
rect 189073 500656 189078 500712
rect 189134 500656 189764 500712
rect 189073 500654 189764 500656
rect 189073 500651 189139 500654
rect 189758 500652 189764 500654
rect 189828 500652 189834 500716
rect 116853 500578 116919 500581
rect 149094 500578 149100 500580
rect 116853 500576 149100 500578
rect 116853 500520 116858 500576
rect 116914 500520 149100 500576
rect 116853 500518 149100 500520
rect 116853 500515 116919 500518
rect 149094 500516 149100 500518
rect 149164 500516 149170 500580
rect 107193 500442 107259 500445
rect 117957 500442 118023 500445
rect 151854 500442 151860 500444
rect 107193 500440 113098 500442
rect 107193 500384 107198 500440
rect 107254 500384 113098 500440
rect 107193 500382 113098 500384
rect 107193 500379 107259 500382
rect 112621 500170 112687 500173
rect 112846 500170 112852 500172
rect 112621 500168 112852 500170
rect 112621 500112 112626 500168
rect 112682 500112 112852 500168
rect 112621 500110 112852 500112
rect 112621 500107 112687 500110
rect 112846 500108 112852 500110
rect 112916 500108 112922 500172
rect 113038 500170 113098 500382
rect 117957 500440 151860 500442
rect 117957 500384 117962 500440
rect 118018 500384 151860 500440
rect 117957 500382 151860 500384
rect 117957 500379 118023 500382
rect 151854 500380 151860 500382
rect 151924 500380 151930 500444
rect 113633 500306 113699 500309
rect 147806 500306 147812 500308
rect 113633 500304 147812 500306
rect 113633 500248 113638 500304
rect 113694 500248 147812 500304
rect 113633 500246 147812 500248
rect 113633 500243 113699 500246
rect 147806 500244 147812 500246
rect 147876 500244 147882 500308
rect 147990 500170 147996 500172
rect 113038 500110 147996 500170
rect 147990 500108 147996 500110
rect 148060 500108 148066 500172
rect 142705 499898 142771 499901
rect 147622 499898 147628 499900
rect 142705 499896 147628 499898
rect 142705 499840 142710 499896
rect 142766 499840 147628 499896
rect 142705 499838 147628 499840
rect 142705 499835 142771 499838
rect 147622 499836 147628 499838
rect 147692 499836 147698 499900
rect 143809 499762 143875 499765
rect 155401 499762 155467 499765
rect 143809 499760 155467 499762
rect 143809 499704 143814 499760
rect 143870 499704 155406 499760
rect 155462 499704 155467 499760
rect 143809 499702 155467 499704
rect 143809 499699 143875 499702
rect 155401 499699 155467 499702
rect 147029 499628 147095 499629
rect 148133 499628 148199 499629
rect 147029 499624 147076 499628
rect 147140 499626 147146 499628
rect 147029 499568 147034 499624
rect 147029 499564 147076 499568
rect 147140 499566 147186 499626
rect 148133 499624 148180 499628
rect 148244 499626 148250 499628
rect 149237 499626 149303 499629
rect 149646 499626 149652 499628
rect 148133 499568 148138 499624
rect 147140 499564 147146 499566
rect 148133 499564 148180 499568
rect 148244 499566 148290 499626
rect 149237 499624 149652 499626
rect 149237 499568 149242 499624
rect 149298 499568 149652 499624
rect 149237 499566 149652 499568
rect 148244 499564 148250 499566
rect 147029 499563 147095 499564
rect 148133 499563 148199 499564
rect 149237 499563 149303 499566
rect 149646 499564 149652 499566
rect 149716 499564 149722 499628
rect 149830 499564 149836 499628
rect 149900 499626 149906 499628
rect 150341 499626 150407 499629
rect 149900 499624 150407 499626
rect 149900 499568 150346 499624
rect 150402 499568 150407 499624
rect 149900 499566 150407 499568
rect 149900 499564 149906 499566
rect 150341 499563 150407 499566
rect 150934 499564 150940 499628
rect 151004 499626 151010 499628
rect 151353 499626 151419 499629
rect 152457 499628 152523 499629
rect 152406 499626 152412 499628
rect 151004 499624 151419 499626
rect 151004 499568 151358 499624
rect 151414 499568 151419 499624
rect 151004 499566 151419 499568
rect 152366 499566 152412 499626
rect 152476 499624 152523 499628
rect 152518 499568 152523 499624
rect 151004 499564 151010 499566
rect 151353 499563 151419 499566
rect 152406 499564 152412 499566
rect 152476 499564 152523 499568
rect 152457 499563 152523 499564
rect 580901 498674 580967 498677
rect 583520 498674 584960 498764
rect 580901 498672 584960 498674
rect 580901 498616 580906 498672
rect 580962 498616 584960 498672
rect 580901 498614 584960 498616
rect 580901 498611 580967 498614
rect 583520 498524 584960 498614
rect 124213 498130 124279 498133
rect 154798 498130 154804 498132
rect 124213 498128 154804 498130
rect 124213 498072 124218 498128
rect 124274 498072 154804 498128
rect 124213 498070 154804 498072
rect 124213 498067 124279 498070
rect 154798 498068 154804 498070
rect 154868 498068 154874 498132
rect 114553 497994 114619 497997
rect 149278 497994 149284 497996
rect 114553 497992 149284 497994
rect 114553 497936 114558 497992
rect 114614 497936 149284 497992
rect 114553 497934 149284 497936
rect 114553 497931 114619 497934
rect 149278 497932 149284 497934
rect 149348 497932 149354 497996
rect 110597 497858 110663 497861
rect 150382 497858 150388 497860
rect 110597 497856 150388 497858
rect 110597 497800 110602 497856
rect 110658 497800 150388 497856
rect 110597 497798 150388 497800
rect 110597 497795 110663 497798
rect 150382 497796 150388 497798
rect 150452 497796 150458 497860
rect 110413 497722 110479 497725
rect 150750 497722 150756 497724
rect 110413 497720 150756 497722
rect 110413 497664 110418 497720
rect 110474 497664 150756 497720
rect 110413 497662 150756 497664
rect 110413 497659 110479 497662
rect 150750 497660 150756 497662
rect 150820 497660 150826 497724
rect 153193 497722 153259 497725
rect 153694 497722 153700 497724
rect 153193 497720 153700 497722
rect 153193 497664 153198 497720
rect 153254 497664 153700 497720
rect 153193 497662 153700 497664
rect 153193 497659 153259 497662
rect 153694 497660 153700 497662
rect 153764 497660 153770 497724
rect 107653 497586 107719 497589
rect 148358 497586 148364 497588
rect 107653 497584 148364 497586
rect 107653 497528 107658 497584
rect 107714 497528 148364 497584
rect 107653 497526 148364 497528
rect 107653 497523 107719 497526
rect 148358 497524 148364 497526
rect 148428 497524 148434 497588
rect 109033 497450 109099 497453
rect 150566 497450 150572 497452
rect 109033 497448 150572 497450
rect 109033 497392 109038 497448
rect 109094 497392 150572 497448
rect 109033 497390 150572 497392
rect 109033 497387 109099 497390
rect 150566 497388 150572 497390
rect 150636 497388 150642 497452
rect 125593 497314 125659 497317
rect 153142 497314 153148 497316
rect 125593 497312 153148 497314
rect 125593 497256 125598 497312
rect 125654 497256 153148 497312
rect 125593 497254 153148 497256
rect 125593 497251 125659 497254
rect 153142 497252 153148 497254
rect 153212 497252 153218 497316
rect 128353 497178 128419 497181
rect 154614 497178 154620 497180
rect 128353 497176 154620 497178
rect 128353 497120 128358 497176
rect 128414 497120 154620 497176
rect 128353 497118 154620 497120
rect 128353 497115 128419 497118
rect 154614 497116 154620 497118
rect 154684 497116 154690 497180
rect -960 495546 480 495636
rect 3509 495546 3575 495549
rect -960 495544 3575 495546
rect -960 495488 3514 495544
rect 3570 495488 3575 495544
rect -960 495486 3575 495488
rect -960 495396 480 495486
rect 3509 495483 3575 495486
rect 146845 492690 146911 492693
rect 154205 492690 154271 492693
rect 146845 492688 154271 492690
rect 146845 492632 146850 492688
rect 146906 492632 154210 492688
rect 154266 492632 154271 492688
rect 146845 492630 154271 492632
rect 146845 492627 146911 492630
rect 154205 492627 154271 492630
rect 496721 487794 496787 487797
rect 550582 487794 550588 487796
rect 496721 487792 550588 487794
rect 496721 487736 496726 487792
rect 496782 487736 550588 487792
rect 496721 487734 550588 487736
rect 496721 487731 496787 487734
rect 550582 487732 550588 487734
rect 550652 487732 550658 487796
rect 583520 486692 584960 486932
rect 147438 485890 147444 485892
rect 147262 485830 147444 485890
rect 147262 485620 147322 485830
rect 147438 485828 147444 485830
rect 147508 485828 147514 485892
rect 147254 485556 147260 485620
rect 147324 485556 147330 485620
rect 155861 483034 155927 483037
rect 156137 483034 156203 483037
rect 155861 483032 156203 483034
rect 155861 482976 155866 483032
rect 155922 482976 156142 483032
rect 156198 482976 156203 483032
rect 155861 482974 156203 482976
rect 155861 482971 155927 482974
rect 156137 482971 156203 482974
rect -960 481130 480 481220
rect 3141 481130 3207 481133
rect -960 481128 3207 481130
rect -960 481072 3146 481128
rect 3202 481072 3207 481128
rect -960 481070 3207 481072
rect -960 480980 480 481070
rect 3141 481067 3207 481070
rect 506381 477186 506447 477189
rect 552238 477186 552244 477188
rect 506381 477184 552244 477186
rect 506381 477128 506386 477184
rect 506442 477128 552244 477184
rect 506381 477126 552244 477128
rect 506381 477123 506447 477126
rect 552238 477124 552244 477126
rect 552308 477124 552314 477188
rect 503529 477050 503595 477053
rect 552790 477050 552796 477052
rect 503529 477048 552796 477050
rect 503529 476992 503534 477048
rect 503590 476992 552796 477048
rect 503529 476990 552796 476992
rect 503529 476987 503595 476990
rect 552790 476988 552796 476990
rect 552860 476988 552866 477052
rect 502241 476914 502307 476917
rect 552606 476914 552612 476916
rect 502241 476912 552612 476914
rect 502241 476856 502246 476912
rect 502302 476856 552612 476912
rect 502241 476854 552612 476856
rect 502241 476851 502307 476854
rect 552606 476852 552612 476854
rect 552676 476852 552682 476916
rect 499389 476778 499455 476781
rect 552422 476778 552428 476780
rect 499389 476776 552428 476778
rect 499389 476720 499394 476776
rect 499450 476720 552428 476776
rect 499389 476718 552428 476720
rect 499389 476715 499455 476718
rect 552422 476716 552428 476718
rect 552492 476716 552498 476780
rect 542905 476236 542971 476237
rect 542854 476234 542860 476236
rect 542814 476174 542860 476234
rect 542924 476232 542971 476236
rect 542966 476176 542971 476232
rect 542854 476172 542860 476174
rect 542924 476172 542971 476176
rect 542905 476171 542971 476172
rect 508497 476100 508563 476101
rect 508446 476098 508452 476100
rect 508406 476038 508452 476098
rect 508516 476096 508563 476100
rect 508558 476040 508563 476096
rect 508446 476036 508452 476038
rect 508516 476036 508563 476040
rect 508497 476035 508563 476036
rect 509141 476098 509207 476101
rect 551134 476098 551140 476100
rect 509141 476096 551140 476098
rect 509141 476040 509146 476096
rect 509202 476040 551140 476096
rect 509141 476038 551140 476040
rect 509141 476035 509207 476038
rect 551134 476036 551140 476038
rect 551204 476036 551210 476100
rect 507761 475962 507827 475965
rect 551686 475962 551692 475964
rect 507761 475960 551692 475962
rect 507761 475904 507766 475960
rect 507822 475904 551692 475960
rect 507761 475902 551692 475904
rect 507761 475899 507827 475902
rect 551686 475900 551692 475902
rect 551756 475900 551762 475964
rect 503621 475826 503687 475829
rect 554998 475826 555004 475828
rect 503621 475824 555004 475826
rect 503621 475768 503626 475824
rect 503682 475768 555004 475824
rect 503621 475766 555004 475768
rect 503621 475763 503687 475766
rect 554998 475764 555004 475766
rect 555068 475764 555074 475828
rect 500861 475690 500927 475693
rect 553342 475690 553348 475692
rect 500861 475688 553348 475690
rect 500861 475632 500866 475688
rect 500922 475632 553348 475688
rect 500861 475630 553348 475632
rect 500861 475627 500927 475630
rect 553342 475628 553348 475630
rect 553412 475628 553418 475692
rect 493961 475554 494027 475557
rect 552473 475554 552539 475557
rect 493961 475552 552539 475554
rect 493961 475496 493966 475552
rect 494022 475496 552478 475552
rect 552534 475496 552539 475552
rect 493961 475494 552539 475496
rect 493961 475491 494027 475494
rect 552473 475491 552539 475494
rect 495341 475418 495407 475421
rect 552054 475418 552060 475420
rect 495341 475416 552060 475418
rect 495341 475360 495346 475416
rect 495402 475360 552060 475416
rect 495341 475358 552060 475360
rect 495341 475355 495407 475358
rect 552054 475356 552060 475358
rect 552124 475356 552130 475420
rect 583520 474996 584960 475236
rect 550582 474540 550588 474604
rect 550652 474602 550658 474604
rect 552289 474602 552355 474605
rect 550652 474600 552355 474602
rect 550652 474544 552294 474600
rect 552350 474544 552355 474600
rect 550652 474542 552355 474544
rect 550652 474540 550658 474542
rect 552289 474539 552355 474542
rect 520181 474330 520247 474333
rect 553526 474330 553532 474332
rect 520181 474328 553532 474330
rect 520181 474272 520186 474328
rect 520242 474272 553532 474328
rect 520181 474270 553532 474272
rect 520181 474267 520247 474270
rect 553526 474268 553532 474270
rect 553596 474268 553602 474332
rect 513281 474194 513347 474197
rect 553710 474194 553716 474196
rect 513281 474192 553716 474194
rect 513281 474136 513286 474192
rect 513342 474136 553716 474192
rect 513281 474134 553716 474136
rect 513281 474131 513347 474134
rect 553710 474132 553716 474134
rect 553780 474132 553786 474196
rect 505001 474058 505067 474061
rect 505001 474056 550098 474058
rect 505001 474000 505006 474056
rect 505062 474000 550098 474056
rect 505001 473998 550098 474000
rect 505001 473995 505067 473998
rect 299422 473860 299428 473924
rect 299492 473922 299498 473924
rect 309041 473922 309107 473925
rect 299492 473920 309107 473922
rect 299492 473864 309046 473920
rect 309102 473864 309107 473920
rect 299492 473862 309107 473864
rect 299492 473860 299498 473862
rect 309041 473859 309107 473862
rect 318742 473860 318748 473924
rect 318812 473922 318818 473924
rect 328310 473922 328316 473924
rect 318812 473862 328316 473922
rect 318812 473860 318818 473862
rect 328310 473860 328316 473862
rect 328380 473860 328386 473924
rect 338062 473860 338068 473924
rect 338132 473922 338138 473924
rect 347630 473922 347636 473924
rect 338132 473862 347636 473922
rect 338132 473860 338138 473862
rect 347630 473860 347636 473862
rect 347700 473860 347706 473924
rect 357382 473860 357388 473924
rect 357452 473922 357458 473924
rect 366950 473922 366956 473924
rect 357452 473862 366956 473922
rect 357452 473860 357458 473862
rect 366950 473860 366956 473862
rect 367020 473860 367026 473924
rect 384982 473860 384988 473924
rect 385052 473922 385058 473924
rect 389817 473922 389883 473925
rect 385052 473920 389883 473922
rect 385052 473864 389822 473920
rect 389878 473864 389883 473920
rect 385052 473862 389883 473864
rect 385052 473860 385058 473862
rect 389817 473859 389883 473862
rect 518014 473860 518020 473924
rect 518084 473922 518090 473924
rect 520733 473922 520799 473925
rect 518084 473920 520799 473922
rect 518084 473864 520738 473920
rect 520794 473864 520799 473920
rect 518084 473862 520799 473864
rect 550038 473922 550098 473998
rect 550214 473996 550220 474060
rect 550284 474058 550290 474060
rect 554078 474058 554084 474060
rect 550284 473998 554084 474058
rect 550284 473996 550290 473998
rect 554078 473996 554084 473998
rect 554148 473996 554154 474060
rect 555366 473922 555372 473924
rect 550038 473862 555372 473922
rect 518084 473860 518090 473862
rect 520733 473859 520799 473862
rect 555366 473860 555372 473862
rect 555436 473860 555442 473924
rect 280654 473724 280660 473788
rect 280724 473786 280730 473788
rect 408585 473786 408651 473789
rect 418153 473786 418219 473789
rect 280724 473726 289738 473786
rect 280724 473724 280730 473726
rect 289678 473378 289738 473726
rect 408585 473784 415410 473786
rect 408585 473728 408590 473784
rect 408646 473728 415410 473784
rect 408585 473726 415410 473728
rect 408585 473723 408651 473726
rect 299422 473650 299428 473652
rect 292622 473590 299428 473650
rect 292622 473378 292682 473590
rect 299422 473588 299428 473590
rect 299492 473588 299498 473652
rect 328310 473588 328316 473652
rect 328380 473650 328386 473652
rect 328380 473590 328562 473650
rect 328380 473588 328386 473590
rect 318742 473514 318748 473516
rect 311942 473454 318748 473514
rect 289678 473318 292682 473378
rect 309041 473378 309107 473381
rect 311942 473378 312002 473454
rect 318742 473452 318748 473454
rect 318812 473452 318818 473516
rect 328502 473514 328562 473590
rect 347630 473588 347636 473652
rect 347700 473650 347706 473652
rect 347700 473590 347882 473650
rect 347700 473588 347706 473590
rect 331070 473514 331076 473516
rect 328502 473454 331076 473514
rect 331070 473452 331076 473454
rect 331140 473452 331146 473516
rect 331254 473452 331260 473516
rect 331324 473514 331330 473516
rect 338062 473514 338068 473516
rect 331324 473454 338068 473514
rect 331324 473452 331330 473454
rect 338062 473452 338068 473454
rect 338132 473452 338138 473516
rect 347822 473514 347882 473590
rect 366950 473588 366956 473652
rect 367020 473650 367026 473652
rect 384982 473650 384988 473652
rect 367020 473590 367202 473650
rect 367020 473588 367026 473590
rect 350390 473514 350396 473516
rect 347822 473454 350396 473514
rect 350390 473452 350396 473454
rect 350460 473452 350466 473516
rect 350574 473452 350580 473516
rect 350644 473514 350650 473516
rect 357382 473514 357388 473516
rect 350644 473454 357388 473514
rect 350644 473452 350650 473454
rect 357382 473452 357388 473454
rect 357452 473452 357458 473516
rect 367142 473514 367202 473590
rect 381494 473590 384988 473650
rect 369710 473514 369716 473516
rect 367142 473454 369716 473514
rect 369710 473452 369716 473454
rect 369780 473452 369786 473516
rect 369894 473452 369900 473516
rect 369964 473514 369970 473516
rect 381494 473514 381554 473590
rect 384982 473588 384988 473590
rect 385052 473588 385058 473652
rect 389817 473650 389883 473653
rect 408401 473650 408467 473653
rect 389817 473648 394618 473650
rect 389817 473592 389822 473648
rect 389878 473592 394618 473648
rect 389817 473590 394618 473592
rect 389817 473587 389883 473590
rect 369964 473454 381554 473514
rect 394558 473514 394618 473590
rect 400814 473648 408467 473650
rect 400814 473592 408406 473648
rect 408462 473592 408467 473648
rect 400814 473590 408467 473592
rect 415350 473650 415410 473726
rect 418153 473784 424978 473786
rect 418153 473728 418158 473784
rect 418214 473728 424978 473784
rect 418153 473726 424978 473728
rect 418153 473723 418219 473726
rect 418061 473650 418127 473653
rect 415350 473648 418127 473650
rect 415350 473592 418066 473648
rect 418122 473592 418127 473648
rect 415350 473590 418127 473592
rect 424918 473650 424978 473726
rect 434662 473724 434668 473788
rect 434732 473786 434738 473788
rect 437381 473786 437447 473789
rect 434732 473784 437447 473786
rect 434732 473728 437386 473784
rect 437442 473728 437447 473784
rect 434732 473726 437447 473728
rect 434732 473724 434738 473726
rect 437381 473723 437447 473726
rect 437565 473786 437631 473789
rect 481633 473786 481699 473789
rect 437565 473784 447058 473786
rect 437565 473728 437570 473784
rect 437626 473728 447058 473784
rect 437565 473726 447058 473728
rect 437565 473723 437631 473726
rect 425094 473650 425100 473652
rect 424918 473590 425100 473650
rect 400814 473514 400874 473590
rect 408401 473587 408467 473590
rect 418061 473587 418127 473590
rect 425094 473588 425100 473590
rect 425164 473588 425170 473652
rect 394558 473454 400874 473514
rect 446998 473514 447058 473726
rect 456750 473726 466378 473786
rect 456750 473514 456810 473726
rect 446998 473454 456810 473514
rect 466318 473514 466378 473726
rect 476070 473784 481699 473786
rect 476070 473728 481638 473784
rect 481694 473728 481699 473784
rect 476070 473726 481699 473728
rect 476070 473514 476130 473726
rect 481633 473723 481699 473726
rect 512637 473786 512703 473789
rect 517462 473786 517468 473788
rect 512637 473784 517468 473786
rect 512637 473728 512642 473784
rect 512698 473728 517468 473784
rect 512637 473726 517468 473728
rect 512637 473723 512703 473726
rect 517462 473724 517468 473726
rect 517532 473724 517538 473788
rect 536782 473786 536788 473788
rect 531822 473726 536788 473786
rect 490649 473650 490715 473653
rect 505001 473650 505067 473653
rect 490649 473648 505067 473650
rect 490649 473592 490654 473648
rect 490710 473592 505006 473648
rect 505062 473592 505067 473648
rect 490649 473590 505067 473592
rect 490649 473587 490715 473590
rect 505001 473587 505067 473590
rect 466318 473454 476130 473514
rect 491845 473516 491911 473517
rect 493133 473516 493199 473517
rect 491845 473512 491892 473516
rect 491956 473514 491962 473516
rect 491845 473456 491850 473512
rect 369964 473452 369970 473454
rect 491845 473452 491892 473456
rect 491956 473454 492002 473514
rect 493133 473512 493180 473516
rect 493244 473514 493250 473516
rect 493133 473456 493138 473512
rect 491956 473452 491962 473454
rect 493133 473452 493180 473456
rect 493244 473454 493290 473514
rect 493244 473452 493250 473454
rect 517462 473452 517468 473516
rect 517532 473514 517538 473516
rect 531822 473514 531882 473726
rect 536782 473724 536788 473726
rect 536852 473724 536858 473788
rect 536966 473588 536972 473652
rect 537036 473650 537042 473652
rect 537036 473590 552122 473650
rect 537036 473588 537042 473590
rect 517532 473454 531882 473514
rect 517532 473452 517538 473454
rect 491845 473451 491911 473452
rect 493133 473451 493199 473452
rect 309041 473376 312002 473378
rect 309041 473320 309046 473376
rect 309102 473320 312002 473376
rect 309041 473318 312002 473320
rect 309041 473315 309107 473318
rect 425094 473316 425100 473380
rect 425164 473378 425170 473380
rect 427721 473378 427787 473381
rect 425164 473376 427787 473378
rect 425164 473320 427726 473376
rect 427782 473320 427787 473376
rect 425164 473318 427787 473320
rect 425164 473316 425170 473318
rect 427721 473315 427787 473318
rect 427905 473378 427971 473381
rect 434662 473378 434668 473380
rect 427905 473376 434668 473378
rect 427905 473320 427910 473376
rect 427966 473320 434668 473376
rect 427905 473318 434668 473320
rect 427905 473315 427971 473318
rect 434662 473316 434668 473318
rect 434732 473316 434738 473380
rect 552062 473348 552122 473590
rect 552062 472565 552122 472804
rect 553025 472698 553091 472701
rect 554814 472698 554820 472700
rect 553025 472696 554820 472698
rect 553025 472640 553030 472696
rect 553086 472640 554820 472696
rect 553025 472638 554820 472640
rect 553025 472635 553091 472638
rect 554814 472636 554820 472638
rect 554884 472636 554890 472700
rect 552062 472560 552171 472565
rect 552062 472504 552110 472560
rect 552166 472504 552171 472560
rect 552062 472502 552171 472504
rect 552105 472499 552171 472502
rect 552197 472426 552263 472429
rect 552197 472424 552306 472426
rect 552197 472368 552202 472424
rect 552258 472368 552306 472424
rect 552197 472363 552306 472368
rect 552246 472124 552306 472363
rect 552473 471882 552539 471885
rect 552430 471880 552539 471882
rect 552430 471824 552478 471880
rect 552534 471824 552539 471880
rect 552430 471819 552539 471824
rect 552430 471580 552490 471819
rect 280153 471338 280219 471341
rect 279956 471336 280219 471338
rect 279956 471280 280158 471336
rect 280214 471280 280219 471336
rect 279956 471278 280219 471280
rect 280153 471275 280219 471278
rect 552054 471276 552060 471340
rect 552124 471276 552130 471340
rect 552062 471036 552122 471276
rect 552289 470794 552355 470797
rect 552246 470792 552355 470794
rect 552246 470736 552294 470792
rect 552350 470736 552355 470792
rect 552246 470731 552355 470736
rect 552246 470356 552306 470731
rect 552381 470114 552447 470117
rect 552381 470112 552490 470114
rect 552381 470056 552386 470112
rect 552442 470056 552490 470112
rect 552381 470051 552490 470056
rect 552430 469812 552490 470051
rect 552565 469570 552631 469573
rect 552565 469568 552674 469570
rect 552565 469512 552570 469568
rect 552626 469512 552674 469568
rect 552565 469507 552674 469512
rect 552614 469268 552674 469507
rect 552422 468964 552428 469028
rect 552492 468964 552498 469028
rect 552430 468588 552490 468964
rect 553342 468074 553348 468076
rect 552644 468014 553348 468074
rect 553342 468012 553348 468014
rect 553412 468012 553418 468076
rect 552606 467740 552612 467804
rect 552676 467740 552682 467804
rect 552614 467500 552674 467740
rect -960 466700 480 466940
rect 554998 466850 555004 466852
rect 552644 466790 555004 466850
rect 554998 466788 555004 466790
rect 555068 466788 555074 466852
rect 552790 466306 552796 466308
rect 552644 466246 552796 466306
rect 552790 466244 552796 466246
rect 552860 466244 552866 466308
rect 555366 465626 555372 465628
rect 552644 465566 555372 465626
rect 555366 465564 555372 465566
rect 555436 465564 555442 465628
rect 156045 465354 156111 465357
rect 153916 465352 156111 465354
rect 153916 465296 156050 465352
rect 156106 465296 156111 465352
rect 153916 465294 156111 465296
rect 156045 465291 156111 465294
rect 552238 465292 552244 465356
rect 552308 465292 552314 465356
rect 552246 465052 552306 465292
rect 552054 464748 552060 464812
rect 552124 464748 552130 464812
rect 552062 464508 552122 464748
rect 554814 463858 554820 463860
rect 552644 463798 554820 463858
rect 554814 463796 554820 463798
rect 554884 463796 554890 463860
rect 155769 463722 155835 463725
rect 156137 463722 156203 463725
rect 155769 463720 156203 463722
rect 155769 463664 155774 463720
rect 155830 463664 156142 463720
rect 156198 463664 156203 463720
rect 155769 463662 156203 463664
rect 155769 463659 155835 463662
rect 156137 463659 156203 463662
rect 552054 463524 552060 463588
rect 552124 463524 552130 463588
rect 552062 463284 552122 463524
rect 580165 463450 580231 463453
rect 583520 463450 584960 463540
rect 580165 463448 584960 463450
rect 580165 463392 580170 463448
rect 580226 463392 584960 463448
rect 580165 463390 584960 463392
rect 580165 463387 580231 463390
rect 583520 463300 584960 463390
rect 312537 462770 312603 462773
rect 553025 462770 553091 462773
rect 312537 462768 316020 462770
rect 312537 462712 312542 462768
rect 312598 462712 316020 462768
rect 312537 462710 316020 462712
rect 552644 462768 553091 462770
rect 552644 462712 553030 462768
rect 553086 462712 553091 462768
rect 552644 462710 553091 462712
rect 312537 462707 312603 462710
rect 553025 462707 553091 462710
rect 555877 462090 555943 462093
rect 552644 462088 555943 462090
rect 552644 462032 555882 462088
rect 555938 462032 555943 462088
rect 552644 462030 555943 462032
rect 555877 462027 555943 462030
rect 553710 461546 553716 461548
rect 552644 461486 553716 461546
rect 553710 461484 553716 461486
rect 553780 461484 553786 461548
rect 555785 461002 555851 461005
rect 552644 461000 555851 461002
rect 552644 460944 555790 461000
rect 555846 460944 555851 461000
rect 552644 460942 555851 460944
rect 555785 460939 555851 460942
rect 552381 460730 552447 460733
rect 552381 460728 552490 460730
rect 552381 460672 552386 460728
rect 552442 460672 552490 460728
rect 552381 460667 552490 460672
rect 552430 460292 552490 460667
rect 552657 460050 552723 460053
rect 552614 460048 552723 460050
rect 552614 459992 552662 460048
rect 552718 459992 552723 460048
rect 552614 459987 552723 459992
rect 552614 459748 552674 459987
rect 552933 459234 552999 459237
rect 552644 459232 552999 459234
rect 552644 459176 552938 459232
rect 552994 459176 552999 459232
rect 552644 459174 552999 459176
rect 552933 459171 552999 459174
rect 555693 458554 555759 458557
rect 552644 458552 555759 458554
rect 552644 458496 555698 458552
rect 555754 458496 555759 458552
rect 552644 458494 555759 458496
rect 555693 458491 555759 458494
rect 552841 458010 552907 458013
rect 552644 458008 552907 458010
rect 552644 457952 552846 458008
rect 552902 457952 552907 458008
rect 552644 457950 552907 457952
rect 552841 457947 552907 457950
rect 553526 457330 553532 457332
rect 552644 457270 553532 457330
rect 553526 457268 553532 457270
rect 553596 457268 553602 457332
rect 552841 456786 552907 456789
rect 552644 456784 552907 456786
rect 552644 456728 552846 456784
rect 552902 456728 552907 456784
rect 552644 456726 552907 456728
rect 552841 456723 552907 456726
rect 555049 456242 555115 456245
rect 552644 456240 555115 456242
rect 552644 456184 555054 456240
rect 555110 456184 555115 456240
rect 552644 456182 555115 456184
rect 555049 456179 555115 456182
rect 554865 455562 554931 455565
rect 552644 455560 554931 455562
rect 552644 455504 554870 455560
rect 554926 455504 554931 455560
rect 552644 455502 554931 455504
rect 554865 455499 554931 455502
rect 554957 455018 555023 455021
rect 552644 455016 555023 455018
rect 552644 454960 554962 455016
rect 555018 454960 555023 455016
rect 552644 454958 555023 454960
rect 554957 454955 555023 454958
rect 552381 454746 552447 454749
rect 552381 454744 552490 454746
rect 552381 454688 552386 454744
rect 552442 454688 552490 454744
rect 552381 454683 552490 454688
rect 552430 454444 552490 454683
rect 552749 454202 552815 454205
rect 552614 454200 552815 454202
rect 552614 454144 552754 454200
rect 552810 454144 552815 454200
rect 552614 454142 552815 454144
rect 282913 454066 282979 454069
rect 283189 454066 283255 454069
rect 282913 454064 283255 454066
rect 282913 454008 282918 454064
rect 282974 454008 283194 454064
rect 283250 454008 283255 454064
rect 282913 454006 283255 454008
rect 282913 454003 282979 454006
rect 283189 454003 283255 454006
rect 552614 453764 552674 454142
rect 552749 454139 552815 454142
rect 552565 453522 552631 453525
rect 552565 453520 552674 453522
rect 552565 453464 552570 453520
rect 552626 453464 552674 453520
rect 552565 453459 552674 453464
rect 552614 453220 552674 453459
rect 552657 452978 552723 452981
rect 552614 452976 552723 452978
rect 552614 452920 552662 452976
rect 552718 452920 552723 452976
rect 552614 452915 552723 452920
rect 552614 452676 552674 452915
rect -960 452434 480 452524
rect 3417 452434 3483 452437
rect -960 452432 3483 452434
rect -960 452376 3422 452432
rect 3478 452376 3483 452432
rect -960 452374 3483 452376
rect -960 452284 480 452374
rect 3417 452371 3483 452374
rect 555601 452026 555667 452029
rect 552644 452024 555667 452026
rect 552644 451968 555606 452024
rect 555662 451968 555667 452024
rect 552644 451966 555667 451968
rect 555601 451963 555667 451966
rect 552013 451754 552079 451757
rect 580901 451754 580967 451757
rect 583520 451754 584960 451844
rect 552013 451752 552122 451754
rect 552013 451696 552018 451752
rect 552074 451696 552122 451752
rect 552013 451691 552122 451696
rect 580901 451752 584960 451754
rect 580901 451696 580906 451752
rect 580962 451696 584960 451752
rect 580901 451694 584960 451696
rect 580901 451691 580967 451694
rect 552062 451452 552122 451691
rect 583520 451604 584960 451694
rect 552013 451210 552079 451213
rect 552013 451208 552122 451210
rect 552013 451152 552018 451208
rect 552074 451152 552122 451208
rect 552013 451147 552122 451152
rect 185577 450938 185643 450941
rect 185577 450936 188140 450938
rect 185577 450880 185582 450936
rect 185638 450880 188140 450936
rect 552062 450908 552122 451147
rect 185577 450878 188140 450880
rect 185577 450875 185643 450878
rect 443637 450666 443703 450669
rect 443637 450664 446108 450666
rect 443637 450608 443642 450664
rect 443698 450608 446108 450664
rect 443637 450606 446108 450608
rect 443637 450603 443703 450606
rect 555417 450258 555483 450261
rect 552644 450256 555483 450258
rect 552644 450200 555422 450256
rect 555478 450200 555483 450256
rect 552644 450198 555483 450200
rect 555417 450195 555483 450198
rect 552381 449986 552447 449989
rect 552381 449984 552490 449986
rect 552381 449928 552386 449984
rect 552442 449928 552490 449984
rect 552381 449923 552490 449928
rect 552430 449684 552490 449923
rect 554037 449034 554103 449037
rect 552644 449032 554103 449034
rect 552644 448976 554042 449032
rect 554098 448976 554103 449032
rect 552644 448974 554103 448976
rect 554037 448971 554103 448974
rect 554313 448490 554379 448493
rect 552644 448488 554379 448490
rect 552644 448432 554318 448488
rect 554374 448432 554379 448488
rect 552644 448430 554379 448432
rect 554313 448427 554379 448430
rect 553945 447946 554011 447949
rect 552644 447944 554011 447946
rect 552644 447888 553950 447944
rect 554006 447888 554011 447944
rect 552644 447886 554011 447888
rect 553945 447883 554011 447886
rect 552013 447674 552079 447677
rect 552013 447672 552122 447674
rect 552013 447616 552018 447672
rect 552074 447616 552122 447672
rect 552013 447611 552122 447616
rect 552062 447236 552122 447611
rect 552197 446994 552263 446997
rect 552197 446992 552306 446994
rect 552197 446936 552202 446992
rect 552258 446936 552306 446992
rect 552197 446931 552306 446936
rect 552246 446692 552306 446931
rect 555325 446178 555391 446181
rect 552644 446176 555391 446178
rect 552644 446120 555330 446176
rect 555386 446120 555391 446176
rect 552644 446118 555391 446120
rect 555325 446115 555391 446118
rect 553853 445498 553919 445501
rect 552644 445496 553919 445498
rect 552644 445440 553858 445496
rect 553914 445440 553919 445496
rect 552644 445438 553919 445440
rect 553853 445435 553919 445438
rect 552565 445226 552631 445229
rect 552565 445224 552674 445226
rect 552565 445168 552570 445224
rect 552626 445168 552674 445224
rect 552565 445163 552674 445168
rect 552614 444924 552674 445163
rect 553761 444410 553827 444413
rect 552644 444408 553827 444410
rect 552644 444352 553766 444408
rect 553822 444352 553827 444408
rect 552644 444350 553827 444352
rect 553761 444347 553827 444350
rect 553393 443730 553459 443733
rect 552644 443728 553459 443730
rect 552644 443672 553398 443728
rect 553454 443672 553459 443728
rect 552644 443670 553459 443672
rect 553393 443667 553459 443670
rect 12617 443594 12683 443597
rect 12617 443592 16100 443594
rect 12617 443536 12622 443592
rect 12678 443536 16100 443592
rect 12617 443534 16100 443536
rect 12617 443531 12683 443534
rect 553669 443186 553735 443189
rect 552644 443184 553735 443186
rect 552644 443128 553674 443184
rect 553730 443128 553735 443184
rect 552644 443126 553735 443128
rect 553669 443123 553735 443126
rect 555233 442506 555299 442509
rect 552644 442504 555299 442506
rect 552644 442448 555238 442504
rect 555294 442448 555299 442504
rect 552644 442446 555299 442448
rect 555233 442443 555299 442446
rect 553577 441962 553643 441965
rect 552644 441960 553643 441962
rect 552644 441904 553582 441960
rect 553638 441904 553643 441960
rect 552644 441902 553643 441904
rect 553577 441899 553643 441902
rect 552105 441690 552171 441693
rect 552062 441688 552171 441690
rect 552062 441632 552110 441688
rect 552166 441632 552171 441688
rect 552062 441627 552171 441632
rect 552062 441388 552122 441627
rect 554078 440738 554084 440740
rect 552644 440678 554084 440738
rect 554078 440676 554084 440678
rect 554148 440676 554154 440740
rect 554129 440194 554195 440197
rect 552644 440192 554195 440194
rect 552644 440136 554134 440192
rect 554190 440136 554195 440192
rect 552644 440134 554195 440136
rect 554129 440131 554195 440134
rect 583520 439772 584960 440012
rect 313273 439650 313339 439653
rect 314653 439650 314719 439653
rect 553485 439650 553551 439653
rect 313273 439648 316020 439650
rect 313273 439592 313278 439648
rect 313334 439592 314658 439648
rect 314714 439592 316020 439648
rect 313273 439590 316020 439592
rect 552644 439648 553551 439650
rect 552644 439592 553490 439648
rect 553546 439592 553551 439648
rect 552644 439590 553551 439592
rect 313273 439587 313339 439590
rect 314653 439587 314719 439590
rect 553485 439587 553551 439590
rect 554221 438970 554287 438973
rect 552644 438968 554287 438970
rect 552644 438912 554226 438968
rect 554282 438912 554287 438968
rect 552644 438910 554287 438912
rect 554221 438907 554287 438910
rect 555141 438426 555207 438429
rect 552644 438424 555207 438426
rect 552644 438368 555146 438424
rect 555202 438368 555207 438424
rect 552644 438366 555207 438368
rect 555141 438363 555207 438366
rect -960 438018 480 438108
rect 3509 438018 3575 438021
rect -960 438016 3575 438018
rect -960 437960 3514 438016
rect 3570 437960 3575 438016
rect -960 437958 3575 437960
rect -960 437868 480 437958
rect 3509 437955 3575 437958
rect 555509 437882 555575 437885
rect 552644 437880 555575 437882
rect 552644 437824 555514 437880
rect 555570 437824 555575 437880
rect 552644 437822 555575 437824
rect 555509 437819 555575 437822
rect 556061 437202 556127 437205
rect 552644 437200 556127 437202
rect 552644 437144 556066 437200
rect 556122 437144 556127 437200
rect 552644 437142 556127 437144
rect 556061 437139 556127 437142
rect 554773 436658 554839 436661
rect 552644 436656 554839 436658
rect 552644 436600 554778 436656
rect 554834 436600 554839 436656
rect 552644 436598 554839 436600
rect 554773 436595 554839 436598
rect 554773 436114 554839 436117
rect 552644 436112 554839 436114
rect 552644 436056 554778 436112
rect 554834 436056 554839 436112
rect 552644 436054 554839 436056
rect 554773 436051 554839 436054
rect 554773 435434 554839 435437
rect 552644 435432 554839 435434
rect 552644 435376 554778 435432
rect 554834 435376 554839 435432
rect 552644 435374 554839 435376
rect 554773 435371 554839 435374
rect 554865 434890 554931 434893
rect 552644 434888 554931 434890
rect 552644 434832 554870 434888
rect 554926 434832 554931 434888
rect 552644 434830 554931 434832
rect 554865 434827 554931 434830
rect 282729 434754 282795 434757
rect 282913 434754 282979 434757
rect 282729 434752 282979 434754
rect 282729 434696 282734 434752
rect 282790 434696 282918 434752
rect 282974 434696 282979 434752
rect 282729 434694 282979 434696
rect 282729 434691 282795 434694
rect 282913 434691 282979 434694
rect 554773 434210 554839 434213
rect 552644 434208 554839 434210
rect 552644 434152 554778 434208
rect 554834 434152 554839 434208
rect 552644 434150 554839 434152
rect 554773 434147 554839 434150
rect 554865 433666 554931 433669
rect 552644 433664 554931 433666
rect 552644 433608 554870 433664
rect 554926 433608 554931 433664
rect 552644 433606 554931 433608
rect 554865 433603 554931 433606
rect 554773 433122 554839 433125
rect 552644 433120 554839 433122
rect 552644 433064 554778 433120
rect 554834 433064 554839 433120
rect 552644 433062 554839 433064
rect 554773 433059 554839 433062
rect 554865 432442 554931 432445
rect 552644 432440 554931 432442
rect 552644 432384 554870 432440
rect 554926 432384 554931 432440
rect 552644 432382 554931 432384
rect 554865 432379 554931 432382
rect 554773 431898 554839 431901
rect 552644 431896 554839 431898
rect 552644 431840 554778 431896
rect 554834 431840 554839 431896
rect 552644 431838 554839 431840
rect 554773 431835 554839 431838
rect 554865 431354 554931 431357
rect 552644 431352 554931 431354
rect 552644 431296 554870 431352
rect 554926 431296 554931 431352
rect 552644 431294 554931 431296
rect 554865 431291 554931 431294
rect 554957 430674 555023 430677
rect 552644 430672 555023 430674
rect 552644 430616 554962 430672
rect 555018 430616 555023 430672
rect 552644 430614 555023 430616
rect 554957 430611 555023 430614
rect 281533 430538 281599 430541
rect 282177 430538 282243 430541
rect 279956 430536 282243 430538
rect 279956 430480 281538 430536
rect 281594 430480 282182 430536
rect 282238 430480 282243 430536
rect 279956 430478 282243 430480
rect 281533 430475 281599 430478
rect 282177 430475 282243 430478
rect 554773 430130 554839 430133
rect 552644 430128 554839 430130
rect 552644 430072 554778 430128
rect 554834 430072 554839 430128
rect 552644 430070 554839 430072
rect 554773 430067 554839 430070
rect 554865 429586 554931 429589
rect 552644 429584 554931 429586
rect 552644 429528 554870 429584
rect 554926 429528 554931 429584
rect 552644 429526 554931 429528
rect 554865 429523 554931 429526
rect 554865 428906 554931 428909
rect 552644 428904 554931 428906
rect 552644 428848 554870 428904
rect 554926 428848 554931 428904
rect 552644 428846 554931 428848
rect 554865 428843 554931 428846
rect 317086 428708 317092 428772
rect 317156 428770 317162 428772
rect 338113 428770 338179 428773
rect 317156 428768 338179 428770
rect 317156 428712 338118 428768
rect 338174 428712 338179 428768
rect 317156 428710 338179 428712
rect 317156 428708 317162 428710
rect 338113 428707 338179 428710
rect 316902 428572 316908 428636
rect 316972 428634 316978 428636
rect 338389 428634 338455 428637
rect 316972 428632 338455 428634
rect 316972 428576 338394 428632
rect 338450 428576 338455 428632
rect 316972 428574 338455 428576
rect 316972 428572 316978 428574
rect 338389 428571 338455 428574
rect 317270 428436 317276 428500
rect 317340 428498 317346 428500
rect 343633 428498 343699 428501
rect 317340 428496 343699 428498
rect 317340 428440 343638 428496
rect 343694 428440 343699 428496
rect 317340 428438 343699 428440
rect 317340 428436 317346 428438
rect 343633 428435 343699 428438
rect 554773 428362 554839 428365
rect 552644 428360 554839 428362
rect 552644 428304 554778 428360
rect 554834 428304 554839 428360
rect 552644 428302 554839 428304
rect 554773 428299 554839 428302
rect 583520 428076 584960 428316
rect 554773 427818 554839 427821
rect 552644 427816 554839 427818
rect 552644 427760 554778 427816
rect 554834 427760 554839 427816
rect 552644 427758 554839 427760
rect 554773 427755 554839 427758
rect -960 423738 480 423828
rect 3417 423738 3483 423741
rect -960 423736 3483 423738
rect -960 423680 3422 423736
rect 3478 423680 3483 423736
rect -960 423678 3483 423680
rect -960 423588 480 423678
rect 3417 423675 3483 423678
rect 153886 421290 153946 421804
rect 281625 421292 281691 421293
rect 155902 421290 155908 421292
rect 153886 421230 155908 421290
rect 155902 421228 155908 421230
rect 155972 421228 155978 421292
rect 281574 421228 281580 421292
rect 281644 421290 281691 421292
rect 281644 421288 281736 421290
rect 281686 421232 281736 421288
rect 281644 421230 281736 421232
rect 281644 421228 281691 421230
rect 281625 421227 281691 421228
rect 580165 416530 580231 416533
rect 583520 416530 584960 416620
rect 580165 416528 584960 416530
rect 580165 416472 580170 416528
rect 580226 416472 584960 416528
rect 580165 416470 584960 416472
rect 580165 416467 580231 416470
rect 583520 416380 584960 416470
rect -960 409172 480 409412
rect 156137 405922 156203 405925
rect 155542 405920 156203 405922
rect 155542 405864 156142 405920
rect 156198 405864 156203 405920
rect 155542 405862 156203 405864
rect 155542 405786 155602 405862
rect 156137 405859 156203 405862
rect 155677 405786 155743 405789
rect 155542 405784 155743 405786
rect 155542 405728 155682 405784
rect 155738 405728 155743 405784
rect 155542 405726 155743 405728
rect 155677 405723 155743 405726
rect 580901 404834 580967 404837
rect 583520 404834 584960 404924
rect 580901 404832 584960 404834
rect 580901 404776 580906 404832
rect 580962 404776 584960 404832
rect 580901 404774 584960 404776
rect 580901 404771 580967 404774
rect 583520 404684 584960 404774
rect 153878 403548 153884 403612
rect 153948 403610 153954 403612
rect 283189 403610 283255 403613
rect 153948 403608 283255 403610
rect 153948 403552 283194 403608
rect 283250 403552 283255 403608
rect 153948 403550 283255 403552
rect 153948 403548 153954 403550
rect 283189 403547 283255 403550
rect 131021 401434 131087 401437
rect 153326 401434 153332 401436
rect 131021 401432 153332 401434
rect 131021 401376 131026 401432
rect 131082 401376 153332 401432
rect 131021 401374 153332 401376
rect 131021 401371 131087 401374
rect 153326 401372 153332 401374
rect 153396 401372 153402 401436
rect 129641 401298 129707 401301
rect 154614 401298 154620 401300
rect 129641 401296 154620 401298
rect 129641 401240 129646 401296
rect 129702 401240 154620 401296
rect 129641 401238 154620 401240
rect 129641 401235 129707 401238
rect 154614 401236 154620 401238
rect 154684 401236 154690 401300
rect 126881 401162 126947 401165
rect 153142 401162 153148 401164
rect 126881 401160 153148 401162
rect 126881 401104 126886 401160
rect 126942 401104 153148 401160
rect 126881 401102 153148 401104
rect 126881 401099 126947 401102
rect 153142 401100 153148 401102
rect 153212 401100 153218 401164
rect 125501 401026 125567 401029
rect 154798 401026 154804 401028
rect 125501 401024 154804 401026
rect 125501 400968 125506 401024
rect 125562 400968 154804 401024
rect 125501 400966 154804 400968
rect 125501 400963 125567 400966
rect 154798 400964 154804 400966
rect 154868 400964 154874 401028
rect 118601 400890 118667 400893
rect 151854 400890 151860 400892
rect 118601 400888 151860 400890
rect 118601 400832 118606 400888
rect 118662 400832 151860 400888
rect 118601 400830 151860 400832
rect 118601 400827 118667 400830
rect 151854 400828 151860 400830
rect 151924 400828 151930 400892
rect 146886 398652 146892 398716
rect 146956 398714 146962 398716
rect 147438 398714 147444 398716
rect 146956 398654 147444 398714
rect 146956 398652 146962 398654
rect 147438 398652 147444 398654
rect 147508 398652 147514 398716
rect -960 395042 480 395132
rect 4797 395042 4863 395045
rect -960 395040 4863 395042
rect -960 394984 4802 395040
rect 4858 394984 4863 395040
rect -960 394982 4863 394984
rect -960 394892 480 394982
rect 4797 394979 4863 394982
rect 583520 392852 584960 393092
rect 284385 392730 284451 392733
rect 282716 392728 284451 392730
rect 282716 392672 284390 392728
rect 284446 392672 284451 392728
rect 282716 392670 284451 392672
rect 284385 392667 284451 392670
rect 147121 389468 147187 389469
rect 147070 389404 147076 389468
rect 147140 389466 147187 389468
rect 147140 389464 147232 389466
rect 147182 389408 147232 389464
rect 147140 389406 147232 389408
rect 147140 389404 147187 389406
rect 147121 389403 147187 389404
rect 146702 386548 146708 386612
rect 146772 386610 146778 386612
rect 147254 386610 147260 386612
rect 146772 386550 147260 386610
rect 146772 386548 146778 386550
rect 147254 386548 147260 386550
rect 147324 386548 147330 386612
rect 147121 386476 147187 386477
rect 147070 386474 147076 386476
rect 147030 386414 147076 386474
rect 147140 386472 147187 386476
rect 147182 386416 147187 386472
rect 147070 386412 147076 386414
rect 147140 386412 147187 386416
rect 147121 386411 147187 386412
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 2773 380626 2839 380629
rect -960 380624 2839 380626
rect -960 380568 2778 380624
rect 2834 380568 2839 380624
rect -960 380566 2839 380568
rect -960 380476 480 380566
rect 2773 380563 2839 380566
rect 78581 377362 78647 377365
rect 75900 377360 78647 377362
rect 75900 377304 78586 377360
rect 78642 377304 78647 377360
rect 75900 377302 78647 377304
rect 78581 377299 78647 377302
rect 155677 376684 155743 376685
rect 155677 376680 155724 376684
rect 155788 376682 155794 376684
rect 155677 376624 155682 376680
rect 155677 376620 155724 376624
rect 155788 376622 155834 376682
rect 155788 376620 155794 376622
rect 155677 376619 155743 376620
rect 155769 369748 155835 369749
rect 155718 369746 155724 369748
rect 155678 369686 155724 369746
rect 155788 369744 155835 369748
rect 155830 369688 155835 369744
rect 155718 369684 155724 369686
rect 155788 369684 155835 369688
rect 155769 369683 155835 369684
rect 284293 369610 284359 369613
rect 282716 369608 284359 369610
rect 282716 369552 284298 369608
rect 284354 369552 284359 369608
rect 282716 369550 284359 369552
rect 284293 369547 284359 369550
rect 580165 369610 580231 369613
rect 583520 369610 584960 369700
rect 580165 369608 584960 369610
rect 580165 369552 580170 369608
rect 580226 369552 584960 369608
rect 580165 369550 584960 369552
rect 580165 369547 580231 369550
rect 583520 369460 584960 369550
rect -960 366210 480 366300
rect 2773 366210 2839 366213
rect -960 366208 2839 366210
rect -960 366152 2778 366208
rect 2834 366152 2839 366208
rect -960 366150 2839 366152
rect -960 366060 480 366150
rect 2773 366147 2839 366150
rect 153878 364306 153884 364308
rect 75870 364246 153884 364306
rect 75870 363732 75930 364246
rect 153878 364244 153884 364246
rect 153948 364244 153954 364308
rect 147254 360498 147260 360500
rect 146894 360438 147260 360498
rect 146894 360092 146954 360438
rect 147254 360436 147260 360438
rect 147324 360436 147330 360500
rect 147070 360300 147076 360364
rect 147140 360300 147146 360364
rect 147078 360092 147138 360300
rect 146886 360028 146892 360092
rect 146956 360028 146962 360092
rect 147070 360028 147076 360092
rect 147140 360028 147146 360092
rect 580901 357914 580967 357917
rect 583520 357914 584960 358004
rect 580901 357912 584960 357914
rect 580901 357856 580906 357912
rect 580962 357856 584960 357912
rect 580901 357854 584960 357856
rect 580901 357851 580967 357854
rect 583520 357764 584960 357854
rect 20478 357308 20484 357372
rect 20548 357370 20554 357372
rect 21357 357370 21423 357373
rect 20548 357368 21423 357370
rect 20548 357312 21362 357368
rect 21418 357312 21423 357368
rect 20548 357310 21423 357312
rect 20548 357308 20554 357310
rect 21357 357307 21423 357310
rect -960 351780 480 352020
rect 147581 351930 147647 351933
rect 147581 351928 147874 351930
rect 147581 351872 147586 351928
rect 147642 351872 147874 351928
rect 147581 351870 147874 351872
rect 147581 351867 147647 351870
rect 114001 351794 114067 351797
rect 122649 351794 122715 351797
rect 114001 351792 122715 351794
rect 114001 351736 114006 351792
rect 114062 351736 122654 351792
rect 122710 351736 122715 351792
rect 114001 351734 122715 351736
rect 114001 351731 114067 351734
rect 122649 351731 122715 351734
rect 146937 351794 147003 351797
rect 147070 351794 147076 351796
rect 146937 351792 147076 351794
rect 146937 351736 146942 351792
rect 146998 351736 147076 351792
rect 146937 351734 147076 351736
rect 146937 351731 147003 351734
rect 147070 351732 147076 351734
rect 147140 351732 147146 351796
rect 147213 351794 147279 351797
rect 147673 351794 147739 351797
rect 147814 351796 147874 351870
rect 147213 351792 147739 351794
rect 147213 351736 147218 351792
rect 147274 351736 147678 351792
rect 147734 351736 147739 351792
rect 147213 351734 147739 351736
rect 147213 351731 147279 351734
rect 147673 351731 147739 351734
rect 147806 351732 147812 351796
rect 147876 351732 147882 351796
rect 148041 351794 148107 351797
rect 148174 351794 148180 351796
rect 148041 351792 148180 351794
rect 148041 351736 148046 351792
rect 148102 351736 148180 351792
rect 148041 351734 148180 351736
rect 148041 351731 148107 351734
rect 148174 351732 148180 351734
rect 148244 351732 148250 351796
rect 149421 351794 149487 351797
rect 149646 351794 149652 351796
rect 149421 351792 149652 351794
rect 149421 351736 149426 351792
rect 149482 351736 149652 351792
rect 149421 351734 149652 351736
rect 149421 351731 149487 351734
rect 149646 351732 149652 351734
rect 149716 351732 149722 351796
rect 149830 351732 149836 351796
rect 149900 351794 149906 351796
rect 150065 351794 150131 351797
rect 149900 351792 150131 351794
rect 149900 351736 150070 351792
rect 150126 351736 150131 351792
rect 149900 351734 150131 351736
rect 149900 351732 149906 351734
rect 150065 351731 150131 351734
rect 150934 351732 150940 351796
rect 151004 351794 151010 351796
rect 151169 351794 151235 351797
rect 152365 351796 152431 351797
rect 152365 351794 152412 351796
rect 151004 351792 151235 351794
rect 151004 351736 151174 351792
rect 151230 351736 151235 351792
rect 151004 351734 151235 351736
rect 152320 351792 152412 351794
rect 152320 351736 152370 351792
rect 152320 351734 152412 351736
rect 151004 351732 151010 351734
rect 151169 351731 151235 351734
rect 152365 351732 152412 351734
rect 152476 351732 152482 351796
rect 189441 351794 189507 351797
rect 189758 351794 189764 351796
rect 189441 351792 189764 351794
rect 189441 351736 189446 351792
rect 189502 351736 189764 351792
rect 189441 351734 189764 351736
rect 152365 351731 152431 351732
rect 189441 351731 189507 351734
rect 189758 351732 189764 351734
rect 189828 351732 189834 351796
rect 191046 351732 191052 351796
rect 191116 351794 191122 351796
rect 191189 351794 191255 351797
rect 191116 351792 191255 351794
rect 191116 351736 191194 351792
rect 191250 351736 191255 351792
rect 191116 351734 191255 351736
rect 191116 351732 191122 351734
rect 191189 351731 191255 351734
rect 111701 351658 111767 351661
rect 150382 351658 150388 351660
rect 111701 351656 150388 351658
rect 111701 351600 111706 351656
rect 111762 351600 150388 351656
rect 111701 351598 150388 351600
rect 111701 351595 111767 351598
rect 150382 351596 150388 351598
rect 150452 351596 150458 351660
rect 189574 351596 189580 351660
rect 189644 351658 189650 351660
rect 189901 351658 189967 351661
rect 189644 351656 189967 351658
rect 189644 351600 189906 351656
rect 189962 351600 189967 351656
rect 189644 351598 189967 351600
rect 189644 351596 189650 351598
rect 189901 351595 189967 351598
rect 110689 351522 110755 351525
rect 147213 351522 147279 351525
rect 110689 351520 147279 351522
rect 110689 351464 110694 351520
rect 110750 351464 147218 351520
rect 147274 351464 147279 351520
rect 110689 351462 147279 351464
rect 110689 351459 110755 351462
rect 147213 351459 147279 351462
rect 147673 351522 147739 351525
rect 150750 351522 150756 351524
rect 147673 351520 150756 351522
rect 147673 351464 147678 351520
rect 147734 351464 150756 351520
rect 147673 351462 150756 351464
rect 147673 351459 147739 351462
rect 150750 351460 150756 351462
rect 150820 351460 150826 351524
rect 108665 351386 108731 351389
rect 148358 351386 148364 351388
rect 108665 351384 148364 351386
rect 108665 351328 108670 351384
rect 108726 351328 148364 351384
rect 108665 351326 148364 351328
rect 108665 351323 108731 351326
rect 148358 351324 148364 351326
rect 148428 351324 148434 351388
rect 153193 351386 153259 351389
rect 153694 351386 153700 351388
rect 153193 351384 153700 351386
rect 153193 351328 153198 351384
rect 153254 351328 153700 351384
rect 153193 351326 153700 351328
rect 153193 351323 153259 351326
rect 153694 351324 153700 351326
rect 153764 351324 153770 351388
rect 109585 351250 109651 351253
rect 142613 351250 142679 351253
rect 109585 351248 142679 351250
rect 109585 351192 109590 351248
rect 109646 351192 142618 351248
rect 142674 351192 142679 351248
rect 109585 351190 142679 351192
rect 109585 351187 109651 351190
rect 142613 351187 142679 351190
rect 142797 351250 142863 351253
rect 149094 351250 149100 351252
rect 142797 351248 149100 351250
rect 142797 351192 142802 351248
rect 142858 351192 149100 351248
rect 142797 351190 149100 351192
rect 142797 351187 142863 351190
rect 149094 351188 149100 351190
rect 149164 351188 149170 351252
rect 107561 351114 107627 351117
rect 147990 351114 147996 351116
rect 107561 351112 147996 351114
rect 107561 351056 107566 351112
rect 107622 351056 147996 351112
rect 107561 351054 147996 351056
rect 107561 351051 107627 351054
rect 147990 351052 147996 351054
rect 148060 351052 148066 351116
rect 117129 350978 117195 350981
rect 142797 350978 142863 350981
rect 117129 350976 142863 350978
rect 117129 350920 117134 350976
rect 117190 350920 142802 350976
rect 142858 350920 142863 350976
rect 117129 350918 142863 350920
rect 117129 350915 117195 350918
rect 142797 350915 142863 350918
rect 146293 350978 146359 350981
rect 146886 350978 146892 350980
rect 146293 350976 146892 350978
rect 146293 350920 146298 350976
rect 146354 350920 146892 350976
rect 146293 350918 146892 350920
rect 146293 350915 146359 350918
rect 146886 350916 146892 350918
rect 146956 350916 146962 350980
rect 115105 350842 115171 350845
rect 147622 350842 147628 350844
rect 115105 350840 147628 350842
rect 115105 350784 115110 350840
rect 115166 350784 147628 350840
rect 115105 350782 147628 350784
rect 115105 350779 115171 350782
rect 147622 350780 147628 350782
rect 147692 350780 147698 350844
rect 149053 350842 149119 350845
rect 149278 350842 149284 350844
rect 149053 350840 149284 350842
rect 149053 350784 149058 350840
rect 149114 350784 149284 350840
rect 149053 350782 149284 350784
rect 149053 350779 149119 350782
rect 149278 350780 149284 350782
rect 149348 350780 149354 350844
rect 122649 350706 122715 350709
rect 142613 350706 142679 350709
rect 150566 350706 150572 350708
rect 122649 350704 122850 350706
rect 122649 350648 122654 350704
rect 122710 350648 122850 350704
rect 122649 350646 122850 350648
rect 122649 350643 122715 350646
rect 122790 350570 122850 350646
rect 142613 350704 150572 350706
rect 142613 350648 142618 350704
rect 142674 350648 150572 350704
rect 142613 350646 150572 350648
rect 142613 350643 142679 350646
rect 150566 350644 150572 350646
rect 150636 350644 150642 350708
rect 147581 350570 147647 350573
rect 122790 350568 147647 350570
rect 122790 350512 147586 350568
rect 147642 350512 147647 350568
rect 122790 350510 147647 350512
rect 147581 350507 147647 350510
rect 583520 345932 584960 346172
rect -960 337514 480 337604
rect 3141 337514 3207 337517
rect -960 337512 3207 337514
rect -960 337456 3146 337512
rect 3202 337456 3207 337512
rect -960 337454 3207 337456
rect -960 337364 480 337454
rect 3141 337451 3207 337454
rect 282177 336018 282243 336021
rect 279006 336016 282243 336018
rect 279006 335960 282182 336016
rect 282238 335960 282243 336016
rect 279006 335958 282243 335960
rect 279006 335920 279066 335958
rect 282177 335955 282243 335958
rect 583520 334236 584960 334476
rect 304257 328266 304323 328269
rect 301668 328264 304323 328266
rect 301668 328208 304262 328264
rect 304318 328208 304323 328264
rect 301668 328206 304323 328208
rect 304257 328203 304323 328206
rect 303613 326362 303679 326365
rect 301668 326360 303679 326362
rect 301668 326304 303618 326360
rect 303674 326304 303679 326360
rect 301668 326302 303679 326304
rect 303613 326299 303679 326302
rect 289721 325274 289787 325277
rect 289721 325272 290812 325274
rect 289721 325216 289726 325272
rect 289782 325216 290812 325272
rect 289721 325214 290812 325216
rect 289721 325211 289787 325214
rect 303613 324458 303679 324461
rect 301668 324456 303679 324458
rect 301668 324400 303618 324456
rect 303674 324400 303679 324456
rect 301668 324398 303679 324400
rect 303613 324395 303679 324398
rect -960 323098 480 323188
rect 2773 323098 2839 323101
rect -960 323096 2839 323098
rect -960 323040 2778 323096
rect 2834 323040 2839 323096
rect -960 323038 2839 323040
rect -960 322948 480 323038
rect 2773 323035 2839 323038
rect 580165 322690 580231 322693
rect 583520 322690 584960 322780
rect 580165 322688 584960 322690
rect 580165 322632 580170 322688
rect 580226 322632 584960 322688
rect 580165 322630 584960 322632
rect 580165 322627 580231 322630
rect 304349 322554 304415 322557
rect 301668 322552 304415 322554
rect 301668 322496 304354 322552
rect 304410 322496 304415 322552
rect 583520 322540 584960 322630
rect 301668 322494 304415 322496
rect 304349 322491 304415 322494
rect 219934 322084 219940 322148
rect 220004 322146 220010 322148
rect 282269 322146 282335 322149
rect 220004 322144 282335 322146
rect 220004 322088 282274 322144
rect 282330 322088 282335 322144
rect 220004 322086 282335 322088
rect 220004 322084 220010 322086
rect 282269 322083 282335 322086
rect 304441 320650 304507 320653
rect 301668 320648 304507 320650
rect 301668 320592 304446 320648
rect 304502 320592 304507 320648
rect 301668 320590 304507 320592
rect 304441 320587 304507 320590
rect 189073 320378 189139 320381
rect 190126 320378 190132 320380
rect 189073 320376 190132 320378
rect 189073 320320 189078 320376
rect 189134 320320 190132 320376
rect 189073 320318 190132 320320
rect 189073 320315 189139 320318
rect 190126 320316 190132 320318
rect 190196 320316 190202 320380
rect 193397 320378 193463 320381
rect 194358 320378 194364 320380
rect 193397 320376 194364 320378
rect 193397 320320 193402 320376
rect 193458 320320 194364 320376
rect 193397 320318 194364 320320
rect 193397 320315 193463 320318
rect 194358 320316 194364 320318
rect 194428 320316 194434 320380
rect 190177 320242 190243 320245
rect 190310 320242 190316 320244
rect 190177 320240 190316 320242
rect 190177 320184 190182 320240
rect 190238 320184 190316 320240
rect 190177 320182 190316 320184
rect 190177 320179 190243 320182
rect 190310 320180 190316 320182
rect 190380 320180 190386 320244
rect 191281 320242 191347 320245
rect 191598 320242 191604 320244
rect 191281 320240 191604 320242
rect 191281 320184 191286 320240
rect 191342 320184 191604 320240
rect 191281 320182 191604 320184
rect 191281 320179 191347 320182
rect 191598 320180 191604 320182
rect 191668 320180 191674 320244
rect 192385 320242 192451 320245
rect 193070 320242 193076 320244
rect 192385 320240 193076 320242
rect 192385 320184 192390 320240
rect 192446 320184 193076 320240
rect 192385 320182 193076 320184
rect 192385 320179 192451 320182
rect 193070 320180 193076 320182
rect 193140 320180 193146 320244
rect 194174 320180 194180 320244
rect 194244 320242 194250 320244
rect 194501 320242 194567 320245
rect 194244 320240 194567 320242
rect 194244 320184 194506 320240
rect 194562 320184 194567 320240
rect 194244 320182 194567 320184
rect 194244 320180 194250 320182
rect 194501 320179 194567 320182
rect 303613 318746 303679 318749
rect 301668 318744 303679 318746
rect 301668 318688 303618 318744
rect 303674 318688 303679 318744
rect 301668 318686 303679 318688
rect 303613 318683 303679 318686
rect 288893 317114 288959 317117
rect 288893 317112 290812 317114
rect 288893 317056 288898 317112
rect 288954 317056 290812 317112
rect 288893 317054 290812 317056
rect 288893 317051 288959 317054
rect 304349 316978 304415 316981
rect 301668 316976 304415 316978
rect 301668 316920 304354 316976
rect 304410 316920 304415 316976
rect 301668 316918 304415 316920
rect 304349 316915 304415 316918
rect 304257 315074 304323 315077
rect 301668 315072 304323 315074
rect 301668 315016 304262 315072
rect 304318 315016 304323 315072
rect 301668 315014 304323 315016
rect 304257 315011 304323 315014
rect 303613 313170 303679 313173
rect 301668 313168 303679 313170
rect 301668 313112 303618 313168
rect 303674 313112 303679 313168
rect 301668 313110 303679 313112
rect 303613 313107 303679 313110
rect 303613 311266 303679 311269
rect 301668 311264 303679 311266
rect 301668 311208 303618 311264
rect 303674 311208 303679 311264
rect 301668 311206 303679 311208
rect 303613 311203 303679 311206
rect 580349 310858 580415 310861
rect 580901 310858 580967 310861
rect 583520 310858 584960 310948
rect 580349 310856 584960 310858
rect 580349 310800 580354 310856
rect 580410 310800 580906 310856
rect 580962 310800 584960 310856
rect 580349 310798 584960 310800
rect 580349 310795 580415 310798
rect 580901 310795 580967 310798
rect 583520 310708 584960 310798
rect 303613 309362 303679 309365
rect 301668 309360 303679 309362
rect 301668 309304 303618 309360
rect 303674 309304 303679 309360
rect 301668 309302 303679 309304
rect 303613 309299 303679 309302
rect 2773 309090 2839 309093
rect 3417 309090 3483 309093
rect 2773 309088 3483 309090
rect 2773 309032 2778 309088
rect 2834 309032 3422 309088
rect 3478 309032 3483 309088
rect 2773 309030 3483 309032
rect 2773 309027 2839 309030
rect 3417 309027 3483 309030
rect 289629 308954 289695 308957
rect 289629 308952 290812 308954
rect -960 308818 480 308908
rect 289629 308896 289634 308952
rect 289690 308896 290812 308952
rect 289629 308894 290812 308896
rect 289629 308891 289695 308894
rect 2773 308818 2839 308821
rect -960 308816 2839 308818
rect -960 308760 2778 308816
rect 2834 308760 2839 308816
rect -960 308758 2839 308760
rect -960 308668 480 308758
rect 2773 308755 2839 308758
rect 303613 307458 303679 307461
rect 301668 307456 303679 307458
rect 301668 307400 303618 307456
rect 303674 307400 303679 307456
rect 301668 307398 303679 307400
rect 303613 307395 303679 307398
rect 300902 305557 300962 305660
rect 300853 305552 300962 305557
rect 300853 305496 300858 305552
rect 300914 305496 300962 305552
rect 300853 305494 300962 305496
rect 300853 305491 300919 305494
rect 292573 302834 292639 302837
rect 332910 302834 332916 302836
rect 292573 302832 332916 302834
rect 292573 302776 292578 302832
rect 292634 302776 332916 302832
rect 292573 302774 332916 302776
rect 292573 302771 292639 302774
rect 332910 302772 332916 302774
rect 332980 302772 332986 302836
rect 583520 299012 584960 299252
rect 280153 295898 280219 295901
rect 279926 295896 280219 295898
rect 279926 295840 280158 295896
rect 280214 295840 280219 295896
rect 279926 295838 280219 295840
rect 113173 295354 113239 295357
rect 111964 295352 113239 295354
rect 111964 295296 113178 295352
rect 113234 295296 113239 295352
rect 279926 295324 279986 295838
rect 280153 295835 280219 295838
rect 111964 295294 113239 295296
rect 113173 295291 113239 295294
rect -960 294402 480 294492
rect 3417 294402 3483 294405
rect -960 294400 3483 294402
rect -960 294344 3422 294400
rect 3478 294344 3483 294400
rect -960 294342 3483 294344
rect -960 294252 480 294342
rect 3417 294339 3483 294342
rect 583520 287316 584960 287556
rect -960 280122 480 280212
rect 2773 280122 2839 280125
rect -960 280120 2839 280122
rect -960 280064 2778 280120
rect 2834 280064 2839 280120
rect -960 280062 2839 280064
rect -960 279972 480 280062
rect 2773 280059 2839 280062
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 17125 274954 17191 274957
rect 185577 274954 185643 274957
rect 17125 274952 20148 274954
rect 17125 274896 17130 274952
rect 17186 274896 20148 274952
rect 17125 274894 20148 274896
rect 185577 274952 188140 274954
rect 185577 274896 185582 274952
rect 185638 274896 188140 274952
rect 185577 274894 188140 274896
rect 17125 274891 17191 274894
rect 185577 274891 185643 274894
rect -960 265706 480 265796
rect 2773 265706 2839 265709
rect -960 265704 2839 265706
rect -960 265648 2778 265704
rect 2834 265648 2839 265704
rect -960 265646 2839 265648
rect -960 265556 480 265646
rect 2773 265643 2839 265646
rect 580349 263938 580415 263941
rect 580901 263938 580967 263941
rect 583520 263938 584960 264028
rect 580349 263936 584960 263938
rect 580349 263880 580354 263936
rect 580410 263880 580906 263936
rect 580962 263880 584960 263936
rect 580349 263878 584960 263880
rect 580349 263875 580415 263878
rect 580901 263875 580967 263878
rect 583520 263788 584960 263878
rect 113909 254554 113975 254557
rect 111964 254552 113975 254554
rect 111964 254496 113914 254552
rect 113970 254496 113975 254552
rect 111964 254494 113975 254496
rect 113909 254491 113975 254494
rect 279926 254010 279986 254524
rect 281533 254010 281599 254013
rect 282177 254010 282243 254013
rect 279926 254008 282243 254010
rect 279926 253952 281538 254008
rect 281594 253952 282182 254008
rect 282238 253952 282243 254008
rect 279926 253950 282243 253952
rect 281533 253947 281599 253950
rect 282177 253947 282243 253950
rect 583520 252092 584960 252332
rect -960 251140 480 251380
rect 583520 240396 584960 240636
rect -960 237010 480 237100
rect 2773 237010 2839 237013
rect -960 237008 2839 237010
rect -960 236952 2778 237008
rect 2834 236952 2839 237008
rect -960 236950 2839 236952
rect -960 236860 480 236950
rect 2773 236947 2839 236950
rect 235257 235242 235323 235245
rect 280102 235242 280108 235244
rect 235257 235240 280108 235242
rect 235257 235184 235262 235240
rect 235318 235184 280108 235240
rect 235257 235182 280108 235184
rect 235257 235179 235323 235182
rect 280102 235180 280108 235182
rect 280172 235180 280178 235244
rect 579981 228850 580047 228853
rect 583520 228850 584960 228940
rect 579981 228848 584960 228850
rect 579981 228792 579986 228848
rect 580042 228792 584960 228848
rect 579981 228790 584960 228792
rect 579981 228787 580047 228790
rect 583520 228700 584960 228790
rect 193070 224844 193076 224908
rect 193140 224906 193146 224908
rect 207749 224906 207815 224909
rect 193140 224904 207815 224906
rect 193140 224848 207754 224904
rect 207810 224848 207815 224904
rect 193140 224846 207815 224848
rect 193140 224844 193146 224846
rect 207749 224843 207815 224846
rect 194358 224708 194364 224772
rect 194428 224770 194434 224772
rect 208853 224770 208919 224773
rect 194428 224768 208919 224770
rect 194428 224712 208858 224768
rect 208914 224712 208919 224768
rect 194428 224710 208919 224712
rect 194428 224708 194434 224710
rect 208853 224707 208919 224710
rect 191598 224572 191604 224636
rect 191668 224634 191674 224636
rect 206645 224634 206711 224637
rect 191668 224632 206711 224634
rect 191668 224576 206650 224632
rect 206706 224576 206711 224632
rect 191668 224574 206711 224576
rect 191668 224572 191674 224574
rect 206645 224571 206711 224574
rect 190126 224436 190132 224500
rect 190196 224498 190202 224500
rect 204529 224498 204595 224501
rect 190196 224496 204595 224498
rect 190196 224440 204534 224496
rect 204590 224440 204595 224496
rect 190196 224438 204595 224440
rect 190196 224436 190202 224438
rect 204529 224435 204595 224438
rect 190310 224300 190316 224364
rect 190380 224362 190386 224364
rect 205633 224362 205699 224365
rect 190380 224360 205699 224362
rect 190380 224304 205638 224360
rect 205694 224304 205699 224360
rect 190380 224302 205699 224304
rect 190380 224300 190386 224302
rect 205633 224299 205699 224302
rect 194174 224164 194180 224228
rect 194244 224226 194250 224228
rect 209865 224226 209931 224229
rect 194244 224224 209931 224226
rect 194244 224168 209870 224224
rect 209926 224168 209931 224224
rect 194244 224166 209931 224168
rect 194244 224164 194250 224166
rect 209865 224163 209931 224166
rect -960 222594 480 222684
rect 2773 222594 2839 222597
rect -960 222592 2839 222594
rect -960 222536 2778 222592
rect 2834 222536 2839 222592
rect -960 222534 2839 222536
rect -960 222444 480 222534
rect 2773 222531 2839 222534
rect 215109 221370 215175 221373
rect 211508 221368 215175 221370
rect 211508 221312 215114 221368
rect 215170 221312 215175 221368
rect 211508 221310 215175 221312
rect 215109 221307 215175 221310
rect 227621 221370 227687 221373
rect 227621 221368 230092 221370
rect 227621 221312 227626 221368
rect 227682 221312 230092 221368
rect 227621 221310 230092 221312
rect 227621 221307 227687 221310
rect 116393 221234 116459 221237
rect 116393 221232 119692 221234
rect 116393 221176 116398 221232
rect 116454 221176 119692 221232
rect 116393 221174 119692 221176
rect 116393 221171 116459 221174
rect 226333 220826 226399 220829
rect 226333 220824 230092 220826
rect 226333 220768 226338 220824
rect 226394 220768 230092 220824
rect 226333 220766 230092 220768
rect 226333 220763 226399 220766
rect 215201 220554 215267 220557
rect 211508 220552 215267 220554
rect 211508 220496 215206 220552
rect 215262 220496 215267 220552
rect 211508 220494 215267 220496
rect 215201 220491 215267 220494
rect 226333 220146 226399 220149
rect 226333 220144 230092 220146
rect 226333 220088 226338 220144
rect 226394 220088 230092 220144
rect 226333 220086 230092 220088
rect 226333 220083 226399 220086
rect 116117 220010 116183 220013
rect 116117 220008 119692 220010
rect 116117 219952 116122 220008
rect 116178 219952 119692 220008
rect 116117 219950 119692 219952
rect 116117 219947 116183 219950
rect 215109 219738 215175 219741
rect 211508 219736 215175 219738
rect 211508 219680 215114 219736
rect 215170 219680 215175 219736
rect 211508 219678 215175 219680
rect 215109 219675 215175 219678
rect 226425 219602 226491 219605
rect 226425 219600 230092 219602
rect 226425 219544 226430 219600
rect 226486 219544 230092 219600
rect 226425 219542 230092 219544
rect 226425 219539 226491 219542
rect 104801 219330 104867 219333
rect 101078 219328 104867 219330
rect 101078 219272 104806 219328
rect 104862 219272 104867 219328
rect 101078 219270 104867 219272
rect 101078 219096 101138 219270
rect 104801 219267 104867 219270
rect 226333 219058 226399 219061
rect 226333 219056 230092 219058
rect 226333 219000 226338 219056
rect 226394 219000 230092 219056
rect 226333 218998 230092 219000
rect 226333 218995 226399 218998
rect 116393 218922 116459 218925
rect 215109 218922 215175 218925
rect 116393 218920 119692 218922
rect 116393 218864 116398 218920
rect 116454 218864 119692 218920
rect 116393 218862 119692 218864
rect 211508 218920 215175 218922
rect 211508 218864 215114 218920
rect 215170 218864 215175 218920
rect 211508 218862 215175 218864
rect 116393 218859 116459 218862
rect 215109 218859 215175 218862
rect 226425 218378 226491 218381
rect 226425 218376 230092 218378
rect 226425 218320 226430 218376
rect 226486 218320 230092 218376
rect 226425 218318 230092 218320
rect 226425 218315 226491 218318
rect 215201 218242 215267 218245
rect 211508 218240 215267 218242
rect 211508 218184 215206 218240
rect 215262 218184 215267 218240
rect 211508 218182 215267 218184
rect 215201 218179 215267 218182
rect 104801 217970 104867 217973
rect 101078 217968 104867 217970
rect 101078 217912 104806 217968
rect 104862 217912 104867 217968
rect 101078 217910 104867 217912
rect 101078 217872 101138 217910
rect 104801 217907 104867 217910
rect 226333 217834 226399 217837
rect 226333 217832 230092 217834
rect 226333 217776 226338 217832
rect 226394 217776 230092 217832
rect 226333 217774 230092 217776
rect 226333 217771 226399 217774
rect 116393 217698 116459 217701
rect 116393 217696 119692 217698
rect 116393 217640 116398 217696
rect 116454 217640 119692 217696
rect 116393 217638 119692 217640
rect 116393 217635 116459 217638
rect 215109 217426 215175 217429
rect 211508 217424 215175 217426
rect 211508 217368 215114 217424
rect 215170 217368 215175 217424
rect 211508 217366 215175 217368
rect 215109 217363 215175 217366
rect 226425 217290 226491 217293
rect 226425 217288 230092 217290
rect 226425 217232 226430 217288
rect 226486 217232 230092 217288
rect 226425 217230 230092 217232
rect 226425 217227 226491 217230
rect 580901 217018 580967 217021
rect 583520 217018 584960 217108
rect 580901 217016 584960 217018
rect 580901 216960 580906 217016
rect 580962 216960 584960 217016
rect 580901 216958 584960 216960
rect 580901 216955 580967 216958
rect 583520 216868 584960 216958
rect 101078 216610 101138 216648
rect 104801 216610 104867 216613
rect 101078 216608 104867 216610
rect 101078 216552 104806 216608
rect 104862 216552 104867 216608
rect 101078 216550 104867 216552
rect 104801 216547 104867 216550
rect 115933 216610 115999 216613
rect 215109 216610 215175 216613
rect 115933 216608 119692 216610
rect 115933 216552 115938 216608
rect 115994 216552 119692 216608
rect 115933 216550 119692 216552
rect 211508 216608 215175 216610
rect 211508 216552 215114 216608
rect 215170 216552 215175 216608
rect 211508 216550 215175 216552
rect 115933 216547 115999 216550
rect 215109 216547 215175 216550
rect 226333 216610 226399 216613
rect 226333 216608 230092 216610
rect 226333 216552 226338 216608
rect 226394 216552 230092 216608
rect 226333 216550 230092 216552
rect 226333 216547 226399 216550
rect 226425 216066 226491 216069
rect 226425 216064 230092 216066
rect 226425 216008 226430 216064
rect 226486 216008 230092 216064
rect 226425 216006 230092 216008
rect 226425 216003 226491 216006
rect 215109 215794 215175 215797
rect 211508 215792 215175 215794
rect 211508 215736 215114 215792
rect 215170 215736 215175 215792
rect 211508 215734 215175 215736
rect 215109 215731 215175 215734
rect 104801 215658 104867 215661
rect 101078 215656 104867 215658
rect 101078 215600 104806 215656
rect 104862 215600 104867 215656
rect 101078 215598 104867 215600
rect 101078 215424 101138 215598
rect 104801 215595 104867 215598
rect 226333 215522 226399 215525
rect 226333 215520 230092 215522
rect 226333 215464 226338 215520
rect 226394 215464 230092 215520
rect 226333 215462 230092 215464
rect 226333 215459 226399 215462
rect 116393 215386 116459 215389
rect 116393 215384 119692 215386
rect 116393 215328 116398 215384
rect 116454 215328 119692 215384
rect 116393 215326 119692 215328
rect 116393 215323 116459 215326
rect 215109 215114 215175 215117
rect 211508 215112 215175 215114
rect 211508 215056 215114 215112
rect 215170 215056 215175 215112
rect 211508 215054 215175 215056
rect 215109 215051 215175 215054
rect 226425 214842 226491 214845
rect 226425 214840 230092 214842
rect 226425 214784 226430 214840
rect 226486 214784 230092 214840
rect 226425 214782 230092 214784
rect 226425 214779 226491 214782
rect 104801 214706 104867 214709
rect 101078 214704 104867 214706
rect 101078 214648 104806 214704
rect 104862 214648 104867 214704
rect 101078 214646 104867 214648
rect 101078 214200 101138 214646
rect 104801 214643 104867 214646
rect 215201 214298 215267 214301
rect 211508 214296 215267 214298
rect 211508 214240 215206 214296
rect 215262 214240 215267 214296
rect 211508 214238 215267 214240
rect 215201 214235 215267 214238
rect 226333 214298 226399 214301
rect 226333 214296 230092 214298
rect 226333 214240 226338 214296
rect 226394 214240 230092 214296
rect 226333 214238 230092 214240
rect 226333 214235 226399 214238
rect 116393 214162 116459 214165
rect 116393 214160 119692 214162
rect 116393 214104 116398 214160
rect 116454 214104 119692 214160
rect 116393 214102 119692 214104
rect 116393 214099 116459 214102
rect 226425 213618 226491 213621
rect 226425 213616 230092 213618
rect 226425 213560 226430 213616
rect 226486 213560 230092 213616
rect 226425 213558 230092 213560
rect 226425 213555 226491 213558
rect 104801 213482 104867 213485
rect 215109 213482 215175 213485
rect 101078 213480 104867 213482
rect 101078 213424 104806 213480
rect 104862 213424 104867 213480
rect 101078 213422 104867 213424
rect 211508 213480 215175 213482
rect 211508 213424 215114 213480
rect 215170 213424 215175 213480
rect 211508 213422 215175 213424
rect 101078 212976 101138 213422
rect 104801 213419 104867 213422
rect 215109 213419 215175 213422
rect 115933 213074 115999 213077
rect 226333 213074 226399 213077
rect 115933 213072 119692 213074
rect 115933 213016 115938 213072
rect 115994 213016 119692 213072
rect 115933 213014 119692 213016
rect 226333 213072 230092 213074
rect 226333 213016 226338 213072
rect 226394 213016 230092 213072
rect 226333 213014 230092 213016
rect 115933 213011 115999 213014
rect 226333 213011 226399 213014
rect 214373 212666 214439 212669
rect 211508 212664 214439 212666
rect 211508 212608 214378 212664
rect 214434 212608 214439 212664
rect 211508 212606 214439 212608
rect 214373 212603 214439 212606
rect 226517 212530 226583 212533
rect 226517 212528 230092 212530
rect 226517 212472 226522 212528
rect 226578 212472 230092 212528
rect 226517 212470 230092 212472
rect 226517 212467 226583 212470
rect 104433 212122 104499 212125
rect 101078 212120 104499 212122
rect 101078 212064 104438 212120
rect 104494 212064 104499 212120
rect 101078 212062 104499 212064
rect 101078 211752 101138 212062
rect 104433 212059 104499 212062
rect 215109 211986 215175 211989
rect 211508 211984 215175 211986
rect 211508 211928 215114 211984
rect 215170 211928 215175 211984
rect 211508 211926 215175 211928
rect 215109 211923 215175 211926
rect 116301 211850 116367 211853
rect 226149 211850 226215 211853
rect 116301 211848 119692 211850
rect 116301 211792 116306 211848
rect 116362 211792 119692 211848
rect 116301 211790 119692 211792
rect 226149 211848 230092 211850
rect 226149 211792 226154 211848
rect 226210 211792 230092 211848
rect 226149 211790 230092 211792
rect 116301 211787 116367 211790
rect 226149 211787 226215 211790
rect 226241 211306 226307 211309
rect 226241 211304 230092 211306
rect 226241 211248 226246 211304
rect 226302 211248 230092 211304
rect 226241 211246 230092 211248
rect 226241 211243 226307 211246
rect 215201 211170 215267 211173
rect 211508 211168 215267 211170
rect 211508 211112 215206 211168
rect 215262 211112 215267 211168
rect 211508 211110 215267 211112
rect 215201 211107 215267 211110
rect 104801 210898 104867 210901
rect 101078 210896 104867 210898
rect 101078 210840 104806 210896
rect 104862 210840 104867 210896
rect 101078 210838 104867 210840
rect 101078 210528 101138 210838
rect 104801 210835 104867 210838
rect 116301 210762 116367 210765
rect 226057 210762 226123 210765
rect 116301 210760 119692 210762
rect 116301 210704 116306 210760
rect 116362 210704 119692 210760
rect 116301 210702 119692 210704
rect 226057 210760 230092 210762
rect 226057 210704 226062 210760
rect 226118 210704 230092 210760
rect 226057 210702 230092 210704
rect 116301 210699 116367 210702
rect 226057 210699 226123 210702
rect 214189 210354 214255 210357
rect 211508 210352 214255 210354
rect 211508 210296 214194 210352
rect 214250 210296 214255 210352
rect 211508 210294 214255 210296
rect 214189 210291 214255 210294
rect 225965 210082 226031 210085
rect 225965 210080 230092 210082
rect 225965 210024 225970 210080
rect 226026 210024 230092 210080
rect 225965 210022 230092 210024
rect 225965 210019 226031 210022
rect 104801 209538 104867 209541
rect 101078 209536 104867 209538
rect 101078 209480 104806 209536
rect 104862 209480 104867 209536
rect 101078 209478 104867 209480
rect 101078 209304 101138 209478
rect 104801 209475 104867 209478
rect 116025 209538 116091 209541
rect 215109 209538 215175 209541
rect 116025 209536 119692 209538
rect 116025 209480 116030 209536
rect 116086 209480 119692 209536
rect 116025 209478 119692 209480
rect 211508 209536 215175 209538
rect 211508 209480 215114 209536
rect 215170 209480 215175 209536
rect 211508 209478 215175 209480
rect 116025 209475 116091 209478
rect 215109 209475 215175 209478
rect 226149 209538 226215 209541
rect 226149 209536 230092 209538
rect 226149 209480 226154 209536
rect 226210 209480 230092 209536
rect 226149 209478 230092 209480
rect 226149 209475 226215 209478
rect 226241 208994 226307 208997
rect 226241 208992 230092 208994
rect 226241 208936 226246 208992
rect 226302 208936 230092 208992
rect 226241 208934 230092 208936
rect 226241 208931 226307 208934
rect 214189 208858 214255 208861
rect 211508 208856 214255 208858
rect 211508 208800 214194 208856
rect 214250 208800 214255 208856
rect 211508 208798 214255 208800
rect 214189 208795 214255 208798
rect 115933 208314 115999 208317
rect 115933 208312 119692 208314
rect -960 208028 480 208268
rect 115933 208256 115938 208312
rect 115994 208256 119692 208312
rect 115933 208254 119692 208256
rect 115933 208251 115999 208254
rect 104801 208178 104867 208181
rect 101078 208176 104867 208178
rect 101078 208120 104806 208176
rect 104862 208120 104867 208176
rect 101078 208118 104867 208120
rect 101078 208080 101138 208118
rect 104801 208115 104867 208118
rect 215109 208042 215175 208045
rect 211508 208040 215175 208042
rect 211508 207984 215114 208040
rect 215170 207984 215175 208040
rect 211508 207982 215175 207984
rect 215109 207979 215175 207982
rect 226149 208042 226215 208045
rect 230062 208042 230122 208284
rect 226149 208040 230122 208042
rect 226149 207984 226154 208040
rect 226210 207984 230122 208040
rect 226149 207982 230122 207984
rect 226149 207979 226215 207982
rect 225873 207770 225939 207773
rect 225873 207768 230092 207770
rect 225873 207712 225878 207768
rect 225934 207712 230092 207768
rect 225873 207710 230092 207712
rect 225873 207707 225939 207710
rect 116025 207226 116091 207229
rect 214281 207226 214347 207229
rect 116025 207224 119692 207226
rect 116025 207168 116030 207224
rect 116086 207168 119692 207224
rect 116025 207166 119692 207168
rect 211508 207224 214347 207226
rect 211508 207168 214286 207224
rect 214342 207168 214347 207224
rect 211508 207166 214347 207168
rect 116025 207163 116091 207166
rect 214281 207163 214347 207166
rect 225965 207226 226031 207229
rect 225965 207224 230092 207226
rect 225965 207168 225970 207224
rect 226026 207168 230092 207224
rect 225965 207166 230092 207168
rect 225965 207163 226031 207166
rect 104801 206954 104867 206957
rect 101078 206952 104867 206954
rect 101078 206896 104806 206952
rect 104862 206896 104867 206952
rect 101078 206894 104867 206896
rect 101078 206856 101138 206894
rect 104801 206891 104867 206894
rect 225781 206546 225847 206549
rect 225781 206544 230092 206546
rect 225781 206488 225786 206544
rect 225842 206488 230092 206544
rect 225781 206486 230092 206488
rect 225781 206483 225847 206486
rect 215109 206410 215175 206413
rect 211508 206408 215175 206410
rect 211508 206352 215114 206408
rect 215170 206352 215175 206408
rect 211508 206350 215175 206352
rect 215109 206347 215175 206350
rect 104709 206274 104775 206277
rect 101078 206272 104775 206274
rect 101078 206216 104714 206272
rect 104770 206216 104775 206272
rect 101078 206214 104775 206216
rect 101078 205632 101138 206214
rect 104709 206211 104775 206214
rect 115933 206002 115999 206005
rect 226057 206002 226123 206005
rect 115933 206000 119692 206002
rect 115933 205944 115938 206000
rect 115994 205944 119692 206000
rect 115933 205942 119692 205944
rect 226057 206000 230092 206002
rect 226057 205944 226062 206000
rect 226118 205944 230092 206000
rect 226057 205942 230092 205944
rect 115933 205939 115999 205942
rect 226057 205939 226123 205942
rect 214373 205730 214439 205733
rect 211508 205728 214439 205730
rect 211508 205672 214378 205728
rect 214434 205672 214439 205728
rect 211508 205670 214439 205672
rect 214373 205667 214439 205670
rect 225597 205322 225663 205325
rect 225597 205320 230092 205322
rect 225597 205264 225602 205320
rect 225658 205264 230092 205320
rect 225597 205262 230092 205264
rect 225597 205259 225663 205262
rect 583520 205172 584960 205412
rect 104801 205050 104867 205053
rect 101078 205048 104867 205050
rect 101078 204992 104806 205048
rect 104862 204992 104867 205048
rect 101078 204990 104867 204992
rect 101078 204408 101138 204990
rect 104801 204987 104867 204990
rect 116393 204914 116459 204917
rect 215109 204914 215175 204917
rect 116393 204912 119692 204914
rect 116393 204856 116398 204912
rect 116454 204856 119692 204912
rect 116393 204854 119692 204856
rect 211508 204912 215175 204914
rect 211508 204856 215114 204912
rect 215170 204856 215175 204912
rect 211508 204854 215175 204856
rect 116393 204851 116459 204854
rect 215109 204851 215175 204854
rect 226149 204778 226215 204781
rect 226149 204776 230092 204778
rect 226149 204720 226154 204776
rect 226210 204720 230092 204776
rect 226149 204718 230092 204720
rect 226149 204715 226215 204718
rect 226241 204234 226307 204237
rect 226241 204232 230092 204234
rect 226241 204176 226246 204232
rect 226302 204176 230092 204232
rect 226241 204174 230092 204176
rect 226241 204171 226307 204174
rect 215109 204098 215175 204101
rect 211508 204096 215175 204098
rect 211508 204040 215114 204096
rect 215170 204040 215175 204096
rect 211508 204038 215175 204040
rect 215109 204035 215175 204038
rect 104801 203690 104867 203693
rect 101078 203688 104867 203690
rect 101078 203632 104806 203688
rect 104862 203632 104867 203688
rect 101078 203630 104867 203632
rect 101078 203184 101138 203630
rect 104801 203627 104867 203630
rect 116301 203690 116367 203693
rect 116301 203688 119692 203690
rect 116301 203632 116306 203688
rect 116362 203632 119692 203688
rect 116301 203630 119692 203632
rect 116301 203627 116367 203630
rect 225965 203554 226031 203557
rect 225965 203552 230092 203554
rect 225965 203496 225970 203552
rect 226026 203496 230092 203552
rect 225965 203494 230092 203496
rect 225965 203491 226031 203494
rect 215201 203282 215267 203285
rect 211508 203280 215267 203282
rect 211508 203224 215206 203280
rect 215262 203224 215267 203280
rect 211508 203222 215267 203224
rect 215201 203219 215267 203222
rect 225689 203010 225755 203013
rect 225689 203008 230092 203010
rect 225689 202952 225694 203008
rect 225750 202952 230092 203008
rect 225689 202950 230092 202952
rect 225689 202947 225755 202950
rect 104801 202466 104867 202469
rect 101078 202464 104867 202466
rect 101078 202408 104806 202464
rect 104862 202408 104867 202464
rect 101078 202406 104867 202408
rect 101078 201960 101138 202406
rect 104801 202403 104867 202406
rect 116117 202466 116183 202469
rect 215109 202466 215175 202469
rect 116117 202464 119692 202466
rect 116117 202408 116122 202464
rect 116178 202408 119692 202464
rect 116117 202406 119692 202408
rect 211508 202464 215175 202466
rect 211508 202408 215114 202464
rect 215170 202408 215175 202464
rect 211508 202406 215175 202408
rect 116117 202403 116183 202406
rect 215109 202403 215175 202406
rect 225873 202466 225939 202469
rect 225873 202464 230092 202466
rect 225873 202408 225878 202464
rect 225934 202408 230092 202464
rect 225873 202406 230092 202408
rect 225873 202403 225939 202406
rect 214281 201786 214347 201789
rect 211508 201784 214347 201786
rect 211508 201728 214286 201784
rect 214342 201728 214347 201784
rect 211508 201726 214347 201728
rect 214281 201723 214347 201726
rect 226149 201786 226215 201789
rect 226149 201784 230092 201786
rect 226149 201728 226154 201784
rect 226210 201728 230092 201784
rect 226149 201726 230092 201728
rect 226149 201723 226215 201726
rect 116117 201378 116183 201381
rect 116117 201376 119692 201378
rect 116117 201320 116122 201376
rect 116178 201320 119692 201376
rect 116117 201318 119692 201320
rect 116117 201315 116183 201318
rect 226333 201242 226399 201245
rect 226333 201240 230092 201242
rect 226333 201184 226338 201240
rect 226394 201184 230092 201240
rect 226333 201182 230092 201184
rect 226333 201179 226399 201182
rect 104801 201106 104867 201109
rect 101078 201104 104867 201106
rect 101078 201048 104806 201104
rect 104862 201048 104867 201104
rect 101078 201046 104867 201048
rect 101078 200736 101138 201046
rect 104801 201043 104867 201046
rect 214373 200970 214439 200973
rect 211508 200968 214439 200970
rect 211508 200912 214378 200968
rect 214434 200912 214439 200968
rect 211508 200910 214439 200912
rect 214373 200907 214439 200910
rect 226057 200698 226123 200701
rect 226057 200696 230092 200698
rect 226057 200640 226062 200696
rect 226118 200640 230092 200696
rect 226057 200638 230092 200640
rect 226057 200635 226123 200638
rect 115933 200154 115999 200157
rect 215109 200154 215175 200157
rect 115933 200152 119692 200154
rect 115933 200096 115938 200152
rect 115994 200096 119692 200152
rect 115933 200094 119692 200096
rect 211508 200152 215175 200154
rect 211508 200096 215114 200152
rect 215170 200096 215175 200152
rect 211508 200094 215175 200096
rect 115933 200091 115999 200094
rect 215109 200091 215175 200094
rect 225781 200018 225847 200021
rect 225781 200016 230092 200018
rect 225781 199960 225786 200016
rect 225842 199960 230092 200016
rect 225781 199958 230092 199960
rect 225781 199955 225847 199958
rect 104801 199882 104867 199885
rect 101078 199880 104867 199882
rect 101078 199824 104806 199880
rect 104862 199824 104867 199880
rect 101078 199822 104867 199824
rect 101078 199512 101138 199822
rect 104801 199819 104867 199822
rect 226425 199474 226491 199477
rect 226425 199472 230092 199474
rect 226425 199416 226430 199472
rect 226486 199416 230092 199472
rect 226425 199414 230092 199416
rect 226425 199411 226491 199414
rect 214097 199338 214163 199341
rect 211508 199336 214163 199338
rect 211508 199280 214102 199336
rect 214158 199280 214163 199336
rect 211508 199278 214163 199280
rect 214097 199275 214163 199278
rect 116393 199066 116459 199069
rect 116393 199064 119692 199066
rect 116393 199008 116398 199064
rect 116454 199008 119692 199064
rect 116393 199006 119692 199008
rect 116393 199003 116459 199006
rect 226333 198930 226399 198933
rect 226333 198928 230092 198930
rect 226333 198872 226338 198928
rect 226394 198872 230092 198928
rect 226333 198870 230092 198872
rect 226333 198867 226399 198870
rect 215109 198658 215175 198661
rect 338113 198658 338179 198661
rect 211508 198656 215175 198658
rect 211508 198600 215114 198656
rect 215170 198600 215175 198656
rect 211508 198598 215175 198600
rect 336628 198656 338179 198658
rect 336628 198600 338118 198656
rect 338174 198600 338179 198656
rect 336628 198598 338179 198600
rect 215109 198595 215175 198598
rect 338113 198595 338179 198598
rect 104801 198522 104867 198525
rect 101078 198520 104867 198522
rect 101078 198464 104806 198520
rect 104862 198464 104867 198520
rect 101078 198462 104867 198464
rect 101078 198288 101138 198462
rect 104801 198459 104867 198462
rect 226425 198250 226491 198253
rect 226425 198248 230092 198250
rect 226425 198192 226430 198248
rect 226486 198192 230092 198248
rect 226425 198190 230092 198192
rect 226425 198187 226491 198190
rect 116393 197842 116459 197845
rect 214097 197842 214163 197845
rect 116393 197840 119692 197842
rect 116393 197784 116398 197840
rect 116454 197784 119692 197840
rect 116393 197782 119692 197784
rect 211508 197840 214163 197842
rect 211508 197784 214102 197840
rect 214158 197784 214163 197840
rect 211508 197782 214163 197784
rect 116393 197779 116459 197782
rect 214097 197779 214163 197782
rect 226333 197706 226399 197709
rect 226333 197704 230092 197706
rect 226333 197648 226338 197704
rect 226394 197648 230092 197704
rect 226333 197646 230092 197648
rect 226333 197643 226399 197646
rect 104801 197298 104867 197301
rect 101078 197296 104867 197298
rect 101078 197240 104806 197296
rect 104862 197240 104867 197296
rect 101078 197238 104867 197240
rect 101078 197200 101138 197238
rect 104801 197235 104867 197238
rect 215109 197026 215175 197029
rect 211508 197024 215175 197026
rect 211508 196968 215114 197024
rect 215170 196968 215175 197024
rect 211508 196966 215175 196968
rect 215109 196963 215175 196966
rect 226609 197026 226675 197029
rect 226609 197024 230092 197026
rect 226609 196968 226614 197024
rect 226670 196968 230092 197024
rect 226609 196966 230092 196968
rect 226609 196963 226675 196966
rect 116393 196754 116459 196757
rect 116393 196752 119692 196754
rect 116393 196696 116398 196752
rect 116454 196696 119692 196752
rect 116393 196694 119692 196696
rect 116393 196691 116459 196694
rect 104525 196618 104591 196621
rect 101078 196616 104591 196618
rect 101078 196560 104530 196616
rect 104586 196560 104591 196616
rect 101078 196558 104591 196560
rect 101078 195976 101138 196558
rect 104525 196555 104591 196558
rect 226701 196482 226767 196485
rect 226701 196480 230092 196482
rect 226701 196424 226706 196480
rect 226762 196424 230092 196480
rect 226701 196422 230092 196424
rect 226701 196419 226767 196422
rect 214373 196210 214439 196213
rect 211508 196208 214439 196210
rect 211508 196152 214378 196208
rect 214434 196152 214439 196208
rect 211508 196150 214439 196152
rect 214373 196147 214439 196150
rect 226333 195938 226399 195941
rect 226333 195936 230092 195938
rect 226333 195880 226338 195936
rect 226394 195880 230092 195936
rect 226333 195878 230092 195880
rect 226333 195875 226399 195878
rect 115933 195530 115999 195533
rect 215109 195530 215175 195533
rect 115933 195528 119692 195530
rect 115933 195472 115938 195528
rect 115994 195472 119692 195528
rect 115933 195470 119692 195472
rect 211508 195528 215175 195530
rect 211508 195472 215114 195528
rect 215170 195472 215175 195528
rect 211508 195470 215175 195472
rect 115933 195467 115999 195470
rect 215109 195467 215175 195470
rect 104801 195394 104867 195397
rect 101078 195392 104867 195394
rect 101078 195336 104806 195392
rect 104862 195336 104867 195392
rect 101078 195334 104867 195336
rect 101078 194752 101138 195334
rect 104801 195331 104867 195334
rect 226609 195258 226675 195261
rect 226609 195256 230092 195258
rect 226609 195200 226614 195256
rect 226670 195200 230092 195256
rect 226609 195198 230092 195200
rect 226609 195195 226675 195198
rect 215201 194714 215267 194717
rect 211508 194712 215267 194714
rect 211508 194656 215206 194712
rect 215262 194656 215267 194712
rect 211508 194654 215267 194656
rect 215201 194651 215267 194654
rect 226977 194714 227043 194717
rect 226977 194712 230092 194714
rect 226977 194656 226982 194712
rect 227038 194656 230092 194712
rect 226977 194654 230092 194656
rect 226977 194651 227043 194654
rect 116117 194306 116183 194309
rect 116117 194304 119692 194306
rect 116117 194248 116122 194304
rect 116178 194248 119692 194304
rect 116117 194246 119692 194248
rect 116117 194243 116183 194246
rect 226425 194170 226491 194173
rect 226425 194168 230092 194170
rect 226425 194112 226430 194168
rect 226486 194112 230092 194168
rect 226425 194110 230092 194112
rect 226425 194107 226491 194110
rect 104801 194034 104867 194037
rect 101078 194032 104867 194034
rect -960 193898 480 193988
rect 101078 193976 104806 194032
rect 104862 193976 104867 194032
rect 101078 193974 104867 193976
rect 2773 193898 2839 193901
rect -960 193896 2839 193898
rect -960 193840 2778 193896
rect 2834 193840 2839 193896
rect -960 193838 2839 193840
rect -960 193748 480 193838
rect 2773 193835 2839 193838
rect 101078 193528 101138 193974
rect 104801 193971 104867 193974
rect 215109 193898 215175 193901
rect 211508 193896 215175 193898
rect 211508 193840 215114 193896
rect 215170 193840 215175 193896
rect 211508 193838 215175 193840
rect 215109 193835 215175 193838
rect 226333 193490 226399 193493
rect 226333 193488 230092 193490
rect 226333 193432 226338 193488
rect 226394 193432 230092 193488
rect 583520 193476 584960 193716
rect 226333 193430 230092 193432
rect 226333 193427 226399 193430
rect 116393 193218 116459 193221
rect 116393 193216 119692 193218
rect 116393 193160 116398 193216
rect 116454 193160 119692 193216
rect 116393 193158 119692 193160
rect 116393 193155 116459 193158
rect 215109 193082 215175 193085
rect 211508 193080 215175 193082
rect 211508 193024 215114 193080
rect 215170 193024 215175 193080
rect 211508 193022 215175 193024
rect 215109 193019 215175 193022
rect 226425 192946 226491 192949
rect 226425 192944 230092 192946
rect 226425 192888 226430 192944
rect 226486 192888 230092 192944
rect 226425 192886 230092 192888
rect 226425 192883 226491 192886
rect 104433 192810 104499 192813
rect 101078 192808 104499 192810
rect 101078 192752 104438 192808
rect 104494 192752 104499 192808
rect 101078 192750 104499 192752
rect 101078 192304 101138 192750
rect 104433 192747 104499 192750
rect 215201 192402 215267 192405
rect 211508 192400 215267 192402
rect 211508 192344 215206 192400
rect 215262 192344 215267 192400
rect 211508 192342 215267 192344
rect 215201 192339 215267 192342
rect 226333 192402 226399 192405
rect 226333 192400 230092 192402
rect 226333 192344 226338 192400
rect 226394 192344 230092 192400
rect 226333 192342 230092 192344
rect 226333 192339 226399 192342
rect 116025 191994 116091 191997
rect 116025 191992 119692 191994
rect 116025 191936 116030 191992
rect 116086 191936 119692 191992
rect 116025 191934 119692 191936
rect 116025 191931 116091 191934
rect 226333 191722 226399 191725
rect 226333 191720 230092 191722
rect 226333 191664 226338 191720
rect 226394 191664 230092 191720
rect 226333 191662 230092 191664
rect 226333 191659 226399 191662
rect 215109 191586 215175 191589
rect 211508 191584 215175 191586
rect 211508 191528 215114 191584
rect 215170 191528 215175 191584
rect 211508 191526 215175 191528
rect 215109 191523 215175 191526
rect 104801 191450 104867 191453
rect 101078 191448 104867 191450
rect 101078 191392 104806 191448
rect 104862 191392 104867 191448
rect 101078 191390 104867 191392
rect 101078 191080 101138 191390
rect 104801 191387 104867 191390
rect 226517 191178 226583 191181
rect 226517 191176 230092 191178
rect 226517 191120 226522 191176
rect 226578 191120 230092 191176
rect 226517 191118 230092 191120
rect 226517 191115 226583 191118
rect 116485 190906 116551 190909
rect 116485 190904 119692 190906
rect 116485 190848 116490 190904
rect 116546 190848 119692 190904
rect 116485 190846 119692 190848
rect 116485 190843 116551 190846
rect 214281 190770 214347 190773
rect 211508 190768 214347 190770
rect 211508 190712 214286 190768
rect 214342 190712 214347 190768
rect 211508 190710 214347 190712
rect 214281 190707 214347 190710
rect 226333 190498 226399 190501
rect 226333 190496 230092 190498
rect 226333 190440 226338 190496
rect 226394 190440 230092 190496
rect 226333 190438 230092 190440
rect 226333 190435 226399 190438
rect 104709 190226 104775 190229
rect 101078 190224 104775 190226
rect 101078 190168 104714 190224
rect 104770 190168 104775 190224
rect 101078 190166 104775 190168
rect 101078 189856 101138 190166
rect 104709 190163 104775 190166
rect 215109 189954 215175 189957
rect 211508 189952 215175 189954
rect 211508 189896 215114 189952
rect 215170 189896 215175 189952
rect 211508 189894 215175 189896
rect 215109 189891 215175 189894
rect 226333 189954 226399 189957
rect 226333 189952 230092 189954
rect 226333 189896 226338 189952
rect 226394 189896 230092 189952
rect 226333 189894 230092 189896
rect 226333 189891 226399 189894
rect 116393 189682 116459 189685
rect 116393 189680 119692 189682
rect 116393 189624 116398 189680
rect 116454 189624 119692 189680
rect 116393 189622 119692 189624
rect 116393 189619 116459 189622
rect 225781 189410 225847 189413
rect 225781 189408 230092 189410
rect 225781 189352 225786 189408
rect 225842 189352 230092 189408
rect 225781 189350 230092 189352
rect 225781 189347 225847 189350
rect 214373 189274 214439 189277
rect 211508 189272 214439 189274
rect 211508 189216 214378 189272
rect 214434 189216 214439 189272
rect 211508 189214 214439 189216
rect 214373 189211 214439 189214
rect 104801 188866 104867 188869
rect 101078 188864 104867 188866
rect 101078 188808 104806 188864
rect 104862 188808 104867 188864
rect 101078 188806 104867 188808
rect 101078 188632 101138 188806
rect 104801 188803 104867 188806
rect 226333 188730 226399 188733
rect 226333 188728 230092 188730
rect 226333 188672 226338 188728
rect 226394 188672 230092 188728
rect 226333 188670 230092 188672
rect 226333 188667 226399 188670
rect 116209 188458 116275 188461
rect 214005 188458 214071 188461
rect 116209 188456 119692 188458
rect 116209 188400 116214 188456
rect 116270 188400 119692 188456
rect 116209 188398 119692 188400
rect 211508 188456 214071 188458
rect 211508 188400 214010 188456
rect 214066 188400 214071 188456
rect 211508 188398 214071 188400
rect 116209 188395 116275 188398
rect 214005 188395 214071 188398
rect 226425 188186 226491 188189
rect 226425 188184 230092 188186
rect 226425 188128 226430 188184
rect 226486 188128 230092 188184
rect 226425 188126 230092 188128
rect 226425 188123 226491 188126
rect 215201 187642 215267 187645
rect 211508 187640 215267 187642
rect 211508 187584 215206 187640
rect 215262 187584 215267 187640
rect 211508 187582 215267 187584
rect 215201 187579 215267 187582
rect 226333 187642 226399 187645
rect 226333 187640 230092 187642
rect 226333 187584 226338 187640
rect 226394 187584 230092 187640
rect 226333 187582 230092 187584
rect 226333 187579 226399 187582
rect 104801 187506 104867 187509
rect 101078 187504 104867 187506
rect 101078 187448 104806 187504
rect 104862 187448 104867 187504
rect 101078 187446 104867 187448
rect 101078 187408 101138 187446
rect 104801 187443 104867 187446
rect 116301 187370 116367 187373
rect 116301 187368 119692 187370
rect 116301 187312 116306 187368
rect 116362 187312 119692 187368
rect 116301 187310 119692 187312
rect 116301 187307 116367 187310
rect 225597 186962 225663 186965
rect 225597 186960 230092 186962
rect 225597 186904 225602 186960
rect 225658 186904 230092 186960
rect 225597 186902 230092 186904
rect 225597 186899 225663 186902
rect 215201 186826 215267 186829
rect 211508 186824 215267 186826
rect 211508 186768 215206 186824
rect 215262 186768 215267 186824
rect 211508 186766 215267 186768
rect 215201 186763 215267 186766
rect 226333 186418 226399 186421
rect 226333 186416 230092 186418
rect 226333 186360 226338 186416
rect 226394 186360 230092 186416
rect 226333 186358 230092 186360
rect 226333 186355 226399 186358
rect 104801 186282 104867 186285
rect 101078 186280 104867 186282
rect 101078 186224 104806 186280
rect 104862 186224 104867 186280
rect 101078 186222 104867 186224
rect 101078 186184 101138 186222
rect 104801 186219 104867 186222
rect 116025 186146 116091 186149
rect 116025 186144 119692 186146
rect 116025 186088 116030 186144
rect 116086 186088 119692 186144
rect 116025 186086 119692 186088
rect 116025 186083 116091 186086
rect 215109 186010 215175 186013
rect 211508 186008 215175 186010
rect 211508 185952 215114 186008
rect 215170 185952 215175 186008
rect 211508 185950 215175 185952
rect 215109 185947 215175 185950
rect 226333 185874 226399 185877
rect 226333 185872 230092 185874
rect 226333 185816 226338 185872
rect 226394 185816 230092 185872
rect 226333 185814 230092 185816
rect 226333 185811 226399 185814
rect 104525 185602 104591 185605
rect 101078 185600 104591 185602
rect 101078 185544 104530 185600
rect 104586 185544 104591 185600
rect 101078 185542 104591 185544
rect 101078 184960 101138 185542
rect 104525 185539 104591 185542
rect 213913 185330 213979 185333
rect 211508 185328 213979 185330
rect 211508 185272 213918 185328
rect 213974 185272 213979 185328
rect 211508 185270 213979 185272
rect 213913 185267 213979 185270
rect 226977 185194 227043 185197
rect 226977 185192 230092 185194
rect 226977 185136 226982 185192
rect 227038 185136 230092 185192
rect 226977 185134 230092 185136
rect 226977 185131 227043 185134
rect 116393 185058 116459 185061
rect 116393 185056 119692 185058
rect 116393 185000 116398 185056
rect 116454 185000 119692 185056
rect 116393 184998 119692 185000
rect 116393 184995 116459 184998
rect 226333 184650 226399 184653
rect 226333 184648 230092 184650
rect 226333 184592 226338 184648
rect 226394 184592 230092 184648
rect 226333 184590 230092 184592
rect 226333 184587 226399 184590
rect 214465 184514 214531 184517
rect 211508 184512 214531 184514
rect 211508 184456 214470 184512
rect 214526 184456 214531 184512
rect 211508 184454 214531 184456
rect 214465 184451 214531 184454
rect 104801 184378 104867 184381
rect 101078 184376 104867 184378
rect 101078 184320 104806 184376
rect 104862 184320 104867 184376
rect 101078 184318 104867 184320
rect 101078 183736 101138 184318
rect 104801 184315 104867 184318
rect 226517 184106 226583 184109
rect 226517 184104 230092 184106
rect 226517 184048 226522 184104
rect 226578 184048 230092 184104
rect 226517 184046 230092 184048
rect 226517 184043 226583 184046
rect 116393 183834 116459 183837
rect 116393 183832 119692 183834
rect 116393 183776 116398 183832
rect 116454 183776 119692 183832
rect 116393 183774 119692 183776
rect 116393 183771 116459 183774
rect 214189 183698 214255 183701
rect 211508 183696 214255 183698
rect 211508 183640 214194 183696
rect 214250 183640 214255 183696
rect 211508 183638 214255 183640
rect 214189 183635 214255 183638
rect 226517 183426 226583 183429
rect 226517 183424 230092 183426
rect 226517 183368 226522 183424
rect 226578 183368 230092 183424
rect 226517 183366 230092 183368
rect 226517 183363 226583 183366
rect 104801 183018 104867 183021
rect 101078 183016 104867 183018
rect 101078 182960 104806 183016
rect 104862 182960 104867 183016
rect 101078 182958 104867 182960
rect 101078 182512 101138 182958
rect 104801 182955 104867 182958
rect 215109 182882 215175 182885
rect 211508 182880 215175 182882
rect 211508 182824 215114 182880
rect 215170 182824 215175 182880
rect 211508 182822 215175 182824
rect 215109 182819 215175 182822
rect 226425 182882 226491 182885
rect 226425 182880 230092 182882
rect 226425 182824 226430 182880
rect 226486 182824 230092 182880
rect 226425 182822 230092 182824
rect 226425 182819 226491 182822
rect 115933 182610 115999 182613
rect 115933 182608 119692 182610
rect 115933 182552 115938 182608
rect 115994 182552 119692 182608
rect 115933 182550 119692 182552
rect 115933 182547 115999 182550
rect 215201 182202 215267 182205
rect 211508 182200 215267 182202
rect 211508 182144 215206 182200
rect 215262 182144 215267 182200
rect 211508 182142 215267 182144
rect 215201 182139 215267 182142
rect 226333 182202 226399 182205
rect 226333 182200 230092 182202
rect 226333 182144 226338 182200
rect 226394 182144 230092 182200
rect 226333 182142 230092 182144
rect 226333 182139 226399 182142
rect 579981 181930 580047 181933
rect 583520 181930 584960 182020
rect 579981 181928 584960 181930
rect 579981 181872 579986 181928
rect 580042 181872 584960 181928
rect 579981 181870 584960 181872
rect 579981 181867 580047 181870
rect 104801 181794 104867 181797
rect 101078 181792 104867 181794
rect 101078 181736 104806 181792
rect 104862 181736 104867 181792
rect 583520 181780 584960 181870
rect 101078 181734 104867 181736
rect 101078 181288 101138 181734
rect 104801 181731 104867 181734
rect 227621 181658 227687 181661
rect 227621 181656 230092 181658
rect 227621 181600 227626 181656
rect 227682 181600 230092 181656
rect 227621 181598 230092 181600
rect 227621 181595 227687 181598
rect 115933 181522 115999 181525
rect 115933 181520 119692 181522
rect 115933 181464 115938 181520
rect 115994 181464 119692 181520
rect 115933 181462 119692 181464
rect 115933 181459 115999 181462
rect 214189 181386 214255 181389
rect 211508 181384 214255 181386
rect 211508 181328 214194 181384
rect 214250 181328 214255 181384
rect 211508 181326 214255 181328
rect 214189 181323 214255 181326
rect 226333 181114 226399 181117
rect 226333 181112 230092 181114
rect 226333 181056 226338 181112
rect 226394 181056 230092 181112
rect 226333 181054 230092 181056
rect 226333 181051 226399 181054
rect 214097 180570 214163 180573
rect 211508 180568 214163 180570
rect 211508 180512 214102 180568
rect 214158 180512 214163 180568
rect 211508 180510 214163 180512
rect 214097 180507 214163 180510
rect 104801 180434 104867 180437
rect 101078 180432 104867 180434
rect 101078 180376 104806 180432
rect 104862 180376 104867 180432
rect 101078 180374 104867 180376
rect 101078 180064 101138 180374
rect 104801 180371 104867 180374
rect 226333 180434 226399 180437
rect 226333 180432 230092 180434
rect 226333 180376 226338 180432
rect 226394 180376 230092 180432
rect 226333 180374 230092 180376
rect 226333 180371 226399 180374
rect 116393 180298 116459 180301
rect 116393 180296 119692 180298
rect 116393 180240 116398 180296
rect 116454 180240 119692 180296
rect 116393 180238 119692 180240
rect 116393 180235 116459 180238
rect 226425 179890 226491 179893
rect 226425 179888 230092 179890
rect 226425 179832 226430 179888
rect 226486 179832 230092 179888
rect 226425 179830 230092 179832
rect 226425 179827 226491 179830
rect 214005 179754 214071 179757
rect 211508 179752 214071 179754
rect 211508 179696 214010 179752
rect 214066 179696 214071 179752
rect 211508 179694 214071 179696
rect 214005 179691 214071 179694
rect -960 179482 480 179572
rect 2773 179482 2839 179485
rect -960 179480 2839 179482
rect -960 179424 2778 179480
rect 2834 179424 2839 179480
rect -960 179422 2839 179424
rect -960 179332 480 179422
rect 2773 179419 2839 179422
rect 227069 179346 227135 179349
rect 227069 179344 230092 179346
rect 227069 179288 227074 179344
rect 227130 179288 230092 179344
rect 227069 179286 230092 179288
rect 227069 179283 227135 179286
rect 115933 179210 115999 179213
rect 115933 179208 119692 179210
rect 115933 179152 115938 179208
rect 115994 179152 119692 179208
rect 115933 179150 119692 179152
rect 115933 179147 115999 179150
rect 104801 179074 104867 179077
rect 213913 179074 213979 179077
rect 101078 179072 104867 179074
rect 101078 179016 104806 179072
rect 104862 179016 104867 179072
rect 101078 179014 104867 179016
rect 211508 179072 213979 179074
rect 211508 179016 213918 179072
rect 213974 179016 213979 179072
rect 211508 179014 213979 179016
rect 101078 178840 101138 179014
rect 104801 179011 104867 179014
rect 213913 179011 213979 179014
rect 226425 178666 226491 178669
rect 226425 178664 230092 178666
rect 226425 178608 226430 178664
rect 226486 178608 230092 178664
rect 226425 178606 230092 178608
rect 226425 178603 226491 178606
rect 214097 178258 214163 178261
rect 211508 178256 214163 178258
rect 211508 178200 214102 178256
rect 214158 178200 214163 178256
rect 211508 178198 214163 178200
rect 214097 178195 214163 178198
rect 226701 178122 226767 178125
rect 226701 178120 230092 178122
rect 226701 178064 226706 178120
rect 226762 178064 230092 178120
rect 226701 178062 230092 178064
rect 226701 178059 226767 178062
rect 115933 177986 115999 177989
rect 115933 177984 119692 177986
rect 115933 177928 115938 177984
rect 115994 177928 119692 177984
rect 115933 177926 119692 177928
rect 115933 177923 115999 177926
rect 104157 177850 104223 177853
rect 101078 177848 104223 177850
rect 101078 177792 104162 177848
rect 104218 177792 104223 177848
rect 101078 177790 104223 177792
rect 101078 177616 101138 177790
rect 104157 177787 104223 177790
rect 226333 177578 226399 177581
rect 226333 177576 230092 177578
rect 226333 177520 226338 177576
rect 226394 177520 230092 177576
rect 226333 177518 230092 177520
rect 226333 177515 226399 177518
rect 215017 177442 215083 177445
rect 211508 177440 215083 177442
rect 211508 177384 215022 177440
rect 215078 177384 215083 177440
rect 211508 177382 215083 177384
rect 215017 177379 215083 177382
rect 116393 176898 116459 176901
rect 227345 176898 227411 176901
rect 116393 176896 119692 176898
rect 116393 176840 116398 176896
rect 116454 176840 119692 176896
rect 116393 176838 119692 176840
rect 227345 176896 230092 176898
rect 227345 176840 227350 176896
rect 227406 176840 230092 176896
rect 227345 176838 230092 176840
rect 116393 176835 116459 176838
rect 227345 176835 227411 176838
rect 215109 176626 215175 176629
rect 211508 176624 215175 176626
rect 211508 176568 215114 176624
rect 215170 176568 215175 176624
rect 211508 176566 215175 176568
rect 215109 176563 215175 176566
rect 104157 176490 104223 176493
rect 101078 176488 104223 176490
rect 101078 176432 104162 176488
rect 104218 176432 104223 176488
rect 101078 176430 104223 176432
rect 101078 176392 101138 176430
rect 104157 176427 104223 176430
rect 227437 176354 227503 176357
rect 227437 176352 230092 176354
rect 227437 176296 227442 176352
rect 227498 176296 230092 176352
rect 227437 176294 230092 176296
rect 227437 176291 227503 176294
rect 215109 175946 215175 175949
rect 211508 175944 215175 175946
rect 211508 175888 215114 175944
rect 215170 175888 215175 175944
rect 211508 175886 215175 175888
rect 215109 175883 215175 175886
rect 226977 175810 227043 175813
rect 226977 175808 230092 175810
rect 226977 175752 226982 175808
rect 227038 175752 230092 175808
rect 226977 175750 230092 175752
rect 226977 175747 227043 175750
rect 116393 175674 116459 175677
rect 116393 175672 119692 175674
rect 116393 175616 116398 175672
rect 116454 175616 119692 175672
rect 116393 175614 119692 175616
rect 116393 175611 116459 175614
rect 101078 175130 101138 175168
rect 104801 175130 104867 175133
rect 215109 175130 215175 175133
rect 101078 175128 104867 175130
rect 101078 175072 104806 175128
rect 104862 175072 104867 175128
rect 101078 175070 104867 175072
rect 211508 175128 215175 175130
rect 211508 175072 215114 175128
rect 215170 175072 215175 175128
rect 211508 175070 215175 175072
rect 104801 175067 104867 175070
rect 215109 175067 215175 175070
rect 104433 174722 104499 174725
rect 101078 174720 104499 174722
rect 101078 174664 104438 174720
rect 104494 174664 104499 174720
rect 101078 174662 104499 174664
rect 101078 174080 101138 174662
rect 104433 174659 104499 174662
rect 115933 174450 115999 174453
rect 115933 174448 119692 174450
rect 115933 174392 115938 174448
rect 115994 174392 119692 174448
rect 115933 174390 119692 174392
rect 115933 174387 115999 174390
rect 214097 174314 214163 174317
rect 211508 174312 214163 174314
rect 211508 174256 214102 174312
rect 214158 174256 214163 174312
rect 211508 174254 214163 174256
rect 214097 174251 214163 174254
rect 283373 173906 283439 173909
rect 332910 173906 332916 173908
rect 283373 173904 332916 173906
rect 283373 173848 283378 173904
rect 283434 173848 332916 173904
rect 283373 173846 332916 173848
rect 283373 173843 283439 173846
rect 332910 173844 332916 173846
rect 332980 173844 332986 173908
rect 4797 173770 4863 173773
rect 4797 173768 9322 173770
rect 4797 173712 4802 173768
rect 4858 173712 9322 173768
rect 4797 173710 9322 173712
rect 4797 173707 4863 173710
rect 9262 173536 9322 173710
rect 215201 173498 215267 173501
rect 211508 173496 215267 173498
rect 211508 173440 215206 173496
rect 215262 173440 215267 173496
rect 211508 173438 215267 173440
rect 215201 173435 215267 173438
rect 104801 173362 104867 173365
rect 101078 173360 104867 173362
rect 101078 173304 104806 173360
rect 104862 173304 104867 173360
rect 101078 173302 104867 173304
rect 101078 172856 101138 173302
rect 104801 173299 104867 173302
rect 116393 173362 116459 173365
rect 116393 173360 119692 173362
rect 116393 173304 116398 173360
rect 116454 173304 119692 173360
rect 116393 173302 119692 173304
rect 116393 173299 116459 173302
rect 232221 173226 232287 173229
rect 283373 173226 283439 173229
rect 232221 173224 283439 173226
rect 232221 173168 232226 173224
rect 232282 173168 283378 173224
rect 283434 173168 283439 173224
rect 232221 173166 283439 173168
rect 232221 173163 232287 173166
rect 283373 173163 283439 173166
rect 214281 172818 214347 172821
rect 211508 172816 214347 172818
rect 211508 172760 214286 172816
rect 214342 172760 214347 172816
rect 211508 172758 214347 172760
rect 214281 172755 214347 172758
rect 104433 172138 104499 172141
rect 101078 172136 104499 172138
rect 101078 172080 104438 172136
rect 104494 172080 104499 172136
rect 101078 172078 104499 172080
rect 101078 171632 101138 172078
rect 104433 172075 104499 172078
rect 116117 172138 116183 172141
rect 116117 172136 119692 172138
rect 116117 172080 116122 172136
rect 116178 172080 119692 172136
rect 116117 172078 119692 172080
rect 116117 172075 116183 172078
rect 214281 172002 214347 172005
rect 211508 172000 214347 172002
rect 211508 171944 214286 172000
rect 214342 171944 214347 172000
rect 211508 171942 214347 171944
rect 214281 171939 214347 171942
rect 215017 171186 215083 171189
rect 211508 171184 215083 171186
rect 211508 171128 215022 171184
rect 215078 171128 215083 171184
rect 211508 171126 215083 171128
rect 215017 171123 215083 171126
rect 116301 171050 116367 171053
rect 116301 171048 119692 171050
rect 116301 170992 116306 171048
rect 116362 170992 119692 171048
rect 116301 170990 119692 170992
rect 116301 170987 116367 170990
rect 104801 170778 104867 170781
rect 101078 170776 104867 170778
rect 101078 170720 104806 170776
rect 104862 170720 104867 170776
rect 101078 170718 104867 170720
rect 101078 170408 101138 170718
rect 104801 170715 104867 170718
rect 214833 170370 214899 170373
rect 211508 170368 214899 170370
rect 211508 170312 214838 170368
rect 214894 170312 214899 170368
rect 211508 170310 214899 170312
rect 214833 170307 214899 170310
rect 580901 170098 580967 170101
rect 583520 170098 584960 170188
rect 580901 170096 584960 170098
rect 580901 170040 580906 170096
rect 580962 170040 584960 170096
rect 580901 170038 584960 170040
rect 580901 170035 580967 170038
rect 583520 169948 584960 170038
rect 116393 169826 116459 169829
rect 116393 169824 119692 169826
rect 116393 169768 116398 169824
rect 116454 169768 119692 169824
rect 116393 169766 119692 169768
rect 116393 169763 116459 169766
rect 215109 169554 215175 169557
rect 211508 169552 215175 169554
rect 211508 169496 215114 169552
rect 215170 169496 215175 169552
rect 211508 169494 215175 169496
rect 215109 169491 215175 169494
rect 104801 169418 104867 169421
rect 101078 169416 104867 169418
rect 101078 169360 104806 169416
rect 104862 169360 104867 169416
rect 101078 169358 104867 169360
rect 101078 169184 101138 169358
rect 104801 169355 104867 169358
rect 215109 168874 215175 168877
rect 211508 168872 215175 168874
rect 211508 168816 215114 168872
rect 215170 168816 215175 168872
rect 211508 168814 215175 168816
rect 215109 168811 215175 168814
rect 116393 168602 116459 168605
rect 116393 168600 119692 168602
rect 116393 168544 116398 168600
rect 116454 168544 119692 168600
rect 116393 168542 119692 168544
rect 116393 168539 116459 168542
rect 104157 168194 104223 168197
rect 101078 168192 104223 168194
rect 101078 168136 104162 168192
rect 104218 168136 104223 168192
rect 101078 168134 104223 168136
rect 101078 167960 101138 168134
rect 104157 168131 104223 168134
rect 213913 168058 213979 168061
rect 211508 168056 213979 168058
rect 211508 168000 213918 168056
rect 213974 168000 213979 168056
rect 211508 167998 213979 168000
rect 213913 167995 213979 167998
rect 115933 167514 115999 167517
rect 115933 167512 119692 167514
rect 115933 167456 115938 167512
rect 115994 167456 119692 167512
rect 115933 167454 119692 167456
rect 115933 167451 115999 167454
rect 214281 167242 214347 167245
rect 211508 167240 214347 167242
rect 211508 167184 214286 167240
rect 214342 167184 214347 167240
rect 211508 167182 214347 167184
rect 214281 167179 214347 167182
rect 104249 166970 104315 166973
rect 101078 166968 104315 166970
rect 101078 166912 104254 166968
rect 104310 166912 104315 166968
rect 101078 166910 104315 166912
rect 101078 166736 101138 166910
rect 104249 166907 104315 166910
rect 215201 166426 215267 166429
rect 211508 166424 215267 166426
rect 211508 166368 215206 166424
rect 215262 166368 215267 166424
rect 211508 166366 215267 166368
rect 215201 166363 215267 166366
rect 115933 166290 115999 166293
rect 115933 166288 119692 166290
rect 115933 166232 115938 166288
rect 115994 166232 119692 166288
rect 115933 166230 119692 166232
rect 115933 166227 115999 166230
rect 214373 165746 214439 165749
rect 211508 165744 214439 165746
rect 211508 165688 214378 165744
rect 214434 165688 214439 165744
rect 211508 165686 214439 165688
rect 214373 165683 214439 165686
rect 104801 165610 104867 165613
rect 101078 165608 104867 165610
rect 101078 165552 104806 165608
rect 104862 165552 104867 165608
rect 101078 165550 104867 165552
rect 101078 165512 101138 165550
rect 104801 165547 104867 165550
rect 116117 165202 116183 165205
rect 116117 165200 119692 165202
rect -960 164916 480 165156
rect 116117 165144 116122 165200
rect 116178 165144 119692 165200
rect 116117 165142 119692 165144
rect 116117 165139 116183 165142
rect 104617 164930 104683 164933
rect 214097 164930 214163 164933
rect 101078 164928 104683 164930
rect 101078 164872 104622 164928
rect 104678 164872 104683 164928
rect 101078 164870 104683 164872
rect 211508 164928 214163 164930
rect 211508 164872 214102 164928
rect 214158 164872 214163 164928
rect 211508 164870 214163 164872
rect 101078 164288 101138 164870
rect 104617 164867 104683 164870
rect 214097 164867 214163 164870
rect 214925 164114 214991 164117
rect 211508 164112 214991 164114
rect 211508 164056 214930 164112
rect 214986 164056 214991 164112
rect 211508 164054 214991 164056
rect 214925 164051 214991 164054
rect 116393 163978 116459 163981
rect 116393 163976 119692 163978
rect 116393 163920 116398 163976
rect 116454 163920 119692 163976
rect 116393 163918 119692 163920
rect 116393 163915 116459 163918
rect 104801 163706 104867 163709
rect 101078 163704 104867 163706
rect 101078 163648 104806 163704
rect 104862 163648 104867 163704
rect 101078 163646 104867 163648
rect 101078 163064 101138 163646
rect 104801 163643 104867 163646
rect 214373 163298 214439 163301
rect 211508 163296 214439 163298
rect 211508 163240 214378 163296
rect 214434 163240 214439 163296
rect 211508 163238 214439 163240
rect 214373 163235 214439 163238
rect 116209 162754 116275 162757
rect 116209 162752 119692 162754
rect 116209 162696 116214 162752
rect 116270 162696 119692 162752
rect 116209 162694 119692 162696
rect 116209 162691 116275 162694
rect 215109 162618 215175 162621
rect 211508 162616 215175 162618
rect 211508 162560 215114 162616
rect 215170 162560 215175 162616
rect 211508 162558 215175 162560
rect 215109 162555 215175 162558
rect 104801 162346 104867 162349
rect 101078 162344 104867 162346
rect 101078 162288 104806 162344
rect 104862 162288 104867 162344
rect 101078 162286 104867 162288
rect 101078 161840 101138 162286
rect 104801 162283 104867 162286
rect 214281 161802 214347 161805
rect 211508 161800 214347 161802
rect 211508 161744 214286 161800
rect 214342 161744 214347 161800
rect 211508 161742 214347 161744
rect 214281 161739 214347 161742
rect 116393 161666 116459 161669
rect 116393 161664 119692 161666
rect 116393 161608 116398 161664
rect 116454 161608 119692 161664
rect 116393 161606 119692 161608
rect 116393 161603 116459 161606
rect 104801 160986 104867 160989
rect 215109 160986 215175 160989
rect 101078 160984 104867 160986
rect 101078 160928 104806 160984
rect 104862 160928 104867 160984
rect 101078 160926 104867 160928
rect 211508 160984 215175 160986
rect 211508 160928 215114 160984
rect 215170 160928 215175 160984
rect 211508 160926 215175 160928
rect 101078 160616 101138 160926
rect 104801 160923 104867 160926
rect 215109 160923 215175 160926
rect 116393 160442 116459 160445
rect 116393 160440 119692 160442
rect 116393 160384 116398 160440
rect 116454 160384 119692 160440
rect 116393 160382 119692 160384
rect 116393 160379 116459 160382
rect 214925 160170 214991 160173
rect 211508 160168 214991 160170
rect 211508 160112 214930 160168
rect 214986 160112 214991 160168
rect 211508 160110 214991 160112
rect 214925 160107 214991 160110
rect 104801 159762 104867 159765
rect 101078 159760 104867 159762
rect 101078 159704 104806 159760
rect 104862 159704 104867 159760
rect 101078 159702 104867 159704
rect 101078 159392 101138 159702
rect 104801 159699 104867 159702
rect 116393 159354 116459 159357
rect 116393 159352 119692 159354
rect 116393 159296 116398 159352
rect 116454 159296 119692 159352
rect 116393 159294 119692 159296
rect 116393 159291 116459 159294
rect 211478 158946 211538 159460
rect 211478 158886 211722 158946
rect 211662 158810 211722 158886
rect 219934 158810 219940 158812
rect 211662 158750 219940 158810
rect 219934 158748 219940 158750
rect 220004 158748 220010 158812
rect 103697 158674 103763 158677
rect 214833 158674 214899 158677
rect 101078 158672 103763 158674
rect 101078 158616 103702 158672
rect 103758 158616 103763 158672
rect 101078 158614 103763 158616
rect 211508 158672 214899 158674
rect 211508 158616 214838 158672
rect 214894 158616 214899 158672
rect 211508 158614 214899 158616
rect 101078 158168 101138 158614
rect 103697 158611 103763 158614
rect 214833 158611 214899 158614
rect 583520 158252 584960 158492
rect 116393 158130 116459 158133
rect 116393 158128 119692 158130
rect 116393 158072 116398 158128
rect 116454 158072 119692 158128
rect 116393 158070 119692 158072
rect 116393 158067 116459 158070
rect 214741 157858 214807 157861
rect 211508 157856 214807 157858
rect 211508 157800 214746 157856
rect 214802 157800 214807 157856
rect 211508 157798 214807 157800
rect 214741 157795 214807 157798
rect 104249 157314 104315 157317
rect 101078 157312 104315 157314
rect 101078 157256 104254 157312
rect 104310 157256 104315 157312
rect 101078 157254 104315 157256
rect 101078 156944 101138 157254
rect 104249 157251 104315 157254
rect 116025 157042 116091 157045
rect 215109 157042 215175 157045
rect 116025 157040 119692 157042
rect 116025 156984 116030 157040
rect 116086 156984 119692 157040
rect 116025 156982 119692 156984
rect 211508 157040 215175 157042
rect 211508 156984 215114 157040
rect 215170 156984 215175 157040
rect 211508 156982 215175 156984
rect 116025 156979 116091 156982
rect 215109 156979 215175 156982
rect 214741 156362 214807 156365
rect 211508 156360 214807 156362
rect 211508 156304 214746 156360
rect 214802 156304 214807 156360
rect 211508 156302 214807 156304
rect 214741 156299 214807 156302
rect 104801 155954 104867 155957
rect 101078 155952 104867 155954
rect 101078 155896 104806 155952
rect 104862 155896 104867 155952
rect 101078 155894 104867 155896
rect 101078 155720 101138 155894
rect 104801 155891 104867 155894
rect 116025 155818 116091 155821
rect 116025 155816 119692 155818
rect 116025 155760 116030 155816
rect 116086 155760 119692 155816
rect 116025 155758 119692 155760
rect 116025 155755 116091 155758
rect 214373 155546 214439 155549
rect 211508 155544 214439 155546
rect 211508 155488 214378 155544
rect 214434 155488 214439 155544
rect 211508 155486 214439 155488
rect 214373 155483 214439 155486
rect 215109 154730 215175 154733
rect 211508 154728 215175 154730
rect 211508 154672 215114 154728
rect 215170 154672 215175 154728
rect 211508 154670 215175 154672
rect 215109 154667 215175 154670
rect 116393 154594 116459 154597
rect 232313 154594 232379 154597
rect 232497 154594 232563 154597
rect 116393 154592 119692 154594
rect 116393 154536 116398 154592
rect 116454 154536 119692 154592
rect 116393 154534 119692 154536
rect 232313 154592 232563 154594
rect 232313 154536 232318 154592
rect 232374 154536 232502 154592
rect 232558 154536 232563 154592
rect 232313 154534 232563 154536
rect 116393 154531 116459 154534
rect 232313 154531 232379 154534
rect 232497 154531 232563 154534
rect 101078 154458 101138 154496
rect 104341 154458 104407 154461
rect 101078 154456 104407 154458
rect 101078 154400 104346 154456
rect 104402 154400 104407 154456
rect 101078 154398 104407 154400
rect 104341 154395 104407 154398
rect 104617 153914 104683 153917
rect 215201 153914 215267 153917
rect 101078 153912 104683 153914
rect 101078 153856 104622 153912
rect 104678 153856 104683 153912
rect 101078 153854 104683 153856
rect 211508 153912 215267 153914
rect 211508 153856 215206 153912
rect 215262 153856 215267 153912
rect 211508 153854 215267 153856
rect 101078 153272 101138 153854
rect 104617 153851 104683 153854
rect 215201 153851 215267 153854
rect 115933 153506 115999 153509
rect 115933 153504 119692 153506
rect 115933 153448 115938 153504
rect 115994 153448 119692 153504
rect 115933 153446 119692 153448
rect 115933 153443 115999 153446
rect 215109 153234 215175 153237
rect 211508 153232 215175 153234
rect 211508 153176 215114 153232
rect 215170 153176 215175 153232
rect 211508 153174 215175 153176
rect 215109 153171 215175 153174
rect 104801 152690 104867 152693
rect 101078 152688 104867 152690
rect 101078 152632 104806 152688
rect 104862 152632 104867 152688
rect 101078 152630 104867 152632
rect 101078 152048 101138 152630
rect 104801 152627 104867 152630
rect 214005 152418 214071 152421
rect 211508 152416 214071 152418
rect 211508 152360 214010 152416
rect 214066 152360 214071 152416
rect 211508 152358 214071 152360
rect 214005 152355 214071 152358
rect 116393 152282 116459 152285
rect 116393 152280 119692 152282
rect 116393 152224 116398 152280
rect 116454 152224 119692 152280
rect 116393 152222 119692 152224
rect 116393 152219 116459 152222
rect 104157 151602 104223 151605
rect 214373 151602 214439 151605
rect 101078 151600 104223 151602
rect 101078 151544 104162 151600
rect 104218 151544 104223 151600
rect 101078 151542 104223 151544
rect 211508 151600 214439 151602
rect 211508 151544 214378 151600
rect 214434 151544 214439 151600
rect 211508 151542 214439 151544
rect 101078 150960 101138 151542
rect 104157 151539 104223 151542
rect 214373 151539 214439 151542
rect 116393 151194 116459 151197
rect 116393 151192 119692 151194
rect 116393 151136 116398 151192
rect 116454 151136 119692 151192
rect 116393 151134 119692 151136
rect 116393 151131 116459 151134
rect -960 150786 480 150876
rect 2773 150786 2839 150789
rect 215109 150786 215175 150789
rect -960 150784 2839 150786
rect -960 150728 2778 150784
rect 2834 150728 2839 150784
rect -960 150726 2839 150728
rect 211508 150784 215175 150786
rect 211508 150728 215114 150784
rect 215170 150728 215175 150784
rect 211508 150726 215175 150728
rect -960 150636 480 150726
rect 2773 150723 2839 150726
rect 215109 150723 215175 150726
rect 103789 150378 103855 150381
rect 101078 150376 103855 150378
rect 101078 150320 103794 150376
rect 103850 150320 103855 150376
rect 101078 150318 103855 150320
rect 101078 149736 101138 150318
rect 103789 150315 103855 150318
rect 116393 149970 116459 149973
rect 214373 149970 214439 149973
rect 116393 149968 119692 149970
rect 116393 149912 116398 149968
rect 116454 149912 119692 149968
rect 116393 149910 119692 149912
rect 211508 149968 214439 149970
rect 211508 149912 214378 149968
rect 214434 149912 214439 149968
rect 211508 149910 214439 149912
rect 116393 149907 116459 149910
rect 214373 149907 214439 149910
rect 227437 149426 227503 149429
rect 227437 149424 230092 149426
rect 227437 149368 227442 149424
rect 227498 149368 230092 149424
rect 227437 149366 230092 149368
rect 227437 149363 227503 149366
rect 215109 149290 215175 149293
rect 211508 149288 215175 149290
rect 211508 149232 215114 149288
rect 215170 149232 215175 149288
rect 211508 149230 215175 149232
rect 215109 149227 215175 149230
rect 103697 149018 103763 149021
rect 101078 149016 103763 149018
rect 101078 148960 103702 149016
rect 103758 148960 103763 149016
rect 101078 148958 103763 148960
rect 101078 148512 101138 148958
rect 103697 148955 103763 148958
rect 227437 148882 227503 148885
rect 227437 148880 230092 148882
rect 227437 148824 227442 148880
rect 227498 148824 230092 148880
rect 227437 148822 230092 148824
rect 227437 148819 227503 148822
rect 116393 148746 116459 148749
rect 116393 148744 119692 148746
rect 116393 148688 116398 148744
rect 116454 148688 119692 148744
rect 116393 148686 119692 148688
rect 116393 148683 116459 148686
rect 215109 148474 215175 148477
rect 211508 148472 215175 148474
rect 211508 148416 215114 148472
rect 215170 148416 215175 148472
rect 211508 148414 215175 148416
rect 215109 148411 215175 148414
rect 227529 148202 227595 148205
rect 227529 148200 230092 148202
rect 227529 148144 227534 148200
rect 227590 148144 230092 148200
rect 227529 148142 230092 148144
rect 227529 148139 227595 148142
rect 104341 147658 104407 147661
rect 101078 147656 104407 147658
rect 101078 147600 104346 147656
rect 104402 147600 104407 147656
rect 101078 147598 104407 147600
rect 101078 147288 101138 147598
rect 104341 147595 104407 147598
rect 115933 147658 115999 147661
rect 214833 147658 214899 147661
rect 115933 147656 119692 147658
rect 115933 147600 115938 147656
rect 115994 147600 119692 147656
rect 115933 147598 119692 147600
rect 211508 147656 214899 147658
rect 211508 147600 214838 147656
rect 214894 147600 214899 147656
rect 211508 147598 214899 147600
rect 115933 147595 115999 147598
rect 214833 147595 214899 147598
rect 225597 147658 225663 147661
rect 225597 147656 230092 147658
rect 225597 147600 225602 147656
rect 225658 147600 230092 147656
rect 225597 147598 230092 147600
rect 225597 147595 225663 147598
rect 226701 146978 226767 146981
rect 226701 146976 230092 146978
rect 226701 146920 226706 146976
rect 226762 146920 230092 146976
rect 226701 146918 230092 146920
rect 226701 146915 226767 146918
rect 215201 146842 215267 146845
rect 211508 146840 215267 146842
rect 211508 146784 215206 146840
rect 215262 146784 215267 146840
rect 211508 146782 215267 146784
rect 215201 146779 215267 146782
rect 583520 146556 584960 146796
rect 116393 146434 116459 146437
rect 226517 146434 226583 146437
rect 116393 146432 119692 146434
rect 116393 146376 116398 146432
rect 116454 146376 119692 146432
rect 116393 146374 119692 146376
rect 226517 146432 230092 146434
rect 226517 146376 226522 146432
rect 226578 146376 230092 146432
rect 226517 146374 230092 146376
rect 116393 146371 116459 146374
rect 226517 146371 226583 146374
rect 104433 146298 104499 146301
rect 101078 146296 104499 146298
rect 101078 146240 104438 146296
rect 104494 146240 104499 146296
rect 101078 146238 104499 146240
rect 101078 146064 101138 146238
rect 104433 146235 104499 146238
rect 215017 146162 215083 146165
rect 211508 146160 215083 146162
rect 211508 146104 215022 146160
rect 215078 146104 215083 146160
rect 211508 146102 215083 146104
rect 215017 146099 215083 146102
rect 227437 145890 227503 145893
rect 227437 145888 230092 145890
rect 227437 145832 227442 145888
rect 227498 145832 230092 145888
rect 227437 145830 230092 145832
rect 227437 145827 227503 145830
rect 116025 145346 116091 145349
rect 215201 145346 215267 145349
rect 116025 145344 119692 145346
rect 116025 145288 116030 145344
rect 116086 145288 119692 145344
rect 116025 145286 119692 145288
rect 211508 145344 215267 145346
rect 211508 145288 215206 145344
rect 215262 145288 215267 145344
rect 211508 145286 215267 145288
rect 116025 145283 116091 145286
rect 215201 145283 215267 145286
rect 226701 145210 226767 145213
rect 226701 145208 230092 145210
rect 226701 145152 226706 145208
rect 226762 145152 230092 145208
rect 226701 145150 230092 145152
rect 226701 145147 226767 145150
rect 101078 144802 101138 144840
rect 104801 144802 104867 144805
rect 101078 144800 104867 144802
rect 101078 144744 104806 144800
rect 104862 144744 104867 144800
rect 101078 144742 104867 144744
rect 104801 144739 104867 144742
rect 227437 144666 227503 144669
rect 227437 144664 230092 144666
rect 227437 144608 227442 144664
rect 227498 144608 230092 144664
rect 227437 144606 230092 144608
rect 227437 144603 227503 144606
rect 214465 144530 214531 144533
rect 211508 144528 214531 144530
rect 211508 144472 214470 144528
rect 214526 144472 214531 144528
rect 211508 144470 214531 144472
rect 214465 144467 214531 144470
rect 104617 144258 104683 144261
rect 101078 144256 104683 144258
rect 101078 144200 104622 144256
rect 104678 144200 104683 144256
rect 101078 144198 104683 144200
rect 101078 143616 101138 144198
rect 104617 144195 104683 144198
rect 116393 144122 116459 144125
rect 116393 144120 119692 144122
rect 116393 144064 116398 144120
rect 116454 144064 119692 144120
rect 116393 144062 119692 144064
rect 116393 144059 116459 144062
rect 226517 143986 226583 143989
rect 226517 143984 230092 143986
rect 226517 143928 226522 143984
rect 226578 143928 230092 143984
rect 226517 143926 230092 143928
rect 226517 143923 226583 143926
rect 215201 143714 215267 143717
rect 211508 143712 215267 143714
rect 211508 143656 215206 143712
rect 215262 143656 215267 143712
rect 211508 143654 215267 143656
rect 215201 143651 215267 143654
rect 227437 143442 227503 143445
rect 227437 143440 230092 143442
rect 227437 143384 227442 143440
rect 227498 143384 230092 143440
rect 227437 143382 230092 143384
rect 227437 143379 227503 143382
rect 104157 143034 104223 143037
rect 215109 143034 215175 143037
rect 101078 143032 104223 143034
rect 101078 142976 104162 143032
rect 104218 142976 104223 143032
rect 101078 142974 104223 142976
rect 211508 143032 215175 143034
rect 211508 142976 215114 143032
rect 215170 142976 215175 143032
rect 211508 142974 215175 142976
rect 101078 142392 101138 142974
rect 104157 142971 104223 142974
rect 215109 142971 215175 142974
rect 116393 142898 116459 142901
rect 226885 142898 226951 142901
rect 116393 142896 119692 142898
rect 116393 142840 116398 142896
rect 116454 142840 119692 142896
rect 116393 142838 119692 142840
rect 226885 142896 230092 142898
rect 226885 142840 226890 142896
rect 226946 142840 230092 142896
rect 226885 142838 230092 142840
rect 116393 142835 116459 142838
rect 226885 142835 226951 142838
rect 215201 142218 215267 142221
rect 211508 142216 215267 142218
rect 211508 142160 215206 142216
rect 215262 142160 215267 142216
rect 211508 142158 215267 142160
rect 215201 142155 215267 142158
rect 227621 142218 227687 142221
rect 227621 142216 230092 142218
rect 227621 142160 227626 142216
rect 227682 142160 230092 142216
rect 227621 142158 230092 142160
rect 227621 142155 227687 142158
rect 104525 141810 104591 141813
rect 101078 141808 104591 141810
rect 101078 141752 104530 141808
rect 104586 141752 104591 141808
rect 101078 141750 104591 141752
rect 101078 141168 101138 141750
rect 104525 141747 104591 141750
rect 116393 141810 116459 141813
rect 116393 141808 119692 141810
rect 116393 141752 116398 141808
rect 116454 141752 119692 141808
rect 116393 141750 119692 141752
rect 116393 141747 116459 141750
rect 226701 141674 226767 141677
rect 226701 141672 230092 141674
rect 226701 141616 226706 141672
rect 226762 141616 230092 141672
rect 226701 141614 230092 141616
rect 226701 141611 226767 141614
rect 215109 141402 215175 141405
rect 211508 141400 215175 141402
rect 211508 141344 215114 141400
rect 215170 141344 215175 141400
rect 211508 141342 215175 141344
rect 215109 141339 215175 141342
rect 227253 140994 227319 140997
rect 227253 140992 230092 140994
rect 227253 140936 227258 140992
rect 227314 140936 230092 140992
rect 227253 140934 230092 140936
rect 227253 140931 227319 140934
rect 103513 140586 103579 140589
rect 101078 140584 103579 140586
rect 101078 140528 103518 140584
rect 103574 140528 103579 140584
rect 101078 140526 103579 140528
rect 101078 139944 101138 140526
rect 103513 140523 103579 140526
rect 116393 140586 116459 140589
rect 215109 140586 215175 140589
rect 116393 140584 119692 140586
rect 116393 140528 116398 140584
rect 116454 140528 119692 140584
rect 116393 140526 119692 140528
rect 211508 140584 215175 140586
rect 211508 140528 215114 140584
rect 215170 140528 215175 140584
rect 211508 140526 215175 140528
rect 116393 140523 116459 140526
rect 215109 140523 215175 140526
rect 227069 140450 227135 140453
rect 227069 140448 230092 140450
rect 227069 140392 227074 140448
rect 227130 140392 230092 140448
rect 227069 140390 230092 140392
rect 227069 140387 227135 140390
rect 214373 139906 214439 139909
rect 211508 139904 214439 139906
rect 211508 139848 214378 139904
rect 214434 139848 214439 139904
rect 211508 139846 214439 139848
rect 214373 139843 214439 139846
rect 227529 139770 227595 139773
rect 227529 139768 230092 139770
rect 227529 139712 227534 139768
rect 227590 139712 230092 139768
rect 227529 139710 230092 139712
rect 227529 139707 227595 139710
rect 116301 139498 116367 139501
rect 116301 139496 119692 139498
rect 116301 139440 116306 139496
rect 116362 139440 119692 139496
rect 116301 139438 119692 139440
rect 116301 139435 116367 139438
rect 103697 139362 103763 139365
rect 101078 139360 103763 139362
rect 101078 139304 103702 139360
rect 103758 139304 103763 139360
rect 101078 139302 103763 139304
rect 101078 138720 101138 139302
rect 103697 139299 103763 139302
rect 227437 139226 227503 139229
rect 227437 139224 230092 139226
rect 227437 139168 227442 139224
rect 227498 139168 230092 139224
rect 227437 139166 230092 139168
rect 227437 139163 227503 139166
rect 214465 139090 214531 139093
rect 211508 139088 214531 139090
rect 211508 139032 214470 139088
rect 214526 139032 214531 139088
rect 211508 139030 214531 139032
rect 214465 139027 214531 139030
rect 227345 138682 227411 138685
rect 227345 138680 230092 138682
rect 227345 138624 227350 138680
rect 227406 138624 230092 138680
rect 227345 138622 230092 138624
rect 227345 138619 227411 138622
rect 115841 138274 115907 138277
rect 215109 138274 215175 138277
rect 115841 138272 119692 138274
rect 115841 138216 115846 138272
rect 115902 138216 119692 138272
rect 115841 138214 119692 138216
rect 211508 138272 215175 138274
rect 211508 138216 215114 138272
rect 215170 138216 215175 138272
rect 211508 138214 215175 138216
rect 115841 138211 115907 138214
rect 215109 138211 215175 138214
rect 104341 138002 104407 138005
rect 101078 138000 104407 138002
rect 101078 137944 104346 138000
rect 104402 137944 104407 138000
rect 101078 137942 104407 137944
rect 101078 137496 101138 137942
rect 104341 137939 104407 137942
rect 227437 138002 227503 138005
rect 227437 138000 230092 138002
rect 227437 137944 227442 138000
rect 227498 137944 230092 138000
rect 227437 137942 230092 137944
rect 227437 137939 227503 137942
rect 214281 137458 214347 137461
rect 211508 137456 214347 137458
rect 211508 137400 214286 137456
rect 214342 137400 214347 137456
rect 211508 137398 214347 137400
rect 214281 137395 214347 137398
rect 226701 137458 226767 137461
rect 226701 137456 230092 137458
rect 226701 137400 226706 137456
rect 226762 137400 230092 137456
rect 226701 137398 230092 137400
rect 226701 137395 226767 137398
rect 116393 137186 116459 137189
rect 116393 137184 119692 137186
rect 116393 137128 116398 137184
rect 116454 137128 119692 137184
rect 116393 137126 119692 137128
rect 116393 137123 116459 137126
rect 215109 136778 215175 136781
rect 211508 136776 215175 136778
rect 211508 136720 215114 136776
rect 215170 136720 215175 136776
rect 211508 136718 215175 136720
rect 215109 136715 215175 136718
rect 226517 136778 226583 136781
rect 226517 136776 230092 136778
rect 226517 136720 226522 136776
rect 226578 136720 230092 136776
rect 226517 136718 230092 136720
rect 226517 136715 226583 136718
rect 104801 136642 104867 136645
rect 101078 136640 104867 136642
rect 101078 136584 104806 136640
rect 104862 136584 104867 136640
rect 101078 136582 104867 136584
rect -960 136370 480 136460
rect 2773 136370 2839 136373
rect -960 136368 2839 136370
rect -960 136312 2778 136368
rect 2834 136312 2839 136368
rect -960 136310 2839 136312
rect -960 136220 480 136310
rect 2773 136307 2839 136310
rect 101078 136272 101138 136582
rect 104801 136579 104867 136582
rect 226609 136234 226675 136237
rect 226609 136232 230092 136234
rect 226609 136176 226614 136232
rect 226670 136176 230092 136232
rect 226609 136174 230092 136176
rect 226609 136171 226675 136174
rect 115933 135962 115999 135965
rect 214189 135962 214255 135965
rect 115933 135960 119692 135962
rect 115933 135904 115938 135960
rect 115994 135904 119692 135960
rect 115933 135902 119692 135904
rect 211508 135960 214255 135962
rect 211508 135904 214194 135960
rect 214250 135904 214255 135960
rect 211508 135902 214255 135904
rect 115933 135899 115999 135902
rect 214189 135899 214255 135902
rect 226425 135690 226491 135693
rect 226425 135688 230092 135690
rect 226425 135632 226430 135688
rect 226486 135632 230092 135688
rect 226425 135630 230092 135632
rect 226425 135627 226491 135630
rect 104801 135146 104867 135149
rect 215201 135146 215267 135149
rect 101078 135144 104867 135146
rect 101078 135088 104806 135144
rect 104862 135088 104867 135144
rect 101078 135086 104867 135088
rect 211508 135144 215267 135146
rect 211508 135088 215206 135144
rect 215262 135088 215267 135144
rect 211508 135086 215267 135088
rect 101078 135048 101138 135086
rect 104801 135083 104867 135086
rect 215201 135083 215267 135086
rect 226793 135010 226859 135013
rect 226793 135008 230092 135010
rect 226793 134952 226798 135008
rect 226854 134952 230092 135008
rect 226793 134950 230092 134952
rect 226793 134947 226859 134950
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 116393 134738 116459 134741
rect 116393 134736 119692 134738
rect 116393 134680 116398 134736
rect 116454 134680 119692 134736
rect 583520 134724 584960 134814
rect 116393 134678 119692 134680
rect 116393 134675 116459 134678
rect 227437 134466 227503 134469
rect 227437 134464 230092 134466
rect 227437 134408 227442 134464
rect 227498 134408 230092 134464
rect 227437 134406 230092 134408
rect 227437 134403 227503 134406
rect 215109 134330 215175 134333
rect 211508 134328 215175 134330
rect 211508 134272 215114 134328
rect 215170 134272 215175 134328
rect 211508 134270 215175 134272
rect 215109 134267 215175 134270
rect 101078 133786 101138 133824
rect 104801 133786 104867 133789
rect 101078 133784 104867 133786
rect 101078 133728 104806 133784
rect 104862 133728 104867 133784
rect 101078 133726 104867 133728
rect 104801 133723 104867 133726
rect 227253 133786 227319 133789
rect 227253 133784 230092 133786
rect 227253 133728 227258 133784
rect 227314 133728 230092 133784
rect 227253 133726 230092 133728
rect 227253 133723 227319 133726
rect 117129 133650 117195 133653
rect 117129 133648 119692 133650
rect 117129 133592 117134 133648
rect 117190 133592 119692 133648
rect 117129 133590 119692 133592
rect 117129 133587 117195 133590
rect 215109 133514 215175 133517
rect 211508 133512 215175 133514
rect 211508 133456 215114 133512
rect 215170 133456 215175 133512
rect 211508 133454 215175 133456
rect 215109 133451 215175 133454
rect 104709 133242 104775 133245
rect 101078 133240 104775 133242
rect 101078 133184 104714 133240
rect 104770 133184 104775 133240
rect 101078 133182 104775 133184
rect 101078 132600 101138 133182
rect 104709 133179 104775 133182
rect 226517 133242 226583 133245
rect 226517 133240 230092 133242
rect 226517 133184 226522 133240
rect 226578 133184 230092 133240
rect 226517 133182 230092 133184
rect 226517 133179 226583 133182
rect 214005 132834 214071 132837
rect 211508 132832 214071 132834
rect 211508 132776 214010 132832
rect 214066 132776 214071 132832
rect 211508 132774 214071 132776
rect 214005 132771 214071 132774
rect 227529 132562 227595 132565
rect 227529 132560 230092 132562
rect 227529 132504 227534 132560
rect 227590 132504 230092 132560
rect 227529 132502 230092 132504
rect 227529 132499 227595 132502
rect 116117 132426 116183 132429
rect 116117 132424 119692 132426
rect 116117 132368 116122 132424
rect 116178 132368 119692 132424
rect 116117 132366 119692 132368
rect 116117 132363 116183 132366
rect 104341 132018 104407 132021
rect 214373 132018 214439 132021
rect 101078 132016 104407 132018
rect 101078 131960 104346 132016
rect 104402 131960 104407 132016
rect 101078 131958 104407 131960
rect 211508 132016 214439 132018
rect 211508 131960 214378 132016
rect 214434 131960 214439 132016
rect 211508 131958 214439 131960
rect 101078 131376 101138 131958
rect 104341 131955 104407 131958
rect 214373 131955 214439 131958
rect 226701 132018 226767 132021
rect 226701 132016 230092 132018
rect 226701 131960 226706 132016
rect 226762 131960 230092 132016
rect 226701 131958 230092 131960
rect 226701 131955 226767 131958
rect 227437 131474 227503 131477
rect 227437 131472 230092 131474
rect 227437 131416 227442 131472
rect 227498 131416 230092 131472
rect 227437 131414 230092 131416
rect 227437 131411 227503 131414
rect 116393 131338 116459 131341
rect 116393 131336 119692 131338
rect 116393 131280 116398 131336
rect 116454 131280 119692 131336
rect 116393 131278 119692 131280
rect 116393 131275 116459 131278
rect 215109 131202 215175 131205
rect 211508 131200 215175 131202
rect 211508 131144 215114 131200
rect 215170 131144 215175 131200
rect 211508 131142 215175 131144
rect 215109 131139 215175 131142
rect 227345 130794 227411 130797
rect 227345 130792 230092 130794
rect 227345 130736 227350 130792
rect 227406 130736 230092 130792
rect 227345 130734 230092 130736
rect 227345 130731 227411 130734
rect 103973 130658 104039 130661
rect 101078 130656 104039 130658
rect 101078 130600 103978 130656
rect 104034 130600 104039 130656
rect 101078 130598 104039 130600
rect 101078 130152 101138 130598
rect 103973 130595 104039 130598
rect 214189 130386 214255 130389
rect 211508 130384 214255 130386
rect 211508 130328 214194 130384
rect 214250 130328 214255 130384
rect 211508 130326 214255 130328
rect 214189 130323 214255 130326
rect 227069 130250 227135 130253
rect 227069 130248 230092 130250
rect 227069 130192 227074 130248
rect 227130 130192 230092 130248
rect 227069 130190 230092 130192
rect 227069 130187 227135 130190
rect 116669 130114 116735 130117
rect 116669 130112 119692 130114
rect 116669 130056 116674 130112
rect 116730 130056 119692 130112
rect 116669 130054 119692 130056
rect 116669 130051 116735 130054
rect 214189 129706 214255 129709
rect 211508 129704 214255 129706
rect 211508 129648 214194 129704
rect 214250 129648 214255 129704
rect 211508 129646 214255 129648
rect 214189 129643 214255 129646
rect 226517 129570 226583 129573
rect 226517 129568 230092 129570
rect 226517 129512 226522 129568
rect 226578 129512 230092 129568
rect 226517 129510 230092 129512
rect 226517 129507 226583 129510
rect 104801 129298 104867 129301
rect 101078 129296 104867 129298
rect 101078 129240 104806 129296
rect 104862 129240 104867 129296
rect 101078 129238 104867 129240
rect 101078 128928 101138 129238
rect 104801 129235 104867 129238
rect 227529 129026 227595 129029
rect 227529 129024 230092 129026
rect 227529 128968 227534 129024
rect 227590 128968 230092 129024
rect 227529 128966 230092 128968
rect 227529 128963 227595 128966
rect 116393 128890 116459 128893
rect 214005 128890 214071 128893
rect 116393 128888 119692 128890
rect 116393 128832 116398 128888
rect 116454 128832 119692 128888
rect 116393 128830 119692 128832
rect 211508 128888 214071 128890
rect 211508 128832 214010 128888
rect 214066 128832 214071 128888
rect 211508 128830 214071 128832
rect 116393 128827 116459 128830
rect 214005 128827 214071 128830
rect 227437 128482 227503 128485
rect 227437 128480 230092 128482
rect 227437 128424 227442 128480
rect 227498 128424 230092 128480
rect 227437 128422 230092 128424
rect 227437 128419 227503 128422
rect 104801 128074 104867 128077
rect 215109 128074 215175 128077
rect 101078 128072 104867 128074
rect 101078 128016 104806 128072
rect 104862 128016 104867 128072
rect 101078 128014 104867 128016
rect 211508 128072 215175 128074
rect 211508 128016 215114 128072
rect 215170 128016 215175 128072
rect 211508 128014 215175 128016
rect 101078 127840 101138 128014
rect 104801 128011 104867 128014
rect 215109 128011 215175 128014
rect 116393 127802 116459 127805
rect 226333 127802 226399 127805
rect 116393 127800 119692 127802
rect 116393 127744 116398 127800
rect 116454 127744 119692 127800
rect 116393 127742 119692 127744
rect 226333 127800 230092 127802
rect 226333 127744 226338 127800
rect 226394 127744 230092 127800
rect 226333 127742 230092 127744
rect 116393 127739 116459 127742
rect 226333 127739 226399 127742
rect 215109 127258 215175 127261
rect 211508 127256 215175 127258
rect 211508 127200 215114 127256
rect 215170 127200 215175 127256
rect 211508 127198 215175 127200
rect 215109 127195 215175 127198
rect 227437 127258 227503 127261
rect 227437 127256 230092 127258
rect 227437 127200 227442 127256
rect 227498 127200 230092 127256
rect 227437 127198 230092 127200
rect 227437 127195 227503 127198
rect 343633 126714 343699 126717
rect 342148 126712 343699 126714
rect 342148 126656 343638 126712
rect 343694 126656 343699 126712
rect 342148 126654 343699 126656
rect 343633 126651 343699 126654
rect 116393 126578 116459 126581
rect 215109 126578 215175 126581
rect 116393 126576 119692 126578
rect 116393 126520 116398 126576
rect 116454 126520 119692 126576
rect 116393 126518 119692 126520
rect 211508 126576 215175 126578
rect 211508 126520 215114 126576
rect 215170 126520 215175 126576
rect 211508 126518 215175 126520
rect 116393 126515 116459 126518
rect 215109 126515 215175 126518
rect 227437 126578 227503 126581
rect 227437 126576 230092 126578
rect 227437 126520 227442 126576
rect 227498 126520 230092 126576
rect 227437 126518 230092 126520
rect 227437 126515 227503 126518
rect 227437 126034 227503 126037
rect 227437 126032 230092 126034
rect 227437 125976 227442 126032
rect 227498 125976 230092 126032
rect 227437 125974 230092 125976
rect 227437 125971 227503 125974
rect 215109 125762 215175 125765
rect 211508 125760 215175 125762
rect 211508 125704 215114 125760
rect 215170 125704 215175 125760
rect 211508 125702 215175 125704
rect 215109 125699 215175 125702
rect 116393 125490 116459 125493
rect 116393 125488 119692 125490
rect 116393 125432 116398 125488
rect 116454 125432 119692 125488
rect 116393 125430 119692 125432
rect 116393 125427 116459 125430
rect 227437 125354 227503 125357
rect 227437 125352 230092 125354
rect 227437 125296 227442 125352
rect 227498 125296 230092 125352
rect 227437 125294 230092 125296
rect 227437 125291 227503 125294
rect 32213 125084 32279 125085
rect 32213 125080 32260 125084
rect 32324 125082 32330 125084
rect 32213 125024 32218 125080
rect 32213 125020 32260 125024
rect 32324 125022 32370 125082
rect 32324 125020 32330 125022
rect 32213 125019 32279 125020
rect 215109 124946 215175 124949
rect 211508 124944 215175 124946
rect 211508 124888 215114 124944
rect 215170 124888 215175 124944
rect 211508 124886 215175 124888
rect 215109 124883 215175 124886
rect 227253 124810 227319 124813
rect 227253 124808 230092 124810
rect 227253 124752 227258 124808
rect 227314 124752 230092 124808
rect 227253 124750 230092 124752
rect 227253 124747 227319 124750
rect 18638 124204 18644 124268
rect 18708 124266 18714 124268
rect 227253 124266 227319 124269
rect 18708 124206 119692 124266
rect 227253 124264 230092 124266
rect 227253 124208 227258 124264
rect 227314 124208 230092 124264
rect 227253 124206 230092 124208
rect 18708 124204 18714 124206
rect 227253 124203 227319 124206
rect 215109 124130 215175 124133
rect 211508 124128 215175 124130
rect 211508 124072 215114 124128
rect 215170 124072 215175 124128
rect 211508 124070 215175 124072
rect 215109 124067 215175 124070
rect 227253 123586 227319 123589
rect 227253 123584 230092 123586
rect 227253 123528 227258 123584
rect 227314 123528 230092 123584
rect 227253 123526 230092 123528
rect 227253 123523 227319 123526
rect 215109 123450 215175 123453
rect 211508 123448 215175 123450
rect 211508 123392 215114 123448
rect 215170 123392 215175 123448
rect 211508 123390 215175 123392
rect 215109 123387 215175 123390
rect 580901 123178 580967 123181
rect 583520 123178 584960 123268
rect 580901 123176 584960 123178
rect 580901 123120 580906 123176
rect 580962 123120 584960 123176
rect 580901 123118 584960 123120
rect 580901 123115 580967 123118
rect 116577 123042 116643 123045
rect 227437 123042 227503 123045
rect 116577 123040 119692 123042
rect 116577 122984 116582 123040
rect 116638 122984 119692 123040
rect 116577 122982 119692 122984
rect 227437 123040 230092 123042
rect 227437 122984 227442 123040
rect 227498 122984 230092 123040
rect 583520 123028 584960 123118
rect 227437 122982 230092 122984
rect 116577 122979 116643 122982
rect 227437 122979 227503 122982
rect 215109 122634 215175 122637
rect 211508 122632 215175 122634
rect 211508 122576 215114 122632
rect 215170 122576 215175 122632
rect 211508 122574 215175 122576
rect 215109 122571 215175 122574
rect 227437 122362 227503 122365
rect 227437 122360 230092 122362
rect 227437 122304 227442 122360
rect 227498 122304 230092 122360
rect 227437 122302 230092 122304
rect 227437 122299 227503 122302
rect -960 121940 480 122180
rect 116393 121954 116459 121957
rect 116393 121952 119692 121954
rect 116393 121896 116398 121952
rect 116454 121896 119692 121952
rect 116393 121894 119692 121896
rect 116393 121891 116459 121894
rect 215109 121818 215175 121821
rect 211508 121816 215175 121818
rect 211508 121760 215114 121816
rect 215170 121760 215175 121816
rect 211508 121758 215175 121760
rect 215109 121755 215175 121758
rect 227437 121818 227503 121821
rect 227437 121816 230092 121818
rect 227437 121760 227442 121816
rect 227498 121760 230092 121816
rect 227437 121758 230092 121760
rect 227437 121755 227503 121758
rect 227437 121274 227503 121277
rect 227437 121272 230092 121274
rect 227437 121216 227442 121272
rect 227498 121216 230092 121272
rect 227437 121214 230092 121216
rect 227437 121211 227503 121214
rect 215109 121002 215175 121005
rect 211508 121000 215175 121002
rect 211508 120944 215114 121000
rect 215170 120944 215175 121000
rect 211508 120942 215175 120944
rect 215109 120939 215175 120942
rect 116393 120730 116459 120733
rect 116393 120728 119692 120730
rect 116393 120672 116398 120728
rect 116454 120672 119692 120728
rect 116393 120670 119692 120672
rect 116393 120667 116459 120670
rect 227437 120594 227503 120597
rect 227437 120592 230092 120594
rect 227437 120536 227442 120592
rect 227498 120536 230092 120592
rect 227437 120534 230092 120536
rect 227437 120531 227503 120534
rect 215109 120322 215175 120325
rect 211508 120320 215175 120322
rect 211508 120264 215114 120320
rect 215170 120264 215175 120320
rect 211508 120262 215175 120264
rect 215109 120259 215175 120262
rect 226425 120050 226491 120053
rect 226425 120048 230092 120050
rect 226425 119992 226430 120048
rect 226486 119992 230092 120048
rect 226425 119990 230092 119992
rect 226425 119987 226491 119990
rect 116393 119642 116459 119645
rect 116393 119640 119692 119642
rect 116393 119584 116398 119640
rect 116454 119584 119692 119640
rect 116393 119582 119692 119584
rect 116393 119579 116459 119582
rect 214189 119506 214255 119509
rect 211508 119504 214255 119506
rect 211508 119448 214194 119504
rect 214250 119448 214255 119504
rect 211508 119446 214255 119448
rect 214189 119443 214255 119446
rect 226333 119370 226399 119373
rect 226333 119368 230092 119370
rect 226333 119312 226338 119368
rect 226394 119312 230092 119368
rect 226333 119310 230092 119312
rect 226333 119307 226399 119310
rect 226241 118826 226307 118829
rect 226241 118824 230092 118826
rect 226241 118768 226246 118824
rect 226302 118768 230092 118824
rect 226241 118766 230092 118768
rect 226241 118763 226307 118766
rect 215109 118690 215175 118693
rect 211508 118688 215175 118690
rect 211508 118632 215114 118688
rect 215170 118632 215175 118688
rect 211508 118630 215175 118632
rect 215109 118627 215175 118630
rect 116393 118418 116459 118421
rect 116393 118416 119692 118418
rect 116393 118360 116398 118416
rect 116454 118360 119692 118416
rect 116393 118358 119692 118360
rect 116393 118355 116459 118358
rect 227437 118146 227503 118149
rect 227437 118144 230092 118146
rect 227437 118088 227442 118144
rect 227498 118088 230092 118144
rect 227437 118086 230092 118088
rect 227437 118083 227503 118086
rect 214281 117874 214347 117877
rect 211508 117872 214347 117874
rect 211508 117816 214286 117872
rect 214342 117816 214347 117872
rect 211508 117814 214347 117816
rect 214281 117811 214347 117814
rect 226149 117602 226215 117605
rect 226149 117600 230092 117602
rect 226149 117544 226154 117600
rect 226210 117544 230092 117600
rect 226149 117542 230092 117544
rect 226149 117539 226215 117542
rect 116301 117194 116367 117197
rect 116301 117192 119692 117194
rect 116301 117136 116306 117192
rect 116362 117136 119692 117192
rect 116301 117134 119692 117136
rect 116301 117131 116367 117134
rect 215109 117058 215175 117061
rect 211508 117056 215175 117058
rect 211508 117000 215114 117056
rect 215170 117000 215175 117056
rect 211508 116998 215175 117000
rect 215109 116995 215175 116998
rect 227437 117058 227503 117061
rect 227437 117056 230092 117058
rect 227437 117000 227442 117056
rect 227498 117000 230092 117056
rect 227437 116998 230092 117000
rect 227437 116995 227503 116998
rect 215201 116378 215267 116381
rect 211508 116376 215267 116378
rect 211508 116320 215206 116376
rect 215262 116320 215267 116376
rect 211508 116318 215267 116320
rect 215201 116315 215267 116318
rect 226241 116378 226307 116381
rect 226241 116376 230092 116378
rect 226241 116320 226246 116376
rect 226302 116320 230092 116376
rect 226241 116318 230092 116320
rect 226241 116315 226307 116318
rect 116393 116106 116459 116109
rect 116393 116104 119692 116106
rect 116393 116048 116398 116104
rect 116454 116048 119692 116104
rect 116393 116046 119692 116048
rect 116393 116043 116459 116046
rect 227069 115834 227135 115837
rect 227069 115832 230092 115834
rect 227069 115776 227074 115832
rect 227130 115776 230092 115832
rect 227069 115774 230092 115776
rect 227069 115771 227135 115774
rect 215109 115562 215175 115565
rect 211508 115560 215175 115562
rect 211508 115504 215114 115560
rect 215170 115504 215175 115560
rect 211508 115502 215175 115504
rect 215109 115499 215175 115502
rect 226149 115154 226215 115157
rect 226149 115152 230092 115154
rect 226149 115096 226154 115152
rect 226210 115096 230092 115152
rect 226149 115094 230092 115096
rect 226149 115091 226215 115094
rect 116393 114882 116459 114885
rect 116393 114880 119692 114882
rect 116393 114824 116398 114880
rect 116454 114824 119692 114880
rect 116393 114822 119692 114824
rect 116393 114819 116459 114822
rect 215201 114746 215267 114749
rect 211508 114744 215267 114746
rect 211508 114688 215206 114744
rect 215262 114688 215267 114744
rect 211508 114686 215267 114688
rect 215201 114683 215267 114686
rect 226057 114610 226123 114613
rect 226057 114608 230092 114610
rect 226057 114552 226062 114608
rect 226118 114552 230092 114608
rect 226057 114550 230092 114552
rect 226057 114547 226123 114550
rect 226241 114066 226307 114069
rect 226241 114064 230092 114066
rect 226241 114008 226246 114064
rect 226302 114008 230092 114064
rect 226241 114006 230092 114008
rect 226241 114003 226307 114006
rect 214005 113930 214071 113933
rect 211508 113928 214071 113930
rect 211508 113872 214010 113928
rect 214066 113872 214071 113928
rect 211508 113870 214071 113872
rect 214005 113867 214071 113870
rect 116393 113794 116459 113797
rect 116393 113792 119692 113794
rect 116393 113736 116398 113792
rect 116454 113736 119692 113792
rect 116393 113734 119692 113736
rect 116393 113731 116459 113734
rect 225965 113386 226031 113389
rect 225965 113384 230092 113386
rect 225965 113328 225970 113384
rect 226026 113328 230092 113384
rect 225965 113326 230092 113328
rect 225965 113323 226031 113326
rect 215109 113250 215175 113253
rect 211508 113248 215175 113250
rect 211508 113192 215114 113248
rect 215170 113192 215175 113248
rect 211508 113190 215175 113192
rect 215109 113187 215175 113190
rect 226149 112842 226215 112845
rect 226149 112840 230092 112842
rect 226149 112784 226154 112840
rect 226210 112784 230092 112840
rect 226149 112782 230092 112784
rect 226149 112779 226215 112782
rect 116393 112570 116459 112573
rect 116393 112568 119692 112570
rect 116393 112512 116398 112568
rect 116454 112512 119692 112568
rect 116393 112510 119692 112512
rect 116393 112507 116459 112510
rect 214373 112434 214439 112437
rect 211508 112432 214439 112434
rect 211508 112376 214378 112432
rect 214434 112376 214439 112432
rect 211508 112374 214439 112376
rect 214373 112371 214439 112374
rect 225781 112162 225847 112165
rect 225781 112160 230092 112162
rect 225781 112104 225786 112160
rect 225842 112104 230092 112160
rect 225781 112102 230092 112104
rect 225781 112099 225847 112102
rect 215109 111618 215175 111621
rect 211508 111616 215175 111618
rect 211508 111560 215114 111616
rect 215170 111560 215175 111616
rect 211508 111558 215175 111560
rect 215109 111555 215175 111558
rect 226241 111618 226307 111621
rect 226241 111616 230092 111618
rect 226241 111560 226246 111616
rect 226302 111560 230092 111616
rect 226241 111558 230092 111560
rect 226241 111555 226307 111558
rect 116393 111482 116459 111485
rect 116393 111480 119692 111482
rect 116393 111424 116398 111480
rect 116454 111424 119692 111480
rect 116393 111422 119692 111424
rect 116393 111419 116459 111422
rect 583520 111332 584960 111572
rect 226057 110938 226123 110941
rect 226057 110936 230092 110938
rect 226057 110880 226062 110936
rect 226118 110880 230092 110936
rect 226057 110878 230092 110880
rect 226057 110875 226123 110878
rect 215201 110802 215267 110805
rect 211508 110800 215267 110802
rect 211508 110744 215206 110800
rect 215262 110744 215267 110800
rect 211508 110742 215267 110744
rect 215201 110739 215267 110742
rect 225689 110394 225755 110397
rect 225689 110392 230092 110394
rect 225689 110336 225694 110392
rect 225750 110336 230092 110392
rect 225689 110334 230092 110336
rect 225689 110331 225755 110334
rect 116393 110258 116459 110261
rect 116393 110256 119692 110258
rect 116393 110200 116398 110256
rect 116454 110200 119692 110256
rect 116393 110198 119692 110200
rect 116393 110195 116459 110198
rect 215109 110122 215175 110125
rect 211508 110120 215175 110122
rect 211508 110064 215114 110120
rect 215170 110064 215175 110120
rect 211508 110062 215175 110064
rect 215109 110059 215175 110062
rect 226149 109850 226215 109853
rect 226149 109848 230092 109850
rect 226149 109792 226154 109848
rect 226210 109792 230092 109848
rect 226149 109790 230092 109792
rect 226149 109787 226215 109790
rect 214465 109306 214531 109309
rect 211508 109304 214531 109306
rect 211508 109248 214470 109304
rect 214526 109248 214531 109304
rect 211508 109246 214531 109248
rect 214465 109243 214531 109246
rect 225597 109170 225663 109173
rect 225597 109168 230092 109170
rect 225597 109112 225602 109168
rect 225658 109112 230092 109168
rect 225597 109110 230092 109112
rect 225597 109107 225663 109110
rect 116301 109034 116367 109037
rect 116301 109032 119692 109034
rect 116301 108976 116306 109032
rect 116362 108976 119692 109032
rect 116301 108974 119692 108976
rect 116301 108971 116367 108974
rect 226241 108626 226307 108629
rect 226241 108624 230092 108626
rect 226241 108568 226246 108624
rect 226302 108568 230092 108624
rect 226241 108566 230092 108568
rect 226241 108563 226307 108566
rect 215109 108490 215175 108493
rect 211508 108488 215175 108490
rect 211508 108432 215114 108488
rect 215170 108432 215175 108488
rect 211508 108430 215175 108432
rect 215109 108427 215175 108430
rect 116393 107946 116459 107949
rect 225781 107946 225847 107949
rect 116393 107944 119692 107946
rect 116393 107888 116398 107944
rect 116454 107888 119692 107944
rect 116393 107886 119692 107888
rect 225781 107944 230092 107946
rect 225781 107888 225786 107944
rect 225842 107888 230092 107944
rect 225781 107886 230092 107888
rect 116393 107883 116459 107886
rect 225781 107883 225847 107886
rect -960 107674 480 107764
rect 2773 107674 2839 107677
rect 215201 107674 215267 107677
rect -960 107672 2839 107674
rect -960 107616 2778 107672
rect 2834 107616 2839 107672
rect -960 107614 2839 107616
rect 211508 107672 215267 107674
rect 211508 107616 215206 107672
rect 215262 107616 215267 107672
rect 211508 107614 215267 107616
rect -960 107524 480 107614
rect 2773 107611 2839 107614
rect 215201 107611 215267 107614
rect 226057 107402 226123 107405
rect 226057 107400 230092 107402
rect 226057 107344 226062 107400
rect 226118 107344 230092 107400
rect 226057 107342 230092 107344
rect 226057 107339 226123 107342
rect 214189 106994 214255 106997
rect 211508 106992 214255 106994
rect 211508 106936 214194 106992
rect 214250 106936 214255 106992
rect 211508 106934 214255 106936
rect 214189 106931 214255 106934
rect 225873 106858 225939 106861
rect 225873 106856 230092 106858
rect 225873 106800 225878 106856
rect 225934 106800 230092 106856
rect 225873 106798 230092 106800
rect 225873 106795 225939 106798
rect 116393 106722 116459 106725
rect 116393 106720 119692 106722
rect 116393 106664 116398 106720
rect 116454 106664 119692 106720
rect 116393 106662 119692 106664
rect 116393 106659 116459 106662
rect 215109 106178 215175 106181
rect 211508 106176 215175 106178
rect 211508 106120 215114 106176
rect 215170 106120 215175 106176
rect 211508 106118 215175 106120
rect 215109 106115 215175 106118
rect 225965 106178 226031 106181
rect 225965 106176 230092 106178
rect 225965 106120 225970 106176
rect 226026 106120 230092 106176
rect 225965 106118 230092 106120
rect 225965 106115 226031 106118
rect 116393 105634 116459 105637
rect 226149 105634 226215 105637
rect 116393 105632 119692 105634
rect 116393 105576 116398 105632
rect 116454 105576 119692 105632
rect 116393 105574 119692 105576
rect 226149 105632 230092 105634
rect 226149 105576 226154 105632
rect 226210 105576 230092 105632
rect 226149 105574 230092 105576
rect 116393 105571 116459 105574
rect 226149 105571 226215 105574
rect 214373 105362 214439 105365
rect 211508 105360 214439 105362
rect 211508 105304 214378 105360
rect 214434 105304 214439 105360
rect 211508 105302 214439 105304
rect 214373 105299 214439 105302
rect 227437 104954 227503 104957
rect 227437 104952 230092 104954
rect 227437 104896 227442 104952
rect 227498 104896 230092 104952
rect 227437 104894 230092 104896
rect 227437 104891 227503 104894
rect 215109 104546 215175 104549
rect 211508 104544 215175 104546
rect 211508 104488 215114 104544
rect 215170 104488 215175 104544
rect 211508 104486 215175 104488
rect 215109 104483 215175 104486
rect 116393 104410 116459 104413
rect 226241 104410 226307 104413
rect 116393 104408 119692 104410
rect 116393 104352 116398 104408
rect 116454 104352 119692 104408
rect 116393 104350 119692 104352
rect 226241 104408 230092 104410
rect 226241 104352 226246 104408
rect 226302 104352 230092 104408
rect 226241 104350 230092 104352
rect 116393 104347 116459 104350
rect 226241 104347 226307 104350
rect 214373 103866 214439 103869
rect 211508 103864 214439 103866
rect 211508 103808 214378 103864
rect 214434 103808 214439 103864
rect 211508 103806 214439 103808
rect 214373 103803 214439 103806
rect 227437 103866 227503 103869
rect 227437 103864 230092 103866
rect 227437 103808 227442 103864
rect 227498 103808 230092 103864
rect 227437 103806 230092 103808
rect 227437 103803 227503 103806
rect 116301 103186 116367 103189
rect 116301 103184 119692 103186
rect 116301 103128 116306 103184
rect 116362 103128 119692 103184
rect 116301 103126 119692 103128
rect 116301 103123 116367 103126
rect 215201 103050 215267 103053
rect 211508 103048 215267 103050
rect 211508 102992 215206 103048
rect 215262 102992 215267 103048
rect 211508 102990 215267 102992
rect 215201 102987 215267 102990
rect 215109 102234 215175 102237
rect 211508 102232 215175 102234
rect 211508 102176 215114 102232
rect 215170 102176 215175 102232
rect 211508 102174 215175 102176
rect 215109 102171 215175 102174
rect 116669 102098 116735 102101
rect 116669 102096 119692 102098
rect 116669 102040 116674 102096
rect 116730 102040 119692 102096
rect 116669 102038 119692 102040
rect 116669 102035 116735 102038
rect 215109 101418 215175 101421
rect 211508 101416 215175 101418
rect 211508 101360 215114 101416
rect 215170 101360 215175 101416
rect 211508 101358 215175 101360
rect 215109 101355 215175 101358
rect 116393 100874 116459 100877
rect 116393 100872 119692 100874
rect 116393 100816 116398 100872
rect 116454 100816 119692 100872
rect 116393 100814 119692 100816
rect 116393 100811 116459 100814
rect 215109 100602 215175 100605
rect 211508 100600 215175 100602
rect 211508 100544 215114 100600
rect 215170 100544 215175 100600
rect 211508 100542 215175 100544
rect 215109 100539 215175 100542
rect 214465 99922 214531 99925
rect 211508 99920 214531 99922
rect 211508 99864 214470 99920
rect 214526 99864 214531 99920
rect 211508 99862 214531 99864
rect 214465 99859 214531 99862
rect 116393 99786 116459 99789
rect 116393 99784 119692 99786
rect 116393 99728 116398 99784
rect 116454 99728 119692 99784
rect 116393 99726 119692 99728
rect 116393 99723 116459 99726
rect 583520 99636 584960 99876
rect 215109 99106 215175 99109
rect 211508 99104 215175 99106
rect 211508 99048 215114 99104
rect 215170 99048 215175 99104
rect 211508 99046 215175 99048
rect 215109 99043 215175 99046
rect 95141 98970 95207 98973
rect 91908 98968 95207 98970
rect 91908 98912 95146 98968
rect 95202 98912 95207 98968
rect 91908 98910 95207 98912
rect 95141 98907 95207 98910
rect 116393 98562 116459 98565
rect 116393 98560 119692 98562
rect 116393 98504 116398 98560
rect 116454 98504 119692 98560
rect 116393 98502 119692 98504
rect 116393 98499 116459 98502
rect 214649 98290 214715 98293
rect 211508 98288 214715 98290
rect 211508 98232 214654 98288
rect 214710 98232 214715 98288
rect 211508 98230 214715 98232
rect 214649 98227 214715 98230
rect 94773 98018 94839 98021
rect 91908 98016 94839 98018
rect 91908 97960 94778 98016
rect 94834 97960 94839 98016
rect 91908 97958 94839 97960
rect 94773 97955 94839 97958
rect 214097 97474 214163 97477
rect 211508 97472 214163 97474
rect 211508 97416 214102 97472
rect 214158 97416 214163 97472
rect 211508 97414 214163 97416
rect 214097 97411 214163 97414
rect 116393 97338 116459 97341
rect 116393 97336 119692 97338
rect 116393 97280 116398 97336
rect 116454 97280 119692 97336
rect 116393 97278 119692 97280
rect 116393 97275 116459 97278
rect 94681 97202 94747 97205
rect 91908 97200 94747 97202
rect 91908 97144 94686 97200
rect 94742 97144 94747 97200
rect 91908 97142 94747 97144
rect 94681 97139 94747 97142
rect 214557 96794 214623 96797
rect 211508 96792 214623 96794
rect 211508 96736 214562 96792
rect 214618 96736 214623 96792
rect 211508 96734 214623 96736
rect 214557 96731 214623 96734
rect 94865 96250 94931 96253
rect 91908 96248 94931 96250
rect 91908 96192 94870 96248
rect 94926 96192 94931 96248
rect 91908 96190 94931 96192
rect 94865 96187 94931 96190
rect 116301 96250 116367 96253
rect 116301 96248 119692 96250
rect 116301 96192 116306 96248
rect 116362 96192 119692 96248
rect 116301 96190 119692 96192
rect 116301 96187 116367 96190
rect 214281 95978 214347 95981
rect 211508 95976 214347 95978
rect 211508 95920 214286 95976
rect 214342 95920 214347 95976
rect 211508 95918 214347 95920
rect 214281 95915 214347 95918
rect 94589 95434 94655 95437
rect 91908 95432 94655 95434
rect 91908 95376 94594 95432
rect 94650 95376 94655 95432
rect 91908 95374 94655 95376
rect 94589 95371 94655 95374
rect 214741 95162 214807 95165
rect 211508 95160 214807 95162
rect 211508 95104 214746 95160
rect 214802 95104 214807 95160
rect 211508 95102 214807 95104
rect 214741 95099 214807 95102
rect 116577 95026 116643 95029
rect 116577 95024 119692 95026
rect 116577 94968 116582 95024
rect 116638 94968 119692 95024
rect 116577 94966 119692 94968
rect 116577 94963 116643 94966
rect 94497 94482 94563 94485
rect 91908 94480 94563 94482
rect 91908 94424 94502 94480
rect 94558 94424 94563 94480
rect 91908 94422 94563 94424
rect 94497 94419 94563 94422
rect 215109 94346 215175 94349
rect 211508 94344 215175 94346
rect 211508 94288 215114 94344
rect 215170 94288 215175 94344
rect 211508 94286 215175 94288
rect 215109 94283 215175 94286
rect 116393 93938 116459 93941
rect 116393 93936 119692 93938
rect 116393 93880 116398 93936
rect 116454 93880 119692 93936
rect 116393 93878 119692 93880
rect 116393 93875 116459 93878
rect 215109 93666 215175 93669
rect 211508 93664 215175 93666
rect 211508 93608 215114 93664
rect 215170 93608 215175 93664
rect 211508 93606 215175 93608
rect 215109 93603 215175 93606
rect 94865 93530 94931 93533
rect 91908 93528 94931 93530
rect 91908 93472 94870 93528
rect 94926 93472 94931 93528
rect 91908 93470 94931 93472
rect 94865 93467 94931 93470
rect -960 93258 480 93348
rect 2773 93258 2839 93261
rect -960 93256 2839 93258
rect -960 93200 2778 93256
rect 2834 93200 2839 93256
rect -960 93198 2839 93200
rect -960 93108 480 93198
rect 2773 93195 2839 93198
rect 215201 92850 215267 92853
rect 211508 92848 215267 92850
rect 211508 92792 215206 92848
rect 215262 92792 215267 92848
rect 211508 92790 215267 92792
rect 215201 92787 215267 92790
rect 94405 92714 94471 92717
rect 91908 92712 94471 92714
rect 91908 92656 94410 92712
rect 94466 92656 94471 92712
rect 91908 92654 94471 92656
rect 94405 92651 94471 92654
rect 116393 92714 116459 92717
rect 116393 92712 119692 92714
rect 116393 92656 116398 92712
rect 116454 92656 119692 92712
rect 116393 92654 119692 92656
rect 116393 92651 116459 92654
rect 214557 92034 214623 92037
rect 211508 92032 214623 92034
rect 211508 91976 214562 92032
rect 214618 91976 214623 92032
rect 211508 91974 214623 91976
rect 214557 91971 214623 91974
rect 95141 91762 95207 91765
rect 91908 91760 95207 91762
rect 91908 91704 95146 91760
rect 95202 91704 95207 91760
rect 91908 91702 95207 91704
rect 95141 91699 95207 91702
rect 116393 91626 116459 91629
rect 116393 91624 119692 91626
rect 116393 91568 116398 91624
rect 116454 91568 119692 91624
rect 116393 91566 119692 91568
rect 116393 91563 116459 91566
rect 214741 91218 214807 91221
rect 211508 91216 214807 91218
rect 211508 91160 214746 91216
rect 214802 91160 214807 91216
rect 211508 91158 214807 91160
rect 214741 91155 214807 91158
rect 94957 90946 95023 90949
rect 91908 90944 95023 90946
rect 91908 90888 94962 90944
rect 95018 90888 95023 90944
rect 91908 90886 95023 90888
rect 94957 90883 95023 90886
rect 214465 90538 214531 90541
rect 211508 90536 214531 90538
rect 211508 90480 214470 90536
rect 214526 90480 214531 90536
rect 211508 90478 214531 90480
rect 214465 90475 214531 90478
rect 116393 90402 116459 90405
rect 116393 90400 119692 90402
rect 116393 90344 116398 90400
rect 116454 90344 119692 90400
rect 116393 90342 119692 90344
rect 116393 90339 116459 90342
rect 95049 89994 95115 89997
rect 91908 89992 95115 89994
rect 91908 89936 95054 89992
rect 95110 89936 95115 89992
rect 91908 89934 95115 89936
rect 95049 89931 95115 89934
rect 215109 89722 215175 89725
rect 211508 89720 215175 89722
rect 211508 89664 215114 89720
rect 215170 89664 215175 89720
rect 211508 89662 215175 89664
rect 215109 89659 215175 89662
rect 95141 89178 95207 89181
rect 91908 89176 95207 89178
rect 91908 89120 95146 89176
rect 95202 89120 95207 89176
rect 91908 89118 95207 89120
rect 95141 89115 95207 89118
rect 115933 89178 115999 89181
rect 115933 89176 119692 89178
rect 115933 89120 115938 89176
rect 115994 89120 119692 89176
rect 115933 89118 119692 89120
rect 115933 89115 115999 89118
rect 214097 88906 214163 88909
rect 211508 88904 214163 88906
rect 211508 88848 214102 88904
rect 214158 88848 214163 88904
rect 211508 88846 214163 88848
rect 214097 88843 214163 88846
rect 95141 88226 95207 88229
rect 91908 88224 95207 88226
rect 91908 88168 95146 88224
rect 95202 88168 95207 88224
rect 91908 88166 95207 88168
rect 95141 88163 95207 88166
rect 116393 88090 116459 88093
rect 215017 88090 215083 88093
rect 116393 88088 119692 88090
rect 116393 88032 116398 88088
rect 116454 88032 119692 88088
rect 116393 88030 119692 88032
rect 211508 88088 215083 88090
rect 211508 88032 215022 88088
rect 215078 88032 215083 88088
rect 211508 88030 215083 88032
rect 116393 88027 116459 88030
rect 215017 88027 215083 88030
rect 580165 87954 580231 87957
rect 583520 87954 584960 88044
rect 580165 87952 584960 87954
rect 580165 87896 580170 87952
rect 580226 87896 584960 87952
rect 580165 87894 584960 87896
rect 580165 87891 580231 87894
rect 583520 87804 584960 87894
rect 215109 87410 215175 87413
rect 211508 87408 215175 87410
rect 211508 87352 215114 87408
rect 215170 87352 215175 87408
rect 211508 87350 215175 87352
rect 215109 87347 215175 87350
rect 94405 87274 94471 87277
rect 91908 87272 94471 87274
rect 91908 87216 94410 87272
rect 94466 87216 94471 87272
rect 91908 87214 94471 87216
rect 94405 87211 94471 87214
rect 116117 86866 116183 86869
rect 116117 86864 119692 86866
rect 116117 86808 116122 86864
rect 116178 86808 119692 86864
rect 116117 86806 119692 86808
rect 116117 86803 116183 86806
rect 215201 86594 215267 86597
rect 211508 86592 215267 86594
rect 211508 86536 215206 86592
rect 215262 86536 215267 86592
rect 211508 86534 215267 86536
rect 215201 86531 215267 86534
rect 94497 86458 94563 86461
rect 91908 86456 94563 86458
rect 91908 86400 94502 86456
rect 94558 86400 94563 86456
rect 91908 86398 94563 86400
rect 94497 86395 94563 86398
rect 116393 85778 116459 85781
rect 215109 85778 215175 85781
rect 116393 85776 119692 85778
rect 116393 85720 116398 85776
rect 116454 85720 119692 85776
rect 116393 85718 119692 85720
rect 211508 85776 215175 85778
rect 211508 85720 215114 85776
rect 215170 85720 215175 85776
rect 211508 85718 215175 85720
rect 116393 85715 116459 85718
rect 215109 85715 215175 85718
rect 94865 85506 94931 85509
rect 91908 85504 94931 85506
rect 91908 85448 94870 85504
rect 94926 85448 94931 85504
rect 91908 85446 94931 85448
rect 94865 85443 94931 85446
rect 214649 84962 214715 84965
rect 211508 84960 214715 84962
rect 211508 84904 214654 84960
rect 214710 84904 214715 84960
rect 211508 84902 214715 84904
rect 214649 84899 214715 84902
rect 95141 84690 95207 84693
rect 91908 84688 95207 84690
rect 91908 84632 95146 84688
rect 95202 84632 95207 84688
rect 91908 84630 95207 84632
rect 95141 84627 95207 84630
rect 117037 84554 117103 84557
rect 117037 84552 119692 84554
rect 117037 84496 117042 84552
rect 117098 84496 119692 84552
rect 117037 84494 119692 84496
rect 117037 84491 117103 84494
rect 215201 84282 215267 84285
rect 211508 84280 215267 84282
rect 211508 84224 215206 84280
rect 215262 84224 215267 84280
rect 211508 84222 215267 84224
rect 215201 84219 215267 84222
rect 94037 83738 94103 83741
rect 91908 83736 94103 83738
rect 91908 83680 94042 83736
rect 94098 83680 94103 83736
rect 91908 83678 94103 83680
rect 94037 83675 94103 83678
rect 214833 83466 214899 83469
rect 211508 83464 214899 83466
rect 211508 83408 214838 83464
rect 214894 83408 214899 83464
rect 211508 83406 214899 83408
rect 214833 83403 214899 83406
rect 116393 83330 116459 83333
rect 116393 83328 119692 83330
rect 116393 83272 116398 83328
rect 116454 83272 119692 83328
rect 116393 83270 119692 83272
rect 116393 83267 116459 83270
rect 94221 82922 94287 82925
rect 91908 82920 94287 82922
rect 91908 82864 94226 82920
rect 94282 82864 94287 82920
rect 91908 82862 94287 82864
rect 94221 82859 94287 82862
rect 214189 82650 214255 82653
rect 211508 82648 214255 82650
rect 211508 82592 214194 82648
rect 214250 82592 214255 82648
rect 211508 82590 214255 82592
rect 214189 82587 214255 82590
rect 115933 82242 115999 82245
rect 115933 82240 119692 82242
rect 115933 82184 115938 82240
rect 115994 82184 119692 82240
rect 115933 82182 119692 82184
rect 115933 82179 115999 82182
rect 95141 81970 95207 81973
rect 91908 81968 95207 81970
rect 91908 81912 95146 81968
rect 95202 81912 95207 81968
rect 91908 81910 95207 81912
rect 95141 81907 95207 81910
rect 214925 81834 214991 81837
rect 211508 81832 214991 81834
rect 211508 81776 214930 81832
rect 214986 81776 214991 81832
rect 211508 81774 214991 81776
rect 214925 81771 214991 81774
rect 227437 81154 227503 81157
rect 227437 81152 230092 81154
rect 227437 81096 227442 81152
rect 227498 81096 230092 81152
rect 227437 81094 230092 81096
rect 227437 81091 227503 81094
rect 94405 81018 94471 81021
rect 91908 81016 94471 81018
rect 91908 80960 94410 81016
rect 94466 80960 94471 81016
rect 91908 80958 94471 80960
rect 94405 80955 94471 80958
rect 116393 81018 116459 81021
rect 214005 81018 214071 81021
rect 116393 81016 119692 81018
rect 116393 80960 116398 81016
rect 116454 80960 119692 81016
rect 116393 80958 119692 80960
rect 211508 81016 214071 81018
rect 211508 80960 214010 81016
rect 214066 80960 214071 81016
rect 211508 80958 214071 80960
rect 116393 80955 116459 80958
rect 214005 80955 214071 80958
rect 227529 80474 227595 80477
rect 227529 80472 230092 80474
rect 227529 80416 227534 80472
rect 227590 80416 230092 80472
rect 227529 80414 230092 80416
rect 227529 80411 227595 80414
rect 215017 80338 215083 80341
rect 211508 80336 215083 80338
rect 211508 80280 215022 80336
rect 215078 80280 215083 80336
rect 211508 80278 215083 80280
rect 215017 80275 215083 80278
rect 94681 80202 94747 80205
rect 91908 80200 94747 80202
rect 91908 80144 94686 80200
rect 94742 80144 94747 80200
rect 91908 80142 94747 80144
rect 94681 80139 94747 80142
rect 116393 79930 116459 79933
rect 116393 79928 119692 79930
rect 116393 79872 116398 79928
rect 116454 79872 119692 79928
rect 116393 79870 119692 79872
rect 116393 79867 116459 79870
rect 227345 79794 227411 79797
rect 227345 79792 230092 79794
rect 227345 79736 227350 79792
rect 227406 79736 230092 79792
rect 227345 79734 230092 79736
rect 227345 79731 227411 79734
rect 215109 79522 215175 79525
rect 211508 79520 215175 79522
rect 211508 79464 215114 79520
rect 215170 79464 215175 79520
rect 211508 79462 215175 79464
rect 215109 79459 215175 79462
rect 95141 79250 95207 79253
rect 91908 79248 95207 79250
rect 91908 79192 95146 79248
rect 95202 79192 95207 79248
rect 91908 79190 95207 79192
rect 95141 79187 95207 79190
rect 227437 79114 227503 79117
rect 227437 79112 230092 79114
rect -960 78828 480 79068
rect 227437 79056 227442 79112
rect 227498 79056 230092 79112
rect 227437 79054 230092 79056
rect 227437 79051 227503 79054
rect 116577 78706 116643 78709
rect 214557 78706 214623 78709
rect 116577 78704 119692 78706
rect 116577 78648 116582 78704
rect 116638 78648 119692 78704
rect 116577 78646 119692 78648
rect 211508 78704 214623 78706
rect 211508 78648 214562 78704
rect 214618 78648 214623 78704
rect 211508 78646 214623 78648
rect 116577 78643 116643 78646
rect 214557 78643 214623 78646
rect 227437 78570 227503 78573
rect 227437 78568 230092 78570
rect 227437 78512 227442 78568
rect 227498 78512 230092 78568
rect 227437 78510 230092 78512
rect 227437 78507 227503 78510
rect 94589 78434 94655 78437
rect 91908 78432 94655 78434
rect 91908 78376 94594 78432
rect 94650 78376 94655 78432
rect 91908 78374 94655 78376
rect 94589 78371 94655 78374
rect 214741 77890 214807 77893
rect 211508 77888 214807 77890
rect 211508 77832 214746 77888
rect 214802 77832 214807 77888
rect 211508 77830 214807 77832
rect 214741 77827 214807 77830
rect 227529 77890 227595 77893
rect 227529 77888 230092 77890
rect 227529 77832 227534 77888
rect 227590 77832 230092 77888
rect 227529 77830 230092 77832
rect 227529 77827 227595 77830
rect 94405 77482 94471 77485
rect 91908 77480 94471 77482
rect 91908 77424 94410 77480
rect 94466 77424 94471 77480
rect 91908 77422 94471 77424
rect 94405 77419 94471 77422
rect 116393 77482 116459 77485
rect 116393 77480 119692 77482
rect 116393 77424 116398 77480
rect 116454 77424 119692 77480
rect 116393 77422 119692 77424
rect 116393 77419 116459 77422
rect 214465 77210 214531 77213
rect 211508 77208 214531 77210
rect 211508 77152 214470 77208
rect 214526 77152 214531 77208
rect 211508 77150 214531 77152
rect 214465 77147 214531 77150
rect 227437 77210 227503 77213
rect 227437 77208 230092 77210
rect 227437 77152 227442 77208
rect 227498 77152 230092 77208
rect 227437 77150 230092 77152
rect 227437 77147 227503 77150
rect 94221 76530 94287 76533
rect 91908 76528 94287 76530
rect 91908 76472 94226 76528
rect 94282 76472 94287 76528
rect 91908 76470 94287 76472
rect 94221 76467 94287 76470
rect 227529 76530 227595 76533
rect 227529 76528 230092 76530
rect 227529 76472 227534 76528
rect 227590 76472 230092 76528
rect 227529 76470 230092 76472
rect 227529 76467 227595 76470
rect 116393 76394 116459 76397
rect 215201 76394 215267 76397
rect 116393 76392 119692 76394
rect 116393 76336 116398 76392
rect 116454 76336 119692 76392
rect 116393 76334 119692 76336
rect 211508 76392 215267 76394
rect 211508 76336 215206 76392
rect 215262 76336 215267 76392
rect 211508 76334 215267 76336
rect 116393 76331 116459 76334
rect 215201 76331 215267 76334
rect 580901 76258 580967 76261
rect 583520 76258 584960 76348
rect 580901 76256 584960 76258
rect 580901 76200 580906 76256
rect 580962 76200 584960 76256
rect 580901 76198 584960 76200
rect 580901 76195 580967 76198
rect 583520 76108 584960 76198
rect 225597 75850 225663 75853
rect 225597 75848 230092 75850
rect 225597 75792 225602 75848
rect 225658 75792 230092 75848
rect 225597 75790 230092 75792
rect 225597 75787 225663 75790
rect 94589 75714 94655 75717
rect 91908 75712 94655 75714
rect 91908 75656 94594 75712
rect 94650 75656 94655 75712
rect 91908 75654 94655 75656
rect 94589 75651 94655 75654
rect 215109 75578 215175 75581
rect 211508 75576 215175 75578
rect 211508 75520 215114 75576
rect 215170 75520 215175 75576
rect 211508 75518 215175 75520
rect 215109 75515 215175 75518
rect 227437 75306 227503 75309
rect 227437 75304 230092 75306
rect 227437 75248 227442 75304
rect 227498 75248 230092 75304
rect 227437 75246 230092 75248
rect 227437 75243 227503 75246
rect 116393 75170 116459 75173
rect 116393 75168 119692 75170
rect 116393 75112 116398 75168
rect 116454 75112 119692 75168
rect 116393 75110 119692 75112
rect 116393 75107 116459 75110
rect 94957 74762 95023 74765
rect 215201 74762 215267 74765
rect 91908 74760 95023 74762
rect 91908 74704 94962 74760
rect 95018 74704 95023 74760
rect 91908 74702 95023 74704
rect 211508 74760 215267 74762
rect 211508 74704 215206 74760
rect 215262 74704 215267 74760
rect 211508 74702 215267 74704
rect 94957 74699 95023 74702
rect 215201 74699 215267 74702
rect 227069 74626 227135 74629
rect 227069 74624 230092 74626
rect 227069 74568 227074 74624
rect 227130 74568 230092 74624
rect 227069 74566 230092 74568
rect 227069 74563 227135 74566
rect 116393 74082 116459 74085
rect 214281 74082 214347 74085
rect 116393 74080 119692 74082
rect 116393 74024 116398 74080
rect 116454 74024 119692 74080
rect 116393 74022 119692 74024
rect 211508 74080 214347 74082
rect 211508 74024 214286 74080
rect 214342 74024 214347 74080
rect 211508 74022 214347 74024
rect 116393 74019 116459 74022
rect 214281 74019 214347 74022
rect 95141 73946 95207 73949
rect 91908 73944 95207 73946
rect 91908 73888 95146 73944
rect 95202 73888 95207 73944
rect 91908 73886 95207 73888
rect 95141 73883 95207 73886
rect 227437 73946 227503 73949
rect 227437 73944 230092 73946
rect 227437 73888 227442 73944
rect 227498 73888 230092 73944
rect 227437 73886 230092 73888
rect 227437 73883 227503 73886
rect 215109 73266 215175 73269
rect 211508 73264 215175 73266
rect 211508 73208 215114 73264
rect 215170 73208 215175 73264
rect 211508 73206 215175 73208
rect 215109 73203 215175 73206
rect 227161 73266 227227 73269
rect 227161 73264 230092 73266
rect 227161 73208 227166 73264
rect 227222 73208 230092 73264
rect 227161 73206 230092 73208
rect 227161 73203 227227 73206
rect 94037 72994 94103 72997
rect 91908 72992 94103 72994
rect 91908 72936 94042 72992
rect 94098 72936 94103 72992
rect 91908 72934 94103 72936
rect 94037 72931 94103 72934
rect 116393 72858 116459 72861
rect 116393 72856 119692 72858
rect 116393 72800 116398 72856
rect 116454 72800 119692 72856
rect 116393 72798 119692 72800
rect 116393 72795 116459 72798
rect 227437 72722 227503 72725
rect 227437 72720 230092 72722
rect 227437 72664 227442 72720
rect 227498 72664 230092 72720
rect 227437 72662 230092 72664
rect 227437 72659 227503 72662
rect 214649 72450 214715 72453
rect 211508 72448 214715 72450
rect 211508 72392 214654 72448
rect 214710 72392 214715 72448
rect 211508 72390 214715 72392
rect 214649 72387 214715 72390
rect 94405 72178 94471 72181
rect 91908 72176 94471 72178
rect 91908 72120 94410 72176
rect 94466 72120 94471 72176
rect 91908 72118 94471 72120
rect 94405 72115 94471 72118
rect 227529 72042 227595 72045
rect 227529 72040 230092 72042
rect 227529 71984 227534 72040
rect 227590 71984 230092 72040
rect 227529 71982 230092 71984
rect 227529 71979 227595 71982
rect 116301 71770 116367 71773
rect 116301 71768 119692 71770
rect 116301 71712 116306 71768
rect 116362 71712 119692 71768
rect 116301 71710 119692 71712
rect 116301 71707 116367 71710
rect 214097 71634 214163 71637
rect 211508 71632 214163 71634
rect 211508 71576 214102 71632
rect 214158 71576 214163 71632
rect 211508 71574 214163 71576
rect 214097 71571 214163 71574
rect 227437 71362 227503 71365
rect 227437 71360 230092 71362
rect 227437 71304 227442 71360
rect 227498 71304 230092 71360
rect 227437 71302 230092 71304
rect 227437 71299 227503 71302
rect 94221 71226 94287 71229
rect 91908 71224 94287 71226
rect 91908 71168 94226 71224
rect 94282 71168 94287 71224
rect 91908 71166 94287 71168
rect 94221 71163 94287 71166
rect 215109 70954 215175 70957
rect 211508 70952 215175 70954
rect 211508 70896 215114 70952
rect 215170 70896 215175 70952
rect 211508 70894 215175 70896
rect 215109 70891 215175 70894
rect 227529 70682 227595 70685
rect 227529 70680 230092 70682
rect 227529 70624 227534 70680
rect 227590 70624 230092 70680
rect 227529 70622 230092 70624
rect 227529 70619 227595 70622
rect 116393 70546 116459 70549
rect 116393 70544 119692 70546
rect 116393 70488 116398 70544
rect 116454 70488 119692 70544
rect 116393 70486 119692 70488
rect 116393 70483 116459 70486
rect 94865 70274 94931 70277
rect 91908 70272 94931 70274
rect 91908 70216 94870 70272
rect 94926 70216 94931 70272
rect 91908 70214 94931 70216
rect 94865 70211 94931 70214
rect 214925 70138 214991 70141
rect 211508 70136 214991 70138
rect 211508 70080 214930 70136
rect 214986 70080 214991 70136
rect 211508 70078 214991 70080
rect 214925 70075 214991 70078
rect 227437 70002 227503 70005
rect 227437 70000 230092 70002
rect 227437 69944 227442 70000
rect 227498 69944 230092 70000
rect 227437 69942 230092 69944
rect 227437 69939 227503 69942
rect 95049 69458 95115 69461
rect 91908 69456 95115 69458
rect 91908 69400 95054 69456
rect 95110 69400 95115 69456
rect 91908 69398 95115 69400
rect 95049 69395 95115 69398
rect 226517 69458 226583 69461
rect 226517 69456 230092 69458
rect 226517 69400 226522 69456
rect 226578 69400 230092 69456
rect 226517 69398 230092 69400
rect 226517 69395 226583 69398
rect 116393 69322 116459 69325
rect 215109 69322 215175 69325
rect 116393 69320 119692 69322
rect 116393 69264 116398 69320
rect 116454 69264 119692 69320
rect 116393 69262 119692 69264
rect 211508 69320 215175 69322
rect 211508 69264 215114 69320
rect 215170 69264 215175 69320
rect 211508 69262 215175 69264
rect 116393 69259 116459 69262
rect 215109 69259 215175 69262
rect 227437 68778 227503 68781
rect 227437 68776 230092 68778
rect 227437 68720 227442 68776
rect 227498 68720 230092 68776
rect 227437 68718 230092 68720
rect 227437 68715 227503 68718
rect 94037 68506 94103 68509
rect 215201 68506 215267 68509
rect 91908 68504 94103 68506
rect 91908 68448 94042 68504
rect 94098 68448 94103 68504
rect 91908 68446 94103 68448
rect 211508 68504 215267 68506
rect 211508 68448 215206 68504
rect 215262 68448 215267 68504
rect 211508 68446 215267 68448
rect 94037 68443 94103 68446
rect 215201 68443 215267 68446
rect 116393 68234 116459 68237
rect 116393 68232 119692 68234
rect 116393 68176 116398 68232
rect 116454 68176 119692 68232
rect 116393 68174 119692 68176
rect 116393 68171 116459 68174
rect 227529 68098 227595 68101
rect 227529 68096 230092 68098
rect 227529 68040 227534 68096
rect 227590 68040 230092 68096
rect 227529 68038 230092 68040
rect 227529 68035 227595 68038
rect 215109 67826 215175 67829
rect 211508 67824 215175 67826
rect 211508 67768 215114 67824
rect 215170 67768 215175 67824
rect 211508 67766 215175 67768
rect 215109 67763 215175 67766
rect 95141 67690 95207 67693
rect 91908 67688 95207 67690
rect 91908 67632 95146 67688
rect 95202 67632 95207 67688
rect 91908 67630 95207 67632
rect 95141 67627 95207 67630
rect 227437 67418 227503 67421
rect 227437 67416 230092 67418
rect 227437 67360 227442 67416
rect 227498 67360 230092 67416
rect 227437 67358 230092 67360
rect 227437 67355 227503 67358
rect 116393 67010 116459 67013
rect 215109 67010 215175 67013
rect 116393 67008 119692 67010
rect 116393 66952 116398 67008
rect 116454 66952 119692 67008
rect 116393 66950 119692 66952
rect 211508 67008 215175 67010
rect 211508 66952 215114 67008
rect 215170 66952 215175 67008
rect 211508 66950 215175 66952
rect 116393 66947 116459 66950
rect 215109 66947 215175 66950
rect 227529 66874 227595 66877
rect 227529 66872 230092 66874
rect 227529 66816 227534 66872
rect 227590 66816 230092 66872
rect 227529 66814 230092 66816
rect 227529 66811 227595 66814
rect 95141 66738 95207 66741
rect 91908 66736 95207 66738
rect 91908 66680 95146 66736
rect 95202 66680 95207 66736
rect 91908 66678 95207 66680
rect 95141 66675 95207 66678
rect 213913 66194 213979 66197
rect 211508 66192 213979 66194
rect 211508 66136 213918 66192
rect 213974 66136 213979 66192
rect 211508 66134 213979 66136
rect 213913 66131 213979 66134
rect 227437 66194 227503 66197
rect 227437 66192 230092 66194
rect 227437 66136 227442 66192
rect 227498 66136 230092 66192
rect 227437 66134 230092 66136
rect 227437 66131 227503 66134
rect 94129 65922 94195 65925
rect 91908 65920 94195 65922
rect 91908 65864 94134 65920
rect 94190 65864 94195 65920
rect 91908 65862 94195 65864
rect 94129 65859 94195 65862
rect 116393 65922 116459 65925
rect 116393 65920 119692 65922
rect 116393 65864 116398 65920
rect 116454 65864 119692 65920
rect 116393 65862 119692 65864
rect 116393 65859 116459 65862
rect 6177 65514 6243 65517
rect 227529 65514 227595 65517
rect 6177 65512 9292 65514
rect 6177 65456 6182 65512
rect 6238 65456 9292 65512
rect 6177 65454 9292 65456
rect 227529 65512 230092 65514
rect 227529 65456 227534 65512
rect 227590 65456 230092 65512
rect 227529 65454 230092 65456
rect 6177 65451 6243 65454
rect 227529 65451 227595 65454
rect 214005 65378 214071 65381
rect 211508 65376 214071 65378
rect 211508 65320 214010 65376
rect 214066 65320 214071 65376
rect 211508 65318 214071 65320
rect 214005 65315 214071 65318
rect 94405 64970 94471 64973
rect 91908 64968 94471 64970
rect 91908 64912 94410 64968
rect 94466 64912 94471 64968
rect 91908 64910 94471 64912
rect 94405 64907 94471 64910
rect 227253 64834 227319 64837
rect 227253 64832 230092 64834
rect 227253 64776 227258 64832
rect 227314 64776 230092 64832
rect 227253 64774 230092 64776
rect 227253 64771 227319 64774
rect 115933 64698 115999 64701
rect 115933 64696 119692 64698
rect -960 64562 480 64652
rect 115933 64640 115938 64696
rect 115994 64640 119692 64696
rect 115933 64638 119692 64640
rect 115933 64635 115999 64638
rect 2773 64562 2839 64565
rect 214097 64562 214163 64565
rect -960 64560 2839 64562
rect -960 64504 2778 64560
rect 2834 64504 2839 64560
rect -960 64502 2839 64504
rect 211508 64560 214163 64562
rect 211508 64504 214102 64560
rect 214158 64504 214163 64560
rect 211508 64502 214163 64504
rect -960 64412 480 64502
rect 2773 64499 2839 64502
rect 214097 64499 214163 64502
rect 583520 64412 584960 64652
rect 227437 64154 227503 64157
rect 227437 64152 230092 64154
rect 227437 64096 227442 64152
rect 227498 64096 230092 64152
rect 227437 64094 230092 64096
rect 227437 64091 227503 64094
rect 94589 64018 94655 64021
rect 91908 64016 94655 64018
rect 91908 63960 94594 64016
rect 94650 63960 94655 64016
rect 91908 63958 94655 63960
rect 94589 63955 94655 63958
rect 215109 63882 215175 63885
rect 211508 63880 215175 63882
rect 211508 63824 215114 63880
rect 215170 63824 215175 63880
rect 211508 63822 215175 63824
rect 215109 63819 215175 63822
rect 227529 63610 227595 63613
rect 227529 63608 230092 63610
rect 227529 63552 227534 63608
rect 227590 63552 230092 63608
rect 227529 63550 230092 63552
rect 227529 63547 227595 63550
rect 116393 63474 116459 63477
rect 116393 63472 119692 63474
rect 116393 63416 116398 63472
rect 116454 63416 119692 63472
rect 116393 63414 119692 63416
rect 116393 63411 116459 63414
rect 95141 63202 95207 63205
rect 91908 63200 95207 63202
rect 91908 63144 95146 63200
rect 95202 63144 95207 63200
rect 91908 63142 95207 63144
rect 95141 63139 95207 63142
rect 214373 63066 214439 63069
rect 211508 63064 214439 63066
rect 211508 63008 214378 63064
rect 214434 63008 214439 63064
rect 211508 63006 214439 63008
rect 214373 63003 214439 63006
rect 227437 62930 227503 62933
rect 227437 62928 230092 62930
rect 227437 62872 227442 62928
rect 227498 62872 230092 62928
rect 227437 62870 230092 62872
rect 227437 62867 227503 62870
rect 116485 62386 116551 62389
rect 116485 62384 119692 62386
rect 116485 62328 116490 62384
rect 116546 62328 119692 62384
rect 116485 62326 119692 62328
rect 116485 62323 116551 62326
rect 94773 62250 94839 62253
rect 215109 62250 215175 62253
rect 91908 62248 94839 62250
rect 91908 62192 94778 62248
rect 94834 62192 94839 62248
rect 91908 62190 94839 62192
rect 211508 62248 215175 62250
rect 211508 62192 215114 62248
rect 215170 62192 215175 62248
rect 211508 62190 215175 62192
rect 94773 62187 94839 62190
rect 215109 62187 215175 62190
rect 227069 62250 227135 62253
rect 227069 62248 230092 62250
rect 227069 62192 227074 62248
rect 227130 62192 230092 62248
rect 227069 62190 230092 62192
rect 227069 62187 227135 62190
rect 227437 61570 227503 61573
rect 227437 61568 230092 61570
rect 227437 61512 227442 61568
rect 227498 61512 230092 61568
rect 227437 61510 230092 61512
rect 227437 61507 227503 61510
rect 94313 61434 94379 61437
rect 214741 61434 214807 61437
rect 91908 61432 94379 61434
rect 91908 61376 94318 61432
rect 94374 61376 94379 61432
rect 91908 61374 94379 61376
rect 211508 61432 214807 61434
rect 211508 61376 214746 61432
rect 214802 61376 214807 61432
rect 211508 61374 214807 61376
rect 94313 61371 94379 61374
rect 214741 61371 214807 61374
rect 116393 61162 116459 61165
rect 116393 61160 119692 61162
rect 116393 61104 116398 61160
rect 116454 61104 119692 61160
rect 116393 61102 119692 61104
rect 116393 61099 116459 61102
rect 226701 61026 226767 61029
rect 226701 61024 230092 61026
rect 226701 60968 226706 61024
rect 226762 60968 230092 61024
rect 226701 60966 230092 60968
rect 226701 60963 226767 60966
rect 215109 60754 215175 60757
rect 211508 60752 215175 60754
rect 211508 60696 215114 60752
rect 215170 60696 215175 60752
rect 211508 60694 215175 60696
rect 215109 60691 215175 60694
rect 94497 60482 94563 60485
rect 91908 60480 94563 60482
rect 91908 60424 94502 60480
rect 94558 60424 94563 60480
rect 91908 60422 94563 60424
rect 94497 60419 94563 60422
rect 227437 60346 227503 60349
rect 227437 60344 230092 60346
rect 227437 60288 227442 60344
rect 227498 60288 230092 60344
rect 227437 60286 230092 60288
rect 227437 60283 227503 60286
rect 116393 60074 116459 60077
rect 116393 60072 119692 60074
rect 116393 60016 116398 60072
rect 116454 60016 119692 60072
rect 116393 60014 119692 60016
rect 116393 60011 116459 60014
rect 214373 59938 214439 59941
rect 211508 59936 214439 59938
rect 211508 59880 214378 59936
rect 214434 59880 214439 59936
rect 211508 59878 214439 59880
rect 214373 59875 214439 59878
rect 227529 59666 227595 59669
rect 227529 59664 230092 59666
rect 227529 59608 227534 59664
rect 227590 59608 230092 59664
rect 227529 59606 230092 59608
rect 227529 59603 227595 59606
rect 94313 59530 94379 59533
rect 91908 59528 94379 59530
rect 91908 59472 94318 59528
rect 94374 59472 94379 59528
rect 91908 59470 94379 59472
rect 94313 59467 94379 59470
rect 214281 59122 214347 59125
rect 211508 59120 214347 59122
rect 211508 59064 214286 59120
rect 214342 59064 214347 59120
rect 211508 59062 214347 59064
rect 214281 59059 214347 59062
rect 227437 58986 227503 58989
rect 227437 58984 230092 58986
rect 227437 58928 227442 58984
rect 227498 58928 230092 58984
rect 227437 58926 230092 58928
rect 227437 58923 227503 58926
rect 116393 58850 116459 58853
rect 116393 58848 119692 58850
rect 116393 58792 116398 58848
rect 116454 58792 119692 58848
rect 116393 58790 119692 58792
rect 116393 58787 116459 58790
rect 94681 58714 94747 58717
rect 91908 58712 94747 58714
rect 91908 58656 94686 58712
rect 94742 58656 94747 58712
rect 91908 58654 94747 58656
rect 94681 58651 94747 58654
rect 214373 58306 214439 58309
rect 211508 58304 214439 58306
rect 211508 58248 214378 58304
rect 214434 58248 214439 58304
rect 211508 58246 214439 58248
rect 214373 58243 214439 58246
rect 227529 58306 227595 58309
rect 227529 58304 230092 58306
rect 227529 58248 227534 58304
rect 227590 58248 230092 58304
rect 227529 58246 230092 58248
rect 227529 58243 227595 58246
rect 94405 57762 94471 57765
rect 91908 57760 94471 57762
rect 91908 57704 94410 57760
rect 94466 57704 94471 57760
rect 91908 57702 94471 57704
rect 94405 57699 94471 57702
rect 227253 57762 227319 57765
rect 227253 57760 230092 57762
rect 227253 57704 227258 57760
rect 227314 57704 230092 57760
rect 227253 57702 230092 57704
rect 227253 57699 227319 57702
rect 116301 57626 116367 57629
rect 213913 57626 213979 57629
rect 116301 57624 119692 57626
rect 116301 57568 116306 57624
rect 116362 57568 119692 57624
rect 116301 57566 119692 57568
rect 211508 57624 213979 57626
rect 211508 57568 213918 57624
rect 213974 57568 213979 57624
rect 211508 57566 213979 57568
rect 116301 57563 116367 57566
rect 213913 57563 213979 57566
rect 227437 57082 227503 57085
rect 227437 57080 230092 57082
rect 227437 57024 227442 57080
rect 227498 57024 230092 57080
rect 227437 57022 230092 57024
rect 227437 57019 227503 57022
rect 94865 56946 94931 56949
rect 91908 56944 94931 56946
rect 91908 56888 94870 56944
rect 94926 56888 94931 56944
rect 91908 56886 94931 56888
rect 94865 56883 94931 56886
rect 214005 56810 214071 56813
rect 211508 56808 214071 56810
rect 211508 56752 214010 56808
rect 214066 56752 214071 56808
rect 211508 56750 214071 56752
rect 214005 56747 214071 56750
rect 116301 56538 116367 56541
rect 116301 56536 119692 56538
rect 116301 56480 116306 56536
rect 116362 56480 119692 56536
rect 116301 56478 119692 56480
rect 116301 56475 116367 56478
rect 227253 56402 227319 56405
rect 227253 56400 230092 56402
rect 227253 56344 227258 56400
rect 227314 56344 230092 56400
rect 227253 56342 230092 56344
rect 227253 56339 227319 56342
rect 95141 55994 95207 55997
rect 215109 55994 215175 55997
rect 91908 55992 95207 55994
rect 91908 55936 95146 55992
rect 95202 55936 95207 55992
rect 91908 55934 95207 55936
rect 211508 55992 215175 55994
rect 211508 55936 215114 55992
rect 215170 55936 215175 55992
rect 211508 55934 215175 55936
rect 95141 55931 95207 55934
rect 215109 55931 215175 55934
rect 227437 55722 227503 55725
rect 227437 55720 230092 55722
rect 227437 55664 227442 55720
rect 227498 55664 230092 55720
rect 227437 55662 230092 55664
rect 227437 55659 227503 55662
rect 116393 55314 116459 55317
rect 116393 55312 119692 55314
rect 116393 55256 116398 55312
rect 116454 55256 119692 55312
rect 116393 55254 119692 55256
rect 116393 55251 116459 55254
rect 94589 55178 94655 55181
rect 214741 55178 214807 55181
rect 91908 55176 94655 55178
rect 91908 55120 94594 55176
rect 94650 55120 94655 55176
rect 91908 55118 94655 55120
rect 211508 55176 214807 55178
rect 211508 55120 214746 55176
rect 214802 55120 214807 55176
rect 211508 55118 214807 55120
rect 94589 55115 94655 55118
rect 214741 55115 214807 55118
rect 227437 55178 227503 55181
rect 227437 55176 230092 55178
rect 227437 55120 227442 55176
rect 227498 55120 230092 55176
rect 227437 55118 230092 55120
rect 227437 55115 227503 55118
rect 215109 54498 215175 54501
rect 211508 54496 215175 54498
rect 211508 54440 215114 54496
rect 215170 54440 215175 54496
rect 211508 54438 215175 54440
rect 215109 54435 215175 54438
rect 226517 54498 226583 54501
rect 226517 54496 230092 54498
rect 226517 54440 226522 54496
rect 226578 54440 230092 54496
rect 226517 54438 230092 54440
rect 226517 54435 226583 54438
rect 94589 54226 94655 54229
rect 91908 54224 94655 54226
rect 91908 54168 94594 54224
rect 94650 54168 94655 54224
rect 91908 54166 94655 54168
rect 94589 54163 94655 54166
rect 116393 54226 116459 54229
rect 116393 54224 119692 54226
rect 116393 54168 116398 54224
rect 116454 54168 119692 54224
rect 116393 54166 119692 54168
rect 116393 54163 116459 54166
rect 227253 53818 227319 53821
rect 227253 53816 230092 53818
rect 227253 53760 227258 53816
rect 227314 53760 230092 53816
rect 227253 53758 230092 53760
rect 227253 53755 227319 53758
rect 214741 53682 214807 53685
rect 211508 53680 214807 53682
rect 211508 53624 214746 53680
rect 214802 53624 214807 53680
rect 211508 53622 214807 53624
rect 214741 53619 214807 53622
rect 94773 53274 94839 53277
rect 91908 53272 94839 53274
rect 91908 53216 94778 53272
rect 94834 53216 94839 53272
rect 91908 53214 94839 53216
rect 94773 53211 94839 53214
rect 227437 53138 227503 53141
rect 227437 53136 230092 53138
rect 227437 53080 227442 53136
rect 227498 53080 230092 53136
rect 227437 53078 230092 53080
rect 227437 53075 227503 53078
rect 116393 53002 116459 53005
rect 116393 53000 119692 53002
rect 116393 52944 116398 53000
rect 116454 52944 119692 53000
rect 116393 52942 119692 52944
rect 116393 52939 116459 52942
rect 215109 52866 215175 52869
rect 211508 52864 215175 52866
rect 211508 52808 215114 52864
rect 215170 52808 215175 52864
rect 211508 52806 215175 52808
rect 215109 52803 215175 52806
rect 583520 52716 584960 52956
rect 95141 52458 95207 52461
rect 91908 52456 95207 52458
rect 91908 52400 95146 52456
rect 95202 52400 95207 52456
rect 91908 52398 95207 52400
rect 95141 52395 95207 52398
rect 227253 52458 227319 52461
rect 227253 52456 230092 52458
rect 227253 52400 227258 52456
rect 227314 52400 230092 52456
rect 227253 52398 230092 52400
rect 227253 52395 227319 52398
rect 214557 52050 214623 52053
rect 211508 52048 214623 52050
rect 211508 51992 214562 52048
rect 214618 51992 214623 52048
rect 211508 51990 214623 51992
rect 214557 51987 214623 51990
rect 115933 51914 115999 51917
rect 227437 51914 227503 51917
rect 115933 51912 119692 51914
rect 115933 51856 115938 51912
rect 115994 51856 119692 51912
rect 115933 51854 119692 51856
rect 227437 51912 230092 51914
rect 227437 51856 227442 51912
rect 227498 51856 230092 51912
rect 227437 51854 230092 51856
rect 115933 51851 115999 51854
rect 227437 51851 227503 51854
rect 94957 51506 95023 51509
rect 91908 51504 95023 51506
rect 91908 51448 94962 51504
rect 95018 51448 95023 51504
rect 91908 51446 95023 51448
rect 94957 51443 95023 51446
rect 215109 51370 215175 51373
rect 211508 51368 215175 51370
rect 211508 51312 215114 51368
rect 215170 51312 215175 51368
rect 211508 51310 215175 51312
rect 215109 51307 215175 51310
rect 227529 51234 227595 51237
rect 227529 51232 230092 51234
rect 227529 51176 227534 51232
rect 227590 51176 230092 51232
rect 227529 51174 230092 51176
rect 227529 51171 227595 51174
rect 95141 50690 95207 50693
rect 91908 50688 95207 50690
rect 91908 50632 95146 50688
rect 95202 50632 95207 50688
rect 91908 50630 95207 50632
rect 95141 50627 95207 50630
rect 116393 50690 116459 50693
rect 116393 50688 119692 50690
rect 116393 50632 116398 50688
rect 116454 50632 119692 50688
rect 116393 50630 119692 50632
rect 116393 50627 116459 50630
rect 214373 50554 214439 50557
rect 211508 50552 214439 50554
rect 211508 50496 214378 50552
rect 214434 50496 214439 50552
rect 211508 50494 214439 50496
rect 214373 50491 214439 50494
rect 226517 50554 226583 50557
rect 226517 50552 230092 50554
rect 226517 50496 226522 50552
rect 226578 50496 230092 50552
rect 226517 50494 230092 50496
rect 226517 50491 226583 50494
rect -960 50146 480 50236
rect 2773 50146 2839 50149
rect -960 50144 2839 50146
rect -960 50088 2778 50144
rect 2834 50088 2839 50144
rect -960 50086 2839 50088
rect -960 49996 480 50086
rect 2773 50083 2839 50086
rect 226977 49874 227043 49877
rect 411989 49874 412055 49877
rect 226977 49872 230092 49874
rect 226977 49816 226982 49872
rect 227038 49816 230092 49872
rect 226977 49814 230092 49816
rect 411989 49872 414092 49874
rect 411989 49816 411994 49872
rect 412050 49816 414092 49872
rect 411989 49814 414092 49816
rect 226977 49811 227043 49814
rect 411989 49811 412055 49814
rect 94037 49738 94103 49741
rect 215109 49738 215175 49741
rect 91908 49736 94103 49738
rect 91908 49680 94042 49736
rect 94098 49680 94103 49736
rect 91908 49678 94103 49680
rect 211508 49736 215175 49738
rect 211508 49680 215114 49736
rect 215170 49680 215175 49736
rect 211508 49678 215175 49680
rect 94037 49675 94103 49678
rect 215109 49675 215175 49678
rect 116393 49466 116459 49469
rect 116393 49464 119692 49466
rect 116393 49408 116398 49464
rect 116454 49408 119692 49464
rect 116393 49406 119692 49408
rect 116393 49403 116459 49406
rect 226701 49330 226767 49333
rect 226701 49328 230092 49330
rect 226701 49272 226706 49328
rect 226762 49272 230092 49328
rect 226701 49270 230092 49272
rect 226701 49267 226767 49270
rect 94129 48922 94195 48925
rect 215109 48922 215175 48925
rect 91908 48920 94195 48922
rect 91908 48864 94134 48920
rect 94190 48864 94195 48920
rect 91908 48862 94195 48864
rect 211508 48920 215175 48922
rect 211508 48864 215114 48920
rect 215170 48864 215175 48920
rect 211508 48862 215175 48864
rect 94129 48859 94195 48862
rect 215109 48859 215175 48862
rect 226793 48650 226859 48653
rect 226793 48648 230092 48650
rect 226793 48592 226798 48648
rect 226854 48592 230092 48648
rect 226793 48590 230092 48592
rect 226793 48587 226859 48590
rect 116117 48378 116183 48381
rect 116117 48376 119692 48378
rect 116117 48320 116122 48376
rect 116178 48320 119692 48376
rect 116117 48318 119692 48320
rect 116117 48315 116183 48318
rect 214741 48106 214807 48109
rect 211508 48104 214807 48106
rect 211508 48048 214746 48104
rect 214802 48048 214807 48104
rect 211508 48046 214807 48048
rect 214741 48043 214807 48046
rect 94865 47970 94931 47973
rect 91908 47968 94931 47970
rect 91908 47912 94870 47968
rect 94926 47912 94931 47968
rect 91908 47910 94931 47912
rect 94865 47907 94931 47910
rect 226333 47970 226399 47973
rect 226333 47968 230092 47970
rect 226333 47912 226338 47968
rect 226394 47912 230092 47968
rect 226333 47910 230092 47912
rect 226333 47907 226399 47910
rect 214005 47426 214071 47429
rect 211508 47424 214071 47426
rect 211508 47368 214010 47424
rect 214066 47368 214071 47424
rect 211508 47366 214071 47368
rect 214005 47363 214071 47366
rect 226609 47290 226675 47293
rect 226609 47288 230092 47290
rect 226609 47232 226614 47288
rect 226670 47232 230092 47288
rect 226609 47230 230092 47232
rect 226609 47227 226675 47230
rect 116393 47154 116459 47157
rect 116393 47152 119692 47154
rect 116393 47096 116398 47152
rect 116454 47096 119692 47152
rect 116393 47094 119692 47096
rect 116393 47091 116459 47094
rect 94773 47018 94839 47021
rect 91908 47016 94839 47018
rect 91908 46960 94778 47016
rect 94834 46960 94839 47016
rect 91908 46958 94839 46960
rect 94773 46955 94839 46958
rect 215201 46610 215267 46613
rect 211508 46608 215267 46610
rect 211508 46552 215206 46608
rect 215262 46552 215267 46608
rect 211508 46550 215267 46552
rect 215201 46547 215267 46550
rect 227345 46610 227411 46613
rect 227345 46608 230092 46610
rect 227345 46552 227350 46608
rect 227406 46552 230092 46608
rect 227345 46550 230092 46552
rect 227345 46547 227411 46550
rect 95049 46202 95115 46205
rect 91908 46200 95115 46202
rect 91908 46144 95054 46200
rect 95110 46144 95115 46200
rect 91908 46142 95115 46144
rect 95049 46139 95115 46142
rect 116393 46066 116459 46069
rect 227069 46066 227135 46069
rect 116393 46064 119692 46066
rect 116393 46008 116398 46064
rect 116454 46008 119692 46064
rect 116393 46006 119692 46008
rect 227069 46064 230092 46066
rect 227069 46008 227074 46064
rect 227130 46008 230092 46064
rect 227069 46006 230092 46008
rect 116393 46003 116459 46006
rect 227069 46003 227135 46006
rect 215109 45794 215175 45797
rect 211508 45792 215175 45794
rect 211508 45736 215114 45792
rect 215170 45736 215175 45792
rect 211508 45734 215175 45736
rect 215109 45731 215175 45734
rect 227529 45386 227595 45389
rect 227529 45384 230092 45386
rect 227529 45328 227534 45384
rect 227590 45328 230092 45384
rect 227529 45326 230092 45328
rect 227529 45323 227595 45326
rect 95141 45250 95207 45253
rect 91908 45248 95207 45250
rect 91908 45192 95146 45248
rect 95202 45192 95207 45248
rect 91908 45190 95207 45192
rect 95141 45187 95207 45190
rect 214465 44978 214531 44981
rect 211508 44976 214531 44978
rect 211508 44920 214470 44976
rect 214526 44920 214531 44976
rect 211508 44918 214531 44920
rect 214465 44915 214531 44918
rect 116393 44842 116459 44845
rect 116393 44840 119692 44842
rect 116393 44784 116398 44840
rect 116454 44784 119692 44840
rect 116393 44782 119692 44784
rect 116393 44779 116459 44782
rect 227437 44706 227503 44709
rect 227437 44704 230092 44706
rect 227437 44648 227442 44704
rect 227498 44648 230092 44704
rect 227437 44646 230092 44648
rect 227437 44643 227503 44646
rect 94405 44434 94471 44437
rect 91908 44432 94471 44434
rect 91908 44376 94410 44432
rect 94466 44376 94471 44432
rect 91908 44374 94471 44376
rect 94405 44371 94471 44374
rect 215109 44298 215175 44301
rect 211508 44296 215175 44298
rect 211508 44240 215114 44296
rect 215170 44240 215175 44296
rect 211508 44238 215175 44240
rect 215109 44235 215175 44238
rect 227621 44026 227687 44029
rect 227621 44024 230092 44026
rect 227621 43968 227626 44024
rect 227682 43968 230092 44024
rect 227621 43966 230092 43968
rect 227621 43963 227687 43966
rect 115933 43618 115999 43621
rect 115933 43616 119692 43618
rect 115933 43560 115938 43616
rect 115994 43560 119692 43616
rect 115933 43558 119692 43560
rect 115933 43555 115999 43558
rect 94957 43482 95023 43485
rect 214373 43482 214439 43485
rect 91908 43480 95023 43482
rect 91908 43424 94962 43480
rect 95018 43424 95023 43480
rect 91908 43422 95023 43424
rect 211508 43480 214439 43482
rect 211508 43424 214378 43480
rect 214434 43424 214439 43480
rect 211508 43422 214439 43424
rect 94957 43419 95023 43422
rect 214373 43419 214439 43422
rect 227069 43482 227135 43485
rect 227069 43480 230092 43482
rect 227069 43424 227074 43480
rect 227130 43424 230092 43480
rect 227069 43422 230092 43424
rect 227069 43419 227135 43422
rect 226701 42802 226767 42805
rect 226701 42800 230092 42802
rect 226701 42744 226706 42800
rect 226762 42744 230092 42800
rect 226701 42742 230092 42744
rect 226701 42739 226767 42742
rect 214097 42666 214163 42669
rect 211508 42664 214163 42666
rect 211508 42608 214102 42664
rect 214158 42608 214163 42664
rect 211508 42606 214163 42608
rect 214097 42603 214163 42606
rect 94129 42530 94195 42533
rect 91908 42528 94195 42530
rect 91908 42472 94134 42528
rect 94190 42472 94195 42528
rect 91908 42470 94195 42472
rect 94129 42467 94195 42470
rect 116393 42530 116459 42533
rect 116393 42528 119692 42530
rect 116393 42472 116398 42528
rect 116454 42472 119692 42528
rect 116393 42470 119692 42472
rect 116393 42467 116459 42470
rect 227437 42122 227503 42125
rect 227437 42120 230092 42122
rect 227437 42064 227442 42120
rect 227498 42064 230092 42120
rect 227437 42062 230092 42064
rect 227437 42059 227503 42062
rect 215109 41850 215175 41853
rect 211508 41848 215175 41850
rect 211508 41792 215114 41848
rect 215170 41792 215175 41848
rect 211508 41790 215175 41792
rect 215109 41787 215175 41790
rect 93945 41714 94011 41717
rect 91908 41712 94011 41714
rect 91908 41656 93950 41712
rect 94006 41656 94011 41712
rect 91908 41654 94011 41656
rect 93945 41651 94011 41654
rect 227345 41442 227411 41445
rect 227345 41440 230092 41442
rect 227345 41384 227350 41440
rect 227406 41384 230092 41440
rect 227345 41382 230092 41384
rect 227345 41379 227411 41382
rect 116301 41306 116367 41309
rect 116301 41304 119692 41306
rect 116301 41248 116306 41304
rect 116362 41248 119692 41304
rect 116301 41246 119692 41248
rect 116301 41243 116367 41246
rect 214649 41170 214715 41173
rect 211508 41168 214715 41170
rect 211508 41112 214654 41168
rect 214710 41112 214715 41168
rect 211508 41110 214715 41112
rect 214649 41107 214715 41110
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect 95049 40762 95115 40765
rect 91908 40760 95115 40762
rect 91908 40704 95054 40760
rect 95110 40704 95115 40760
rect 91908 40702 95115 40704
rect 95049 40699 95115 40702
rect 226425 40762 226491 40765
rect 226425 40760 230092 40762
rect 226425 40704 226430 40760
rect 226486 40704 230092 40760
rect 226425 40702 230092 40704
rect 226425 40699 226491 40702
rect 215109 40354 215175 40357
rect 211508 40352 215175 40354
rect 211508 40296 215114 40352
rect 215170 40296 215175 40352
rect 211508 40294 215175 40296
rect 215109 40291 215175 40294
rect 116393 40218 116459 40221
rect 226333 40218 226399 40221
rect 116393 40216 119692 40218
rect 116393 40160 116398 40216
rect 116454 40160 119692 40216
rect 116393 40158 119692 40160
rect 226333 40216 230092 40218
rect 226333 40160 226338 40216
rect 226394 40160 230092 40216
rect 226333 40158 230092 40160
rect 116393 40155 116459 40158
rect 226333 40155 226399 40158
rect 94589 39946 94655 39949
rect 91908 39944 94655 39946
rect 91908 39888 94594 39944
rect 94650 39888 94655 39944
rect 91908 39886 94655 39888
rect 94589 39883 94655 39886
rect 214465 39538 214531 39541
rect 211508 39536 214531 39538
rect 211508 39480 214470 39536
rect 214526 39480 214531 39536
rect 211508 39478 214531 39480
rect 214465 39475 214531 39478
rect 226609 39538 226675 39541
rect 226609 39536 230092 39538
rect 226609 39480 226614 39536
rect 226670 39480 230092 39536
rect 226609 39478 230092 39480
rect 226609 39475 226675 39478
rect 95141 38994 95207 38997
rect 91908 38992 95207 38994
rect 91908 38936 95146 38992
rect 95202 38936 95207 38992
rect 91908 38934 95207 38936
rect 95141 38931 95207 38934
rect 116393 38994 116459 38997
rect 116393 38992 119692 38994
rect 116393 38936 116398 38992
rect 116454 38936 119692 38992
rect 116393 38934 119692 38936
rect 116393 38931 116459 38934
rect 227069 38858 227135 38861
rect 227069 38856 230092 38858
rect 227069 38800 227074 38856
rect 227130 38800 230092 38856
rect 227069 38798 230092 38800
rect 227069 38795 227135 38798
rect 215109 38722 215175 38725
rect 563697 38722 563763 38725
rect 211508 38720 215175 38722
rect 211508 38664 215114 38720
rect 215170 38664 215175 38720
rect 211508 38662 215175 38664
rect 561108 38720 563763 38722
rect 561108 38664 563702 38720
rect 563758 38664 563763 38720
rect 561108 38662 563763 38664
rect 215109 38659 215175 38662
rect 563697 38659 563763 38662
rect 94497 38178 94563 38181
rect 91908 38176 94563 38178
rect 91908 38120 94502 38176
rect 94558 38120 94563 38176
rect 91908 38118 94563 38120
rect 94497 38115 94563 38118
rect 226885 38178 226951 38181
rect 226885 38176 230092 38178
rect 226885 38120 226890 38176
rect 226946 38120 230092 38176
rect 226885 38118 230092 38120
rect 226885 38115 226951 38118
rect 215109 38042 215175 38045
rect 211508 38040 215175 38042
rect 211508 37984 215114 38040
rect 215170 37984 215175 38040
rect 211508 37982 215175 37984
rect 215109 37979 215175 37982
rect 116393 37770 116459 37773
rect 116393 37768 119692 37770
rect 116393 37712 116398 37768
rect 116454 37712 119692 37768
rect 116393 37710 119692 37712
rect 116393 37707 116459 37710
rect 227437 37634 227503 37637
rect 227437 37632 230092 37634
rect 227437 37576 227442 37632
rect 227498 37576 230092 37632
rect 227437 37574 230092 37576
rect 227437 37571 227503 37574
rect 95049 37226 95115 37229
rect 215109 37226 215175 37229
rect 91908 37224 95115 37226
rect 91908 37168 95054 37224
rect 95110 37168 95115 37224
rect 91908 37166 95115 37168
rect 211508 37224 215175 37226
rect 211508 37168 215114 37224
rect 215170 37168 215175 37224
rect 211508 37166 215175 37168
rect 95049 37163 95115 37166
rect 215109 37163 215175 37166
rect 227529 36954 227595 36957
rect 227529 36952 230092 36954
rect 227529 36896 227534 36952
rect 227590 36896 230092 36952
rect 227529 36894 230092 36896
rect 227529 36891 227595 36894
rect 116393 36682 116459 36685
rect 116393 36680 119692 36682
rect 116393 36624 116398 36680
rect 116454 36624 119692 36680
rect 116393 36622 119692 36624
rect 116393 36619 116459 36622
rect 214557 36410 214623 36413
rect 211508 36408 214623 36410
rect 211508 36352 214562 36408
rect 214618 36352 214623 36408
rect 211508 36350 214623 36352
rect 214557 36347 214623 36350
rect 94589 36274 94655 36277
rect 91908 36272 94655 36274
rect 91908 36216 94594 36272
rect 94650 36216 94655 36272
rect 91908 36214 94655 36216
rect 94589 36211 94655 36214
rect 227437 36274 227503 36277
rect 227437 36272 230092 36274
rect 227437 36216 227442 36272
rect 227498 36216 230092 36272
rect 227437 36214 230092 36216
rect 227437 36211 227503 36214
rect -960 35866 480 35956
rect 3417 35866 3483 35869
rect -960 35864 3483 35866
rect -960 35808 3422 35864
rect 3478 35808 3483 35864
rect -960 35806 3483 35808
rect -960 35716 480 35806
rect 3417 35803 3483 35806
rect 214649 35594 214715 35597
rect 211508 35592 214715 35594
rect 211508 35536 214654 35592
rect 214710 35536 214715 35592
rect 211508 35534 214715 35536
rect 214649 35531 214715 35534
rect 227437 35594 227503 35597
rect 227437 35592 230092 35594
rect 227437 35536 227442 35592
rect 227498 35536 230092 35592
rect 227437 35534 230092 35536
rect 227437 35531 227503 35534
rect 93853 35458 93919 35461
rect 91908 35456 93919 35458
rect 91908 35400 93858 35456
rect 93914 35400 93919 35456
rect 91908 35398 93919 35400
rect 93853 35395 93919 35398
rect 116393 35458 116459 35461
rect 116393 35456 119692 35458
rect 116393 35400 116398 35456
rect 116454 35400 119692 35456
rect 116393 35398 119692 35400
rect 116393 35395 116459 35398
rect 215109 34914 215175 34917
rect 211508 34912 215175 34914
rect 211508 34856 215114 34912
rect 215170 34856 215175 34912
rect 211508 34854 215175 34856
rect 215109 34851 215175 34854
rect 227529 34914 227595 34917
rect 227529 34912 230092 34914
rect 227529 34856 227534 34912
rect 227590 34856 230092 34912
rect 227529 34854 230092 34856
rect 227529 34851 227595 34854
rect 93945 34506 94011 34509
rect 91908 34504 94011 34506
rect 91908 34448 93950 34504
rect 94006 34448 94011 34504
rect 91908 34446 94011 34448
rect 93945 34443 94011 34446
rect 116301 34370 116367 34373
rect 227437 34370 227503 34373
rect 116301 34368 119692 34370
rect 116301 34312 116306 34368
rect 116362 34312 119692 34368
rect 116301 34310 119692 34312
rect 227437 34368 230092 34370
rect 227437 34312 227442 34368
rect 227498 34312 230092 34368
rect 227437 34310 230092 34312
rect 116301 34307 116367 34310
rect 227437 34307 227503 34310
rect 214557 34098 214623 34101
rect 211508 34096 214623 34098
rect 211508 34040 214562 34096
rect 214618 34040 214623 34096
rect 211508 34038 214623 34040
rect 214557 34035 214623 34038
rect 95141 33690 95207 33693
rect 91908 33688 95207 33690
rect 91908 33632 95146 33688
rect 95202 33632 95207 33688
rect 91908 33630 95207 33632
rect 95141 33627 95207 33630
rect 227345 33690 227411 33693
rect 227345 33688 230092 33690
rect 227345 33632 227350 33688
rect 227406 33632 230092 33688
rect 227345 33630 230092 33632
rect 227345 33627 227411 33630
rect 215109 33282 215175 33285
rect 211508 33280 215175 33282
rect 211508 33224 215114 33280
rect 215170 33224 215175 33280
rect 211508 33222 215175 33224
rect 215109 33219 215175 33222
rect 116393 33146 116459 33149
rect 116393 33144 119692 33146
rect 116393 33088 116398 33144
rect 116454 33088 119692 33144
rect 116393 33086 119692 33088
rect 116393 33083 116459 33086
rect 227437 33010 227503 33013
rect 227437 33008 230092 33010
rect 227437 32952 227442 33008
rect 227498 32952 230092 33008
rect 227437 32950 230092 32952
rect 227437 32947 227503 32950
rect 95141 32738 95207 32741
rect 91908 32736 95207 32738
rect 91908 32680 95146 32736
rect 95202 32680 95207 32736
rect 91908 32678 95207 32680
rect 95141 32675 95207 32678
rect 215109 32466 215175 32469
rect 211508 32464 215175 32466
rect 211508 32408 215114 32464
rect 215170 32408 215175 32464
rect 211508 32406 215175 32408
rect 215109 32403 215175 32406
rect 227529 32330 227595 32333
rect 227529 32328 230092 32330
rect 227529 32272 227534 32328
rect 227590 32272 230092 32328
rect 227529 32270 230092 32272
rect 227529 32267 227595 32270
rect 116393 32058 116459 32061
rect 116393 32056 119692 32058
rect 116393 32000 116398 32056
rect 116454 32000 119692 32056
rect 116393 31998 119692 32000
rect 116393 31995 116459 31998
rect 95141 31922 95207 31925
rect 91908 31920 95207 31922
rect 91908 31864 95146 31920
rect 95202 31864 95207 31920
rect 91908 31862 95207 31864
rect 95141 31859 95207 31862
rect 213913 31786 213979 31789
rect 211508 31784 213979 31786
rect 211508 31728 213918 31784
rect 213974 31728 213979 31784
rect 211508 31726 213979 31728
rect 213913 31723 213979 31726
rect 227437 31786 227503 31789
rect 227437 31784 230092 31786
rect 227437 31728 227442 31784
rect 227498 31728 230092 31784
rect 227437 31726 230092 31728
rect 227437 31723 227503 31726
rect 32305 30292 32371 30293
rect 32254 30290 32260 30292
rect 32214 30230 32260 30290
rect 32324 30288 32371 30292
rect 32366 30232 32371 30288
rect 32254 30228 32260 30230
rect 32324 30228 32371 30232
rect 32305 30227 32371 30228
rect 580901 29338 580967 29341
rect 583520 29338 584960 29428
rect 580901 29336 584960 29338
rect 580901 29280 580906 29336
rect 580962 29280 584960 29336
rect 580901 29278 584960 29280
rect 580901 29275 580967 29278
rect 583520 29188 584960 29278
rect 411897 27570 411963 27573
rect 411897 27568 414092 27570
rect 411897 27512 411902 27568
rect 411958 27512 414092 27568
rect 411897 27510 414092 27512
rect 411897 27507 411963 27510
rect -960 21450 480 21540
rect 2773 21450 2839 21453
rect -960 21448 2839 21450
rect -960 21392 2778 21448
rect 2834 21392 2839 21448
rect -960 21390 2839 21392
rect -960 21300 480 21390
rect 2773 21387 2839 21390
rect 583520 17492 584960 17732
rect 406469 16962 406535 16965
rect 414657 16962 414723 16965
rect 406469 16960 414723 16962
rect 406469 16904 406474 16960
rect 406530 16904 414662 16960
rect 414718 16904 414723 16960
rect 406469 16902 414723 16904
rect 406469 16899 406535 16902
rect 414657 16899 414723 16902
rect 424593 16962 424659 16965
rect 435357 16962 435423 16965
rect 424593 16960 435423 16962
rect 424593 16904 424598 16960
rect 424654 16904 435362 16960
rect 435418 16904 435423 16960
rect 424593 16902 435423 16904
rect 424593 16899 424659 16902
rect 435357 16899 435423 16902
rect 439405 16962 439471 16965
rect 452561 16962 452627 16965
rect 439405 16960 452627 16962
rect 439405 16904 439410 16960
rect 439466 16904 452566 16960
rect 452622 16904 452627 16960
rect 439405 16902 452627 16904
rect 439405 16899 439471 16902
rect 452561 16899 452627 16902
rect 250437 15602 250503 15605
rect 429101 15602 429167 15605
rect 250437 15600 429167 15602
rect 250437 15544 250442 15600
rect 250498 15544 429106 15600
rect 429162 15544 429167 15600
rect 250437 15542 429167 15544
rect 250437 15539 250503 15542
rect 429101 15539 429167 15542
rect 246297 15466 246363 15469
rect 426801 15466 426867 15469
rect 246297 15464 426867 15466
rect 246297 15408 246302 15464
rect 246358 15408 426806 15464
rect 426862 15408 426867 15464
rect 246297 15406 426867 15408
rect 246297 15403 246363 15406
rect 426801 15403 426867 15406
rect 131021 15330 131087 15333
rect 415301 15330 415367 15333
rect 131021 15328 415367 15330
rect 131021 15272 131026 15328
rect 131082 15272 415306 15328
rect 415362 15272 415367 15328
rect 131021 15270 415367 15272
rect 131021 15267 131087 15270
rect 415301 15267 415367 15270
rect 307201 14922 307267 14925
rect 472433 14922 472499 14925
rect 307201 14920 472499 14922
rect 307201 14864 307206 14920
rect 307262 14864 472438 14920
rect 472494 14864 472499 14920
rect 307201 14862 472499 14864
rect 307201 14859 307267 14862
rect 472433 14859 472499 14862
rect 158621 14786 158687 14789
rect 424133 14786 424199 14789
rect 158621 14784 424199 14786
rect 158621 14728 158626 14784
rect 158682 14728 424138 14784
rect 424194 14728 424199 14784
rect 158621 14726 424199 14728
rect 158621 14723 158687 14726
rect 424133 14723 424199 14726
rect 151721 14650 151787 14653
rect 421833 14650 421899 14653
rect 151721 14648 421899 14650
rect 151721 14592 151726 14648
rect 151782 14592 421838 14648
rect 421894 14592 421899 14648
rect 151721 14590 421899 14592
rect 151721 14587 151787 14590
rect 421833 14587 421899 14590
rect 126881 14514 126947 14517
rect 414197 14514 414263 14517
rect 126881 14512 414263 14514
rect 126881 14456 126886 14512
rect 126942 14456 414202 14512
rect 414258 14456 414263 14512
rect 126881 14454 414263 14456
rect 126881 14451 126947 14454
rect 414197 14451 414263 14454
rect 215201 13426 215267 13429
rect 442533 13426 442599 13429
rect 215201 13424 442599 13426
rect 215201 13368 215206 13424
rect 215262 13368 442538 13424
rect 442594 13368 442599 13424
rect 215201 13366 442599 13368
rect 215201 13363 215267 13366
rect 442533 13363 442599 13366
rect 201401 13290 201467 13293
rect 437933 13290 437999 13293
rect 201401 13288 437999 13290
rect 201401 13232 201406 13288
rect 201462 13232 437938 13288
rect 437994 13232 437999 13288
rect 201401 13230 437999 13232
rect 201401 13227 201467 13230
rect 437933 13227 437999 13230
rect 172421 13154 172487 13157
rect 425053 13154 425119 13157
rect 172421 13152 425119 13154
rect 172421 13096 172426 13152
rect 172482 13096 425058 13152
rect 425114 13096 425119 13152
rect 172421 13094 425119 13096
rect 172421 13091 172487 13094
rect 425053 13091 425119 13094
rect 136541 13018 136607 13021
rect 417233 13018 417299 13021
rect 136541 13016 417299 13018
rect 136541 12960 136546 13016
rect 136602 12960 417238 13016
rect 417294 12960 417299 13016
rect 136541 12958 417299 12960
rect 136541 12955 136607 12958
rect 417233 12955 417299 12958
rect 422293 12610 422359 12613
rect 422753 12610 422819 12613
rect 422293 12608 422819 12610
rect 422293 12552 422298 12608
rect 422354 12552 422758 12608
rect 422814 12552 422819 12608
rect 422293 12550 422819 12552
rect 422293 12547 422359 12550
rect 422753 12547 422819 12550
rect 466177 12610 466243 12613
rect 471881 12610 471947 12613
rect 466177 12608 471947 12610
rect 466177 12552 466182 12608
rect 466238 12552 471886 12608
rect 471942 12552 471947 12608
rect 466177 12550 471947 12552
rect 466177 12547 466243 12550
rect 471881 12547 471947 12550
rect 340137 12066 340203 12069
rect 440233 12066 440299 12069
rect 340137 12064 440299 12066
rect 340137 12008 340142 12064
rect 340198 12008 440238 12064
rect 440294 12008 440299 12064
rect 340137 12006 440299 12008
rect 340137 12003 340203 12006
rect 440233 12003 440299 12006
rect 244181 11930 244247 11933
rect 451733 11930 451799 11933
rect 244181 11928 451799 11930
rect 244181 11872 244186 11928
rect 244242 11872 451738 11928
rect 451794 11872 451799 11928
rect 244181 11870 451799 11872
rect 244181 11867 244247 11870
rect 451733 11867 451799 11870
rect 165521 11794 165587 11797
rect 423121 11794 423187 11797
rect 165521 11792 423187 11794
rect 165521 11736 165526 11792
rect 165582 11736 423126 11792
rect 423182 11736 423187 11792
rect 165521 11734 423187 11736
rect 165521 11731 165587 11734
rect 423121 11731 423187 11734
rect 142061 11658 142127 11661
rect 419165 11658 419231 11661
rect 142061 11656 419231 11658
rect 142061 11600 142066 11656
rect 142122 11600 419170 11656
rect 419226 11600 419231 11656
rect 142061 11598 419231 11600
rect 142061 11595 142127 11598
rect 419165 11595 419231 11598
rect 393221 10706 393287 10709
rect 419901 10706 419967 10709
rect 393221 10704 419967 10706
rect 393221 10648 393226 10704
rect 393282 10648 419906 10704
rect 419962 10648 419967 10704
rect 393221 10646 419967 10648
rect 393221 10643 393287 10646
rect 419901 10643 419967 10646
rect 242801 10570 242867 10573
rect 451365 10570 451431 10573
rect 242801 10568 451431 10570
rect 242801 10512 242806 10568
rect 242862 10512 451370 10568
rect 451426 10512 451431 10568
rect 242801 10510 451431 10512
rect 242801 10507 242867 10510
rect 451365 10507 451431 10510
rect 238661 10434 238727 10437
rect 450169 10434 450235 10437
rect 238661 10432 450235 10434
rect 238661 10376 238666 10432
rect 238722 10376 450174 10432
rect 450230 10376 450235 10432
rect 238661 10374 450235 10376
rect 238661 10371 238727 10374
rect 450169 10371 450235 10374
rect 224861 10298 224927 10301
rect 445569 10298 445635 10301
rect 224861 10296 445635 10298
rect 224861 10240 224866 10296
rect 224922 10240 445574 10296
rect 445630 10240 445635 10296
rect 224861 10238 445635 10240
rect 224861 10235 224927 10238
rect 445569 10235 445635 10238
rect 307753 9346 307819 9349
rect 440969 9346 441035 9349
rect 307753 9344 441035 9346
rect 307753 9288 307758 9344
rect 307814 9288 440974 9344
rect 441030 9288 441035 9344
rect 307753 9286 441035 9288
rect 307753 9283 307819 9286
rect 440969 9283 441035 9286
rect 273161 9210 273227 9213
rect 429193 9210 429259 9213
rect 273161 9208 429259 9210
rect 273161 9152 273166 9208
rect 273222 9152 429198 9208
rect 429254 9152 429259 9208
rect 273161 9150 429259 9152
rect 273161 9147 273227 9150
rect 429193 9147 429259 9150
rect 177757 9074 177823 9077
rect 430665 9074 430731 9077
rect 177757 9072 430731 9074
rect 177757 9016 177762 9072
rect 177818 9016 430670 9072
rect 430726 9016 430731 9072
rect 177757 9014 430731 9016
rect 177757 9011 177823 9014
rect 430665 9011 430731 9014
rect 138473 8938 138539 8941
rect 417969 8938 418035 8941
rect 138473 8936 418035 8938
rect 138473 8880 138478 8936
rect 138534 8880 417974 8936
rect 418030 8880 418035 8936
rect 138473 8878 418035 8880
rect 138473 8875 138539 8878
rect 417969 8875 418035 8878
rect 232497 8122 232563 8125
rect 448237 8122 448303 8125
rect 232497 8120 448303 8122
rect 232497 8064 232502 8120
rect 232558 8064 448242 8120
rect 448298 8064 448303 8120
rect 232497 8062 448303 8064
rect 232497 8059 232563 8062
rect 448237 8059 448303 8062
rect 211061 7986 211127 7989
rect 441337 7986 441403 7989
rect 211061 7984 441403 7986
rect 211061 7928 211066 7984
rect 211122 7928 441342 7984
rect 441398 7928 441403 7984
rect 211061 7926 441403 7928
rect 211061 7923 211127 7926
rect 441337 7923 441403 7926
rect 193305 7850 193371 7853
rect 426709 7850 426775 7853
rect 193305 7848 426775 7850
rect 193305 7792 193310 7848
rect 193366 7792 426714 7848
rect 426770 7792 426775 7848
rect 193305 7790 426775 7792
rect 193305 7787 193371 7790
rect 426709 7787 426775 7790
rect 145649 7714 145715 7717
rect 420269 7714 420335 7717
rect 145649 7712 420335 7714
rect 145649 7656 145654 7712
rect 145710 7656 420274 7712
rect 420330 7656 420335 7712
rect 145649 7654 420335 7656
rect 145649 7651 145715 7654
rect 420269 7651 420335 7654
rect 127801 7578 127867 7581
rect 414565 7578 414631 7581
rect 127801 7576 414631 7578
rect 127801 7520 127806 7576
rect 127862 7520 414570 7576
rect 414626 7520 414631 7576
rect 127801 7518 414631 7520
rect 127801 7515 127867 7518
rect 414565 7515 414631 7518
rect -960 7170 480 7260
rect 2773 7170 2839 7173
rect -960 7168 2839 7170
rect -960 7112 2778 7168
rect 2834 7112 2839 7168
rect -960 7110 2839 7112
rect -960 7020 480 7110
rect 2773 7107 2839 7110
rect 272885 6490 272951 6493
rect 461301 6490 461367 6493
rect 272885 6488 461367 6490
rect 272885 6432 272890 6488
rect 272946 6432 461306 6488
rect 461362 6432 461367 6488
rect 272885 6430 461367 6432
rect 272885 6427 272951 6430
rect 461301 6427 461367 6430
rect 191741 6354 191807 6357
rect 418245 6354 418311 6357
rect 191741 6352 418311 6354
rect 191741 6296 191746 6352
rect 191802 6296 418250 6352
rect 418306 6296 418311 6352
rect 191741 6294 418311 6296
rect 191741 6291 191807 6294
rect 418245 6291 418311 6294
rect 175365 6218 175431 6221
rect 429285 6218 429351 6221
rect 175365 6216 429351 6218
rect 175365 6160 175370 6216
rect 175426 6160 429290 6216
rect 429346 6160 429351 6216
rect 175365 6158 429351 6160
rect 175365 6155 175431 6158
rect 429285 6155 429351 6158
rect 583520 5796 584960 6036
rect 289813 5266 289879 5269
rect 440509 5266 440575 5269
rect 289813 5264 440575 5266
rect 289813 5208 289818 5264
rect 289874 5208 440514 5264
rect 440570 5208 440575 5264
rect 289813 5206 440575 5208
rect 289813 5203 289879 5206
rect 440509 5203 440575 5206
rect 198181 5130 198247 5133
rect 417509 5130 417575 5133
rect 198181 5128 417575 5130
rect 198181 5072 198186 5128
rect 198242 5072 417514 5128
rect 417570 5072 417575 5128
rect 198181 5070 417575 5072
rect 198181 5067 198247 5070
rect 417509 5067 417575 5070
rect 222929 4994 222995 4997
rect 445017 4994 445083 4997
rect 222929 4992 445083 4994
rect 222929 4936 222934 4992
rect 222990 4936 445022 4992
rect 445078 4936 445083 4992
rect 222929 4934 445083 4936
rect 222929 4931 222995 4934
rect 445017 4931 445083 4934
rect 212257 4858 212323 4861
rect 441981 4858 442047 4861
rect 212257 4856 442047 4858
rect 212257 4800 212262 4856
rect 212318 4800 441986 4856
rect 442042 4800 442047 4856
rect 212257 4798 442047 4800
rect 212257 4795 212323 4798
rect 441981 4795 442047 4798
rect 296713 3770 296779 3773
rect 442993 3770 443059 3773
rect 296713 3768 443059 3770
rect 296713 3712 296718 3768
rect 296774 3712 442998 3768
rect 443054 3712 443059 3768
rect 296713 3710 443059 3712
rect 296713 3707 296779 3710
rect 442993 3707 443059 3710
rect 483013 3770 483079 3773
rect 484393 3770 484459 3773
rect 483013 3768 484459 3770
rect 483013 3712 483018 3768
rect 483074 3712 484398 3768
rect 484454 3712 484459 3768
rect 483013 3710 484459 3712
rect 483013 3707 483079 3710
rect 484393 3707 484459 3710
rect 289537 3634 289603 3637
rect 436737 3634 436803 3637
rect 446397 3634 446463 3637
rect 289537 3632 436803 3634
rect 289537 3576 289542 3632
rect 289598 3576 436742 3632
rect 436798 3576 436803 3632
rect 289537 3574 436803 3576
rect 289537 3571 289603 3574
rect 436737 3571 436803 3574
rect 436878 3632 446463 3634
rect 436878 3576 446402 3632
rect 446458 3576 446463 3632
rect 436878 3574 446463 3576
rect 275277 3498 275343 3501
rect 427077 3498 427143 3501
rect 275277 3496 427143 3498
rect 275277 3440 275282 3496
rect 275338 3440 427082 3496
rect 427138 3440 427143 3496
rect 275277 3438 427143 3440
rect 275277 3435 275343 3438
rect 427077 3435 427143 3438
rect 434713 3498 434779 3501
rect 436878 3498 436938 3574
rect 446397 3571 446463 3574
rect 455965 3634 456031 3637
rect 469029 3634 469095 3637
rect 455965 3632 469095 3634
rect 455965 3576 455970 3632
rect 456026 3576 469034 3632
rect 469090 3576 469095 3632
rect 455965 3574 469095 3576
rect 455965 3571 456031 3574
rect 469029 3571 469095 3574
rect 434713 3496 436938 3498
rect 434713 3440 434718 3496
rect 434774 3440 436938 3496
rect 434713 3438 436938 3440
rect 439497 3498 439563 3501
rect 444281 3498 444347 3501
rect 439497 3496 444347 3498
rect 439497 3440 439502 3496
rect 439558 3440 444286 3496
rect 444342 3440 444347 3496
rect 439497 3438 444347 3440
rect 434713 3435 434779 3438
rect 439497 3435 439563 3438
rect 444281 3435 444347 3438
rect 483197 3498 483263 3501
rect 483381 3498 483447 3501
rect 483197 3496 483447 3498
rect 483197 3440 483202 3496
rect 483258 3440 483386 3496
rect 483442 3440 483447 3496
rect 483197 3438 483447 3440
rect 483197 3435 483263 3438
rect 483381 3435 483447 3438
rect 282453 3362 282519 3365
rect 433333 3362 433399 3365
rect 282453 3360 433399 3362
rect 282453 3304 282458 3360
rect 282514 3304 433338 3360
rect 433394 3304 433399 3360
rect 282453 3302 433399 3304
rect 282453 3299 282519 3302
rect 433333 3299 433399 3302
rect 483013 3362 483079 3365
rect 483565 3362 483631 3365
rect 483013 3360 483631 3362
rect 483013 3304 483018 3360
rect 483074 3304 483570 3360
rect 483626 3304 483631 3360
rect 483013 3302 483631 3304
rect 483013 3299 483079 3302
rect 483565 3299 483631 3302
rect 412633 3090 412699 3093
rect 414197 3090 414263 3093
rect 412633 3088 414263 3090
rect 412633 3032 412638 3088
rect 412694 3032 414202 3088
rect 414258 3032 414263 3088
rect 412633 3030 414263 3032
rect 412633 3027 412699 3030
rect 414197 3027 414263 3030
rect 356053 2954 356119 2957
rect 369117 2954 369183 2957
rect 356053 2952 369183 2954
rect 356053 2896 356058 2952
rect 356114 2896 369122 2952
rect 369178 2896 369183 2952
rect 356053 2894 369183 2896
rect 356053 2891 356119 2894
rect 369117 2891 369183 2894
rect 374085 2954 374151 2957
rect 378961 2954 379027 2957
rect 374085 2952 379027 2954
rect 374085 2896 374090 2952
rect 374146 2896 378966 2952
rect 379022 2896 379027 2952
rect 374085 2894 379027 2896
rect 374085 2891 374151 2894
rect 378961 2891 379027 2894
rect 256693 2682 256759 2685
rect 432045 2682 432111 2685
rect 256693 2680 432111 2682
rect 256693 2624 256698 2680
rect 256754 2624 432050 2680
rect 432106 2624 432111 2680
rect 256693 2622 432111 2624
rect 256693 2619 256759 2622
rect 432045 2619 432111 2622
rect 176561 2138 176627 2141
rect 429469 2138 429535 2141
rect 176561 2136 429535 2138
rect 176561 2080 176566 2136
rect 176622 2080 429474 2136
rect 429530 2080 429535 2136
rect 176561 2078 429535 2080
rect 176561 2075 176627 2078
rect 429469 2075 429535 2078
rect 169385 2002 169451 2005
rect 427905 2002 427971 2005
rect 169385 2000 427971 2002
rect 169385 1944 169390 2000
rect 169446 1944 427910 2000
rect 427966 1944 427971 2000
rect 169385 1942 427971 1944
rect 169385 1939 169451 1942
rect 427905 1939 427971 1942
<< via3 >>
rect 317092 700572 317156 700636
rect 317276 700436 317340 700500
rect 18644 700300 18708 700364
rect 316908 700300 316972 700364
rect 283052 684448 283116 684452
rect 283052 684392 283066 684448
rect 283066 684392 283116 684448
rect 283052 684388 283116 684392
rect 219020 679144 219084 679148
rect 219020 679088 219070 679144
rect 219070 679088 219084 679144
rect 219020 679084 219084 679088
rect 283052 678872 283116 678876
rect 283052 678816 283102 678872
rect 283102 678816 283116 678872
rect 283052 678812 283116 678816
rect 219020 676288 219084 676292
rect 219020 676232 219034 676288
rect 219034 676232 219084 676288
rect 219020 676228 219084 676232
rect 280660 667932 280724 667996
rect 492444 663852 492508 663916
rect 493916 662084 493980 662148
rect 551324 660044 551388 660108
rect 553348 659364 553412 659428
rect 551324 657868 551388 657932
rect 553532 656916 553596 656980
rect 552060 655556 552124 655620
rect 553900 654468 553964 654532
rect 553716 653244 553780 653308
rect 554084 652020 554148 652084
rect 551324 650524 551388 650588
rect 551508 646580 551572 646644
rect 551324 645764 551388 645828
rect 552244 641004 552308 641068
rect 552428 636244 552492 636308
rect 552796 631348 552860 631412
rect 551692 630804 551756 630868
rect 551508 630668 551572 630732
rect 551692 630532 551756 630596
rect 551324 627948 551388 628012
rect 552612 626452 552676 626516
rect 280108 619516 280172 619580
rect 31156 617748 31220 617812
rect 31340 617612 31404 617676
rect 30788 617476 30852 617540
rect 31524 617536 31588 617540
rect 31524 617480 31538 617536
rect 31538 617480 31588 617536
rect 31524 617476 31588 617480
rect 551692 616252 551756 616316
rect 27476 614892 27540 614956
rect 27292 614348 27356 614412
rect 28580 613260 28644 613324
rect 27660 613124 27724 613188
rect 551508 612716 551572 612780
rect 26924 612580 26988 612644
rect 24900 611900 24964 611964
rect 27108 611356 27172 611420
rect 27844 610812 27908 610876
rect 26740 610132 26804 610196
rect 28028 609044 28092 609108
rect 26004 608364 26068 608428
rect 28212 606732 28276 606796
rect 28396 605644 28460 605708
rect 25636 604692 25700 604756
rect 551738 604284 551802 604348
rect 25820 602924 25884 602988
rect 551324 602788 551388 602852
rect 551692 602788 551756 602852
rect 25268 601156 25332 601220
rect 28626 598360 28690 598364
rect 28626 598304 28630 598360
rect 28630 598304 28686 598360
rect 28686 598304 28690 598360
rect 28626 598300 28690 598304
rect 28580 597620 28644 597684
rect 28580 596668 28644 596732
rect 28580 594628 28644 594692
rect 551876 593948 551940 594012
rect 28580 593464 28644 593468
rect 28580 593408 28594 593464
rect 28594 593408 28644 593464
rect 28580 593404 28644 593408
rect 551324 593404 551388 593468
rect 551692 593404 551756 593468
rect 25268 592180 25332 592244
rect 25084 591908 25148 591972
rect 28580 591908 28644 591972
rect 28580 591288 28644 591292
rect 28580 591232 28594 591288
rect 28594 591232 28644 591288
rect 28580 591228 28644 591232
rect 551324 588508 551388 588572
rect 25084 587828 25148 587892
rect 551692 582524 551756 582588
rect 551876 582252 551940 582316
rect 551324 576948 551388 577012
rect 551692 576948 551756 577012
rect 25636 576540 25700 576604
rect 26372 576540 26436 576604
rect 551508 573412 551572 573476
rect 551876 573412 551940 573476
rect 20484 571916 20548 571980
rect 29500 571372 29564 571436
rect 30420 571372 30484 571436
rect 550772 570420 550836 570484
rect 551692 570420 551756 570484
rect 551508 570012 551572 570076
rect 551876 570012 551940 570076
rect 29316 567836 29380 567900
rect 29868 567836 29932 567900
rect 551876 567700 551940 567764
rect 550588 567564 550652 567628
rect 551876 567564 551940 567628
rect 29132 567488 29196 567492
rect 29132 567432 29146 567488
rect 29146 567432 29196 567488
rect 29132 567428 29196 567432
rect 29684 565660 29748 565724
rect 29132 565388 29196 565452
rect 551324 563212 551388 563276
rect 551324 562940 551388 563004
rect 29316 560764 29380 560828
rect 29868 560764 29932 560828
rect 551508 558996 551572 559060
rect 28948 558452 29012 558516
rect 29500 558452 29564 558516
rect 29500 558316 29564 558380
rect 550588 558180 550652 558244
rect 551692 558180 551756 558244
rect 30052 557424 30116 557428
rect 30052 557368 30066 557424
rect 30066 557368 30116 557424
rect 30052 557364 30116 557368
rect 30236 557092 30300 557156
rect 550772 553964 550836 554028
rect 551508 553964 551572 554028
rect 28948 547708 29012 547772
rect 25820 547028 25884 547092
rect 552796 547028 552860 547092
rect 29132 545804 29196 545868
rect 29684 545804 29748 545868
rect 551140 543764 551204 543828
rect 551876 543764 551940 543828
rect 551140 543628 551204 543692
rect 551508 543628 551572 543692
rect 30052 540908 30116 540972
rect 29316 538324 29380 538388
rect 29500 538188 29564 538252
rect 28028 534924 28092 534988
rect 26004 534788 26068 534852
rect 27844 534652 27908 534716
rect 28396 533836 28460 533900
rect 28212 533700 28276 533764
rect 30236 533564 30300 533628
rect 31156 533564 31220 533628
rect 551508 533564 551572 533628
rect 31340 533428 31404 533492
rect 554084 533428 554148 533492
rect 31524 533292 31588 533356
rect 553900 533292 553964 533356
rect 26740 532612 26804 532676
rect 550956 532612 551020 532676
rect 27108 532476 27172 532540
rect 550772 532476 550836 532540
rect 26924 532340 26988 532404
rect 552060 532340 552124 532404
rect 29500 532204 29564 532268
rect 553716 532204 553780 532268
rect 27292 532068 27356 532132
rect 550588 532068 550652 532132
rect 27476 531932 27540 531996
rect 553532 531932 553596 531996
rect 29684 531796 29748 531860
rect 552244 531796 552308 531860
rect 29868 531660 29932 531724
rect 552428 531660 552492 531724
rect 29132 531388 29196 531452
rect 95188 531252 95252 531316
rect 104940 531252 105004 531316
rect 493916 531252 493980 531316
rect 492444 531116 492508 531180
rect 30236 530844 30300 530908
rect 552612 530844 552676 530908
rect 29132 530708 29196 530772
rect 551324 530708 551388 530772
rect 27660 530572 27724 530636
rect 553348 530572 553412 530636
rect 493548 529892 493612 529956
rect 574876 527716 574940 527780
rect 574876 502692 574940 502756
rect 130700 500788 130764 500852
rect 189580 500788 189644 500852
rect 191052 500788 191116 500852
rect 491892 500848 491956 500852
rect 491892 500792 491906 500848
rect 491906 500792 491956 500848
rect 491892 500788 491956 500792
rect 493180 500848 493244 500852
rect 493180 500792 493194 500848
rect 493194 500792 493244 500848
rect 493180 500788 493244 500792
rect 508452 500788 508516 500852
rect 518020 500848 518084 500852
rect 518020 500792 518034 500848
rect 518034 500792 518084 500848
rect 518020 500788 518084 500792
rect 542860 500788 542924 500852
rect 550220 500788 550284 500852
rect 189764 500652 189828 500716
rect 149100 500516 149164 500580
rect 112852 500108 112916 500172
rect 151860 500380 151924 500444
rect 147812 500244 147876 500308
rect 147996 500108 148060 500172
rect 147628 499836 147692 499900
rect 147076 499624 147140 499628
rect 147076 499568 147090 499624
rect 147090 499568 147140 499624
rect 147076 499564 147140 499568
rect 148180 499624 148244 499628
rect 148180 499568 148194 499624
rect 148194 499568 148244 499624
rect 148180 499564 148244 499568
rect 149652 499564 149716 499628
rect 149836 499564 149900 499628
rect 150940 499564 151004 499628
rect 152412 499624 152476 499628
rect 152412 499568 152462 499624
rect 152462 499568 152476 499624
rect 152412 499564 152476 499568
rect 154804 498068 154868 498132
rect 149284 497932 149348 497996
rect 150388 497796 150452 497860
rect 150756 497660 150820 497724
rect 153700 497660 153764 497724
rect 148364 497524 148428 497588
rect 150572 497388 150636 497452
rect 153148 497252 153212 497316
rect 154620 497116 154684 497180
rect 550588 487732 550652 487796
rect 147444 485828 147508 485892
rect 147260 485556 147324 485620
rect 552244 477124 552308 477188
rect 552796 476988 552860 477052
rect 552612 476852 552676 476916
rect 552428 476716 552492 476780
rect 542860 476232 542924 476236
rect 542860 476176 542910 476232
rect 542910 476176 542924 476232
rect 542860 476172 542924 476176
rect 508452 476096 508516 476100
rect 508452 476040 508502 476096
rect 508502 476040 508516 476096
rect 508452 476036 508516 476040
rect 551140 476036 551204 476100
rect 551692 475900 551756 475964
rect 555004 475764 555068 475828
rect 553348 475628 553412 475692
rect 552060 475356 552124 475420
rect 550588 474540 550652 474604
rect 553532 474268 553596 474332
rect 553716 474132 553780 474196
rect 299428 473860 299492 473924
rect 318748 473860 318812 473924
rect 328316 473860 328380 473924
rect 338068 473860 338132 473924
rect 347636 473860 347700 473924
rect 357388 473860 357452 473924
rect 366956 473860 367020 473924
rect 384988 473860 385052 473924
rect 518020 473860 518084 473924
rect 550220 473996 550284 474060
rect 554084 473996 554148 474060
rect 555372 473860 555436 473924
rect 280660 473724 280724 473788
rect 299428 473588 299492 473652
rect 328316 473588 328380 473652
rect 318748 473452 318812 473516
rect 347636 473588 347700 473652
rect 331076 473452 331140 473516
rect 331260 473452 331324 473516
rect 338068 473452 338132 473516
rect 366956 473588 367020 473652
rect 350396 473452 350460 473516
rect 350580 473452 350644 473516
rect 357388 473452 357452 473516
rect 369716 473452 369780 473516
rect 369900 473452 369964 473516
rect 384988 473588 385052 473652
rect 434668 473724 434732 473788
rect 425100 473588 425164 473652
rect 517468 473724 517532 473788
rect 491892 473512 491956 473516
rect 491892 473456 491906 473512
rect 491906 473456 491956 473512
rect 491892 473452 491956 473456
rect 493180 473512 493244 473516
rect 493180 473456 493194 473512
rect 493194 473456 493244 473512
rect 493180 473452 493244 473456
rect 517468 473452 517532 473516
rect 536788 473724 536852 473788
rect 536972 473588 537036 473652
rect 425100 473316 425164 473380
rect 434668 473316 434732 473380
rect 554820 472636 554884 472700
rect 552060 471276 552124 471340
rect 552428 468964 552492 469028
rect 553348 468012 553412 468076
rect 552612 467740 552676 467804
rect 555004 466788 555068 466852
rect 552796 466244 552860 466308
rect 555372 465564 555436 465628
rect 552244 465292 552308 465356
rect 552060 464748 552124 464812
rect 554820 463796 554884 463860
rect 552060 463524 552124 463588
rect 553716 461484 553780 461548
rect 553532 457268 553596 457332
rect 554084 440676 554148 440740
rect 317092 428708 317156 428772
rect 316908 428572 316972 428636
rect 317276 428436 317340 428500
rect 155908 421228 155972 421292
rect 281580 421288 281644 421292
rect 281580 421232 281630 421288
rect 281630 421232 281644 421288
rect 281580 421228 281644 421232
rect 153884 403548 153948 403612
rect 153332 401372 153396 401436
rect 154620 401236 154684 401300
rect 153148 401100 153212 401164
rect 154804 400964 154868 401028
rect 151860 400828 151924 400892
rect 146892 398652 146956 398716
rect 147444 398652 147508 398716
rect 147076 389464 147140 389468
rect 147076 389408 147126 389464
rect 147126 389408 147140 389464
rect 147076 389404 147140 389408
rect 146708 386548 146772 386612
rect 147260 386548 147324 386612
rect 147076 386472 147140 386476
rect 147076 386416 147126 386472
rect 147126 386416 147140 386472
rect 147076 386412 147140 386416
rect 155724 376680 155788 376684
rect 155724 376624 155738 376680
rect 155738 376624 155788 376680
rect 155724 376620 155788 376624
rect 155724 369744 155788 369748
rect 155724 369688 155774 369744
rect 155774 369688 155788 369744
rect 155724 369684 155788 369688
rect 153884 364244 153948 364308
rect 147260 360436 147324 360500
rect 147076 360300 147140 360364
rect 146892 360028 146956 360092
rect 147076 360028 147140 360092
rect 20484 357308 20548 357372
rect 147076 351732 147140 351796
rect 147812 351732 147876 351796
rect 148180 351732 148244 351796
rect 149652 351732 149716 351796
rect 149836 351732 149900 351796
rect 150940 351732 151004 351796
rect 152412 351792 152476 351796
rect 152412 351736 152426 351792
rect 152426 351736 152476 351792
rect 152412 351732 152476 351736
rect 189764 351732 189828 351796
rect 191052 351732 191116 351796
rect 150388 351596 150452 351660
rect 189580 351596 189644 351660
rect 150756 351460 150820 351524
rect 148364 351324 148428 351388
rect 153700 351324 153764 351388
rect 149100 351188 149164 351252
rect 147996 351052 148060 351116
rect 146892 350916 146956 350980
rect 147628 350780 147692 350844
rect 149284 350780 149348 350844
rect 150572 350644 150636 350708
rect 219940 322084 220004 322148
rect 190132 320316 190196 320380
rect 194364 320316 194428 320380
rect 190316 320180 190380 320244
rect 191604 320180 191668 320244
rect 193076 320180 193140 320244
rect 194180 320180 194244 320244
rect 332916 302772 332980 302836
rect 280108 235180 280172 235244
rect 193076 224844 193140 224908
rect 194364 224708 194428 224772
rect 191604 224572 191668 224636
rect 190132 224436 190196 224500
rect 190316 224300 190380 224364
rect 194180 224164 194244 224228
rect 332916 173844 332980 173908
rect 219940 158748 220004 158812
rect 32260 125080 32324 125084
rect 32260 125024 32274 125080
rect 32274 125024 32324 125080
rect 32260 125020 32324 125024
rect 18644 124204 18708 124268
rect 32260 30288 32324 30292
rect 32260 30232 32310 30288
rect 32310 30232 32324 30288
rect 32260 30228 32324 30232
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 -6926 -7976 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 -5986 -7036 709922
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 -5046 -6096 708982
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 -4106 -5156 708042
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 -3166 -4216 707102
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 -2226 -3276 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18643 700364 18709 700365
rect 18643 700300 18644 700364
rect 18708 700300 18709 700364
rect 18643 700299 18709 700300
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 13408 182454 13728 182476
rect 13408 182218 13450 182454
rect 13686 182218 13728 182454
rect 13408 182134 13728 182218
rect 13408 181898 13450 182134
rect 13686 181898 13728 182134
rect 13408 181876 13728 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 13408 146454 13728 146476
rect 13408 146218 13450 146454
rect 13686 146218 13728 146454
rect 13408 146134 13728 146218
rect 13408 145898 13450 146134
rect 13686 145898 13728 146134
rect 13408 145876 13728 145898
rect 18646 124269 18706 700299
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 31155 617812 31221 617813
rect 31155 617748 31156 617812
rect 31220 617748 31221 617812
rect 31155 617747 31221 617748
rect 30787 617540 30853 617541
rect 30787 617476 30788 617540
rect 30852 617476 30853 617540
rect 30787 617475 30853 617476
rect 30790 615770 30850 617475
rect 30790 615710 31034 615770
rect 27475 614956 27541 614957
rect 27475 614892 27476 614956
rect 27540 614892 27541 614956
rect 27475 614891 27541 614892
rect 27291 614412 27357 614413
rect 27291 614348 27292 614412
rect 27356 614348 27357 614412
rect 27291 614347 27357 614348
rect 26923 612644 26989 612645
rect 26923 612580 26924 612644
rect 26988 612580 26989 612644
rect 26923 612579 26989 612580
rect 24899 611964 24965 611965
rect 24899 611900 24900 611964
rect 24964 611900 24965 611964
rect 24899 611899 24965 611900
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 20483 571980 20549 571981
rect 20483 571916 20484 571980
rect 20548 571916 20549 571980
rect 20483 571915 20549 571916
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 487040 19404 487898
rect 18804 380454 19404 400000
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 20486 357373 20546 571915
rect 24902 571658 24962 611899
rect 26739 610196 26805 610197
rect 26739 610132 26740 610196
rect 26804 610132 26805 610196
rect 26739 610131 26805 610132
rect 26003 608428 26069 608429
rect 26003 608364 26004 608428
rect 26068 608364 26069 608428
rect 26003 608363 26069 608364
rect 25635 604756 25701 604757
rect 25635 604692 25636 604756
rect 25700 604692 25701 604756
rect 25635 604691 25701 604692
rect 25267 601220 25333 601221
rect 25267 601156 25268 601220
rect 25332 601156 25333 601220
rect 25267 601155 25333 601156
rect 25270 592245 25330 601155
rect 25267 592244 25333 592245
rect 25267 592180 25268 592244
rect 25332 592180 25333 592244
rect 25267 592179 25333 592180
rect 25083 591972 25149 591973
rect 25083 591908 25084 591972
rect 25148 591908 25149 591972
rect 25083 591907 25149 591908
rect 25086 587893 25146 591907
rect 25083 587892 25149 587893
rect 25083 587828 25084 587892
rect 25148 587828 25149 587892
rect 25083 587827 25149 587828
rect 25638 576605 25698 604691
rect 25819 602988 25885 602989
rect 25819 602924 25820 602988
rect 25884 602924 25885 602988
rect 25819 602923 25885 602924
rect 25635 576604 25701 576605
rect 25635 576540 25636 576604
rect 25700 576540 25701 576604
rect 25635 576539 25701 576540
rect 25822 547093 25882 602923
rect 25819 547092 25885 547093
rect 25819 547028 25820 547092
rect 25884 547028 25885 547092
rect 25819 547027 25885 547028
rect 26006 534853 26066 608363
rect 26371 576604 26437 576605
rect 26371 576540 26372 576604
rect 26436 576540 26437 576604
rect 26371 576539 26437 576540
rect 26374 573018 26434 576539
rect 26003 534852 26069 534853
rect 26003 534788 26004 534852
rect 26068 534788 26069 534852
rect 26003 534787 26069 534788
rect 26742 532677 26802 610131
rect 26739 532676 26805 532677
rect 26739 532612 26740 532676
rect 26804 532612 26805 532676
rect 26739 532611 26805 532612
rect 26926 532405 26986 612579
rect 27107 611420 27173 611421
rect 27107 611356 27108 611420
rect 27172 611356 27173 611420
rect 27107 611355 27173 611356
rect 27110 532541 27170 611355
rect 27107 532540 27173 532541
rect 27107 532476 27108 532540
rect 27172 532476 27173 532540
rect 27107 532475 27173 532476
rect 26923 532404 26989 532405
rect 26923 532340 26924 532404
rect 26988 532340 26989 532404
rect 26923 532339 26989 532340
rect 27294 532133 27354 614347
rect 27291 532132 27357 532133
rect 27291 532068 27292 532132
rect 27356 532068 27357 532132
rect 27291 532067 27357 532068
rect 27478 531997 27538 614891
rect 28579 613324 28645 613325
rect 28579 613260 28580 613324
rect 28644 613260 28645 613324
rect 28579 613259 28645 613260
rect 28950 613262 29378 613322
rect 27659 613188 27725 613189
rect 27659 613124 27660 613188
rect 27724 613124 27725 613188
rect 27659 613123 27725 613124
rect 27475 531996 27541 531997
rect 27475 531932 27476 531996
rect 27540 531932 27541 531996
rect 27475 531931 27541 531932
rect 27662 530637 27722 613123
rect 28582 613050 28642 613259
rect 28950 613050 29010 613262
rect 28582 612990 29010 613050
rect 27843 610876 27909 610877
rect 27843 610812 27844 610876
rect 27908 610812 27909 610876
rect 27843 610811 27909 610812
rect 27846 534717 27906 610811
rect 28027 609108 28093 609109
rect 28027 609044 28028 609108
rect 28092 609044 28093 609108
rect 28027 609043 28093 609044
rect 28030 534989 28090 609043
rect 29318 608970 29378 613262
rect 29318 608910 29930 608970
rect 28211 606796 28277 606797
rect 28211 606732 28212 606796
rect 28276 606732 28277 606796
rect 28211 606731 28277 606732
rect 28027 534988 28093 534989
rect 28027 534924 28028 534988
rect 28092 534924 28093 534988
rect 28027 534923 28093 534924
rect 27843 534716 27909 534717
rect 27843 534652 27844 534716
rect 27908 534652 27909 534716
rect 27843 534651 27909 534652
rect 28214 533765 28274 606731
rect 28395 605708 28461 605709
rect 28395 605644 28396 605708
rect 28460 605644 28461 605708
rect 28395 605643 28461 605644
rect 28398 533901 28458 605643
rect 28625 598364 28691 598365
rect 28625 598300 28626 598364
rect 28690 598362 28691 598364
rect 29870 598362 29930 608910
rect 28690 598302 29930 598362
rect 28690 598300 28691 598302
rect 28625 598299 28691 598300
rect 28579 597684 28645 597685
rect 28579 597620 28580 597684
rect 28644 597620 28645 597684
rect 28579 597619 28645 597620
rect 28582 597410 28642 597619
rect 28582 597350 29746 597410
rect 28579 596732 28645 596733
rect 28579 596668 28580 596732
rect 28644 596730 28645 596732
rect 28644 596670 29378 596730
rect 28644 596668 28645 596670
rect 28579 596667 28645 596668
rect 29318 596050 29378 596670
rect 29134 595990 29378 596050
rect 29686 596050 29746 597350
rect 29686 595990 30482 596050
rect 28579 594692 28645 594693
rect 28579 594628 28580 594692
rect 28644 594690 28645 594692
rect 29134 594690 29194 595990
rect 28644 594630 29194 594690
rect 28644 594628 28645 594630
rect 28579 594627 28645 594628
rect 28579 593468 28645 593469
rect 28579 593404 28580 593468
rect 28644 593404 28645 593468
rect 28579 593403 28645 593404
rect 28582 592650 28642 593403
rect 28582 592590 29930 592650
rect 28950 592182 29378 592242
rect 28579 591972 28645 591973
rect 28579 591908 28580 591972
rect 28644 591970 28645 591972
rect 28950 591970 29010 592182
rect 28644 591910 29010 591970
rect 28644 591908 28645 591910
rect 28579 591907 28645 591908
rect 28579 591292 28645 591293
rect 28579 591228 28580 591292
rect 28644 591290 28645 591292
rect 28644 591230 28826 591290
rect 28644 591228 28645 591230
rect 28579 591227 28645 591228
rect 28766 585170 28826 591230
rect 28766 585110 29010 585170
rect 28950 583130 29010 585110
rect 28582 583070 29010 583130
rect 28582 577690 28642 583070
rect 28582 577630 28826 577690
rect 28766 571570 28826 577630
rect 29318 573610 29378 592182
rect 29318 573550 29746 573610
rect 28766 571510 29194 571570
rect 29134 567493 29194 571510
rect 29499 571436 29565 571437
rect 29499 571372 29500 571436
rect 29564 571372 29565 571436
rect 29499 571371 29565 571372
rect 29315 567900 29381 567901
rect 29315 567836 29316 567900
rect 29380 567836 29381 567900
rect 29315 567835 29381 567836
rect 29131 567492 29197 567493
rect 29131 567428 29132 567492
rect 29196 567428 29197 567492
rect 29131 567427 29197 567428
rect 29131 565452 29197 565453
rect 29131 565388 29132 565452
rect 29196 565388 29197 565452
rect 29131 565387 29197 565388
rect 28947 558516 29013 558517
rect 28947 558452 28948 558516
rect 29012 558452 29013 558516
rect 28947 558451 29013 558452
rect 28950 547773 29010 558451
rect 28947 547772 29013 547773
rect 28947 547708 28948 547772
rect 29012 547708 29013 547772
rect 28947 547707 29013 547708
rect 29134 545869 29194 565387
rect 29318 560829 29378 567835
rect 29315 560828 29381 560829
rect 29315 560764 29316 560828
rect 29380 560764 29381 560828
rect 29315 560763 29381 560764
rect 29502 558517 29562 571371
rect 29686 565725 29746 573550
rect 29870 567901 29930 592590
rect 30422 591290 30482 595990
rect 30054 591230 30482 591290
rect 29867 567900 29933 567901
rect 29867 567836 29868 567900
rect 29932 567836 29933 567900
rect 29867 567835 29933 567836
rect 29683 565724 29749 565725
rect 29683 565660 29684 565724
rect 29748 565660 29749 565724
rect 29683 565659 29749 565660
rect 29867 560828 29933 560829
rect 29867 560764 29868 560828
rect 29932 560764 29933 560828
rect 29867 560763 29933 560764
rect 29499 558516 29565 558517
rect 29499 558452 29500 558516
rect 29564 558452 29565 558516
rect 29499 558451 29565 558452
rect 29499 558380 29565 558381
rect 29499 558316 29500 558380
rect 29564 558316 29565 558380
rect 29499 558315 29565 558316
rect 29502 547770 29562 558315
rect 29318 547710 29562 547770
rect 29131 545868 29197 545869
rect 29131 545804 29132 545868
rect 29196 545804 29197 545868
rect 29131 545803 29197 545804
rect 29318 538389 29378 547710
rect 29683 545868 29749 545869
rect 29683 545804 29684 545868
rect 29748 545804 29749 545868
rect 29683 545803 29749 545804
rect 29315 538388 29381 538389
rect 29315 538324 29316 538388
rect 29380 538324 29381 538388
rect 29315 538323 29381 538324
rect 29499 538252 29565 538253
rect 29499 538188 29500 538252
rect 29564 538188 29565 538252
rect 29499 538187 29565 538188
rect 28395 533900 28461 533901
rect 28395 533836 28396 533900
rect 28460 533836 28461 533900
rect 28395 533835 28461 533836
rect 28211 533764 28277 533765
rect 28211 533700 28212 533764
rect 28276 533700 28277 533764
rect 28211 533699 28277 533700
rect 29502 532269 29562 538187
rect 29499 532268 29565 532269
rect 29499 532204 29500 532268
rect 29564 532204 29565 532268
rect 29499 532203 29565 532204
rect 29686 531861 29746 545803
rect 29683 531860 29749 531861
rect 29683 531796 29684 531860
rect 29748 531796 29749 531860
rect 29683 531795 29749 531796
rect 29870 531725 29930 560763
rect 30054 557429 30114 591230
rect 30422 571437 30482 572102
rect 30419 571436 30485 571437
rect 30419 571372 30420 571436
rect 30484 571372 30485 571436
rect 30419 571371 30485 571372
rect 30051 557428 30117 557429
rect 30051 557364 30052 557428
rect 30116 557364 30117 557428
rect 30051 557363 30117 557364
rect 30235 557156 30301 557157
rect 30235 557092 30236 557156
rect 30300 557092 30301 557156
rect 30235 557091 30301 557092
rect 30238 545050 30298 557091
rect 30054 544990 30298 545050
rect 30054 540973 30114 544990
rect 30051 540972 30117 540973
rect 30051 540908 30052 540972
rect 30116 540908 30117 540972
rect 30051 540907 30117 540908
rect 30235 533628 30301 533629
rect 30235 533564 30236 533628
rect 30300 533564 30301 533628
rect 30235 533563 30301 533564
rect 29867 531724 29933 531725
rect 29867 531660 29868 531724
rect 29932 531660 29933 531724
rect 29867 531659 29933 531660
rect 29131 531452 29197 531453
rect 29131 531388 29132 531452
rect 29196 531388 29197 531452
rect 29131 531387 29197 531388
rect 29134 530773 29194 531387
rect 30238 530909 30298 533563
rect 30974 531538 31034 615710
rect 31158 533629 31218 617747
rect 36804 617680 37404 649898
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 617680 55404 631898
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 617680 73404 649898
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 617680 91404 631898
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 617680 109404 649898
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 617680 127404 631898
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 31339 617676 31405 617677
rect 31339 617612 31340 617676
rect 31404 617612 31405 617676
rect 31339 617611 31405 617612
rect 31155 533628 31221 533629
rect 31155 533564 31156 533628
rect 31220 533564 31221 533628
rect 31155 533563 31221 533564
rect 31342 533493 31402 617611
rect 31523 617540 31589 617541
rect 31523 617476 31524 617540
rect 31588 617476 31589 617540
rect 31523 617475 31589 617476
rect 31339 533492 31405 533493
rect 31339 533428 31340 533492
rect 31404 533428 31405 533492
rect 31339 533427 31405 533428
rect 31526 533357 31586 617475
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 36804 542454 37404 571440
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 31523 533356 31589 533357
rect 31523 533292 31524 533356
rect 31588 533292 31589 533356
rect 31523 533291 31589 533292
rect 30235 530908 30301 530909
rect 30235 530844 30236 530908
rect 30300 530844 30301 530908
rect 30235 530843 30301 530844
rect 29131 530772 29197 530773
rect 29131 530708 29132 530772
rect 29196 530708 29197 530772
rect 29131 530707 29197 530708
rect 27659 530636 27725 530637
rect 27659 530572 27660 530636
rect 27724 530572 27725 530636
rect 27659 530571 27725 530572
rect 36804 528912 37404 541898
rect 54804 560454 55404 571440
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 528912 55404 559898
rect 72804 542454 73404 571440
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 528912 73404 541898
rect 90804 560454 91404 571440
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 528912 91404 559898
rect 95190 531317 95250 571422
rect 108804 542454 109404 571440
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 95187 531316 95253 531317
rect 95187 531252 95188 531316
rect 95252 531252 95253 531316
rect 95187 531251 95253 531252
rect 104939 531252 104940 531302
rect 105004 531252 105005 531302
rect 104939 531251 105005 531252
rect 108804 528912 109404 541898
rect 126804 560454 127404 571440
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 528912 127404 559898
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 528912 145404 541898
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 528912 163404 559898
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 618224 199404 631898
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 219019 679148 219085 679149
rect 219019 679084 219020 679148
rect 219084 679084 219085 679148
rect 219019 679083 219085 679084
rect 219022 676293 219082 679083
rect 219019 676292 219085 676293
rect 219019 676228 219020 676292
rect 219084 676228 219085 676292
rect 219019 676227 219085 676228
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 618224 217404 649898
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 618224 235404 631898
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 618224 253404 649898
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 283051 684452 283117 684453
rect 283051 684388 283052 684452
rect 283116 684388 283117 684452
rect 283051 684387 283117 684388
rect 283054 678877 283114 684387
rect 283051 678876 283117 678877
rect 283051 678812 283052 678876
rect 283116 678812 283117 678876
rect 283051 678811 283117 678812
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 280659 667996 280725 667997
rect 280659 667932 280660 667996
rect 280724 667932 280725 667996
rect 280659 667931 280725 667932
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 618224 271404 631898
rect 280107 619580 280173 619581
rect 280107 619516 280108 619580
rect 280172 619516 280173 619580
rect 280107 619515 280173 619516
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 528912 181404 541898
rect 198804 560454 199404 574112
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 528912 199404 559898
rect 216804 542454 217404 574112
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 528912 217404 541898
rect 234804 560454 235404 574112
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 528912 235404 559898
rect 252804 542454 253404 574112
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 528912 253404 541898
rect 270804 560454 271404 574112
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 528912 271404 559898
rect 107675 524454 107995 524476
rect 107675 524218 107717 524454
rect 107953 524218 107995 524454
rect 107675 524134 107995 524218
rect 107675 523898 107717 524134
rect 107953 523898 107995 524134
rect 107675 523876 107995 523898
rect 192805 524454 193125 524476
rect 192805 524218 192847 524454
rect 193083 524218 193125 524454
rect 192805 524134 193125 524218
rect 192805 523898 192847 524134
rect 193083 523898 193125 524134
rect 192805 523876 193125 523898
rect 65109 506454 65429 506476
rect 65109 506218 65151 506454
rect 65387 506218 65429 506454
rect 65109 506134 65429 506218
rect 65109 505898 65151 506134
rect 65387 505898 65429 506134
rect 65109 505876 65429 505898
rect 150240 506454 150560 506476
rect 150240 506218 150282 506454
rect 150518 506218 150560 506454
rect 150240 506134 150560 506218
rect 150240 505898 150282 506134
rect 150518 505898 150560 506134
rect 150240 505876 150560 505898
rect 235370 506454 235690 506476
rect 235370 506218 235412 506454
rect 235648 506218 235690 506454
rect 235370 506134 235690 506218
rect 235370 505898 235412 506134
rect 235648 505898 235690 506134
rect 235370 505876 235690 505898
rect 36804 487040 37404 502800
rect 54804 488454 55404 502800
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 487040 55404 487898
rect 72804 487040 73404 502800
rect 90804 488454 91404 502800
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 487040 91404 487898
rect 108804 487040 109404 502800
rect 126804 488454 127404 502800
rect 130699 500852 130765 500853
rect 130699 500788 130700 500852
rect 130764 500788 130765 500852
rect 130699 500787 130765 500788
rect 130702 498218 130762 500787
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 487040 127404 487898
rect 144804 487040 145404 502800
rect 149099 500580 149165 500581
rect 149099 500516 149100 500580
rect 149164 500516 149165 500580
rect 149099 500515 149165 500516
rect 147811 500308 147877 500309
rect 147811 500244 147812 500308
rect 147876 500244 147877 500308
rect 147811 500243 147877 500244
rect 147075 499628 147141 499629
rect 147075 499564 147076 499628
rect 147140 499564 147141 499628
rect 147075 499563 147141 499564
rect 23684 470454 24004 470476
rect 23684 470218 23726 470454
rect 23962 470218 24004 470454
rect 23684 470134 24004 470218
rect 23684 469898 23726 470134
rect 23962 469898 24004 470134
rect 23684 469876 24004 469898
rect 54404 470454 54724 470476
rect 54404 470218 54446 470454
rect 54682 470218 54724 470454
rect 54404 470134 54724 470218
rect 54404 469898 54446 470134
rect 54682 469898 54724 470134
rect 54404 469876 54724 469898
rect 85124 470454 85444 470476
rect 85124 470218 85166 470454
rect 85402 470218 85444 470454
rect 85124 470134 85444 470218
rect 85124 469898 85166 470134
rect 85402 469898 85444 470134
rect 85124 469876 85444 469898
rect 115844 470454 116164 470476
rect 115844 470218 115886 470454
rect 116122 470218 116164 470454
rect 115844 470134 116164 470218
rect 115844 469898 115886 470134
rect 116122 469898 116164 470134
rect 115844 469876 116164 469898
rect 146564 470454 146884 470476
rect 146564 470218 146606 470454
rect 146842 470218 146884 470454
rect 146564 470134 146884 470218
rect 146564 469898 146606 470134
rect 146842 469898 146884 470134
rect 146564 469876 146884 469898
rect 39044 452454 39364 452476
rect 39044 452218 39086 452454
rect 39322 452218 39364 452454
rect 39044 452134 39364 452218
rect 39044 451898 39086 452134
rect 39322 451898 39364 452134
rect 39044 451876 39364 451898
rect 69764 452454 70084 452476
rect 69764 452218 69806 452454
rect 70042 452218 70084 452454
rect 69764 452134 70084 452218
rect 69764 451898 69806 452134
rect 70042 451898 70084 452134
rect 69764 451876 70084 451898
rect 100484 452454 100804 452476
rect 100484 452218 100526 452454
rect 100762 452218 100804 452454
rect 100484 452134 100804 452218
rect 100484 451898 100526 452134
rect 100762 451898 100804 452134
rect 100484 451876 100804 451898
rect 131204 452454 131524 452476
rect 131204 452218 131246 452454
rect 131482 452218 131524 452454
rect 131204 452134 131524 452218
rect 131204 451898 131246 452134
rect 131482 451898 131524 452134
rect 131204 451876 131524 451898
rect 23684 434454 24004 434476
rect 23684 434218 23726 434454
rect 23962 434218 24004 434454
rect 23684 434134 24004 434218
rect 23684 433898 23726 434134
rect 23962 433898 24004 434134
rect 23684 433876 24004 433898
rect 54404 434454 54724 434476
rect 54404 434218 54446 434454
rect 54682 434218 54724 434454
rect 54404 434134 54724 434218
rect 54404 433898 54446 434134
rect 54682 433898 54724 434134
rect 54404 433876 54724 433898
rect 85124 434454 85444 434476
rect 85124 434218 85166 434454
rect 85402 434218 85444 434454
rect 85124 434134 85444 434218
rect 85124 433898 85166 434134
rect 85402 433898 85444 434134
rect 85124 433876 85444 433898
rect 115844 434454 116164 434476
rect 115844 434218 115886 434454
rect 116122 434218 116164 434454
rect 115844 434134 116164 434218
rect 115844 433898 115886 434134
rect 116122 433898 116164 434134
rect 115844 433876 116164 433898
rect 146564 434454 146884 434476
rect 146564 434218 146606 434454
rect 146842 434218 146884 434454
rect 146564 434134 146884 434218
rect 146564 433898 146606 434134
rect 146842 433898 146884 434134
rect 146564 433876 146884 433898
rect 39044 416454 39364 416476
rect 39044 416218 39086 416454
rect 39322 416218 39364 416454
rect 39044 416134 39364 416218
rect 39044 415898 39086 416134
rect 39322 415898 39364 416134
rect 39044 415876 39364 415898
rect 69764 416454 70084 416476
rect 69764 416218 69806 416454
rect 70042 416218 70084 416454
rect 69764 416134 70084 416218
rect 69764 415898 69806 416134
rect 70042 415898 70084 416134
rect 69764 415876 70084 415898
rect 100484 416454 100804 416476
rect 100484 416218 100526 416454
rect 100762 416218 100804 416454
rect 100484 416134 100804 416218
rect 100484 415898 100526 416134
rect 100762 415898 100804 416134
rect 100484 415876 100804 415898
rect 131204 416454 131524 416476
rect 131204 416218 131246 416454
rect 131482 416218 131524 416454
rect 131204 416134 131524 416218
rect 131204 415898 131246 416134
rect 131482 415898 131524 416134
rect 131204 415876 131524 415898
rect 36804 398454 37404 400000
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 384200 37404 397898
rect 54804 384200 55404 400000
rect 72804 398454 73404 400000
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 384200 73404 397898
rect 38875 380454 39195 380476
rect 38875 380218 38917 380454
rect 39153 380218 39195 380454
rect 38875 380134 39195 380218
rect 38875 379898 38917 380134
rect 39153 379898 39195 380134
rect 38875 379876 39195 379898
rect 56805 380454 57125 380476
rect 56805 380218 56847 380454
rect 57083 380218 57125 380454
rect 56805 380134 57125 380218
rect 56805 379898 56847 380134
rect 57083 379898 57125 380134
rect 56805 379876 57125 379898
rect 90804 380454 91404 400000
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 29909 362454 30229 362476
rect 29909 362218 29951 362454
rect 30187 362218 30229 362454
rect 29909 362134 30229 362218
rect 29909 361898 29951 362134
rect 30187 361898 30229 362134
rect 29909 361876 30229 361898
rect 47840 362454 48160 362476
rect 47840 362218 47882 362454
rect 48118 362218 48160 362454
rect 47840 362134 48160 362218
rect 47840 361898 47882 362134
rect 48118 361898 48160 362134
rect 47840 361876 48160 361898
rect 65770 362454 66090 362476
rect 65770 362218 65812 362454
rect 66048 362218 66090 362454
rect 65770 362134 66090 362218
rect 65770 361898 65812 362134
rect 66048 361898 66090 362134
rect 65770 361876 66090 361898
rect 20483 357372 20549 357373
rect 20483 357308 20484 357372
rect 20548 357308 20549 357372
rect 20483 357307 20549 357308
rect 36804 348912 37404 357000
rect 54804 348912 55404 357000
rect 72804 348912 73404 357000
rect 90804 348912 91404 379898
rect 108804 398454 109404 400000
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 348912 109404 361898
rect 126804 380454 127404 400000
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 348912 127404 379898
rect 144804 398454 145404 400000
rect 146891 398716 146957 398717
rect 146891 398652 146892 398716
rect 146956 398652 146957 398716
rect 146891 398651 146957 398652
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 146894 391370 146954 398651
rect 146710 391310 146954 391370
rect 146710 386613 146770 391310
rect 147078 389469 147138 499563
rect 147446 485893 147506 500022
rect 147627 499900 147693 499901
rect 147627 499836 147628 499900
rect 147692 499836 147693 499900
rect 147627 499835 147693 499836
rect 147443 485892 147509 485893
rect 147443 485828 147444 485892
rect 147508 485828 147509 485892
rect 147443 485827 147509 485828
rect 147259 485620 147325 485621
rect 147259 485556 147260 485620
rect 147324 485556 147325 485620
rect 147259 485555 147325 485556
rect 147262 417890 147322 485555
rect 147262 417830 147506 417890
rect 147446 398717 147506 417830
rect 147443 398716 147509 398717
rect 147443 398652 147444 398716
rect 147508 398652 147509 398716
rect 147443 398651 147509 398652
rect 147075 389468 147141 389469
rect 147075 389404 147076 389468
rect 147140 389404 147141 389468
rect 147075 389403 147141 389404
rect 146707 386612 146773 386613
rect 146707 386548 146708 386612
rect 146772 386548 146773 386612
rect 146707 386547 146773 386548
rect 147259 386612 147325 386613
rect 147259 386548 147260 386612
rect 147324 386548 147325 386612
rect 147259 386547 147325 386548
rect 147075 386476 147141 386477
rect 147075 386412 147076 386476
rect 147140 386412 147141 386476
rect 147075 386411 147141 386412
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 348912 145404 361898
rect 147078 360365 147138 386411
rect 147262 360501 147322 386547
rect 147259 360500 147325 360501
rect 147259 360436 147260 360500
rect 147324 360436 147325 360500
rect 147259 360435 147325 360436
rect 147075 360364 147141 360365
rect 147075 360300 147076 360364
rect 147140 360300 147141 360364
rect 147075 360299 147141 360300
rect 146891 360092 146957 360093
rect 146891 360028 146892 360092
rect 146956 360028 146957 360092
rect 146891 360027 146957 360028
rect 147075 360092 147141 360093
rect 147075 360028 147076 360092
rect 147140 360028 147141 360092
rect 147075 360027 147141 360028
rect 146894 350981 146954 360027
rect 147078 351797 147138 360027
rect 147075 351796 147141 351797
rect 147075 351732 147076 351796
rect 147140 351732 147141 351796
rect 147075 351731 147141 351732
rect 146891 350980 146957 350981
rect 146891 350916 146892 350980
rect 146956 350916 146957 350980
rect 146891 350915 146957 350916
rect 147630 350845 147690 499835
rect 147814 351797 147874 500243
rect 147995 500172 148061 500173
rect 147995 500108 147996 500172
rect 148060 500108 148061 500172
rect 147995 500107 148061 500108
rect 147811 351796 147877 351797
rect 147811 351732 147812 351796
rect 147876 351732 147877 351796
rect 147811 351731 147877 351732
rect 147998 351117 148058 500107
rect 148179 499628 148245 499629
rect 148179 499564 148180 499628
rect 148244 499564 148245 499628
rect 148179 499563 148245 499564
rect 148182 351797 148242 499563
rect 148363 497588 148429 497589
rect 148363 497524 148364 497588
rect 148428 497524 148429 497588
rect 148363 497523 148429 497524
rect 148179 351796 148245 351797
rect 148179 351732 148180 351796
rect 148244 351732 148245 351796
rect 148179 351731 148245 351732
rect 148366 351389 148426 497523
rect 148363 351388 148429 351389
rect 148363 351324 148364 351388
rect 148428 351324 148429 351388
rect 148363 351323 148429 351324
rect 149102 351253 149162 500515
rect 151859 500444 151925 500445
rect 151859 500380 151860 500444
rect 151924 500380 151925 500444
rect 151859 500379 151925 500380
rect 149651 499628 149717 499629
rect 149651 499564 149652 499628
rect 149716 499564 149717 499628
rect 149651 499563 149717 499564
rect 149835 499628 149901 499629
rect 149835 499564 149836 499628
rect 149900 499564 149901 499628
rect 149835 499563 149901 499564
rect 150939 499628 151005 499629
rect 150939 499564 150940 499628
rect 151004 499564 151005 499628
rect 150939 499563 151005 499564
rect 149283 497996 149349 497997
rect 149283 497932 149284 497996
rect 149348 497932 149349 497996
rect 149283 497931 149349 497932
rect 149099 351252 149165 351253
rect 149099 351188 149100 351252
rect 149164 351188 149165 351252
rect 149099 351187 149165 351188
rect 147995 351116 148061 351117
rect 147995 351052 147996 351116
rect 148060 351052 148061 351116
rect 147995 351051 148061 351052
rect 149286 350845 149346 497931
rect 149654 351797 149714 499563
rect 149838 351797 149898 499563
rect 150387 497860 150453 497861
rect 150387 497796 150388 497860
rect 150452 497796 150453 497860
rect 150387 497795 150453 497796
rect 149651 351796 149717 351797
rect 149651 351732 149652 351796
rect 149716 351732 149717 351796
rect 149651 351731 149717 351732
rect 149835 351796 149901 351797
rect 149835 351732 149836 351796
rect 149900 351732 149901 351796
rect 149835 351731 149901 351732
rect 150390 351661 150450 497795
rect 150755 497724 150821 497725
rect 150755 497660 150756 497724
rect 150820 497660 150821 497724
rect 150755 497659 150821 497660
rect 150571 497452 150637 497453
rect 150571 497388 150572 497452
rect 150636 497388 150637 497452
rect 150571 497387 150637 497388
rect 150387 351660 150453 351661
rect 150387 351596 150388 351660
rect 150452 351596 150453 351660
rect 150387 351595 150453 351596
rect 147627 350844 147693 350845
rect 147627 350780 147628 350844
rect 147692 350780 147693 350844
rect 147627 350779 147693 350780
rect 149283 350844 149349 350845
rect 149283 350780 149284 350844
rect 149348 350780 149349 350844
rect 149283 350779 149349 350780
rect 150574 350709 150634 497387
rect 150758 351525 150818 497659
rect 150942 351797 151002 499563
rect 151862 400893 151922 500379
rect 152411 499628 152477 499629
rect 152411 499564 152412 499628
rect 152476 499564 152477 499628
rect 152411 499563 152477 499564
rect 151859 400892 151925 400893
rect 151859 400828 151860 400892
rect 151924 400828 151925 400892
rect 151859 400827 151925 400828
rect 152414 351797 152474 499563
rect 154803 498132 154869 498133
rect 154803 498068 154804 498132
rect 154868 498068 154869 498132
rect 154803 498067 154869 498068
rect 153147 497316 153213 497317
rect 153147 497252 153148 497316
rect 153212 497252 153213 497316
rect 153147 497251 153213 497252
rect 153150 401165 153210 497251
rect 153334 401437 153394 497982
rect 153699 497724 153765 497725
rect 153699 497660 153700 497724
rect 153764 497660 153765 497724
rect 153699 497659 153765 497660
rect 153331 401436 153397 401437
rect 153331 401372 153332 401436
rect 153396 401372 153397 401436
rect 153331 401371 153397 401372
rect 153147 401164 153213 401165
rect 153147 401100 153148 401164
rect 153212 401100 153213 401164
rect 153147 401099 153213 401100
rect 150939 351796 151005 351797
rect 150939 351732 150940 351796
rect 151004 351732 151005 351796
rect 150939 351731 151005 351732
rect 152411 351796 152477 351797
rect 152411 351732 152412 351796
rect 152476 351732 152477 351796
rect 152411 351731 152477 351732
rect 150755 351524 150821 351525
rect 150755 351460 150756 351524
rect 150820 351460 150821 351524
rect 150755 351459 150821 351460
rect 153702 351389 153762 497659
rect 154619 497180 154685 497181
rect 154619 497116 154620 497180
rect 154684 497116 154685 497180
rect 154619 497115 154685 497116
rect 153883 403612 153949 403613
rect 153883 403548 153884 403612
rect 153948 403548 153949 403612
rect 153883 403547 153949 403548
rect 153886 364309 153946 403547
rect 154622 401301 154682 497115
rect 154619 401300 154685 401301
rect 154619 401236 154620 401300
rect 154684 401236 154685 401300
rect 154619 401235 154685 401236
rect 154806 401029 154866 498067
rect 162804 488454 163404 502800
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 154803 401028 154869 401029
rect 154803 400964 154804 401028
rect 154868 400964 154869 401028
rect 154803 400963 154869 400964
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 155723 376684 155789 376685
rect 155723 376620 155724 376684
rect 155788 376620 155789 376684
rect 155723 376619 155789 376620
rect 155726 369749 155786 376619
rect 155723 369748 155789 369749
rect 155723 369684 155724 369748
rect 155788 369684 155789 369748
rect 155723 369683 155789 369684
rect 153883 364308 153949 364309
rect 153883 364244 153884 364308
rect 153948 364244 153949 364308
rect 153883 364243 153949 364244
rect 153699 351388 153765 351389
rect 153699 351324 153700 351388
rect 153764 351324 153765 351388
rect 153699 351323 153765 351324
rect 150571 350708 150637 350709
rect 150571 350644 150572 350708
rect 150636 350644 150637 350708
rect 150571 350643 150637 350644
rect 162804 348912 163404 379898
rect 180804 470454 181404 502800
rect 189579 500852 189645 500853
rect 189579 500788 189580 500852
rect 189644 500788 189645 500852
rect 189579 500787 189645 500788
rect 191051 500852 191117 500853
rect 191051 500788 191052 500852
rect 191116 500788 191117 500852
rect 191051 500787 191117 500788
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 348912 181404 361898
rect 189582 351661 189642 500787
rect 189763 500716 189829 500717
rect 189763 500652 189764 500716
rect 189828 500652 189829 500716
rect 189763 500651 189829 500652
rect 189766 351797 189826 500651
rect 191054 351797 191114 500787
rect 198804 491600 199404 502800
rect 216804 491600 217404 502800
rect 234804 491600 235404 502800
rect 252804 491600 253404 502800
rect 270804 491600 271404 502800
rect 207614 488454 207934 488476
rect 207614 488218 207656 488454
rect 207892 488218 207934 488454
rect 207614 488134 207934 488218
rect 207614 487898 207656 488134
rect 207892 487898 207934 488134
rect 207614 487876 207934 487898
rect 238334 488454 238654 488476
rect 238334 488218 238376 488454
rect 238612 488218 238654 488454
rect 238334 488134 238654 488218
rect 238334 487898 238376 488134
rect 238612 487898 238654 488134
rect 238334 487876 238654 487898
rect 269054 488454 269374 488476
rect 269054 488218 269096 488454
rect 269332 488218 269374 488454
rect 269054 488134 269374 488218
rect 269054 487898 269096 488134
rect 269332 487898 269374 488134
rect 269054 487876 269374 487898
rect 192254 470454 192574 470476
rect 192254 470218 192296 470454
rect 192532 470218 192574 470454
rect 192254 470134 192574 470218
rect 192254 469898 192296 470134
rect 192532 469898 192574 470134
rect 192254 469876 192574 469898
rect 222974 470454 223294 470476
rect 222974 470218 223016 470454
rect 223252 470218 223294 470454
rect 222974 470134 223294 470218
rect 222974 469898 223016 470134
rect 223252 469898 223294 470134
rect 222974 469876 223294 469898
rect 253694 470454 254014 470476
rect 253694 470218 253736 470454
rect 253972 470218 254014 470454
rect 253694 470134 254014 470218
rect 253694 469898 253736 470134
rect 253972 469898 254014 470134
rect 253694 469876 254014 469898
rect 207614 452454 207934 452476
rect 207614 452218 207656 452454
rect 207892 452218 207934 452454
rect 207614 452134 207934 452218
rect 207614 451898 207656 452134
rect 207892 451898 207934 452134
rect 207614 451876 207934 451898
rect 238334 452454 238654 452476
rect 238334 452218 238376 452454
rect 238612 452218 238654 452454
rect 238334 452134 238654 452218
rect 238334 451898 238376 452134
rect 238612 451898 238654 452134
rect 238334 451876 238654 451898
rect 269054 452454 269374 452476
rect 269054 452218 269096 452454
rect 269332 452218 269374 452454
rect 269054 452134 269374 452218
rect 269054 451898 269096 452134
rect 269332 451898 269374 452134
rect 269054 451876 269374 451898
rect 192254 434454 192574 434476
rect 192254 434218 192296 434454
rect 192532 434218 192574 434454
rect 192254 434134 192574 434218
rect 192254 433898 192296 434134
rect 192532 433898 192574 434134
rect 192254 433876 192574 433898
rect 222974 434454 223294 434476
rect 222974 434218 223016 434454
rect 223252 434218 223294 434454
rect 222974 434134 223294 434218
rect 222974 433898 223016 434134
rect 223252 433898 223294 434134
rect 222974 433876 223294 433898
rect 253694 434454 254014 434476
rect 253694 434218 253736 434454
rect 253972 434218 254014 434454
rect 253694 434134 254014 434218
rect 253694 433898 253736 434134
rect 253972 433898 254014 434134
rect 253694 433876 254014 433898
rect 207614 416454 207934 416476
rect 207614 416218 207656 416454
rect 207892 416218 207934 416454
rect 207614 416134 207934 416218
rect 207614 415898 207656 416134
rect 207892 415898 207934 416134
rect 207614 415876 207934 415898
rect 238334 416454 238654 416476
rect 238334 416218 238376 416454
rect 238612 416218 238654 416454
rect 238334 416134 238654 416218
rect 238334 415898 238376 416134
rect 238612 415898 238654 416134
rect 238334 415876 238654 415898
rect 269054 416454 269374 416476
rect 269054 416218 269096 416454
rect 269332 416218 269374 416454
rect 269054 416134 269374 416218
rect 269054 415898 269096 416134
rect 269332 415898 269374 416134
rect 269054 415876 269374 415898
rect 198804 402224 199404 410000
rect 216804 402224 217404 410000
rect 234804 402224 235404 410000
rect 252804 402224 253404 410000
rect 270804 402224 271404 410000
rect 189763 351796 189829 351797
rect 189763 351732 189764 351796
rect 189828 351732 189829 351796
rect 189763 351731 189829 351732
rect 191051 351796 191117 351797
rect 191051 351732 191052 351796
rect 191116 351732 191117 351796
rect 191051 351731 191117 351732
rect 189579 351660 189645 351661
rect 189579 351596 189580 351660
rect 189644 351596 189645 351660
rect 189579 351595 189645 351596
rect 198804 348912 199404 358112
rect 216804 348912 217404 358112
rect 234804 348912 235404 358112
rect 252804 348912 253404 358112
rect 270804 348912 271404 358112
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 107675 344454 107995 344476
rect 107675 344218 107717 344454
rect 107953 344218 107995 344454
rect 107675 344134 107995 344218
rect 107675 343898 107717 344134
rect 107953 343898 107995 344134
rect 107675 343876 107995 343898
rect 192805 344454 193125 344476
rect 192805 344218 192847 344454
rect 193083 344218 193125 344454
rect 192805 344134 193125 344218
rect 192805 343898 192847 344134
rect 193083 343898 193125 344134
rect 192805 343876 193125 343898
rect 65109 326454 65429 326476
rect 65109 326218 65151 326454
rect 65387 326218 65429 326454
rect 65109 326134 65429 326218
rect 65109 325898 65151 326134
rect 65387 325898 65429 326134
rect 65109 325876 65429 325898
rect 150240 326454 150560 326476
rect 150240 326218 150282 326454
rect 150518 326218 150560 326454
rect 150240 326134 150560 326218
rect 150240 325898 150282 326134
rect 150518 325898 150560 326134
rect 150240 325876 150560 325898
rect 235370 326454 235690 326476
rect 235370 326218 235412 326454
rect 235648 326218 235690 326454
rect 235370 326134 235690 326218
rect 235370 325898 235412 326134
rect 235648 325898 235690 326134
rect 235370 325876 235690 325898
rect 36804 315600 37404 322800
rect 54804 315600 55404 322800
rect 72804 315600 73404 322800
rect 90804 315600 91404 322800
rect 108804 315600 109404 322800
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 39614 308454 39934 308476
rect 39614 308218 39656 308454
rect 39892 308218 39934 308454
rect 39614 308134 39934 308218
rect 39614 307898 39656 308134
rect 39892 307898 39934 308134
rect 39614 307876 39934 307898
rect 70334 308454 70654 308476
rect 70334 308218 70376 308454
rect 70612 308218 70654 308454
rect 70334 308134 70654 308218
rect 70334 307898 70376 308134
rect 70612 307898 70654 308134
rect 70334 307876 70654 307898
rect 101054 308454 101374 308476
rect 101054 308218 101096 308454
rect 101332 308218 101374 308454
rect 101054 308134 101374 308218
rect 101054 307898 101096 308134
rect 101332 307898 101374 308134
rect 101054 307876 101374 307898
rect 126804 308454 127404 322800
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 24254 290454 24574 290476
rect 24254 290218 24296 290454
rect 24532 290218 24574 290454
rect 24254 290134 24574 290218
rect 24254 289898 24296 290134
rect 24532 289898 24574 290134
rect 24254 289876 24574 289898
rect 54974 290454 55294 290476
rect 54974 290218 55016 290454
rect 55252 290218 55294 290454
rect 54974 290134 55294 290218
rect 54974 289898 55016 290134
rect 55252 289898 55294 290134
rect 54974 289876 55294 289898
rect 85694 290454 86014 290476
rect 85694 290218 85736 290454
rect 85972 290218 86014 290454
rect 85694 290134 86014 290218
rect 85694 289898 85736 290134
rect 85972 289898 86014 290134
rect 85694 289876 86014 289898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 39614 272454 39934 272476
rect 39614 272218 39656 272454
rect 39892 272218 39934 272454
rect 39614 272134 39934 272218
rect 39614 271898 39656 272134
rect 39892 271898 39934 272134
rect 39614 271876 39934 271898
rect 70334 272454 70654 272476
rect 70334 272218 70376 272454
rect 70612 272218 70654 272454
rect 70334 272134 70654 272218
rect 70334 271898 70376 272134
rect 70612 271898 70654 272134
rect 70334 271876 70654 271898
rect 101054 272454 101374 272476
rect 101054 272218 101096 272454
rect 101332 272218 101374 272454
rect 101054 272134 101374 272218
rect 101054 271898 101096 272134
rect 101332 271898 101374 272134
rect 101054 271876 101374 271898
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 24254 254454 24574 254476
rect 24254 254218 24296 254454
rect 24532 254218 24574 254454
rect 24254 254134 24574 254218
rect 24254 253898 24296 254134
rect 24532 253898 24574 254134
rect 24254 253876 24574 253898
rect 54974 254454 55294 254476
rect 54974 254218 55016 254454
rect 55252 254218 55294 254454
rect 54974 254134 55294 254218
rect 54974 253898 55016 254134
rect 55252 253898 55294 254134
rect 54974 253876 55294 253898
rect 85694 254454 86014 254476
rect 85694 254218 85736 254454
rect 85972 254218 86014 254454
rect 85694 254134 86014 254218
rect 85694 253898 85736 254134
rect 85972 253898 86014 254134
rect 85694 253876 86014 253898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 219708 19404 235898
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 36804 219708 37404 234000
rect 54804 219708 55404 234000
rect 72804 219708 73404 234000
rect 90804 219708 91404 234000
rect 108804 218454 109404 234000
rect 126804 221840 127404 235898
rect 144804 290454 145404 322800
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 221840 145404 253898
rect 162804 308454 163404 322800
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 221840 163404 235898
rect 180804 290454 181404 322800
rect 190131 320380 190197 320381
rect 190131 320316 190132 320380
rect 190196 320316 190197 320380
rect 190131 320315 190197 320316
rect 194363 320380 194429 320381
rect 194363 320316 194364 320380
rect 194428 320316 194429 320380
rect 194363 320315 194429 320316
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 221840 181404 253898
rect 190134 224501 190194 320315
rect 190315 320244 190381 320245
rect 190315 320180 190316 320244
rect 190380 320180 190381 320244
rect 190315 320179 190381 320180
rect 191603 320244 191669 320245
rect 191603 320180 191604 320244
rect 191668 320180 191669 320244
rect 191603 320179 191669 320180
rect 193075 320244 193141 320245
rect 193075 320180 193076 320244
rect 193140 320180 193141 320244
rect 193075 320179 193141 320180
rect 194179 320244 194245 320245
rect 194179 320180 194180 320244
rect 194244 320180 194245 320244
rect 194179 320179 194245 320180
rect 190131 224500 190197 224501
rect 190131 224436 190132 224500
rect 190196 224436 190197 224500
rect 190131 224435 190197 224436
rect 190318 224365 190378 320179
rect 191606 224637 191666 320179
rect 192208 290454 192528 290476
rect 192208 290218 192250 290454
rect 192486 290218 192528 290454
rect 192208 290134 192528 290218
rect 192208 289898 192250 290134
rect 192486 289898 192528 290134
rect 192208 289876 192528 289898
rect 192208 254454 192528 254476
rect 192208 254218 192250 254454
rect 192486 254218 192528 254454
rect 192208 254134 192528 254218
rect 192208 253898 192250 254134
rect 192486 253898 192528 254134
rect 192208 253876 192528 253898
rect 193078 224909 193138 320179
rect 193075 224908 193141 224909
rect 193075 224844 193076 224908
rect 193140 224844 193141 224908
rect 193075 224843 193141 224844
rect 191603 224636 191669 224637
rect 191603 224572 191604 224636
rect 191668 224572 191669 224636
rect 191603 224571 191669 224572
rect 190315 224364 190381 224365
rect 190315 224300 190316 224364
rect 190380 224300 190381 224364
rect 190315 224299 190381 224300
rect 194182 224229 194242 320179
rect 194366 224773 194426 320315
rect 198804 315600 199404 322800
rect 216804 315600 217404 322800
rect 219939 322148 220005 322149
rect 219939 322084 219940 322148
rect 220004 322084 220005 322148
rect 219939 322083 220005 322084
rect 207568 308454 207888 308476
rect 207568 308218 207610 308454
rect 207846 308218 207888 308454
rect 207568 308134 207888 308218
rect 207568 307898 207610 308134
rect 207846 307898 207888 308134
rect 207568 307876 207888 307898
rect 207568 272454 207888 272476
rect 207568 272218 207610 272454
rect 207846 272218 207888 272454
rect 207568 272134 207888 272218
rect 207568 271898 207610 272134
rect 207846 271898 207888 272134
rect 207568 271876 207888 271898
rect 194363 224772 194429 224773
rect 194363 224708 194364 224772
rect 194428 224708 194429 224772
rect 194363 224707 194429 224708
rect 194179 224228 194245 224229
rect 194179 224164 194180 224228
rect 194244 224164 194245 224228
rect 194179 224163 194245 224164
rect 198804 221840 199404 234000
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 28768 200454 29088 200476
rect 28768 200218 28810 200454
rect 29046 200218 29088 200454
rect 28768 200134 29088 200218
rect 28768 199898 28810 200134
rect 29046 199898 29088 200134
rect 28768 199876 29088 199898
rect 59488 200454 59808 200476
rect 59488 200218 59530 200454
rect 59766 200218 59808 200454
rect 59488 200134 59808 200218
rect 59488 199898 59530 200134
rect 59766 199898 59808 200134
rect 59488 199876 59808 199898
rect 90208 200454 90528 200476
rect 90208 200218 90250 200454
rect 90486 200218 90528 200454
rect 90208 200134 90528 200218
rect 90208 199898 90250 200134
rect 90486 199898 90528 200134
rect 90208 199876 90528 199898
rect 44128 182454 44448 182476
rect 44128 182218 44170 182454
rect 44406 182218 44448 182454
rect 44128 182134 44448 182218
rect 44128 181898 44170 182134
rect 44406 181898 44448 182134
rect 44128 181876 44448 181898
rect 74848 182454 75168 182476
rect 74848 182218 74890 182454
rect 75126 182218 75168 182454
rect 74848 182134 75168 182218
rect 74848 181898 74890 182134
rect 75126 181898 75168 182134
rect 74848 181876 75168 181898
rect 108804 182454 109404 217898
rect 123808 218454 124128 218476
rect 123808 218218 123850 218454
rect 124086 218218 124128 218454
rect 123808 218134 124128 218218
rect 123808 217898 123850 218134
rect 124086 217898 124128 218134
rect 123808 217876 124128 217898
rect 154528 218454 154848 218476
rect 154528 218218 154570 218454
rect 154806 218218 154848 218454
rect 154528 218134 154848 218218
rect 154528 217898 154570 218134
rect 154806 217898 154848 218134
rect 154528 217876 154848 217898
rect 185248 218454 185568 218476
rect 185248 218218 185290 218454
rect 185526 218218 185568 218454
rect 185248 218134 185568 218218
rect 185248 217898 185290 218134
rect 185526 217898 185568 218134
rect 185248 217876 185568 217898
rect 216804 218454 217404 234000
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 139168 200454 139488 200476
rect 139168 200218 139210 200454
rect 139446 200218 139488 200454
rect 139168 200134 139488 200218
rect 139168 199898 139210 200134
rect 139446 199898 139488 200134
rect 139168 199876 139488 199898
rect 169888 200454 170208 200476
rect 169888 200218 169930 200454
rect 170166 200218 170208 200454
rect 169888 200134 170208 200218
rect 169888 199898 169930 200134
rect 170166 199898 170208 200134
rect 169888 199876 170208 199898
rect 200608 200454 200928 200476
rect 200608 200218 200650 200454
rect 200886 200218 200928 200454
rect 200608 200134 200928 200218
rect 200608 199898 200650 200134
rect 200886 199898 200928 200134
rect 200608 199876 200928 199898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 28768 164454 29088 164476
rect 28768 164218 28810 164454
rect 29046 164218 29088 164454
rect 28768 164134 29088 164218
rect 28768 163898 28810 164134
rect 29046 163898 29088 164134
rect 28768 163876 29088 163898
rect 59488 164454 59808 164476
rect 59488 164218 59530 164454
rect 59766 164218 59808 164454
rect 59488 164134 59808 164218
rect 59488 163898 59530 164134
rect 59766 163898 59808 164134
rect 59488 163876 59808 163898
rect 90208 164454 90528 164476
rect 90208 164218 90250 164454
rect 90486 164218 90528 164454
rect 90208 164134 90528 164218
rect 90208 163898 90250 164134
rect 90486 163898 90528 164134
rect 90208 163876 90528 163898
rect 44128 146454 44448 146476
rect 44128 146218 44170 146454
rect 44406 146218 44448 146454
rect 44128 146134 44448 146218
rect 44128 145898 44170 146134
rect 44406 145898 44448 146134
rect 44128 145876 44448 145898
rect 74848 146454 75168 146476
rect 74848 146218 74890 146454
rect 75126 146218 75168 146454
rect 74848 146134 75168 146218
rect 74848 145898 74890 146134
rect 75126 145898 75168 146134
rect 74848 145876 75168 145898
rect 108804 146454 109404 181898
rect 123808 182454 124128 182476
rect 123808 182218 123850 182454
rect 124086 182218 124128 182454
rect 123808 182134 124128 182218
rect 123808 181898 123850 182134
rect 124086 181898 124128 182134
rect 123808 181876 124128 181898
rect 154528 182454 154848 182476
rect 154528 182218 154570 182454
rect 154806 182218 154848 182454
rect 154528 182134 154848 182218
rect 154528 181898 154570 182134
rect 154806 181898 154848 182134
rect 154528 181876 154848 181898
rect 185248 182454 185568 182476
rect 185248 182218 185290 182454
rect 185526 182218 185568 182454
rect 185248 182134 185568 182218
rect 185248 181898 185290 182134
rect 185526 181898 185568 182134
rect 185248 181876 185568 181898
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 139168 164454 139488 164476
rect 139168 164218 139210 164454
rect 139446 164218 139488 164454
rect 139168 164134 139488 164218
rect 139168 163898 139210 164134
rect 139446 163898 139488 164134
rect 139168 163876 139488 163898
rect 169888 164454 170208 164476
rect 169888 164218 169930 164454
rect 170166 164218 170208 164454
rect 169888 164134 170208 164218
rect 169888 163898 169930 164134
rect 170166 163898 170208 164134
rect 169888 163876 170208 163898
rect 200608 164454 200928 164476
rect 200608 164218 200650 164454
rect 200886 164218 200928 164454
rect 200608 164134 200928 164218
rect 200608 163898 200650 164134
rect 200886 163898 200928 164134
rect 200608 163876 200928 163898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 18643 124268 18709 124269
rect 18643 124204 18644 124268
rect 18708 124204 18709 124268
rect 18643 124203 18709 124204
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 18804 99440 19404 127228
rect 32259 125084 32325 125085
rect 32259 125020 32260 125084
rect 32324 125020 32325 125084
rect 32259 125019 32325 125020
rect 28768 92454 29088 92476
rect 28768 92218 28810 92454
rect 29046 92218 29088 92454
rect 28768 92134 29088 92218
rect 28768 91898 28810 92134
rect 29046 91898 29088 92134
rect 28768 91876 29088 91898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 13408 74454 13728 74476
rect 13408 74218 13450 74454
rect 13686 74218 13728 74454
rect 13408 74134 13728 74218
rect 13408 73898 13450 74134
rect 13686 73898 13728 74134
rect 13408 73876 13728 73898
rect 28768 56454 29088 56476
rect 28768 56218 28810 56454
rect 29046 56218 29088 56454
rect 28768 56134 29088 56218
rect 28768 55898 28810 56134
rect 29046 55898 29088 56134
rect 28768 55876 29088 55898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 13408 38454 13728 38476
rect 13408 38218 13450 38454
rect 13686 38218 13728 38454
rect 13408 38134 13728 38218
rect 13408 37898 13450 38134
rect 13686 37898 13728 38134
rect 13408 37876 13728 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 18804 20454 19404 31440
rect 32262 30293 32322 125019
rect 36804 110454 37404 127228
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 99440 37404 109898
rect 54804 99440 55404 127228
rect 72804 110454 73404 127228
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 99440 73404 109898
rect 90804 99440 91404 127228
rect 108804 110454 109404 145898
rect 123808 146454 124128 146476
rect 123808 146218 123850 146454
rect 124086 146218 124128 146454
rect 123808 146134 124128 146218
rect 123808 145898 123850 146134
rect 124086 145898 124128 146134
rect 123808 145876 124128 145898
rect 154528 146454 154848 146476
rect 154528 146218 154570 146454
rect 154806 146218 154848 146454
rect 154528 146134 154848 146218
rect 154528 145898 154570 146134
rect 154806 145898 154848 146134
rect 154528 145876 154848 145898
rect 185248 146454 185568 146476
rect 185248 146218 185290 146454
rect 185526 146218 185568 146454
rect 185248 146134 185568 146218
rect 185248 145898 185290 146134
rect 185526 145898 185568 146134
rect 185248 145876 185568 145898
rect 216804 146454 217404 181898
rect 219942 158813 220002 322083
rect 234804 315600 235404 322800
rect 252804 315600 253404 322800
rect 270804 315600 271404 322800
rect 238288 308454 238608 308476
rect 238288 308218 238330 308454
rect 238566 308218 238608 308454
rect 238288 308134 238608 308218
rect 238288 307898 238330 308134
rect 238566 307898 238608 308134
rect 238288 307876 238608 307898
rect 269008 308454 269328 308476
rect 269008 308218 269050 308454
rect 269286 308218 269328 308454
rect 269008 308134 269328 308218
rect 269008 307898 269050 308134
rect 269286 307898 269328 308134
rect 269008 307876 269328 307898
rect 222928 290454 223248 290476
rect 222928 290218 222970 290454
rect 223206 290218 223248 290454
rect 222928 290134 223248 290218
rect 222928 289898 222970 290134
rect 223206 289898 223248 290134
rect 222928 289876 223248 289898
rect 253648 290454 253968 290476
rect 253648 290218 253690 290454
rect 253926 290218 253968 290454
rect 253648 290134 253968 290218
rect 253648 289898 253690 290134
rect 253926 289898 253968 290134
rect 253648 289876 253968 289898
rect 238288 272454 238608 272476
rect 238288 272218 238330 272454
rect 238566 272218 238608 272454
rect 238288 272134 238608 272218
rect 238288 271898 238330 272134
rect 238566 271898 238608 272134
rect 238288 271876 238608 271898
rect 269008 272454 269328 272476
rect 269008 272218 269050 272454
rect 269286 272218 269328 272454
rect 269008 272134 269328 272218
rect 269008 271898 269050 272134
rect 269286 271898 269328 272134
rect 269008 271876 269328 271898
rect 222928 254454 223248 254476
rect 222928 254218 222970 254454
rect 223206 254218 223248 254454
rect 222928 254134 223248 254218
rect 222928 253898 222970 254134
rect 223206 253898 223248 254134
rect 222928 253876 223248 253898
rect 253648 254454 253968 254476
rect 253648 254218 253690 254454
rect 253926 254218 253968 254454
rect 253648 254134 253968 254218
rect 253648 253898 253690 254134
rect 253926 253898 253968 254134
rect 253648 253876 253968 253898
rect 280110 235245 280170 619515
rect 280662 473789 280722 667931
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 280659 473788 280725 473789
rect 280659 473724 280660 473788
rect 280724 473724 280725 473788
rect 280659 473723 280725 473724
rect 288804 470454 289404 505898
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 317091 700636 317157 700637
rect 317091 700572 317092 700636
rect 317156 700572 317157 700636
rect 317091 700571 317157 700572
rect 316907 700364 316973 700365
rect 316907 700300 316908 700364
rect 316972 700300 316973 700364
rect 316907 700299 316973 700300
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 299427 473924 299493 473925
rect 299427 473860 299428 473924
rect 299492 473860 299493 473924
rect 299427 473859 299493 473860
rect 299430 473653 299490 473859
rect 299427 473652 299493 473653
rect 299427 473588 299428 473652
rect 299492 473588 299493 473652
rect 299427 473587 299493 473588
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 326454 289404 361898
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 316910 428637 316970 700299
rect 317094 428773 317154 700571
rect 317275 700500 317341 700501
rect 317275 700436 317276 700500
rect 317340 700436 317341 700500
rect 317275 700435 317341 700436
rect 317091 428772 317157 428773
rect 317091 428708 317092 428772
rect 317156 428708 317157 428772
rect 317091 428707 317157 428708
rect 316907 428636 316973 428637
rect 316907 428572 316908 428636
rect 316972 428572 316973 428636
rect 316907 428571 316973 428572
rect 317278 428501 317338 700435
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 657040 325404 685898
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 657040 343404 667898
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 657040 361404 685898
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 657040 379404 667898
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 657040 397404 685898
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 657040 415404 667898
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 657040 433404 685898
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 657040 451404 667898
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 662480 469404 685898
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 662480 487404 667898
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 492443 663916 492509 663917
rect 492443 663852 492444 663916
rect 492508 663852 492509 663916
rect 492443 663851 492509 663852
rect 323730 650454 324050 650476
rect 323730 650218 323772 650454
rect 324008 650218 324050 650454
rect 323730 650134 324050 650218
rect 323730 649898 323772 650134
rect 324008 649898 324050 650134
rect 323730 649876 324050 649898
rect 354450 650454 354770 650476
rect 354450 650218 354492 650454
rect 354728 650218 354770 650454
rect 354450 650134 354770 650218
rect 354450 649898 354492 650134
rect 354728 649898 354770 650134
rect 354450 649876 354770 649898
rect 385170 650454 385490 650476
rect 385170 650218 385212 650454
rect 385448 650218 385490 650454
rect 385170 650134 385490 650218
rect 385170 649898 385212 650134
rect 385448 649898 385490 650134
rect 385170 649876 385490 649898
rect 415890 650454 416210 650476
rect 415890 650218 415932 650454
rect 416168 650218 416210 650454
rect 415890 650134 416210 650218
rect 415890 649898 415932 650134
rect 416168 649898 416210 650134
rect 415890 649876 416210 649898
rect 446610 650454 446930 650476
rect 446610 650218 446652 650454
rect 446888 650218 446930 650454
rect 446610 650134 446930 650218
rect 446610 649898 446652 650134
rect 446888 649898 446930 650134
rect 446610 649876 446930 649898
rect 464208 650454 464528 650476
rect 464208 650218 464250 650454
rect 464486 650218 464528 650454
rect 464208 650134 464528 650218
rect 464208 649898 464250 650134
rect 464486 649898 464528 650134
rect 464208 649876 464528 649898
rect 339090 632454 339410 632476
rect 339090 632218 339132 632454
rect 339368 632218 339410 632454
rect 339090 632134 339410 632218
rect 339090 631898 339132 632134
rect 339368 631898 339410 632134
rect 339090 631876 339410 631898
rect 369810 632454 370130 632476
rect 369810 632218 369852 632454
rect 370088 632218 370130 632454
rect 369810 632134 370130 632218
rect 369810 631898 369852 632134
rect 370088 631898 370130 632134
rect 369810 631876 370130 631898
rect 400530 632454 400850 632476
rect 400530 632218 400572 632454
rect 400808 632218 400850 632454
rect 400530 632134 400850 632218
rect 400530 631898 400572 632134
rect 400808 631898 400850 632134
rect 400530 631876 400850 631898
rect 431250 632454 431570 632476
rect 431250 632218 431292 632454
rect 431528 632218 431570 632454
rect 431250 632134 431570 632218
rect 431250 631898 431292 632134
rect 431528 631898 431570 632134
rect 431250 631876 431570 631898
rect 479568 632454 479888 632476
rect 479568 632218 479610 632454
rect 479846 632218 479888 632454
rect 479568 632134 479888 632218
rect 479568 631898 479610 632134
rect 479846 631898 479888 632134
rect 479568 631876 479888 631898
rect 323730 614454 324050 614476
rect 323730 614218 323772 614454
rect 324008 614218 324050 614454
rect 323730 614134 324050 614218
rect 323730 613898 323772 614134
rect 324008 613898 324050 614134
rect 323730 613876 324050 613898
rect 354450 614454 354770 614476
rect 354450 614218 354492 614454
rect 354728 614218 354770 614454
rect 354450 614134 354770 614218
rect 354450 613898 354492 614134
rect 354728 613898 354770 614134
rect 354450 613876 354770 613898
rect 385170 614454 385490 614476
rect 385170 614218 385212 614454
rect 385448 614218 385490 614454
rect 385170 614134 385490 614218
rect 385170 613898 385212 614134
rect 385448 613898 385490 614134
rect 385170 613876 385490 613898
rect 415890 614454 416210 614476
rect 415890 614218 415932 614454
rect 416168 614218 416210 614454
rect 415890 614134 416210 614218
rect 415890 613898 415932 614134
rect 416168 613898 416210 614134
rect 415890 613876 416210 613898
rect 446610 614454 446930 614476
rect 446610 614218 446652 614454
rect 446888 614218 446930 614454
rect 446610 614134 446930 614218
rect 446610 613898 446652 614134
rect 446888 613898 446930 614134
rect 446610 613876 446930 613898
rect 464208 614454 464528 614476
rect 464208 614218 464250 614454
rect 464486 614218 464528 614454
rect 464208 614134 464528 614218
rect 464208 613898 464250 614134
rect 464486 613898 464528 614134
rect 464208 613876 464528 613898
rect 339090 596454 339410 596476
rect 339090 596218 339132 596454
rect 339368 596218 339410 596454
rect 339090 596134 339410 596218
rect 339090 595898 339132 596134
rect 339368 595898 339410 596134
rect 339090 595876 339410 595898
rect 369810 596454 370130 596476
rect 369810 596218 369852 596454
rect 370088 596218 370130 596454
rect 369810 596134 370130 596218
rect 369810 595898 369852 596134
rect 370088 595898 370130 596134
rect 369810 595876 370130 595898
rect 400530 596454 400850 596476
rect 400530 596218 400572 596454
rect 400808 596218 400850 596454
rect 400530 596134 400850 596218
rect 400530 595898 400572 596134
rect 400808 595898 400850 596134
rect 400530 595876 400850 595898
rect 431250 596454 431570 596476
rect 431250 596218 431292 596454
rect 431528 596218 431570 596454
rect 431250 596134 431570 596218
rect 431250 595898 431292 596134
rect 431528 595898 431570 596134
rect 431250 595876 431570 595898
rect 479568 596454 479888 596476
rect 479568 596218 479610 596454
rect 479846 596218 479888 596454
rect 479568 596134 479888 596218
rect 479568 595898 479610 596134
rect 479846 595898 479888 596134
rect 479568 595876 479888 595898
rect 323730 578454 324050 578476
rect 323730 578218 323772 578454
rect 324008 578218 324050 578454
rect 323730 578134 324050 578218
rect 323730 577898 323772 578134
rect 324008 577898 324050 578134
rect 323730 577876 324050 577898
rect 354450 578454 354770 578476
rect 354450 578218 354492 578454
rect 354728 578218 354770 578454
rect 354450 578134 354770 578218
rect 354450 577898 354492 578134
rect 354728 577898 354770 578134
rect 354450 577876 354770 577898
rect 385170 578454 385490 578476
rect 385170 578218 385212 578454
rect 385448 578218 385490 578454
rect 385170 578134 385490 578218
rect 385170 577898 385212 578134
rect 385448 577898 385490 578134
rect 385170 577876 385490 577898
rect 415890 578454 416210 578476
rect 415890 578218 415932 578454
rect 416168 578218 416210 578454
rect 415890 578134 416210 578218
rect 415890 577898 415932 578134
rect 416168 577898 416210 578134
rect 415890 577876 416210 577898
rect 446610 578454 446930 578476
rect 446610 578218 446652 578454
rect 446888 578218 446930 578454
rect 446610 578134 446930 578218
rect 446610 577898 446652 578134
rect 446888 577898 446930 578134
rect 446610 577876 446930 577898
rect 464208 578454 464528 578476
rect 464208 578218 464250 578454
rect 464486 578218 464528 578454
rect 464208 578134 464528 578218
rect 464208 577898 464250 578134
rect 464486 577898 464528 578134
rect 464208 577876 464528 577898
rect 324804 542454 325404 570000
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 528912 325404 541898
rect 342804 560454 343404 570000
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 528912 343404 559898
rect 360804 542454 361404 570000
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 528912 361404 541898
rect 378804 560454 379404 570000
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 528912 379404 559898
rect 396804 542454 397404 570000
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 528912 397404 541898
rect 414804 560454 415404 570000
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 528912 415404 559898
rect 432804 542454 433404 570000
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 528912 433404 541898
rect 450804 560454 451404 570000
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 528912 451404 559898
rect 468804 542454 469404 570000
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 528912 469404 541898
rect 486804 560454 487404 570000
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 528912 487404 559898
rect 492446 531181 492506 663851
rect 504804 662480 505404 685898
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 662480 523404 667898
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 662480 541404 685898
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 493915 662148 493981 662149
rect 493915 662084 493916 662148
rect 493980 662084 493981 662148
rect 493915 662083 493981 662084
rect 493918 531317 493978 662083
rect 551323 660108 551389 660109
rect 551323 660044 551324 660108
rect 551388 660044 551389 660108
rect 551323 660043 551389 660044
rect 551326 659970 551386 660043
rect 549854 659910 551386 659970
rect 494928 650454 495248 650476
rect 494928 650218 494970 650454
rect 495206 650218 495248 650454
rect 494928 650134 495248 650218
rect 494928 649898 494970 650134
rect 495206 649898 495248 650134
rect 494928 649876 495248 649898
rect 525648 650454 525968 650476
rect 525648 650218 525690 650454
rect 525926 650218 525968 650454
rect 525648 650134 525968 650218
rect 525648 649898 525690 650134
rect 525926 649898 525968 650134
rect 525648 649876 525968 649898
rect 510288 632454 510608 632476
rect 510288 632218 510330 632454
rect 510566 632218 510608 632454
rect 510288 632134 510608 632218
rect 510288 631898 510330 632134
rect 510566 631898 510608 632134
rect 510288 631876 510608 631898
rect 541008 632454 541328 632476
rect 541008 632218 541050 632454
rect 541286 632218 541328 632454
rect 541008 632134 541328 632218
rect 541008 631898 541050 632134
rect 541286 631898 541328 632134
rect 541008 631876 541328 631898
rect 494928 614454 495248 614476
rect 494928 614218 494970 614454
rect 495206 614218 495248 614454
rect 494928 614134 495248 614218
rect 494928 613898 494970 614134
rect 495206 613898 495248 614134
rect 494928 613876 495248 613898
rect 525648 614454 525968 614476
rect 525648 614218 525690 614454
rect 525926 614218 525968 614454
rect 525648 614134 525968 614218
rect 525648 613898 525690 614134
rect 525926 613898 525968 614134
rect 525648 613876 525968 613898
rect 510288 596454 510608 596476
rect 510288 596218 510330 596454
rect 510566 596218 510608 596454
rect 510288 596134 510608 596218
rect 510288 595898 510330 596134
rect 510566 595898 510608 596134
rect 510288 595876 510608 595898
rect 541008 596454 541328 596476
rect 541008 596218 541050 596454
rect 541286 596218 541328 596454
rect 541008 596134 541328 596218
rect 541008 595898 541050 596134
rect 541286 595898 541328 596134
rect 541008 595876 541328 595898
rect 494928 578454 495248 578476
rect 494928 578218 494970 578454
rect 495206 578218 495248 578454
rect 494928 578134 495248 578218
rect 494928 577898 494970 578134
rect 495206 577898 495248 578134
rect 494928 577876 495248 577898
rect 525648 578454 525968 578476
rect 525648 578218 525690 578454
rect 525926 578218 525968 578454
rect 525648 578134 525968 578218
rect 525648 577898 525690 578134
rect 525926 577898 525968 578134
rect 525648 577876 525968 577898
rect 549486 573474 549546 588422
rect 549854 574378 549914 659910
rect 553347 659428 553413 659429
rect 553347 659364 553348 659428
rect 553412 659364 553413 659428
rect 553347 659363 553413 659364
rect 551323 657932 551389 657933
rect 551323 657930 551324 657932
rect 551142 657870 551324 657930
rect 551142 651130 551202 657870
rect 551323 657868 551324 657870
rect 551388 657868 551389 657932
rect 551323 657867 551389 657868
rect 552059 655620 552125 655621
rect 552059 655556 552060 655620
rect 552124 655556 552125 655620
rect 552059 655555 552125 655556
rect 550774 651070 551202 651130
rect 550774 640930 550834 651070
rect 551323 650588 551389 650589
rect 551323 650524 551324 650588
rect 551388 650524 551389 650588
rect 551323 650523 551389 650524
rect 551326 650450 551386 650523
rect 551142 650390 551386 650450
rect 551142 647050 551202 650390
rect 551142 646990 551754 647050
rect 551507 646644 551573 646645
rect 551507 646580 551508 646644
rect 551572 646580 551573 646644
rect 551507 646579 551573 646580
rect 551323 645828 551389 645829
rect 551323 645764 551324 645828
rect 551388 645764 551389 645828
rect 551323 645763 551389 645764
rect 551326 642970 551386 645763
rect 550406 640870 550834 640930
rect 550958 642910 551386 642970
rect 550406 640250 550466 640870
rect 550406 640190 550650 640250
rect 550590 629370 550650 640190
rect 550590 629310 550834 629370
rect 550774 602170 550834 629310
rect 550222 602110 550834 602170
rect 550222 598090 550282 602110
rect 550222 598030 550650 598090
rect 550590 577690 550650 598030
rect 550958 585170 551018 642910
rect 551510 630733 551570 646579
rect 551694 630869 551754 646990
rect 551691 630868 551757 630869
rect 551691 630804 551692 630868
rect 551756 630804 551757 630868
rect 551691 630803 551757 630804
rect 551507 630732 551573 630733
rect 551507 630668 551508 630732
rect 551572 630668 551573 630732
rect 551507 630667 551573 630668
rect 551691 630596 551757 630597
rect 551691 630532 551692 630596
rect 551756 630532 551757 630596
rect 551691 630531 551757 630532
rect 551323 628012 551389 628013
rect 551323 628010 551324 628012
rect 551142 627950 551324 628010
rect 551142 602850 551202 627950
rect 551323 627948 551324 627950
rect 551388 627948 551389 628012
rect 551323 627947 551389 627948
rect 551694 616317 551754 630531
rect 551691 616316 551757 616317
rect 551691 616252 551692 616316
rect 551756 616252 551757 616316
rect 551691 616251 551757 616252
rect 551507 612780 551573 612781
rect 551507 612716 551508 612780
rect 551572 612716 551573 612780
rect 551507 612715 551573 612716
rect 551510 604890 551570 612715
rect 551510 604830 551800 604890
rect 551740 604349 551800 604830
rect 551737 604348 551803 604349
rect 551737 604284 551738 604348
rect 551802 604284 551803 604348
rect 551737 604283 551803 604284
rect 551323 602852 551389 602853
rect 551323 602850 551324 602852
rect 551142 602790 551324 602850
rect 551323 602788 551324 602790
rect 551388 602788 551389 602852
rect 551323 602787 551389 602788
rect 551691 602852 551757 602853
rect 551691 602788 551692 602852
rect 551756 602788 551757 602852
rect 551691 602787 551757 602788
rect 551694 593469 551754 602787
rect 551875 594012 551941 594013
rect 551875 593948 551876 594012
rect 551940 593948 551941 594012
rect 551875 593947 551941 593948
rect 551323 593468 551389 593469
rect 551323 593404 551324 593468
rect 551388 593404 551389 593468
rect 551323 593403 551389 593404
rect 551691 593468 551757 593469
rect 551691 593404 551692 593468
rect 551756 593404 551757 593468
rect 551691 593403 551757 593404
rect 551326 593330 551386 593403
rect 551326 593270 551754 593330
rect 550958 585110 551386 585170
rect 551326 583810 551386 585110
rect 550958 583750 551386 583810
rect 550958 578370 551018 583750
rect 551694 582589 551754 593270
rect 551691 582588 551757 582589
rect 551691 582524 551692 582588
rect 551756 582524 551757 582588
rect 551691 582523 551757 582524
rect 551878 582450 551938 593947
rect 550406 577630 550650 577690
rect 550774 578310 551018 578370
rect 551694 582390 551938 582450
rect 550406 576330 550466 577630
rect 550774 577010 550834 578310
rect 551694 577013 551754 582390
rect 551875 582316 551941 582317
rect 551875 582252 551876 582316
rect 551940 582252 551941 582316
rect 551875 582251 551941 582252
rect 551323 577012 551389 577013
rect 550774 576950 551018 577010
rect 550406 576270 550834 576330
rect 549486 573414 550650 573474
rect 504804 542454 505404 570000
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 493915 531316 493981 531317
rect 492443 531180 492509 531181
rect 492443 531116 492444 531180
rect 492508 531116 492509 531180
rect 492443 531115 492509 531116
rect 493550 529957 493610 531302
rect 493915 531252 493916 531316
rect 493980 531252 493981 531316
rect 493915 531251 493981 531252
rect 493547 529956 493613 529957
rect 493547 529892 493548 529956
rect 493612 529892 493613 529956
rect 493547 529891 493613 529892
rect 504804 528912 505404 541898
rect 522804 560454 523404 570000
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 528912 523404 559898
rect 540804 542454 541404 570000
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 528912 541404 541898
rect 549854 531538 549914 572782
rect 550590 567629 550650 573414
rect 550774 570485 550834 576270
rect 550771 570484 550837 570485
rect 550771 570420 550772 570484
rect 550836 570420 550837 570484
rect 550771 570419 550837 570420
rect 550587 567628 550653 567629
rect 550587 567564 550588 567628
rect 550652 567564 550653 567628
rect 550587 567563 550653 567564
rect 550587 558244 550653 558245
rect 550587 558180 550588 558244
rect 550652 558180 550653 558244
rect 550587 558179 550653 558180
rect 550590 532133 550650 558179
rect 550771 554028 550837 554029
rect 550771 553964 550772 554028
rect 550836 553964 550837 554028
rect 550771 553963 550837 553964
rect 550774 532541 550834 553963
rect 550958 532677 551018 576950
rect 551323 576948 551324 577012
rect 551388 576948 551389 577012
rect 551323 576947 551389 576948
rect 551691 577012 551757 577013
rect 551691 576948 551692 577012
rect 551756 576948 551757 577012
rect 551691 576947 551757 576948
rect 551326 563277 551386 576947
rect 551878 573477 551938 582251
rect 551507 573476 551573 573477
rect 551507 573412 551508 573476
rect 551572 573412 551573 573476
rect 551507 573411 551573 573412
rect 551875 573476 551941 573477
rect 551875 573412 551876 573476
rect 551940 573412 551941 573476
rect 551875 573411 551941 573412
rect 551510 570077 551570 573411
rect 551691 570484 551757 570485
rect 551691 570420 551692 570484
rect 551756 570420 551757 570484
rect 551691 570419 551757 570420
rect 551507 570076 551573 570077
rect 551507 570012 551508 570076
rect 551572 570012 551573 570076
rect 551507 570011 551573 570012
rect 551323 563276 551389 563277
rect 551323 563212 551324 563276
rect 551388 563212 551389 563276
rect 551323 563211 551389 563212
rect 551323 563004 551389 563005
rect 551323 562940 551324 563004
rect 551388 562940 551389 563004
rect 551323 562939 551389 562940
rect 551139 543828 551205 543829
rect 551139 543764 551140 543828
rect 551204 543764 551205 543828
rect 551139 543763 551205 543764
rect 551142 543693 551202 543763
rect 551139 543692 551205 543693
rect 551139 543628 551140 543692
rect 551204 543628 551205 543692
rect 551139 543627 551205 543628
rect 550955 532676 551021 532677
rect 550955 532612 550956 532676
rect 551020 532612 551021 532676
rect 550955 532611 551021 532612
rect 550771 532540 550837 532541
rect 550771 532476 550772 532540
rect 550836 532476 550837 532540
rect 550771 532475 550837 532476
rect 550587 532132 550653 532133
rect 550587 532068 550588 532132
rect 550652 532068 550653 532132
rect 550587 532067 550653 532068
rect 551326 530773 551386 562939
rect 551507 559060 551573 559061
rect 551507 558996 551508 559060
rect 551572 558996 551573 559060
rect 551507 558995 551573 558996
rect 551510 554029 551570 558995
rect 551694 558245 551754 570419
rect 551875 570076 551941 570077
rect 551875 570012 551876 570076
rect 551940 570012 551941 570076
rect 551875 570011 551941 570012
rect 551878 567765 551938 570011
rect 551875 567764 551941 567765
rect 551875 567700 551876 567764
rect 551940 567700 551941 567764
rect 551875 567699 551941 567700
rect 551875 567628 551941 567629
rect 551875 567564 551876 567628
rect 551940 567564 551941 567628
rect 551875 567563 551941 567564
rect 551691 558244 551757 558245
rect 551691 558180 551692 558244
rect 551756 558180 551757 558244
rect 551691 558179 551757 558180
rect 551507 554028 551573 554029
rect 551507 553964 551508 554028
rect 551572 553964 551573 554028
rect 551507 553963 551573 553964
rect 551878 543829 551938 567563
rect 551875 543828 551941 543829
rect 551875 543764 551876 543828
rect 551940 543764 551941 543828
rect 551875 543763 551941 543764
rect 551507 543692 551573 543693
rect 551507 543628 551508 543692
rect 551572 543628 551573 543692
rect 551507 543627 551573 543628
rect 551510 533629 551570 543627
rect 551507 533628 551573 533629
rect 551507 533564 551508 533628
rect 551572 533564 551573 533628
rect 551507 533563 551573 533564
rect 552062 532405 552122 655555
rect 552243 641068 552309 641069
rect 552243 641004 552244 641068
rect 552308 641004 552309 641068
rect 552243 641003 552309 641004
rect 552059 532404 552125 532405
rect 552059 532340 552060 532404
rect 552124 532340 552125 532404
rect 552059 532339 552125 532340
rect 552246 531861 552306 641003
rect 552427 636308 552493 636309
rect 552427 636244 552428 636308
rect 552492 636244 552493 636308
rect 552427 636243 552493 636244
rect 552243 531860 552309 531861
rect 552243 531796 552244 531860
rect 552308 531796 552309 531860
rect 552243 531795 552309 531796
rect 552430 531725 552490 636243
rect 552795 631412 552861 631413
rect 552795 631348 552796 631412
rect 552860 631348 552861 631412
rect 552795 631347 552861 631348
rect 552611 626516 552677 626517
rect 552611 626452 552612 626516
rect 552676 626452 552677 626516
rect 552611 626451 552677 626452
rect 552427 531724 552493 531725
rect 552427 531660 552428 531724
rect 552492 531660 552493 531724
rect 552427 531659 552493 531660
rect 552614 530909 552674 626451
rect 552798 547093 552858 631347
rect 552795 547092 552861 547093
rect 552795 547028 552796 547092
rect 552860 547028 552861 547092
rect 552795 547027 552861 547028
rect 552611 530908 552677 530909
rect 552611 530844 552612 530908
rect 552676 530844 552677 530908
rect 552611 530843 552677 530844
rect 551323 530772 551389 530773
rect 551323 530708 551324 530772
rect 551388 530708 551389 530772
rect 551323 530707 551389 530708
rect 553350 530637 553410 659363
rect 553531 656980 553597 656981
rect 553531 656916 553532 656980
rect 553596 656916 553597 656980
rect 553531 656915 553597 656916
rect 553534 531997 553594 656915
rect 553899 654532 553965 654533
rect 553899 654468 553900 654532
rect 553964 654468 553965 654532
rect 553899 654467 553965 654468
rect 553715 653308 553781 653309
rect 553715 653244 553716 653308
rect 553780 653244 553781 653308
rect 553715 653243 553781 653244
rect 553718 532269 553778 653243
rect 553902 533357 553962 654467
rect 554083 652084 554149 652085
rect 554083 652020 554084 652084
rect 554148 652020 554149 652084
rect 554083 652019 554149 652020
rect 554086 533493 554146 652019
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 554083 533492 554149 533493
rect 554083 533428 554084 533492
rect 554148 533428 554149 533492
rect 554083 533427 554149 533428
rect 553899 533356 553965 533357
rect 553899 533292 553900 533356
rect 553964 533292 553965 533356
rect 553899 533291 553965 533292
rect 553715 532268 553781 532269
rect 553715 532204 553716 532268
rect 553780 532204 553781 532268
rect 553715 532203 553781 532204
rect 553531 531996 553597 531997
rect 553531 531932 553532 531996
rect 553596 531932 553597 531996
rect 553531 531931 553597 531932
rect 553347 530636 553413 530637
rect 553347 530572 553348 530636
rect 553412 530572 553413 530636
rect 553347 530571 553413 530572
rect 558804 528912 559404 559898
rect 576804 704838 577404 705800
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 574875 527780 574941 527781
rect 574875 527716 574876 527780
rect 574940 527716 574941 527780
rect 574875 527715 574941 527716
rect 403721 524454 404041 524476
rect 403721 524218 403763 524454
rect 403999 524218 404041 524454
rect 403721 524134 404041 524218
rect 403721 523898 403763 524134
rect 403999 523898 404041 524134
rect 403721 523876 404041 523898
rect 488851 524454 489171 524476
rect 488851 524218 488893 524454
rect 489129 524218 489171 524454
rect 488851 524134 489171 524218
rect 488851 523898 488893 524134
rect 489129 523898 489171 524134
rect 488851 523876 489171 523898
rect 361155 506454 361475 506476
rect 361155 506218 361197 506454
rect 361433 506218 361475 506454
rect 361155 506134 361475 506218
rect 361155 505898 361197 506134
rect 361433 505898 361475 506134
rect 361155 505876 361475 505898
rect 446286 506454 446606 506476
rect 446286 506218 446328 506454
rect 446564 506218 446606 506454
rect 446286 506134 446606 506218
rect 446286 505898 446328 506134
rect 446564 505898 446606 506134
rect 446286 505876 446606 505898
rect 531417 506454 531737 506476
rect 531417 506218 531459 506454
rect 531695 506218 531737 506454
rect 531417 506134 531737 506218
rect 531417 505898 531459 506134
rect 531695 505898 531737 506134
rect 531417 505876 531737 505898
rect 324804 474240 325404 502800
rect 342804 488454 343404 502800
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 474240 343404 487898
rect 360804 474240 361404 502800
rect 378804 488454 379404 502800
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 474240 379404 487898
rect 396804 474240 397404 502800
rect 414804 488454 415404 502800
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 318747 473924 318813 473925
rect 318747 473860 318748 473924
rect 318812 473860 318813 473924
rect 318747 473859 318813 473860
rect 328315 473924 328381 473925
rect 328315 473860 328316 473924
rect 328380 473860 328381 473924
rect 328315 473859 328381 473860
rect 338067 473924 338133 473925
rect 338067 473860 338068 473924
rect 338132 473860 338133 473924
rect 338067 473859 338133 473860
rect 347635 473924 347701 473925
rect 347635 473860 347636 473924
rect 347700 473860 347701 473924
rect 347635 473859 347701 473860
rect 357387 473924 357453 473925
rect 357387 473860 357388 473924
rect 357452 473860 357453 473924
rect 357387 473859 357453 473860
rect 366955 473924 367021 473925
rect 366955 473860 366956 473924
rect 367020 473860 367021 473924
rect 366955 473859 367021 473860
rect 384987 473924 385053 473925
rect 384987 473860 384988 473924
rect 385052 473860 385053 473924
rect 384987 473859 385053 473860
rect 318750 473517 318810 473859
rect 328318 473653 328378 473859
rect 328315 473652 328381 473653
rect 328315 473588 328316 473652
rect 328380 473588 328381 473652
rect 328315 473587 328381 473588
rect 331078 473590 331322 473650
rect 331078 473517 331138 473590
rect 331262 473517 331322 473590
rect 338070 473517 338130 473859
rect 347638 473653 347698 473859
rect 347635 473652 347701 473653
rect 347635 473588 347636 473652
rect 347700 473588 347701 473652
rect 347635 473587 347701 473588
rect 350398 473590 350642 473650
rect 350398 473517 350458 473590
rect 350582 473517 350642 473590
rect 357390 473517 357450 473859
rect 366958 473653 367018 473859
rect 384990 473653 385050 473859
rect 366955 473652 367021 473653
rect 366955 473588 366956 473652
rect 367020 473588 367021 473652
rect 384987 473652 385053 473653
rect 366955 473587 367021 473588
rect 369718 473590 369962 473650
rect 369718 473517 369778 473590
rect 369902 473517 369962 473590
rect 384987 473588 384988 473652
rect 385052 473588 385053 473652
rect 384987 473587 385053 473588
rect 318747 473516 318813 473517
rect 318747 473452 318748 473516
rect 318812 473452 318813 473516
rect 318747 473451 318813 473452
rect 331075 473516 331141 473517
rect 331075 473452 331076 473516
rect 331140 473452 331141 473516
rect 331075 473451 331141 473452
rect 331259 473516 331325 473517
rect 331259 473452 331260 473516
rect 331324 473452 331325 473516
rect 331259 473451 331325 473452
rect 338067 473516 338133 473517
rect 338067 473452 338068 473516
rect 338132 473452 338133 473516
rect 338067 473451 338133 473452
rect 350395 473516 350461 473517
rect 350395 473452 350396 473516
rect 350460 473452 350461 473516
rect 350395 473451 350461 473452
rect 350579 473516 350645 473517
rect 350579 473452 350580 473516
rect 350644 473452 350645 473516
rect 350579 473451 350645 473452
rect 357387 473516 357453 473517
rect 357387 473452 357388 473516
rect 357452 473452 357453 473516
rect 357387 473451 357453 473452
rect 369715 473516 369781 473517
rect 369715 473452 369716 473516
rect 369780 473452 369781 473516
rect 369715 473451 369781 473452
rect 369899 473516 369965 473517
rect 369899 473452 369900 473516
rect 369964 473452 369965 473516
rect 369899 473451 369965 473452
rect 414804 452454 415404 487898
rect 425099 473652 425165 473653
rect 425099 473588 425100 473652
rect 425164 473588 425165 473652
rect 425099 473587 425165 473588
rect 425102 473381 425162 473587
rect 425099 473380 425165 473381
rect 425099 473316 425100 473380
rect 425164 473316 425165 473380
rect 425099 473315 425165 473316
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 317275 428500 317341 428501
rect 317275 428436 317276 428500
rect 317340 428436 317341 428500
rect 317275 428435 317341 428436
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 288804 290454 289404 325898
rect 293189 326454 293509 326476
rect 293189 326218 293231 326454
rect 293467 326218 293509 326454
rect 293189 326134 293509 326218
rect 293189 325898 293231 326134
rect 293467 325898 293509 326134
rect 293189 325876 293509 325898
rect 294635 308454 294955 308476
rect 294635 308218 294677 308454
rect 294913 308218 294955 308454
rect 294635 308134 294955 308218
rect 294635 307898 294677 308134
rect 294913 307898 294955 308134
rect 294635 307876 294955 307898
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 280107 235244 280173 235245
rect 280107 235180 280108 235244
rect 280172 235180 280173 235244
rect 280107 235179 280173 235180
rect 234804 221680 235404 234000
rect 252804 221680 253404 234000
rect 270804 221680 271404 234000
rect 288804 221680 289404 253898
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 221680 307404 235898
rect 324804 398454 325404 430128
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 342804 416454 343404 430128
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 380454 343404 415898
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 332915 302836 332981 302837
rect 332915 302772 332916 302836
rect 332980 302772 332981 302836
rect 332915 302771 332981 302772
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 221680 325404 253898
rect 234804 164454 235404 175440
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 219939 158812 220005 158813
rect 219939 158748 219940 158812
rect 220004 158748 220005 158812
rect 219939 158747 220005 158748
rect 234804 149680 235404 163898
rect 252804 149680 253404 175440
rect 270804 164454 271404 175440
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 149680 271404 163898
rect 288804 149680 289404 175440
rect 306804 164454 307404 175440
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 149680 307404 163898
rect 324804 149680 325404 175440
rect 332918 173909 332978 302771
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 332915 173908 332981 173909
rect 332915 173844 332916 173908
rect 332980 173844 332981 173908
rect 332915 173843 332981 173844
rect 342804 164454 343404 199898
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 139168 128454 139488 128476
rect 139168 128218 139210 128454
rect 139446 128218 139488 128454
rect 139168 128134 139488 128218
rect 139168 127898 139210 128134
rect 139446 127898 139488 128134
rect 139168 127876 139488 127898
rect 169888 128454 170208 128476
rect 169888 128218 169930 128454
rect 170166 128218 170208 128454
rect 169888 128134 170208 128218
rect 169888 127898 169930 128134
rect 170166 127898 170208 128134
rect 169888 127876 170208 127898
rect 200608 128454 200928 128476
rect 200608 128218 200650 128454
rect 200886 128218 200928 128454
rect 200608 128134 200928 128218
rect 200608 127898 200650 128134
rect 200886 127898 200928 128134
rect 200608 127876 200928 127898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 59488 92454 59808 92476
rect 59488 92218 59530 92454
rect 59766 92218 59808 92454
rect 59488 92134 59808 92218
rect 59488 91898 59530 92134
rect 59766 91898 59808 92134
rect 59488 91876 59808 91898
rect 90208 92454 90528 92476
rect 90208 92218 90250 92454
rect 90486 92218 90528 92454
rect 90208 92134 90528 92218
rect 90208 91898 90250 92134
rect 90486 91898 90528 92134
rect 90208 91876 90528 91898
rect 44128 74454 44448 74476
rect 44128 74218 44170 74454
rect 44406 74218 44448 74454
rect 44128 74134 44448 74218
rect 44128 73898 44170 74134
rect 44406 73898 44448 74134
rect 44128 73876 44448 73898
rect 74848 74454 75168 74476
rect 74848 74218 74890 74454
rect 75126 74218 75168 74454
rect 74848 74134 75168 74218
rect 74848 73898 74890 74134
rect 75126 73898 75168 74134
rect 74848 73876 75168 73898
rect 108804 74454 109404 109898
rect 123808 110454 124128 110476
rect 123808 110218 123850 110454
rect 124086 110218 124128 110454
rect 123808 110134 124128 110218
rect 123808 109898 123850 110134
rect 124086 109898 124128 110134
rect 123808 109876 124128 109898
rect 154528 110454 154848 110476
rect 154528 110218 154570 110454
rect 154806 110218 154848 110454
rect 154528 110134 154848 110218
rect 154528 109898 154570 110134
rect 154806 109898 154848 110134
rect 154528 109876 154848 109898
rect 185248 110454 185568 110476
rect 185248 110218 185290 110454
rect 185526 110218 185568 110454
rect 185248 110134 185568 110218
rect 185248 109898 185290 110134
rect 185526 109898 185568 110134
rect 185248 109876 185568 109898
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 139168 92454 139488 92476
rect 139168 92218 139210 92454
rect 139446 92218 139488 92454
rect 139168 92134 139488 92218
rect 139168 91898 139210 92134
rect 139446 91898 139488 92134
rect 139168 91876 139488 91898
rect 169888 92454 170208 92476
rect 169888 92218 169930 92454
rect 170166 92218 170208 92454
rect 169888 92134 170208 92218
rect 169888 91898 169930 92134
rect 170166 91898 170208 92134
rect 169888 91876 170208 91898
rect 200608 92454 200928 92476
rect 200608 92218 200650 92454
rect 200886 92218 200928 92454
rect 200608 92134 200928 92218
rect 200608 91898 200650 92134
rect 200886 91898 200928 92134
rect 200608 91876 200928 91898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 59488 56454 59808 56476
rect 59488 56218 59530 56454
rect 59766 56218 59808 56454
rect 59488 56134 59808 56218
rect 59488 55898 59530 56134
rect 59766 55898 59808 56134
rect 59488 55876 59808 55898
rect 90208 56454 90528 56476
rect 90208 56218 90250 56454
rect 90486 56218 90528 56454
rect 90208 56134 90528 56218
rect 90208 55898 90250 56134
rect 90486 55898 90528 56134
rect 90208 55876 90528 55898
rect 44128 38454 44448 38476
rect 44128 38218 44170 38454
rect 44406 38218 44448 38454
rect 44128 38134 44448 38218
rect 44128 37898 44170 38134
rect 44406 37898 44448 38134
rect 44128 37876 44448 37898
rect 74848 38454 75168 38476
rect 74848 38218 74890 38454
rect 75126 38218 75168 38454
rect 74848 38134 75168 38218
rect 74848 37898 74890 38134
rect 75126 37898 75168 38134
rect 74848 37876 75168 37898
rect 108804 38454 109404 73898
rect 123808 74454 124128 74476
rect 123808 74218 123850 74454
rect 124086 74218 124128 74454
rect 123808 74134 124128 74218
rect 123808 73898 123850 74134
rect 124086 73898 124128 74134
rect 123808 73876 124128 73898
rect 154528 74454 154848 74476
rect 154528 74218 154570 74454
rect 154806 74218 154848 74454
rect 154528 74134 154848 74218
rect 154528 73898 154570 74134
rect 154806 73898 154848 74134
rect 154528 73876 154848 73898
rect 185248 74454 185568 74476
rect 185248 74218 185290 74454
rect 185526 74218 185568 74454
rect 185248 74134 185568 74218
rect 185248 73898 185290 74134
rect 185526 73898 185568 74134
rect 185248 73876 185568 73898
rect 216804 74454 217404 109898
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 234804 92454 235404 103440
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 81488 235404 91898
rect 252804 81488 253404 103440
rect 270804 92454 271404 103440
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 81488 271404 91898
rect 288804 81488 289404 103440
rect 306804 92454 307404 103440
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 81488 307404 91898
rect 324804 81488 325404 103440
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 139168 56454 139488 56476
rect 139168 56218 139210 56454
rect 139446 56218 139488 56454
rect 139168 56134 139488 56218
rect 139168 55898 139210 56134
rect 139446 55898 139488 56134
rect 139168 55876 139488 55898
rect 169888 56454 170208 56476
rect 169888 56218 169930 56454
rect 170166 56218 170208 56454
rect 169888 56134 170208 56218
rect 169888 55898 169930 56134
rect 170166 55898 170208 56134
rect 169888 55876 170208 55898
rect 200608 56454 200928 56476
rect 200608 56218 200650 56454
rect 200886 56218 200928 56454
rect 200608 56134 200928 56218
rect 200608 55898 200650 56134
rect 200886 55898 200928 56134
rect 200608 55876 200928 55898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 32259 30292 32325 30293
rect 32259 30228 32260 30292
rect 32324 30228 32325 30292
rect 32259 30227 32325 30228
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 36804 2454 37404 31440
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 54804 20454 55404 31440
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 72804 2454 73404 31440
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 90804 20454 91404 31440
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 108804 2454 109404 37898
rect 123808 38454 124128 38476
rect 123808 38218 123850 38454
rect 124086 38218 124128 38454
rect 123808 38134 124128 38218
rect 123808 37898 123850 38134
rect 124086 37898 124128 38134
rect 123808 37876 124128 37898
rect 154528 38454 154848 38476
rect 154528 38218 154570 38454
rect 154806 38218 154848 38454
rect 154528 38134 154848 38218
rect 154528 37898 154570 38134
rect 154806 37898 154848 38134
rect 154528 37876 154848 37898
rect 185248 38454 185568 38476
rect 185248 38218 185290 38454
rect 185526 38218 185568 38454
rect 185248 38134 185568 38218
rect 185248 37898 185290 38134
rect 185526 37898 185568 38134
rect 185248 37876 185568 37898
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 126804 20454 127404 31440
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 144804 2454 145404 31440
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 162804 20454 163404 31440
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 180804 2454 181404 31440
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 198804 20454 199404 31440
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 216804 2454 217404 37898
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 234804 20454 235404 31440
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 252804 2454 253404 31440
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 270804 20454 271404 31440
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 288804 2454 289404 31440
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 306804 20454 307404 31440
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 324804 2454 325404 31440
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 360804 398454 361404 430128
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 362454 361404 397898
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 182454 361404 217898
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 378804 416454 379404 430128
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 380454 379404 415898
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 396804 398454 397404 430128
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 362454 397404 397898
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 60928 415404 91898
rect 432804 470454 433404 502800
rect 450804 488454 451404 502800
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 434667 473788 434733 473789
rect 434667 473724 434668 473788
rect 434732 473724 434733 473788
rect 434667 473723 434733 473724
rect 434670 473381 434730 473723
rect 450804 473680 451404 487898
rect 468804 473680 469404 502800
rect 486804 488454 487404 502800
rect 491891 500852 491957 500853
rect 491891 500788 491892 500852
rect 491956 500788 491957 500852
rect 491891 500787 491957 500788
rect 493179 500852 493245 500853
rect 493179 500788 493180 500852
rect 493244 500788 493245 500852
rect 493179 500787 493245 500788
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 473680 487404 487898
rect 491894 473517 491954 500787
rect 493182 473517 493242 500787
rect 504804 473680 505404 502800
rect 508451 500852 508517 500853
rect 508451 500788 508452 500852
rect 508516 500788 508517 500852
rect 508451 500787 508517 500788
rect 518019 500852 518085 500853
rect 518019 500788 518020 500852
rect 518084 500788 518085 500852
rect 518019 500787 518085 500788
rect 508454 476101 508514 500787
rect 508451 476100 508517 476101
rect 508451 476036 508452 476100
rect 508516 476036 508517 476100
rect 508451 476035 508517 476036
rect 518022 473925 518082 500787
rect 522804 488454 523404 502800
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 518019 473924 518085 473925
rect 518019 473860 518020 473924
rect 518084 473860 518085 473924
rect 518019 473859 518085 473860
rect 517467 473788 517533 473789
rect 517467 473724 517468 473788
rect 517532 473724 517533 473788
rect 517467 473723 517533 473724
rect 517470 473517 517530 473723
rect 522804 473680 523404 487898
rect 536787 473788 536853 473789
rect 536787 473724 536788 473788
rect 536852 473724 536853 473788
rect 536787 473723 536853 473724
rect 536790 473650 536850 473723
rect 540804 473680 541404 502800
rect 542859 500852 542925 500853
rect 542859 500788 542860 500852
rect 542924 500788 542925 500852
rect 542859 500787 542925 500788
rect 550219 500852 550285 500853
rect 550219 500788 550220 500852
rect 550284 500788 550285 500852
rect 550219 500787 550285 500788
rect 542862 476237 542922 500787
rect 542859 476236 542925 476237
rect 542859 476172 542860 476236
rect 542924 476172 542925 476236
rect 542859 476171 542925 476172
rect 550222 474061 550282 500787
rect 558804 488454 559404 502800
rect 574878 502757 574938 527715
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 574875 502756 574941 502757
rect 574875 502692 574876 502756
rect 574940 502692 574941 502756
rect 574875 502691 574941 502692
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 550587 487796 550653 487797
rect 550587 487732 550588 487796
rect 550652 487732 550653 487796
rect 550587 487731 550653 487732
rect 550590 474605 550650 487731
rect 552243 477188 552309 477189
rect 552243 477124 552244 477188
rect 552308 477124 552309 477188
rect 552243 477123 552309 477124
rect 551139 476100 551205 476101
rect 551139 476036 551140 476100
rect 551204 476036 551205 476100
rect 551139 476035 551205 476036
rect 550587 474604 550653 474605
rect 550587 474540 550588 474604
rect 550652 474540 550653 474604
rect 550587 474539 550653 474540
rect 550219 474060 550285 474061
rect 550219 473996 550220 474060
rect 550284 473996 550285 474060
rect 550219 473995 550285 473996
rect 536971 473652 537037 473653
rect 536971 473650 536972 473652
rect 536790 473590 536972 473650
rect 536971 473588 536972 473590
rect 537036 473588 537037 473652
rect 536971 473587 537037 473588
rect 491891 473516 491957 473517
rect 491891 473452 491892 473516
rect 491956 473452 491957 473516
rect 491891 473451 491957 473452
rect 493179 473516 493245 473517
rect 493179 473452 493180 473516
rect 493244 473452 493245 473516
rect 493179 473451 493245 473452
rect 517467 473516 517533 473517
rect 517467 473452 517468 473516
rect 517532 473452 517533 473516
rect 517467 473451 517533 473452
rect 434667 473380 434733 473381
rect 434667 473316 434668 473380
rect 434732 473316 434733 473380
rect 434667 473315 434733 473316
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 551142 463450 551202 476035
rect 551691 475964 551757 475965
rect 551691 475900 551692 475964
rect 551756 475900 551757 475964
rect 551691 475899 551757 475900
rect 551694 464810 551754 475899
rect 552059 475420 552125 475421
rect 552059 475356 552060 475420
rect 552124 475356 552125 475420
rect 552059 475355 552125 475356
rect 552062 471341 552122 475355
rect 552059 471340 552125 471341
rect 552059 471276 552060 471340
rect 552124 471276 552125 471340
rect 552059 471275 552125 471276
rect 552246 465357 552306 477123
rect 552795 477052 552861 477053
rect 552795 476988 552796 477052
rect 552860 476988 552861 477052
rect 552795 476987 552861 476988
rect 552611 476916 552677 476917
rect 552611 476852 552612 476916
rect 552676 476852 552677 476916
rect 552611 476851 552677 476852
rect 552427 476780 552493 476781
rect 552427 476716 552428 476780
rect 552492 476716 552493 476780
rect 552427 476715 552493 476716
rect 552430 469029 552490 476715
rect 552427 469028 552493 469029
rect 552427 468964 552428 469028
rect 552492 468964 552493 469028
rect 552427 468963 552493 468964
rect 552614 467805 552674 476851
rect 552611 467804 552677 467805
rect 552611 467740 552612 467804
rect 552676 467740 552677 467804
rect 552611 467739 552677 467740
rect 552798 466309 552858 476987
rect 555003 475828 555069 475829
rect 555003 475764 555004 475828
rect 555068 475764 555069 475828
rect 555003 475763 555069 475764
rect 553347 475692 553413 475693
rect 553347 475628 553348 475692
rect 553412 475628 553413 475692
rect 553347 475627 553413 475628
rect 553350 468077 553410 475627
rect 553531 474332 553597 474333
rect 553531 474268 553532 474332
rect 553596 474268 553597 474332
rect 553531 474267 553597 474268
rect 553347 468076 553413 468077
rect 553347 468012 553348 468076
rect 553412 468012 553413 468076
rect 553347 468011 553413 468012
rect 552795 466308 552861 466309
rect 552795 466244 552796 466308
rect 552860 466244 552861 466308
rect 552795 466243 552861 466244
rect 552243 465356 552309 465357
rect 552243 465292 552244 465356
rect 552308 465292 552309 465356
rect 552243 465291 552309 465292
rect 552059 464812 552125 464813
rect 552059 464810 552060 464812
rect 551694 464750 552060 464810
rect 552059 464748 552060 464750
rect 552124 464748 552125 464812
rect 552059 464747 552125 464748
rect 552059 463588 552125 463589
rect 552059 463524 552060 463588
rect 552124 463524 552125 463588
rect 552059 463523 552125 463524
rect 552062 463450 552122 463523
rect 551142 463390 552122 463450
rect 553534 457333 553594 474267
rect 553715 474196 553781 474197
rect 553715 474132 553716 474196
rect 553780 474132 553781 474196
rect 553715 474131 553781 474132
rect 553718 461549 553778 474131
rect 554083 474060 554149 474061
rect 554083 473996 554084 474060
rect 554148 473996 554149 474060
rect 554083 473995 554149 473996
rect 553715 461548 553781 461549
rect 553715 461484 553716 461548
rect 553780 461484 553781 461548
rect 553715 461483 553781 461484
rect 553531 457332 553597 457333
rect 553531 457268 553532 457332
rect 553596 457268 553597 457332
rect 553531 457267 553597 457268
rect 554086 440741 554146 473995
rect 554819 472700 554885 472701
rect 554819 472636 554820 472700
rect 554884 472636 554885 472700
rect 554819 472635 554885 472636
rect 554822 463861 554882 472635
rect 555006 466853 555066 475763
rect 555371 473924 555437 473925
rect 555371 473860 555372 473924
rect 555436 473860 555437 473924
rect 555371 473859 555437 473860
rect 555003 466852 555069 466853
rect 555003 466788 555004 466852
rect 555068 466788 555069 466852
rect 555003 466787 555069 466788
rect 555374 465629 555434 473859
rect 555371 465628 555437 465629
rect 555371 465564 555372 465628
rect 555436 465564 555437 465628
rect 555371 465563 555437 465564
rect 554819 463860 554885 463861
rect 554819 463796 554820 463860
rect 554884 463796 554885 463860
rect 554819 463795 554885 463796
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 554083 440740 554149 440741
rect 554083 440676 554084 440740
rect 554148 440676 554149 440740
rect 554083 440675 554149 440676
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 60928 433404 73898
rect 450804 416454 451404 427440
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 60928 451404 91898
rect 468804 398454 469404 427440
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 60928 469404 73898
rect 486804 416454 487404 427440
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 60928 487404 91898
rect 504804 398454 505404 427440
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 60928 505404 73898
rect 522804 416454 523404 427440
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 60928 523404 91898
rect 540804 398454 541404 427440
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 60928 541404 73898
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 60928 559404 91898
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 433568 56454 433888 56476
rect 433568 56218 433610 56454
rect 433846 56218 433888 56454
rect 433568 56134 433888 56218
rect 433568 55898 433610 56134
rect 433846 55898 433888 56134
rect 433568 55876 433888 55898
rect 464288 56454 464608 56476
rect 464288 56218 464330 56454
rect 464566 56218 464608 56454
rect 464288 56134 464608 56218
rect 464288 55898 464330 56134
rect 464566 55898 464608 56134
rect 464288 55876 464608 55898
rect 495008 56454 495328 56476
rect 495008 56218 495050 56454
rect 495286 56218 495328 56454
rect 495008 56134 495328 56218
rect 495008 55898 495050 56134
rect 495286 55898 495328 56134
rect 495008 55876 495328 55898
rect 525728 56454 526048 56476
rect 525728 56218 525770 56454
rect 526006 56218 526048 56454
rect 525728 56134 526048 56218
rect 525728 55898 525770 56134
rect 526006 55898 526048 56134
rect 525728 55876 526048 55898
rect 556448 56454 556768 56476
rect 556448 56218 556490 56454
rect 556726 56218 556768 56454
rect 556448 56134 556768 56218
rect 556448 55898 556490 56134
rect 556726 55898 556768 56134
rect 556448 55876 556768 55898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 418208 38454 418528 38476
rect 418208 38218 418250 38454
rect 418486 38218 418528 38454
rect 418208 38134 418528 38218
rect 418208 37898 418250 38134
rect 418486 37898 418528 38134
rect 418208 37876 418528 37898
rect 448928 38454 449248 38476
rect 448928 38218 448970 38454
rect 449206 38218 449248 38454
rect 448928 38134 449248 38218
rect 448928 37898 448970 38134
rect 449206 37898 449248 38134
rect 448928 37876 449248 37898
rect 479648 38454 479968 38476
rect 479648 38218 479690 38454
rect 479926 38218 479968 38454
rect 479648 38134 479968 38218
rect 479648 37898 479690 38134
rect 479926 37898 479968 38134
rect 479648 37876 479968 37898
rect 510368 38454 510688 38476
rect 510368 38218 510410 38454
rect 510646 38218 510688 38454
rect 510368 38134 510688 38218
rect 510368 37898 510410 38134
rect 510646 37898 510688 38134
rect 510368 37876 510688 37898
rect 541088 38454 541408 38476
rect 541088 38218 541130 38454
rect 541366 38218 541408 38454
rect 541088 38134 541408 38218
rect 541088 37898 541130 38134
rect 541366 37898 541408 38134
rect 541088 37876 541408 37898
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 433568 20454 433888 20476
rect 433568 20218 433610 20454
rect 433846 20218 433888 20454
rect 433568 20134 433888 20218
rect 433568 19898 433610 20134
rect 433846 19898 433888 20134
rect 433568 19876 433888 19898
rect 464288 20454 464608 20476
rect 464288 20218 464330 20454
rect 464566 20218 464608 20454
rect 464288 20134 464608 20218
rect 464288 19898 464330 20134
rect 464566 19898 464608 20134
rect 464288 19876 464608 19898
rect 495008 20454 495328 20476
rect 495008 20218 495050 20454
rect 495286 20218 495328 20454
rect 495008 20134 495328 20218
rect 495008 19898 495050 20134
rect 495286 19898 495328 20134
rect 495008 19876 495328 19898
rect 525728 20454 526048 20476
rect 525728 20218 525770 20454
rect 526006 20218 526048 20454
rect 525728 20134 526048 20218
rect 525728 19898 525770 20134
rect 526006 19898 526048 20134
rect 525728 19876 526048 19898
rect 556448 20454 556768 20476
rect 556448 20218 556490 20454
rect 556726 20218 556768 20454
rect 556448 20134 556768 20218
rect 556448 19898 556490 20134
rect 556726 19898 556768 20134
rect 556448 19876 556768 19898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 414804 -1286 415404 16320
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 432804 2454 433404 16320
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 450804 -1286 451404 16320
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 468804 2454 469404 16320
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 486804 -1286 487404 16320
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 504804 2454 505404 16320
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 522804 -1286 523404 16320
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 540804 2454 541404 16320
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 558804 -1286 559404 16320
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 587200 -2226 587800 706162
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 588140 -3166 588740 707102
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 589080 -4106 589680 708042
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 590020 -5046 590620 708982
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 590960 -5986 591560 709922
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 591900 -6926 592500 710862
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 13450 182218 13686 182454
rect 13450 181898 13686 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 13450 146218 13686 146454
rect 13450 145898 13686 146134
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 24814 571422 25050 571658
rect 26286 572782 26522 573018
rect 30334 572102 30570 572338
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 30886 531302 31122 531538
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 95102 571422 95338 571658
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 104854 531316 105090 531538
rect 104854 531302 104940 531316
rect 104940 531302 105004 531316
rect 105004 531302 105090 531316
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 107717 524218 107953 524454
rect 107717 523898 107953 524134
rect 192847 524218 193083 524454
rect 192847 523898 193083 524134
rect 65151 506218 65387 506454
rect 65151 505898 65387 506134
rect 150282 506218 150518 506454
rect 150282 505898 150518 506134
rect 235412 506218 235648 506454
rect 235412 505898 235648 506134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 112766 500172 113002 500258
rect 112766 500108 112852 500172
rect 112852 500108 112916 500172
rect 112916 500108 113002 500172
rect 112766 500022 113002 500108
rect 130614 497982 130850 498218
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 147358 500022 147594 500258
rect 23726 470218 23962 470454
rect 23726 469898 23962 470134
rect 54446 470218 54682 470454
rect 54446 469898 54682 470134
rect 85166 470218 85402 470454
rect 85166 469898 85402 470134
rect 115886 470218 116122 470454
rect 115886 469898 116122 470134
rect 146606 470218 146842 470454
rect 146606 469898 146842 470134
rect 39086 452218 39322 452454
rect 39086 451898 39322 452134
rect 69806 452218 70042 452454
rect 69806 451898 70042 452134
rect 100526 452218 100762 452454
rect 100526 451898 100762 452134
rect 131246 452218 131482 452454
rect 131246 451898 131482 452134
rect 23726 434218 23962 434454
rect 23726 433898 23962 434134
rect 54446 434218 54682 434454
rect 54446 433898 54682 434134
rect 85166 434218 85402 434454
rect 85166 433898 85402 434134
rect 115886 434218 116122 434454
rect 115886 433898 116122 434134
rect 146606 434218 146842 434454
rect 146606 433898 146842 434134
rect 39086 416218 39322 416454
rect 39086 415898 39322 416134
rect 69806 416218 70042 416454
rect 69806 415898 70042 416134
rect 100526 416218 100762 416454
rect 100526 415898 100762 416134
rect 131246 416218 131482 416454
rect 131246 415898 131482 416134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 38917 380218 39153 380454
rect 38917 379898 39153 380134
rect 56847 380218 57083 380454
rect 56847 379898 57083 380134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 29951 362218 30187 362454
rect 29951 361898 30187 362134
rect 47882 362218 48118 362454
rect 47882 361898 48118 362134
rect 65812 362218 66048 362454
rect 65812 361898 66048 362134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 153246 497982 153482 498218
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 155822 421292 156058 421378
rect 155822 421228 155908 421292
rect 155908 421228 155972 421292
rect 155972 421228 156058 421292
rect 155822 421142 156058 421228
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 207656 488218 207892 488454
rect 207656 487898 207892 488134
rect 238376 488218 238612 488454
rect 238376 487898 238612 488134
rect 269096 488218 269332 488454
rect 269096 487898 269332 488134
rect 192296 470218 192532 470454
rect 192296 469898 192532 470134
rect 223016 470218 223252 470454
rect 223016 469898 223252 470134
rect 253736 470218 253972 470454
rect 253736 469898 253972 470134
rect 207656 452218 207892 452454
rect 207656 451898 207892 452134
rect 238376 452218 238612 452454
rect 238376 451898 238612 452134
rect 269096 452218 269332 452454
rect 269096 451898 269332 452134
rect 192296 434218 192532 434454
rect 192296 433898 192532 434134
rect 223016 434218 223252 434454
rect 223016 433898 223252 434134
rect 253736 434218 253972 434454
rect 253736 433898 253972 434134
rect 207656 416218 207892 416454
rect 207656 415898 207892 416134
rect 238376 416218 238612 416454
rect 238376 415898 238612 416134
rect 269096 416218 269332 416454
rect 269096 415898 269332 416134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 107717 344218 107953 344454
rect 107717 343898 107953 344134
rect 192847 344218 193083 344454
rect 192847 343898 193083 344134
rect 65151 326218 65387 326454
rect 65151 325898 65387 326134
rect 150282 326218 150518 326454
rect 150282 325898 150518 326134
rect 235412 326218 235648 326454
rect 235412 325898 235648 326134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 39656 308218 39892 308454
rect 39656 307898 39892 308134
rect 70376 308218 70612 308454
rect 70376 307898 70612 308134
rect 101096 308218 101332 308454
rect 101096 307898 101332 308134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 24296 290218 24532 290454
rect 24296 289898 24532 290134
rect 55016 290218 55252 290454
rect 55016 289898 55252 290134
rect 85736 290218 85972 290454
rect 85736 289898 85972 290134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 39656 272218 39892 272454
rect 39656 271898 39892 272134
rect 70376 272218 70612 272454
rect 70376 271898 70612 272134
rect 101096 272218 101332 272454
rect 101096 271898 101332 272134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 24296 254218 24532 254454
rect 24296 253898 24532 254134
rect 55016 254218 55252 254454
rect 55016 253898 55252 254134
rect 85736 254218 85972 254454
rect 85736 253898 85972 254134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 192250 290218 192486 290454
rect 192250 289898 192486 290134
rect 192250 254218 192486 254454
rect 192250 253898 192486 254134
rect 207610 308218 207846 308454
rect 207610 307898 207846 308134
rect 207610 272218 207846 272454
rect 207610 271898 207846 272134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 28810 200218 29046 200454
rect 28810 199898 29046 200134
rect 59530 200218 59766 200454
rect 59530 199898 59766 200134
rect 90250 200218 90486 200454
rect 90250 199898 90486 200134
rect 44170 182218 44406 182454
rect 44170 181898 44406 182134
rect 74890 182218 75126 182454
rect 74890 181898 75126 182134
rect 123850 218218 124086 218454
rect 123850 217898 124086 218134
rect 154570 218218 154806 218454
rect 154570 217898 154806 218134
rect 185290 218218 185526 218454
rect 185290 217898 185526 218134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 139210 200218 139446 200454
rect 139210 199898 139446 200134
rect 169930 200218 170166 200454
rect 169930 199898 170166 200134
rect 200650 200218 200886 200454
rect 200650 199898 200886 200134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 28810 164218 29046 164454
rect 28810 163898 29046 164134
rect 59530 164218 59766 164454
rect 59530 163898 59766 164134
rect 90250 164218 90486 164454
rect 90250 163898 90486 164134
rect 44170 146218 44406 146454
rect 44170 145898 44406 146134
rect 74890 146218 75126 146454
rect 74890 145898 75126 146134
rect 123850 182218 124086 182454
rect 123850 181898 124086 182134
rect 154570 182218 154806 182454
rect 154570 181898 154806 182134
rect 185290 182218 185526 182454
rect 185290 181898 185526 182134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 139210 164218 139446 164454
rect 139210 163898 139446 164134
rect 169930 164218 170166 164454
rect 169930 163898 170166 164134
rect 200650 164218 200886 164454
rect 200650 163898 200886 164134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 28810 92218 29046 92454
rect 28810 91898 29046 92134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 13450 74218 13686 74454
rect 13450 73898 13686 74134
rect 28810 56218 29046 56454
rect 28810 55898 29046 56134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 13450 38218 13686 38454
rect 13450 37898 13686 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 123850 146218 124086 146454
rect 123850 145898 124086 146134
rect 154570 146218 154806 146454
rect 154570 145898 154806 146134
rect 185290 146218 185526 146454
rect 185290 145898 185526 146134
rect 238330 308218 238566 308454
rect 238330 307898 238566 308134
rect 269050 308218 269286 308454
rect 269050 307898 269286 308134
rect 222970 290218 223206 290454
rect 222970 289898 223206 290134
rect 253690 290218 253926 290454
rect 253690 289898 253926 290134
rect 238330 272218 238566 272454
rect 238330 271898 238566 272134
rect 269050 272218 269286 272454
rect 269050 271898 269286 272134
rect 222970 254218 223206 254454
rect 222970 253898 223206 254134
rect 253690 254218 253926 254454
rect 253690 253898 253926 254134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 281494 421292 281730 421378
rect 281494 421228 281580 421292
rect 281580 421228 281644 421292
rect 281644 421228 281730 421292
rect 281494 421142 281730 421228
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 323772 650218 324008 650454
rect 323772 649898 324008 650134
rect 354492 650218 354728 650454
rect 354492 649898 354728 650134
rect 385212 650218 385448 650454
rect 385212 649898 385448 650134
rect 415932 650218 416168 650454
rect 415932 649898 416168 650134
rect 446652 650218 446888 650454
rect 446652 649898 446888 650134
rect 464250 650218 464486 650454
rect 464250 649898 464486 650134
rect 339132 632218 339368 632454
rect 339132 631898 339368 632134
rect 369852 632218 370088 632454
rect 369852 631898 370088 632134
rect 400572 632218 400808 632454
rect 400572 631898 400808 632134
rect 431292 632218 431528 632454
rect 431292 631898 431528 632134
rect 479610 632218 479846 632454
rect 479610 631898 479846 632134
rect 323772 614218 324008 614454
rect 323772 613898 324008 614134
rect 354492 614218 354728 614454
rect 354492 613898 354728 614134
rect 385212 614218 385448 614454
rect 385212 613898 385448 614134
rect 415932 614218 416168 614454
rect 415932 613898 416168 614134
rect 446652 614218 446888 614454
rect 446652 613898 446888 614134
rect 464250 614218 464486 614454
rect 464250 613898 464486 614134
rect 339132 596218 339368 596454
rect 339132 595898 339368 596134
rect 369852 596218 370088 596454
rect 369852 595898 370088 596134
rect 400572 596218 400808 596454
rect 400572 595898 400808 596134
rect 431292 596218 431528 596454
rect 431292 595898 431528 596134
rect 479610 596218 479846 596454
rect 479610 595898 479846 596134
rect 323772 578218 324008 578454
rect 323772 577898 324008 578134
rect 354492 578218 354728 578454
rect 354492 577898 354728 578134
rect 385212 578218 385448 578454
rect 385212 577898 385448 578134
rect 415932 578218 416168 578454
rect 415932 577898 416168 578134
rect 446652 578218 446888 578454
rect 446652 577898 446888 578134
rect 464250 578218 464486 578454
rect 464250 577898 464486 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 493462 531302 493698 531538
rect 494970 650218 495206 650454
rect 494970 649898 495206 650134
rect 525690 650218 525926 650454
rect 525690 649898 525926 650134
rect 510330 632218 510566 632454
rect 510330 631898 510566 632134
rect 541050 632218 541286 632454
rect 541050 631898 541286 632134
rect 494970 614218 495206 614454
rect 494970 613898 495206 614134
rect 525690 614218 525926 614454
rect 525690 613898 525926 614134
rect 510330 596218 510566 596454
rect 510330 595898 510566 596134
rect 541050 596218 541286 596454
rect 541050 595898 541286 596134
rect 549398 588422 549634 588658
rect 494970 578218 495206 578454
rect 494970 577898 495206 578134
rect 525690 578218 525926 578454
rect 525690 577898 525926 578134
rect 551238 588572 551474 588658
rect 551238 588508 551324 588572
rect 551324 588508 551388 588572
rect 551388 588508 551474 588572
rect 551238 588422 551474 588508
rect 549766 574142 550002 574378
rect 549766 572782 550002 573018
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 549766 531302 550002 531538
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 403763 524218 403999 524454
rect 403763 523898 403999 524134
rect 488893 524218 489129 524454
rect 488893 523898 489129 524134
rect 361197 506218 361433 506454
rect 361197 505898 361433 506134
rect 446328 506218 446564 506454
rect 446328 505898 446564 506134
rect 531459 506218 531695 506454
rect 531459 505898 531695 506134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 293231 326218 293467 326454
rect 293231 325898 293467 326134
rect 294677 308218 294913 308454
rect 294677 307898 294913 308134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 139210 128218 139446 128454
rect 139210 127898 139446 128134
rect 169930 128218 170166 128454
rect 169930 127898 170166 128134
rect 200650 128218 200886 128454
rect 200650 127898 200886 128134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 59530 92218 59766 92454
rect 59530 91898 59766 92134
rect 90250 92218 90486 92454
rect 90250 91898 90486 92134
rect 44170 74218 44406 74454
rect 44170 73898 44406 74134
rect 74890 74218 75126 74454
rect 74890 73898 75126 74134
rect 123850 110218 124086 110454
rect 123850 109898 124086 110134
rect 154570 110218 154806 110454
rect 154570 109898 154806 110134
rect 185290 110218 185526 110454
rect 185290 109898 185526 110134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 139210 92218 139446 92454
rect 139210 91898 139446 92134
rect 169930 92218 170166 92454
rect 169930 91898 170166 92134
rect 200650 92218 200886 92454
rect 200650 91898 200886 92134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 59530 56218 59766 56454
rect 59530 55898 59766 56134
rect 90250 56218 90486 56454
rect 90250 55898 90486 56134
rect 44170 38218 44406 38454
rect 44170 37898 44406 38134
rect 74890 38218 75126 38454
rect 74890 37898 75126 38134
rect 123850 74218 124086 74454
rect 123850 73898 124086 74134
rect 154570 74218 154806 74454
rect 154570 73898 154806 74134
rect 185290 74218 185526 74454
rect 185290 73898 185526 74134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 139210 56218 139446 56454
rect 139210 55898 139446 56134
rect 169930 56218 170166 56454
rect 169930 55898 170166 56134
rect 200650 56218 200886 56454
rect 200650 55898 200886 56134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 123850 38218 124086 38454
rect 123850 37898 124086 38134
rect 154570 38218 154806 38454
rect 154570 37898 154806 38134
rect 185290 38218 185526 38454
rect 185290 37898 185526 38134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 433610 56218 433846 56454
rect 433610 55898 433846 56134
rect 464330 56218 464566 56454
rect 464330 55898 464566 56134
rect 495050 56218 495286 56454
rect 495050 55898 495286 56134
rect 525770 56218 526006 56454
rect 525770 55898 526006 56134
rect 556490 56218 556726 56454
rect 556490 55898 556726 56134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 418250 38218 418486 38454
rect 418250 37898 418486 38134
rect 448970 38218 449206 38454
rect 448970 37898 449206 38134
rect 479690 38218 479926 38454
rect 479690 37898 479926 38134
rect 510410 38218 510646 38454
rect 510410 37898 510646 38134
rect 541130 38218 541366 38454
rect 541130 37898 541366 38134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 433610 20218 433846 20454
rect 433610 19898 433846 20134
rect 464330 20218 464566 20454
rect 464330 19898 464566 20134
rect 495050 20218 495286 20454
rect 495050 19898 495286 20134
rect 525770 20218 526006 20454
rect 525770 19898 526006 20134
rect 556490 20218 556726 20454
rect 556490 19898 556726 20134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 323730 650476 324050 650478
rect 354450 650476 354770 650478
rect 385170 650476 385490 650478
rect 415890 650476 416210 650478
rect 446610 650476 446930 650478
rect 464208 650476 464528 650478
rect 494928 650476 495248 650478
rect 525648 650476 525968 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 323772 650454
rect 324008 650218 354492 650454
rect 354728 650218 385212 650454
rect 385448 650218 415932 650454
rect 416168 650218 446652 650454
rect 446888 650218 464250 650454
rect 464486 650218 494970 650454
rect 495206 650218 525690 650454
rect 525926 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 323772 650134
rect 324008 649898 354492 650134
rect 354728 649898 385212 650134
rect 385448 649898 415932 650134
rect 416168 649898 446652 650134
rect 446888 649898 464250 650134
rect 464486 649898 494970 650134
rect 495206 649898 525690 650134
rect 525926 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 323730 649874 324050 649876
rect 354450 649874 354770 649876
rect 385170 649874 385490 649876
rect 415890 649874 416210 649876
rect 446610 649874 446930 649876
rect 464208 649874 464528 649876
rect 494928 649874 495248 649876
rect 525648 649874 525968 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 339090 632476 339410 632478
rect 369810 632476 370130 632478
rect 400530 632476 400850 632478
rect 431250 632476 431570 632478
rect 479568 632476 479888 632478
rect 510288 632476 510608 632478
rect 541008 632476 541328 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 339132 632454
rect 339368 632218 369852 632454
rect 370088 632218 400572 632454
rect 400808 632218 431292 632454
rect 431528 632218 479610 632454
rect 479846 632218 510330 632454
rect 510566 632218 541050 632454
rect 541286 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 339132 632134
rect 339368 631898 369852 632134
rect 370088 631898 400572 632134
rect 400808 631898 431292 632134
rect 431528 631898 479610 632134
rect 479846 631898 510330 632134
rect 510566 631898 541050 632134
rect 541286 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 339090 631874 339410 631876
rect 369810 631874 370130 631876
rect 400530 631874 400850 631876
rect 431250 631874 431570 631876
rect 479568 631874 479888 631876
rect 510288 631874 510608 631876
rect 541008 631874 541328 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 288804 614476 289404 614478
rect 323730 614476 324050 614478
rect 354450 614476 354770 614478
rect 385170 614476 385490 614478
rect 415890 614476 416210 614478
rect 446610 614476 446930 614478
rect 464208 614476 464528 614478
rect 494928 614476 495248 614478
rect 525648 614476 525968 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 288986 614454
rect 289222 614218 323772 614454
rect 324008 614218 354492 614454
rect 354728 614218 385212 614454
rect 385448 614218 415932 614454
rect 416168 614218 446652 614454
rect 446888 614218 464250 614454
rect 464486 614218 494970 614454
rect 495206 614218 525690 614454
rect 525926 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 288986 614134
rect 289222 613898 323772 614134
rect 324008 613898 354492 614134
rect 354728 613898 385212 614134
rect 385448 613898 415932 614134
rect 416168 613898 446652 614134
rect 446888 613898 464250 614134
rect 464486 613898 494970 614134
rect 495206 613898 525690 614134
rect 525926 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 288804 613874 289404 613876
rect 323730 613874 324050 613876
rect 354450 613874 354770 613876
rect 385170 613874 385490 613876
rect 415890 613874 416210 613876
rect 446610 613874 446930 613876
rect 464208 613874 464528 613876
rect 494928 613874 495248 613876
rect 525648 613874 525968 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 162804 596476 163404 596478
rect 306804 596476 307404 596478
rect 339090 596476 339410 596478
rect 369810 596476 370130 596478
rect 400530 596476 400850 596478
rect 431250 596476 431570 596478
rect 479568 596476 479888 596478
rect 510288 596476 510608 596478
rect 541008 596476 541328 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 162986 596454
rect 163222 596218 306986 596454
rect 307222 596218 339132 596454
rect 339368 596218 369852 596454
rect 370088 596218 400572 596454
rect 400808 596218 431292 596454
rect 431528 596218 479610 596454
rect 479846 596218 510330 596454
rect 510566 596218 541050 596454
rect 541286 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 162986 596134
rect 163222 595898 306986 596134
rect 307222 595898 339132 596134
rect 339368 595898 369852 596134
rect 370088 595898 400572 596134
rect 400808 595898 431292 596134
rect 431528 595898 479610 596134
rect 479846 595898 510330 596134
rect 510566 595898 541050 596134
rect 541286 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 162804 595874 163404 595876
rect 306804 595874 307404 595876
rect 339090 595874 339410 595876
rect 369810 595874 370130 595876
rect 400530 595874 400850 595876
rect 431250 595874 431570 595876
rect 479568 595874 479888 595876
rect 510288 595874 510608 595876
rect 541008 595874 541328 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect 549356 588658 551516 588700
rect 549356 588422 549398 588658
rect 549634 588422 551238 588658
rect 551474 588422 551516 588658
rect 549356 588380 551516 588422
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 288804 578476 289404 578478
rect 323730 578476 324050 578478
rect 354450 578476 354770 578478
rect 385170 578476 385490 578478
rect 415890 578476 416210 578478
rect 446610 578476 446930 578478
rect 464208 578476 464528 578478
rect 494928 578476 495248 578478
rect 525648 578476 525968 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 288986 578454
rect 289222 578218 323772 578454
rect 324008 578218 354492 578454
rect 354728 578218 385212 578454
rect 385448 578218 415932 578454
rect 416168 578218 446652 578454
rect 446888 578218 464250 578454
rect 464486 578218 494970 578454
rect 495206 578218 525690 578454
rect 525926 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 288986 578134
rect 289222 577898 323772 578134
rect 324008 577898 354492 578134
rect 354728 577898 385212 578134
rect 385448 577898 415932 578134
rect 416168 577898 446652 578134
rect 446888 577898 464250 578134
rect 464486 577898 494970 578134
rect 495206 577898 525690 578134
rect 525926 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 288804 577874 289404 577876
rect 323730 577874 324050 577876
rect 354450 577874 354770 577876
rect 385170 577874 385490 577876
rect 415890 577874 416210 577876
rect 446610 577874 446930 577876
rect 464208 577874 464528 577876
rect 494928 577874 495248 577876
rect 525648 577874 525968 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect 549724 574378 550044 574420
rect 549724 574142 549766 574378
rect 550002 574142 550044 574378
rect 26244 573018 29508 573060
rect 26244 572782 26286 573018
rect 26522 572782 29508 573018
rect 26244 572740 29508 572782
rect 549724 573018 550044 574142
rect 549724 572782 549766 573018
rect 550002 572782 550044 573018
rect 549724 572740 550044 572782
rect 29188 572380 29508 572740
rect 29188 572338 30612 572380
rect 29188 572102 30334 572338
rect 30570 572102 30612 572338
rect 29188 572060 30612 572102
rect 24772 571658 95380 571700
rect 24772 571422 24814 571658
rect 25050 571422 95102 571658
rect 95338 571422 95380 571658
rect 24772 571380 95380 571422
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586260 559874 586860 559876
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect 30844 531538 105132 531580
rect 30844 531302 30886 531538
rect 31122 531302 104854 531538
rect 105090 531302 105132 531538
rect 30844 531260 105132 531302
rect 493420 531538 550044 531580
rect 493420 531302 493462 531538
rect 493698 531302 549766 531538
rect 550002 531302 550044 531538
rect 493420 531260 550044 531302
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 107675 524476 107995 524478
rect 192805 524476 193125 524478
rect 306804 524476 307404 524478
rect 403721 524476 404041 524478
rect 488851 524476 489171 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 107717 524454
rect 107953 524218 192847 524454
rect 193083 524218 306986 524454
rect 307222 524218 403763 524454
rect 403999 524218 488893 524454
rect 489129 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 107717 524134
rect 107953 523898 192847 524134
rect 193083 523898 306986 524134
rect 307222 523898 403763 524134
rect 403999 523898 488893 524134
rect 489129 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 107675 523874 107995 523876
rect 192805 523874 193125 523876
rect 306804 523874 307404 523876
rect 403721 523874 404041 523876
rect 488851 523874 489171 523876
rect 586260 523874 586860 523876
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 65109 506476 65429 506478
rect 150240 506476 150560 506478
rect 235370 506476 235690 506478
rect 288804 506476 289404 506478
rect 361155 506476 361475 506478
rect 446286 506476 446606 506478
rect 531417 506476 531737 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 65151 506454
rect 65387 506218 150282 506454
rect 150518 506218 235412 506454
rect 235648 506218 288986 506454
rect 289222 506218 361197 506454
rect 361433 506218 446328 506454
rect 446564 506218 531459 506454
rect 531695 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 65151 506134
rect 65387 505898 150282 506134
rect 150518 505898 235412 506134
rect 235648 505898 288986 506134
rect 289222 505898 361197 506134
rect 361433 505898 446328 506134
rect 446564 505898 531459 506134
rect 531695 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 65109 505874 65429 505876
rect 150240 505874 150560 505876
rect 235370 505874 235690 505876
rect 288804 505874 289404 505876
rect 361155 505874 361475 505876
rect 446286 505874 446606 505876
rect 531417 505874 531737 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect 112724 500258 147636 500300
rect 112724 500022 112766 500258
rect 113002 500022 147358 500258
rect 147594 500022 147636 500258
rect 112724 499980 147636 500022
rect 130572 498218 153524 498260
rect 130572 497982 130614 498218
rect 130850 497982 153246 498218
rect 153482 497982 153524 498218
rect 130572 497940 153524 497982
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 207614 488476 207934 488478
rect 238334 488476 238654 488478
rect 269054 488476 269374 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 207656 488454
rect 207892 488218 238376 488454
rect 238612 488218 269096 488454
rect 269332 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 207656 488134
rect 207892 487898 238376 488134
rect 238612 487898 269096 488134
rect 269332 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 207614 487874 207934 487876
rect 238334 487874 238654 487876
rect 269054 487874 269374 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586260 487874 586860 487876
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 23684 470476 24004 470478
rect 54404 470476 54724 470478
rect 85124 470476 85444 470478
rect 115844 470476 116164 470478
rect 146564 470476 146884 470478
rect 180804 470476 181404 470478
rect 192254 470476 192574 470478
rect 222974 470476 223294 470478
rect 253694 470476 254014 470478
rect 288804 470476 289404 470478
rect 432804 470476 433404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 23726 470454
rect 23962 470218 54446 470454
rect 54682 470218 85166 470454
rect 85402 470218 115886 470454
rect 116122 470218 146606 470454
rect 146842 470218 180986 470454
rect 181222 470218 192296 470454
rect 192532 470218 223016 470454
rect 223252 470218 253736 470454
rect 253972 470218 288986 470454
rect 289222 470218 432986 470454
rect 433222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 23726 470134
rect 23962 469898 54446 470134
rect 54682 469898 85166 470134
rect 85402 469898 115886 470134
rect 116122 469898 146606 470134
rect 146842 469898 180986 470134
rect 181222 469898 192296 470134
rect 192532 469898 223016 470134
rect 223252 469898 253736 470134
rect 253972 469898 288986 470134
rect 289222 469898 432986 470134
rect 433222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 23684 469874 24004 469876
rect 54404 469874 54724 469876
rect 85124 469874 85444 469876
rect 115844 469874 116164 469876
rect 146564 469874 146884 469876
rect 180804 469874 181404 469876
rect 192254 469874 192574 469876
rect 222974 469874 223294 469876
rect 253694 469874 254014 469876
rect 288804 469874 289404 469876
rect 432804 469874 433404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -2936 452476 -2336 452478
rect 39044 452476 39364 452478
rect 69764 452476 70084 452478
rect 100484 452476 100804 452478
rect 131204 452476 131524 452478
rect 162804 452476 163404 452478
rect 207614 452476 207934 452478
rect 238334 452476 238654 452478
rect 269054 452476 269374 452478
rect 306804 452476 307404 452478
rect 414804 452476 415404 452478
rect 558804 452476 559404 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 39086 452454
rect 39322 452218 69806 452454
rect 70042 452218 100526 452454
rect 100762 452218 131246 452454
rect 131482 452218 162986 452454
rect 163222 452218 207656 452454
rect 207892 452218 238376 452454
rect 238612 452218 269096 452454
rect 269332 452218 306986 452454
rect 307222 452218 414986 452454
rect 415222 452218 558986 452454
rect 559222 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 39086 452134
rect 39322 451898 69806 452134
rect 70042 451898 100526 452134
rect 100762 451898 131246 452134
rect 131482 451898 162986 452134
rect 163222 451898 207656 452134
rect 207892 451898 238376 452134
rect 238612 451898 269096 452134
rect 269332 451898 306986 452134
rect 307222 451898 414986 452134
rect 415222 451898 558986 452134
rect 559222 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 39044 451874 39364 451876
rect 69764 451874 70084 451876
rect 100484 451874 100804 451876
rect 131204 451874 131524 451876
rect 162804 451874 163404 451876
rect 207614 451874 207934 451876
rect 238334 451874 238654 451876
rect 269054 451874 269374 451876
rect 306804 451874 307404 451876
rect 414804 451874 415404 451876
rect 558804 451874 559404 451876
rect 586260 451874 586860 451876
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 23684 434476 24004 434478
rect 54404 434476 54724 434478
rect 85124 434476 85444 434478
rect 115844 434476 116164 434478
rect 146564 434476 146884 434478
rect 180804 434476 181404 434478
rect 192254 434476 192574 434478
rect 222974 434476 223294 434478
rect 253694 434476 254014 434478
rect 288804 434476 289404 434478
rect 432804 434476 433404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 23726 434454
rect 23962 434218 54446 434454
rect 54682 434218 85166 434454
rect 85402 434218 115886 434454
rect 116122 434218 146606 434454
rect 146842 434218 180986 434454
rect 181222 434218 192296 434454
rect 192532 434218 223016 434454
rect 223252 434218 253736 434454
rect 253972 434218 288986 434454
rect 289222 434218 432986 434454
rect 433222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 23726 434134
rect 23962 433898 54446 434134
rect 54682 433898 85166 434134
rect 85402 433898 115886 434134
rect 116122 433898 146606 434134
rect 146842 433898 180986 434134
rect 181222 433898 192296 434134
rect 192532 433898 223016 434134
rect 223252 433898 253736 434134
rect 253972 433898 288986 434134
rect 289222 433898 432986 434134
rect 433222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 23684 433874 24004 433876
rect 54404 433874 54724 433876
rect 85124 433874 85444 433876
rect 115844 433874 116164 433876
rect 146564 433874 146884 433876
rect 180804 433874 181404 433876
rect 192254 433874 192574 433876
rect 222974 433874 223294 433876
rect 253694 433874 254014 433876
rect 288804 433874 289404 433876
rect 432804 433874 433404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect 155780 421378 281772 421420
rect 155780 421142 155822 421378
rect 156058 421142 281494 421378
rect 281730 421142 281772 421378
rect 155780 421100 281772 421142
rect -2936 416476 -2336 416478
rect 39044 416476 39364 416478
rect 69764 416476 70084 416478
rect 100484 416476 100804 416478
rect 131204 416476 131524 416478
rect 162804 416476 163404 416478
rect 207614 416476 207934 416478
rect 238334 416476 238654 416478
rect 269054 416476 269374 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 39086 416454
rect 39322 416218 69806 416454
rect 70042 416218 100526 416454
rect 100762 416218 131246 416454
rect 131482 416218 162986 416454
rect 163222 416218 207656 416454
rect 207892 416218 238376 416454
rect 238612 416218 269096 416454
rect 269332 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 39086 416134
rect 39322 415898 69806 416134
rect 70042 415898 100526 416134
rect 100762 415898 131246 416134
rect 131482 415898 162986 416134
rect 163222 415898 207656 416134
rect 207892 415898 238376 416134
rect 238612 415898 269096 416134
rect 269332 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 39044 415874 39364 415876
rect 69764 415874 70084 415876
rect 100484 415874 100804 415876
rect 131204 415874 131524 415876
rect 162804 415874 163404 415876
rect 207614 415874 207934 415876
rect 238334 415874 238654 415876
rect 269054 415874 269374 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586260 415874 586860 415876
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 38875 380476 39195 380478
rect 56805 380476 57125 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 38917 380454
rect 39153 380218 56847 380454
rect 57083 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 38917 380134
rect 39153 379898 56847 380134
rect 57083 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 38875 379874 39195 379876
rect 56805 379874 57125 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 29909 362476 30229 362478
rect 47840 362476 48160 362478
rect 65770 362476 66090 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 29951 362454
rect 30187 362218 47882 362454
rect 48118 362218 65812 362454
rect 66048 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 29951 362134
rect 30187 361898 47882 362134
rect 48118 361898 65812 362134
rect 66048 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 29909 361874 30229 361876
rect 47840 361874 48160 361876
rect 65770 361874 66090 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 107675 344476 107995 344478
rect 192805 344476 193125 344478
rect 306804 344476 307404 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 107717 344454
rect 107953 344218 192847 344454
rect 193083 344218 306986 344454
rect 307222 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 107717 344134
rect 107953 343898 192847 344134
rect 193083 343898 306986 344134
rect 307222 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 107675 343874 107995 343876
rect 192805 343874 193125 343876
rect 306804 343874 307404 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 65109 326476 65429 326478
rect 150240 326476 150560 326478
rect 235370 326476 235690 326478
rect 288804 326476 289404 326478
rect 293189 326476 293509 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 65151 326454
rect 65387 326218 150282 326454
rect 150518 326218 235412 326454
rect 235648 326218 288986 326454
rect 289222 326218 293231 326454
rect 293467 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 65151 326134
rect 65387 325898 150282 326134
rect 150518 325898 235412 326134
rect 235648 325898 288986 326134
rect 289222 325898 293231 326134
rect 293467 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 65109 325874 65429 325876
rect 150240 325874 150560 325876
rect 235370 325874 235690 325876
rect 288804 325874 289404 325876
rect 293189 325874 293509 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 39614 308476 39934 308478
rect 70334 308476 70654 308478
rect 101054 308476 101374 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 207568 308476 207888 308478
rect 238288 308476 238608 308478
rect 269008 308476 269328 308478
rect 294635 308476 294955 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 39656 308454
rect 39892 308218 70376 308454
rect 70612 308218 101096 308454
rect 101332 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 207610 308454
rect 207846 308218 238330 308454
rect 238566 308218 269050 308454
rect 269286 308218 294677 308454
rect 294913 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 39656 308134
rect 39892 307898 70376 308134
rect 70612 307898 101096 308134
rect 101332 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 207610 308134
rect 207846 307898 238330 308134
rect 238566 307898 269050 308134
rect 269286 307898 294677 308134
rect 294913 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 39614 307874 39934 307876
rect 70334 307874 70654 307876
rect 101054 307874 101374 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 207568 307874 207888 307876
rect 238288 307874 238608 307876
rect 269008 307874 269328 307876
rect 294635 307874 294955 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 24254 290476 24574 290478
rect 54974 290476 55294 290478
rect 85694 290476 86014 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 192208 290476 192528 290478
rect 222928 290476 223248 290478
rect 253648 290476 253968 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 24296 290454
rect 24532 290218 55016 290454
rect 55252 290218 85736 290454
rect 85972 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 192250 290454
rect 192486 290218 222970 290454
rect 223206 290218 253690 290454
rect 253926 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 24296 290134
rect 24532 289898 55016 290134
rect 55252 289898 85736 290134
rect 85972 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 192250 290134
rect 192486 289898 222970 290134
rect 223206 289898 253690 290134
rect 253926 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 24254 289874 24574 289876
rect 54974 289874 55294 289876
rect 85694 289874 86014 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 192208 289874 192528 289876
rect 222928 289874 223248 289876
rect 253648 289874 253968 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 39614 272476 39934 272478
rect 70334 272476 70654 272478
rect 101054 272476 101374 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 207568 272476 207888 272478
rect 238288 272476 238608 272478
rect 269008 272476 269328 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 39656 272454
rect 39892 272218 70376 272454
rect 70612 272218 101096 272454
rect 101332 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 207610 272454
rect 207846 272218 238330 272454
rect 238566 272218 269050 272454
rect 269286 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 39656 272134
rect 39892 271898 70376 272134
rect 70612 271898 101096 272134
rect 101332 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 207610 272134
rect 207846 271898 238330 272134
rect 238566 271898 269050 272134
rect 269286 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 39614 271874 39934 271876
rect 70334 271874 70654 271876
rect 101054 271874 101374 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 207568 271874 207888 271876
rect 238288 271874 238608 271876
rect 269008 271874 269328 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586260 271874 586860 271876
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 24254 254476 24574 254478
rect 54974 254476 55294 254478
rect 85694 254476 86014 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 192208 254476 192528 254478
rect 222928 254476 223248 254478
rect 253648 254476 253968 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 24296 254454
rect 24532 254218 55016 254454
rect 55252 254218 85736 254454
rect 85972 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 192250 254454
rect 192486 254218 222970 254454
rect 223206 254218 253690 254454
rect 253926 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 24296 254134
rect 24532 253898 55016 254134
rect 55252 253898 85736 254134
rect 85972 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 192250 254134
rect 192486 253898 222970 254134
rect 223206 253898 253690 254134
rect 253926 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 24254 253874 24574 253876
rect 54974 253874 55294 253876
rect 85694 253874 86014 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 192208 253874 192528 253876
rect 222928 253874 223248 253876
rect 253648 253874 253968 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586260 235874 586860 235876
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 108804 218476 109404 218478
rect 123808 218476 124128 218478
rect 154528 218476 154848 218478
rect 185248 218476 185568 218478
rect 216804 218476 217404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 108986 218454
rect 109222 218218 123850 218454
rect 124086 218218 154570 218454
rect 154806 218218 185290 218454
rect 185526 218218 216986 218454
rect 217222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 108986 218134
rect 109222 217898 123850 218134
rect 124086 217898 154570 218134
rect 154806 217898 185290 218134
rect 185526 217898 216986 218134
rect 217222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 108804 217874 109404 217876
rect 123808 217874 124128 217876
rect 154528 217874 154848 217876
rect 185248 217874 185568 217876
rect 216804 217874 217404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -2936 200476 -2336 200478
rect 28768 200476 29088 200478
rect 59488 200476 59808 200478
rect 90208 200476 90528 200478
rect 139168 200476 139488 200478
rect 169888 200476 170208 200478
rect 200608 200476 200928 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 28810 200454
rect 29046 200218 59530 200454
rect 59766 200218 90250 200454
rect 90486 200218 139210 200454
rect 139446 200218 169930 200454
rect 170166 200218 200650 200454
rect 200886 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 28810 200134
rect 29046 199898 59530 200134
rect 59766 199898 90250 200134
rect 90486 199898 139210 200134
rect 139446 199898 169930 200134
rect 170166 199898 200650 200134
rect 200886 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 28768 199874 29088 199876
rect 59488 199874 59808 199876
rect 90208 199874 90528 199876
rect 139168 199874 139488 199876
rect 169888 199874 170208 199876
rect 200608 199874 200928 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586260 199874 586860 199876
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 13408 182476 13728 182478
rect 44128 182476 44448 182478
rect 74848 182476 75168 182478
rect 108804 182476 109404 182478
rect 123808 182476 124128 182478
rect 154528 182476 154848 182478
rect 185248 182476 185568 182478
rect 216804 182476 217404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 13450 182454
rect 13686 182218 44170 182454
rect 44406 182218 74890 182454
rect 75126 182218 108986 182454
rect 109222 182218 123850 182454
rect 124086 182218 154570 182454
rect 154806 182218 185290 182454
rect 185526 182218 216986 182454
rect 217222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 13450 182134
rect 13686 181898 44170 182134
rect 44406 181898 74890 182134
rect 75126 181898 108986 182134
rect 109222 181898 123850 182134
rect 124086 181898 154570 182134
rect 154806 181898 185290 182134
rect 185526 181898 216986 182134
rect 217222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 13408 181874 13728 181876
rect 44128 181874 44448 181876
rect 74848 181874 75168 181876
rect 108804 181874 109404 181876
rect 123808 181874 124128 181876
rect 154528 181874 154848 181876
rect 185248 181874 185568 181876
rect 216804 181874 217404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -2936 164476 -2336 164478
rect 28768 164476 29088 164478
rect 59488 164476 59808 164478
rect 90208 164476 90528 164478
rect 139168 164476 139488 164478
rect 169888 164476 170208 164478
rect 200608 164476 200928 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 28810 164454
rect 29046 164218 59530 164454
rect 59766 164218 90250 164454
rect 90486 164218 139210 164454
rect 139446 164218 169930 164454
rect 170166 164218 200650 164454
rect 200886 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 28810 164134
rect 29046 163898 59530 164134
rect 59766 163898 90250 164134
rect 90486 163898 139210 164134
rect 139446 163898 169930 164134
rect 170166 163898 200650 164134
rect 200886 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 28768 163874 29088 163876
rect 59488 163874 59808 163876
rect 90208 163874 90528 163876
rect 139168 163874 139488 163876
rect 169888 163874 170208 163876
rect 200608 163874 200928 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586260 163874 586860 163876
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 13408 146476 13728 146478
rect 44128 146476 44448 146478
rect 74848 146476 75168 146478
rect 108804 146476 109404 146478
rect 123808 146476 124128 146478
rect 154528 146476 154848 146478
rect 185248 146476 185568 146478
rect 216804 146476 217404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 13450 146454
rect 13686 146218 44170 146454
rect 44406 146218 74890 146454
rect 75126 146218 108986 146454
rect 109222 146218 123850 146454
rect 124086 146218 154570 146454
rect 154806 146218 185290 146454
rect 185526 146218 216986 146454
rect 217222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 13450 146134
rect 13686 145898 44170 146134
rect 44406 145898 74890 146134
rect 75126 145898 108986 146134
rect 109222 145898 123850 146134
rect 124086 145898 154570 146134
rect 154806 145898 185290 146134
rect 185526 145898 216986 146134
rect 217222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 13408 145874 13728 145876
rect 44128 145874 44448 145876
rect 74848 145874 75168 145876
rect 108804 145874 109404 145876
rect 123808 145874 124128 145876
rect 154528 145874 154848 145876
rect 185248 145874 185568 145876
rect 216804 145874 217404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -2936 128476 -2336 128478
rect 139168 128476 139488 128478
rect 169888 128476 170208 128478
rect 200608 128476 200928 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 139210 128454
rect 139446 128218 169930 128454
rect 170166 128218 200650 128454
rect 200886 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 139210 128134
rect 139446 127898 169930 128134
rect 170166 127898 200650 128134
rect 200886 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 139168 127874 139488 127876
rect 169888 127874 170208 127876
rect 200608 127874 200928 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586260 127874 586860 127876
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 123808 110476 124128 110478
rect 154528 110476 154848 110478
rect 185248 110476 185568 110478
rect 216804 110476 217404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 123850 110454
rect 124086 110218 154570 110454
rect 154806 110218 185290 110454
rect 185526 110218 216986 110454
rect 217222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 123850 110134
rect 124086 109898 154570 110134
rect 154806 109898 185290 110134
rect 185526 109898 216986 110134
rect 217222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 123808 109874 124128 109876
rect 154528 109874 154848 109876
rect 185248 109874 185568 109876
rect 216804 109874 217404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -2936 92476 -2336 92478
rect 28768 92476 29088 92478
rect 59488 92476 59808 92478
rect 90208 92476 90528 92478
rect 139168 92476 139488 92478
rect 169888 92476 170208 92478
rect 200608 92476 200928 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 28810 92454
rect 29046 92218 59530 92454
rect 59766 92218 90250 92454
rect 90486 92218 139210 92454
rect 139446 92218 169930 92454
rect 170166 92218 200650 92454
rect 200886 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 28810 92134
rect 29046 91898 59530 92134
rect 59766 91898 90250 92134
rect 90486 91898 139210 92134
rect 139446 91898 169930 92134
rect 170166 91898 200650 92134
rect 200886 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 28768 91874 29088 91876
rect 59488 91874 59808 91876
rect 90208 91874 90528 91876
rect 139168 91874 139488 91876
rect 169888 91874 170208 91876
rect 200608 91874 200928 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586260 91874 586860 91876
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 13408 74476 13728 74478
rect 44128 74476 44448 74478
rect 74848 74476 75168 74478
rect 108804 74476 109404 74478
rect 123808 74476 124128 74478
rect 154528 74476 154848 74478
rect 185248 74476 185568 74478
rect 216804 74476 217404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 13450 74454
rect 13686 74218 44170 74454
rect 44406 74218 74890 74454
rect 75126 74218 108986 74454
rect 109222 74218 123850 74454
rect 124086 74218 154570 74454
rect 154806 74218 185290 74454
rect 185526 74218 216986 74454
rect 217222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 13450 74134
rect 13686 73898 44170 74134
rect 44406 73898 74890 74134
rect 75126 73898 108986 74134
rect 109222 73898 123850 74134
rect 124086 73898 154570 74134
rect 154806 73898 185290 74134
rect 185526 73898 216986 74134
rect 217222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 13408 73874 13728 73876
rect 44128 73874 44448 73876
rect 74848 73874 75168 73876
rect 108804 73874 109404 73876
rect 123808 73874 124128 73876
rect 154528 73874 154848 73876
rect 185248 73874 185568 73876
rect 216804 73874 217404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -2936 56476 -2336 56478
rect 28768 56476 29088 56478
rect 59488 56476 59808 56478
rect 90208 56476 90528 56478
rect 139168 56476 139488 56478
rect 169888 56476 170208 56478
rect 200608 56476 200928 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 433568 56476 433888 56478
rect 464288 56476 464608 56478
rect 495008 56476 495328 56478
rect 525728 56476 526048 56478
rect 556448 56476 556768 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 28810 56454
rect 29046 56218 59530 56454
rect 59766 56218 90250 56454
rect 90486 56218 139210 56454
rect 139446 56218 169930 56454
rect 170166 56218 200650 56454
rect 200886 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 433610 56454
rect 433846 56218 464330 56454
rect 464566 56218 495050 56454
rect 495286 56218 525770 56454
rect 526006 56218 556490 56454
rect 556726 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 28810 56134
rect 29046 55898 59530 56134
rect 59766 55898 90250 56134
rect 90486 55898 139210 56134
rect 139446 55898 169930 56134
rect 170166 55898 200650 56134
rect 200886 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 433610 56134
rect 433846 55898 464330 56134
rect 464566 55898 495050 56134
rect 495286 55898 525770 56134
rect 526006 55898 556490 56134
rect 556726 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 28768 55874 29088 55876
rect 59488 55874 59808 55876
rect 90208 55874 90528 55876
rect 139168 55874 139488 55876
rect 169888 55874 170208 55876
rect 200608 55874 200928 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 433568 55874 433888 55876
rect 464288 55874 464608 55876
rect 495008 55874 495328 55876
rect 525728 55874 526048 55876
rect 556448 55874 556768 55876
rect 586260 55874 586860 55876
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 13408 38476 13728 38478
rect 44128 38476 44448 38478
rect 74848 38476 75168 38478
rect 108804 38476 109404 38478
rect 123808 38476 124128 38478
rect 154528 38476 154848 38478
rect 185248 38476 185568 38478
rect 216804 38476 217404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 418208 38476 418528 38478
rect 448928 38476 449248 38478
rect 479648 38476 479968 38478
rect 510368 38476 510688 38478
rect 541088 38476 541408 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 13450 38454
rect 13686 38218 44170 38454
rect 44406 38218 74890 38454
rect 75126 38218 108986 38454
rect 109222 38218 123850 38454
rect 124086 38218 154570 38454
rect 154806 38218 185290 38454
rect 185526 38218 216986 38454
rect 217222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 418250 38454
rect 418486 38218 448970 38454
rect 449206 38218 479690 38454
rect 479926 38218 510410 38454
rect 510646 38218 541130 38454
rect 541366 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 13450 38134
rect 13686 37898 44170 38134
rect 44406 37898 74890 38134
rect 75126 37898 108986 38134
rect 109222 37898 123850 38134
rect 124086 37898 154570 38134
rect 154806 37898 185290 38134
rect 185526 37898 216986 38134
rect 217222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 418250 38134
rect 418486 37898 448970 38134
rect 449206 37898 479690 38134
rect 479926 37898 510410 38134
rect 510646 37898 541130 38134
rect 541366 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 13408 37874 13728 37876
rect 44128 37874 44448 37876
rect 74848 37874 75168 37876
rect 108804 37874 109404 37876
rect 123808 37874 124128 37876
rect 154528 37874 154848 37876
rect 185248 37874 185568 37876
rect 216804 37874 217404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 418208 37874 418528 37876
rect 448928 37874 449248 37876
rect 479648 37874 479968 37876
rect 510368 37874 510688 37876
rect 541088 37874 541408 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 433568 20476 433888 20478
rect 464288 20476 464608 20478
rect 495008 20476 495328 20478
rect 525728 20476 526048 20478
rect 556448 20476 556768 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 433610 20454
rect 433846 20218 464330 20454
rect 464566 20218 495050 20454
rect 495286 20218 525770 20454
rect 526006 20218 556490 20454
rect 556726 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 433610 20134
rect 433846 19898 464330 20134
rect 464566 19898 495050 20134
rect 495286 19898 525770 20134
rect 526006 19898 556490 20134
rect 556726 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 433568 19874 433888 19876
rect 464288 19874 464608 19876
rect 495008 19874 495328 19876
rect 525728 19874 526048 19876
rect 556448 19874 556768 19876
rect 586260 19874 586860 19876
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 591900 -7506 592500 -7504
use fd_hd  i_fd0_1
timestamp 1608318970
transform 1 0 230000 0 1 31440
box 0 0 108256 50048
use fd_hs  i_fd0_2
timestamp 1608318970
transform 1 0 230000 0 1 103440
box 0 0 112240 46240
use fd_ms  i_fd0_3
timestamp 1608318970
transform 1 0 230000 0 1 175440
box 0 0 106720 46240
use wb_interface  i_itf0
timestamp 1608318970
transform 1 0 119600 0 1 31440
box 0 0 92000 190400
use tdc_inline_1  i_tdc0_1
timestamp 1608318970
transform 1 0 9200 0 1 31440
box 0 0 82800 68000
use tdc_inline_2  i_tdc0_2
timestamp 1608318970
transform 1 0 9200 0 1 127228
box 0 0 92000 92480
use rescue_top  inst_rescue
timestamp 1608318970
transform 1 0 414000 0 1 16320
box 0 0 147200 44608
use fd_inline_1  i_fd2_2
timestamp 1608318970
transform 1 0 20000 0 -1 384200
box 290 2042 56000 27200
use fd_hd_25_1  i_fd2_3
timestamp 1608318970
transform 1 0 188000 0 -1 402224
box 0 0 94746 44112
use wb_extender  i_itf2
timestamp 1608318970
transform 1 0 21600 0 1 322800
box 474 0 257600 26112
use tdc_inline_3  i_tdc2_0
timestamp 1608318970
transform 1 0 20046 0 1 234000
box 0 2128 92000 81600
use tdc_inline_3  i_tdc2_1
timestamp 1608318970
transform 1 0 188000 0 1 234000
box 0 2128 92000 81600
use zero  b_zero.i_zero
timestamp 1608318970
transform 1 0 290800 0 1 304800
box 0 0 10880 24480
use fd_hs  i_fd3_2
timestamp 1608318970
transform 1 0 28000 0 1 571440
box 0 0 112240 46240
use fd_hd_25_1  i_fd3_3
timestamp 1608318970
transform 1 0 188000 0 -1 618224
box 0 0 94746 44112
use wb_extender  i_itf3
timestamp 1608318970
transform 1 0 21600 0 1 502800
box 474 0 257600 26112
use tdc_hd_cbuf2_x4  i_tdc3_0
timestamp 1608318970
transform 1 0 16000 0 1 400000
box 0 2128 138000 87040
use tdc_inline_3  i_tdc3_1
timestamp 1608318970
transform 1 0 188046 0 1 410000
box 0 2128 92000 81600
use fd_ms  i_fd4_2
timestamp 1608318970
transform -1 0 552720 0 1 427440
box 0 0 106720 46240
use fd_hd_25_1  i_fd4_3
timestamp 1608318970
transform -1 0 410746 0 1 430128
box 0 0 94746 44112
use wb_extender  i_itf4
timestamp 1608318970
transform -1 0 575246 0 -1 528912
box 474 0 257600 26112
use tdc_inline_2  i_tdc4_0
timestamp 1608318970
transform 1 0 460000 0 1 570000
box 0 0 92000 92480
use tdc_hd_cbuf2_x4  i_tdc4_1
timestamp 1608318970
transform 1 0 316046 0 -1 657040
box 0 2128 138000 87040
<< labels >>
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 0 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 1 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 2 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 3 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 4 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 5 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 6 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 7 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 8 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 9 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 10 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 11 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 12 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 13 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 14 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 15 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 16 nsew default tristate
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 17 nsew default input
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 18 nsew default input
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 19 nsew default input
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 20 nsew default input
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 21 nsew default input
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 22 nsew default input
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 23 nsew default input
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 24 nsew default input
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 25 nsew default input
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 26 nsew default input
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 27 nsew default input
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 28 nsew default input
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 29 nsew default input
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 30 nsew default input
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 31 nsew default input
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 32 nsew default input
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 33 nsew default input
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 34 nsew default input
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 35 nsew default input
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 36 nsew default input
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 37 nsew default input
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 38 nsew default input
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 39 nsew default input
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 40 nsew default input
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 41 nsew default input
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 42 nsew default input
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 43 nsew default input
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 44 nsew default input
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 45 nsew default input
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 46 nsew default input
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 47 nsew default input
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 48 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 49 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 50 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 51 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 52 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 53 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 54 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 55 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 56 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 57 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 58 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 59 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 60 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 61 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 62 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 63 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 64 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 65 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 66 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 67 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 68 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 69 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 70 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 71 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 72 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 73 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 74 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 75 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 76 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 77 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 78 nsew default tristate
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 79 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 80 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 81 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 82 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 83 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 84 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 85 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 86 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 87 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 88 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 89 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 90 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 91 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 92 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 93 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 94 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 95 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 96 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 97 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 98 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 99 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 100 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 101 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 102 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 103 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 104 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 105 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 106 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 107 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 108 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 109 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 110 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 111 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 112 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 113 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 114 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 115 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 116 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 117 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 118 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 119 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 120 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 121 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 122 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 123 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 124 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 125 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 126 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 127 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 128 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 129 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 130 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 131 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 132 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 133 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 134 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 135 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 136 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 137 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 138 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 139 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 140 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 141 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 142 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 143 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 638 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 639 nsew default input
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 640 nsew default input
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 641 nsew default input
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 642 nsew default input
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
