magic
tech sky130A
magscale 1 2
timestamp 1607421480
<< locali >>
rect 41245 5559 41279 5797
rect 87797 5559 87831 5797
rect 50721 2907 50755 3009
rect 102609 2363 102643 2533
<< viali >>
rect 1133 7293 1167 7327
rect 1409 7293 1443 7327
rect 3249 7293 3283 7327
rect 3525 7293 3559 7327
rect 5365 7293 5399 7327
rect 5641 7293 5675 7327
rect 7481 7293 7515 7327
rect 7757 7293 7791 7327
rect 9597 7293 9631 7327
rect 9873 7293 9907 7327
rect 11713 7293 11747 7327
rect 11989 7293 12023 7327
rect 13829 7293 13863 7327
rect 14105 7293 14139 7327
rect 15945 7293 15979 7327
rect 16221 7293 16255 7327
rect 18061 7293 18095 7327
rect 18337 7293 18371 7327
rect 20177 7293 20211 7327
rect 20453 7293 20487 7327
rect 22293 7293 22327 7327
rect 22569 7293 22603 7327
rect 24409 7293 24443 7327
rect 24685 7293 24719 7327
rect 26525 7293 26559 7327
rect 26801 7293 26835 7327
rect 28641 7293 28675 7327
rect 28917 7293 28951 7327
rect 30757 7293 30791 7327
rect 31033 7293 31067 7327
rect 32873 7293 32907 7327
rect 33149 7293 33183 7327
rect 34989 7293 35023 7327
rect 35265 7293 35299 7327
rect 37105 7293 37139 7327
rect 37381 7293 37415 7327
rect 39221 7293 39255 7327
rect 39497 7293 39531 7327
rect 41337 7293 41371 7327
rect 41613 7293 41647 7327
rect 43453 7293 43487 7327
rect 43729 7293 43763 7327
rect 45569 7293 45603 7327
rect 45845 7293 45879 7327
rect 47685 7293 47719 7327
rect 47961 7293 47995 7327
rect 49801 7293 49835 7327
rect 50077 7293 50111 7327
rect 51917 7293 51951 7327
rect 52193 7293 52227 7327
rect 54033 7293 54067 7327
rect 54309 7293 54343 7327
rect 56149 7293 56183 7327
rect 56425 7293 56459 7327
rect 58265 7293 58299 7327
rect 58541 7293 58575 7327
rect 60381 7293 60415 7327
rect 60657 7293 60691 7327
rect 62497 7293 62531 7327
rect 62773 7293 62807 7327
rect 64613 7293 64647 7327
rect 64889 7293 64923 7327
rect 66729 7293 66763 7327
rect 67005 7293 67039 7327
rect 68845 7293 68879 7327
rect 69121 7293 69155 7327
rect 70961 7293 70995 7327
rect 71237 7293 71271 7327
rect 73077 7293 73111 7327
rect 73353 7293 73387 7327
rect 75193 7293 75227 7327
rect 75469 7293 75503 7327
rect 77309 7293 77343 7327
rect 77585 7293 77619 7327
rect 79425 7293 79459 7327
rect 79701 7293 79735 7327
rect 81541 7293 81575 7327
rect 81817 7293 81851 7327
rect 83657 7293 83691 7327
rect 83933 7293 83967 7327
rect 85773 7293 85807 7327
rect 86049 7293 86083 7327
rect 87889 7293 87923 7327
rect 88165 7293 88199 7327
rect 90005 7293 90039 7327
rect 90281 7293 90315 7327
rect 92121 7293 92155 7327
rect 92397 7293 92431 7327
rect 94237 7293 94271 7327
rect 94513 7293 94547 7327
rect 96353 7293 96387 7327
rect 96629 7293 96663 7327
rect 98469 7293 98503 7327
rect 98745 7293 98779 7327
rect 100585 7293 100619 7327
rect 100861 7293 100895 7327
rect 102701 7293 102735 7327
rect 102977 7293 103011 7327
rect 104817 7293 104851 7327
rect 105093 7293 105127 7327
rect 11253 7225 11287 7259
rect 13369 7225 13403 7259
rect 23949 7225 23983 7259
rect 30297 7225 30331 7259
rect 47225 7225 47259 7259
rect 64153 7225 64187 7259
rect 78965 7225 78999 7259
rect 81081 7225 81115 7259
rect 95893 7225 95927 7259
rect 98009 7225 98043 7259
rect 2513 7157 2547 7191
rect 4629 7157 4663 7191
rect 6745 7157 6779 7191
rect 9045 7157 9079 7191
rect 15209 7157 15243 7191
rect 17325 7157 17359 7191
rect 19441 7157 19475 7191
rect 21557 7157 21591 7191
rect 25973 7157 26007 7191
rect 28089 7157 28123 7191
rect 32137 7157 32171 7191
rect 34253 7157 34287 7191
rect 36369 7157 36403 7191
rect 38485 7157 38519 7191
rect 40601 7157 40635 7191
rect 42901 7157 42935 7191
rect 45017 7157 45051 7191
rect 49065 7157 49099 7191
rect 51181 7157 51215 7191
rect 53297 7157 53331 7191
rect 55413 7157 55447 7191
rect 57529 7157 57563 7191
rect 59829 7157 59863 7191
rect 61945 7157 61979 7191
rect 65993 7157 66027 7191
rect 68109 7157 68143 7191
rect 70225 7157 70259 7191
rect 72341 7157 72375 7191
rect 74457 7157 74491 7191
rect 76757 7157 76791 7191
rect 82921 7157 82955 7191
rect 85221 7157 85255 7191
rect 87153 7157 87187 7191
rect 89269 7157 89303 7191
rect 91385 7157 91419 7191
rect 93685 7157 93719 7191
rect 99849 7157 99883 7191
rect 101965 7157 101999 7191
rect 104081 7157 104115 7191
rect 106197 7157 106231 7191
rect 2513 6953 2547 6987
rect 4629 6953 4663 6987
rect 6745 6953 6779 6987
rect 8861 6953 8895 6987
rect 10977 6953 11011 6987
rect 13093 6953 13127 6987
rect 15209 6953 15243 6987
rect 17325 6953 17359 6987
rect 19441 6953 19475 6987
rect 21557 6953 21591 6987
rect 23673 6953 23707 6987
rect 25789 6953 25823 6987
rect 27905 6953 27939 6987
rect 30021 6953 30055 6987
rect 32137 6953 32171 6987
rect 34253 6953 34287 6987
rect 36369 6953 36403 6987
rect 38485 6953 38519 6987
rect 40601 6953 40635 6987
rect 42717 6953 42751 6987
rect 44833 6953 44867 6987
rect 46949 6953 46983 6987
rect 49065 6953 49099 6987
rect 51181 6953 51215 6987
rect 53297 6953 53331 6987
rect 55413 6953 55447 6987
rect 57529 6953 57563 6987
rect 59645 6953 59679 6987
rect 61761 6953 61795 6987
rect 63877 6953 63911 6987
rect 65993 6953 66027 6987
rect 68109 6953 68143 6987
rect 70225 6953 70259 6987
rect 72341 6953 72375 6987
rect 74457 6953 74491 6987
rect 76573 6953 76607 6987
rect 78689 6953 78723 6987
rect 80805 6953 80839 6987
rect 82921 6953 82955 6987
rect 85037 6953 85071 6987
rect 87153 6953 87187 6987
rect 89269 6953 89303 6987
rect 91385 6953 91419 6987
rect 93501 6953 93535 6987
rect 95617 6953 95651 6987
rect 97733 6953 97767 6987
rect 99849 6953 99883 6987
rect 101965 6953 101999 6987
rect 104081 6953 104115 6987
rect 106197 6953 106231 6987
rect 1133 6817 1167 6851
rect 3249 6817 3283 6851
rect 5365 6817 5399 6851
rect 7481 6817 7515 6851
rect 9597 6817 9631 6851
rect 11713 6817 11747 6851
rect 13829 6817 13863 6851
rect 15945 6817 15979 6851
rect 18061 6817 18095 6851
rect 20177 6817 20211 6851
rect 22293 6817 22327 6851
rect 24409 6817 24443 6851
rect 26525 6817 26559 6851
rect 28641 6817 28675 6851
rect 30757 6817 30791 6851
rect 32873 6817 32907 6851
rect 34989 6817 35023 6851
rect 37105 6817 37139 6851
rect 39221 6817 39255 6851
rect 41337 6817 41371 6851
rect 43453 6817 43487 6851
rect 45569 6817 45603 6851
rect 47685 6817 47719 6851
rect 49801 6817 49835 6851
rect 51917 6817 51951 6851
rect 54033 6817 54067 6851
rect 56149 6817 56183 6851
rect 58265 6817 58299 6851
rect 62497 6817 62531 6851
rect 64613 6817 64647 6851
rect 66729 6817 66763 6851
rect 68845 6817 68879 6851
rect 70961 6817 70995 6851
rect 73077 6817 73111 6851
rect 75193 6817 75227 6851
rect 79425 6817 79459 6851
rect 81541 6817 81575 6851
rect 83657 6817 83691 6851
rect 85773 6817 85807 6851
rect 87889 6817 87923 6851
rect 90005 6817 90039 6851
rect 92121 6817 92155 6851
rect 94237 6817 94271 6851
rect 96353 6817 96387 6851
rect 98469 6817 98503 6851
rect 100585 6817 100619 6851
rect 102701 6817 102735 6851
rect 104817 6817 104851 6851
rect 1409 6749 1443 6783
rect 3525 6749 3559 6783
rect 5641 6749 5675 6783
rect 7757 6749 7791 6783
rect 9873 6749 9907 6783
rect 11989 6749 12023 6783
rect 14105 6749 14139 6783
rect 16221 6749 16255 6783
rect 18337 6749 18371 6783
rect 20453 6749 20487 6783
rect 22569 6749 22603 6783
rect 24685 6749 24719 6783
rect 26801 6749 26835 6783
rect 28917 6749 28951 6783
rect 31033 6749 31067 6783
rect 33149 6749 33183 6783
rect 35265 6749 35299 6783
rect 37381 6749 37415 6783
rect 39497 6749 39531 6783
rect 41613 6749 41647 6783
rect 43729 6749 43763 6783
rect 45845 6749 45879 6783
rect 47961 6749 47995 6783
rect 50077 6749 50111 6783
rect 52193 6749 52227 6783
rect 54309 6749 54343 6783
rect 56425 6749 56459 6783
rect 58541 6749 58575 6783
rect 60381 6749 60415 6783
rect 60657 6749 60691 6783
rect 62773 6749 62807 6783
rect 64889 6749 64923 6783
rect 67005 6749 67039 6783
rect 69121 6749 69155 6783
rect 71237 6749 71271 6783
rect 73353 6749 73387 6783
rect 75469 6749 75503 6783
rect 77309 6749 77343 6783
rect 77585 6749 77619 6783
rect 79701 6749 79735 6783
rect 81817 6749 81851 6783
rect 83933 6749 83967 6783
rect 86049 6749 86083 6783
rect 88165 6749 88199 6783
rect 90281 6749 90315 6783
rect 92397 6749 92431 6783
rect 94513 6749 94547 6783
rect 96629 6749 96663 6783
rect 98745 6749 98779 6783
rect 100861 6749 100895 6783
rect 102977 6749 103011 6783
rect 105093 6749 105127 6783
rect 3249 6341 3283 6375
rect 3433 6205 3467 6239
rect 5549 6205 5583 6239
rect 7481 6205 7515 6239
rect 7665 6205 7699 6239
rect 9597 6205 9631 6239
rect 9781 6205 9815 6239
rect 11713 6205 11747 6239
rect 11897 6205 11931 6239
rect 13829 6205 13863 6239
rect 14013 6205 14047 6239
rect 15945 6205 15979 6239
rect 16129 6205 16163 6239
rect 18061 6205 18095 6239
rect 18245 6205 18279 6239
rect 20177 6205 20211 6239
rect 20361 6205 20395 6239
rect 22293 6205 22327 6239
rect 22477 6205 22511 6239
rect 24409 6205 24443 6239
rect 24593 6205 24627 6239
rect 26525 6205 26559 6239
rect 26709 6205 26743 6239
rect 28641 6205 28675 6239
rect 28825 6205 28859 6239
rect 30757 6205 30791 6239
rect 30941 6205 30975 6239
rect 32873 6205 32907 6239
rect 33057 6205 33091 6239
rect 34989 6205 35023 6239
rect 35173 6205 35207 6239
rect 37105 6205 37139 6239
rect 37289 6205 37323 6239
rect 39221 6205 39255 6239
rect 41521 6205 41555 6239
rect 43453 6205 43487 6239
rect 43637 6205 43671 6239
rect 45569 6205 45603 6239
rect 45753 6205 45787 6239
rect 47685 6205 47719 6239
rect 47869 6205 47903 6239
rect 49801 6205 49835 6239
rect 49985 6205 50019 6239
rect 52101 6205 52135 6239
rect 54033 6205 54067 6239
rect 54217 6205 54251 6239
rect 56149 6205 56183 6239
rect 56333 6205 56367 6239
rect 58265 6205 58299 6239
rect 58449 6205 58483 6239
rect 60381 6205 60415 6239
rect 60565 6205 60599 6239
rect 62497 6205 62531 6239
rect 62681 6205 62715 6239
rect 64613 6205 64647 6239
rect 64797 6205 64831 6239
rect 66729 6205 66763 6239
rect 66913 6205 66947 6239
rect 68845 6205 68879 6239
rect 69029 6205 69063 6239
rect 70961 6205 70995 6239
rect 71145 6205 71179 6239
rect 73077 6205 73111 6239
rect 73261 6205 73295 6239
rect 75193 6205 75227 6239
rect 77493 6205 77527 6239
rect 79425 6205 79459 6239
rect 79609 6205 79643 6239
rect 81541 6205 81575 6239
rect 81725 6205 81759 6239
rect 83657 6205 83691 6239
rect 83841 6205 83875 6239
rect 85773 6205 85807 6239
rect 88073 6205 88107 6239
rect 90005 6205 90039 6239
rect 90189 6205 90223 6239
rect 92121 6205 92155 6239
rect 92305 6205 92339 6239
rect 94237 6205 94271 6239
rect 94421 6205 94455 6239
rect 96353 6205 96387 6239
rect 96537 6205 96571 6239
rect 98469 6205 98503 6239
rect 98653 6205 98687 6239
rect 100585 6205 100619 6239
rect 100769 6205 100803 6239
rect 102701 6205 102735 6239
rect 102885 6205 102919 6239
rect 104817 6205 104851 6239
rect 105001 6205 105035 6239
rect 5365 6137 5399 6171
rect 39405 6137 39439 6171
rect 41337 6137 41371 6171
rect 75377 6137 75411 6171
rect 77309 6137 77343 6171
rect 85957 6137 85991 6171
rect 87889 6137 87923 6171
rect 52009 6069 52043 6103
rect 20361 5865 20395 5899
rect 22477 5865 22511 5899
rect 30941 5865 30975 5899
rect 35173 5865 35207 5899
rect 41521 5865 41555 5899
rect 60565 5865 60599 5899
rect 71145 5865 71179 5899
rect 77493 5865 77527 5899
rect 81725 5865 81759 5899
rect 102885 5865 102919 5899
rect 9873 5797 9907 5831
rect 11805 5797 11839 5831
rect 11989 5797 12023 5831
rect 13921 5797 13955 5831
rect 22385 5797 22419 5831
rect 24501 5797 24535 5831
rect 32965 5797 32999 5831
rect 37197 5797 37231 5831
rect 41245 5797 41279 5831
rect 41429 5797 41463 5831
rect 43545 5797 43579 5831
rect 45845 5797 45879 5831
rect 47777 5797 47811 5831
rect 56425 5797 56459 5831
rect 58357 5797 58391 5831
rect 58541 5797 58575 5831
rect 60473 5797 60507 5831
rect 62589 5797 62623 5831
rect 73169 5797 73203 5831
rect 77401 5797 77435 5831
rect 79517 5797 79551 5831
rect 83749 5797 83783 5831
rect 87797 5797 87831 5831
rect 87981 5797 88015 5831
rect 88165 5797 88199 5831
rect 90097 5797 90131 5831
rect 92397 5797 92431 5831
rect 94329 5797 94363 5831
rect 94513 5797 94547 5831
rect 96445 5797 96479 5831
rect 104909 5797 104943 5831
rect 105093 5797 105127 5831
rect 1225 5729 1259 5763
rect 1409 5729 1443 5763
rect 3341 5729 3375 5763
rect 5457 5729 5491 5763
rect 5641 5729 5675 5763
rect 7573 5729 7607 5763
rect 9689 5729 9723 5763
rect 16037 5729 16071 5763
rect 18153 5729 18187 5763
rect 18337 5729 18371 5763
rect 20269 5729 20303 5763
rect 26617 5729 26651 5763
rect 28733 5729 28767 5763
rect 28917 5729 28951 5763
rect 30849 5729 30883 5763
rect 33149 5729 33183 5763
rect 35081 5729 35115 5763
rect 39313 5729 39347 5763
rect 7757 5661 7791 5695
rect 14105 5661 14139 5695
rect 24685 5661 24719 5695
rect 26801 5661 26835 5695
rect 37381 5661 37415 5695
rect 16221 5593 16255 5627
rect 45661 5729 45695 5763
rect 47961 5729 47995 5763
rect 49893 5729 49927 5763
rect 52009 5729 52043 5763
rect 52193 5729 52227 5763
rect 54125 5729 54159 5763
rect 56241 5729 56275 5763
rect 64705 5729 64739 5763
rect 64889 5729 64923 5763
rect 66821 5729 66855 5763
rect 68937 5729 68971 5763
rect 69121 5729 69155 5763
rect 71053 5729 71087 5763
rect 75285 5729 75319 5763
rect 79701 5729 79735 5763
rect 81633 5729 81667 5763
rect 85865 5729 85899 5763
rect 43729 5661 43763 5695
rect 54309 5661 54343 5695
rect 62773 5661 62807 5695
rect 73353 5661 73387 5695
rect 83933 5661 83967 5695
rect 50077 5593 50111 5627
rect 67005 5593 67039 5627
rect 92213 5729 92247 5763
rect 96629 5729 96663 5763
rect 98561 5729 98595 5763
rect 100677 5729 100711 5763
rect 100861 5729 100895 5763
rect 102793 5729 102827 5763
rect 90281 5661 90315 5695
rect 98745 5661 98779 5695
rect 3433 5525 3467 5559
rect 39405 5525 39439 5559
rect 41245 5525 41279 5559
rect 75377 5525 75411 5559
rect 85957 5525 85991 5559
rect 87797 5525 87831 5559
rect 1133 5185 1167 5219
rect 1409 5185 1443 5219
rect 3249 5185 3283 5219
rect 3525 5185 3559 5219
rect 5365 5185 5399 5219
rect 5641 5185 5675 5219
rect 7481 5185 7515 5219
rect 7757 5185 7791 5219
rect 9597 5185 9631 5219
rect 9873 5185 9907 5219
rect 11713 5185 11747 5219
rect 11989 5185 12023 5219
rect 13829 5185 13863 5219
rect 14105 5185 14139 5219
rect 15945 5185 15979 5219
rect 16221 5185 16255 5219
rect 18061 5185 18095 5219
rect 18337 5185 18371 5219
rect 20177 5185 20211 5219
rect 20453 5185 20487 5219
rect 22293 5185 22327 5219
rect 22569 5185 22603 5219
rect 24409 5185 24443 5219
rect 24685 5185 24719 5219
rect 26525 5185 26559 5219
rect 26801 5185 26835 5219
rect 28641 5185 28675 5219
rect 28917 5185 28951 5219
rect 30757 5185 30791 5219
rect 31033 5185 31067 5219
rect 32873 5185 32907 5219
rect 33149 5185 33183 5219
rect 35265 5185 35299 5219
rect 37105 5185 37139 5219
rect 37381 5185 37415 5219
rect 39221 5185 39255 5219
rect 39497 5185 39531 5219
rect 41337 5185 41371 5219
rect 41613 5185 41647 5219
rect 43453 5185 43487 5219
rect 43729 5185 43763 5219
rect 45569 5185 45603 5219
rect 45845 5185 45879 5219
rect 47685 5185 47719 5219
rect 47961 5185 47995 5219
rect 49801 5185 49835 5219
rect 50077 5185 50111 5219
rect 51917 5185 51951 5219
rect 52193 5185 52227 5219
rect 54033 5185 54067 5219
rect 54309 5185 54343 5219
rect 56149 5185 56183 5219
rect 56425 5185 56459 5219
rect 58265 5185 58299 5219
rect 58541 5185 58575 5219
rect 60657 5185 60691 5219
rect 62497 5185 62531 5219
rect 62773 5185 62807 5219
rect 64613 5185 64647 5219
rect 64889 5185 64923 5219
rect 66729 5185 66763 5219
rect 67005 5185 67039 5219
rect 68845 5185 68879 5219
rect 69121 5185 69155 5219
rect 70961 5185 70995 5219
rect 71237 5185 71271 5219
rect 73077 5185 73111 5219
rect 73353 5185 73387 5219
rect 75193 5185 75227 5219
rect 75469 5185 75503 5219
rect 77585 5185 77619 5219
rect 79425 5185 79459 5219
rect 79701 5185 79735 5219
rect 81541 5185 81575 5219
rect 81817 5185 81851 5219
rect 83657 5185 83691 5219
rect 83933 5185 83967 5219
rect 85773 5185 85807 5219
rect 86049 5185 86083 5219
rect 87889 5185 87923 5219
rect 88165 5185 88199 5219
rect 90005 5185 90039 5219
rect 90281 5185 90315 5219
rect 92121 5185 92155 5219
rect 92397 5185 92431 5219
rect 94237 5185 94271 5219
rect 94513 5185 94547 5219
rect 96353 5185 96387 5219
rect 96629 5185 96663 5219
rect 98469 5185 98503 5219
rect 98745 5185 98779 5219
rect 100585 5185 100619 5219
rect 100861 5185 100895 5219
rect 102701 5185 102735 5219
rect 102977 5185 103011 5219
rect 104817 5185 104851 5219
rect 105093 5185 105127 5219
rect 34989 5117 35023 5151
rect 60381 5117 60415 5151
rect 77309 5117 77343 5151
rect 2513 4981 2547 5015
rect 4629 4981 4663 5015
rect 6745 4981 6779 5015
rect 8861 4981 8895 5015
rect 10977 4981 11011 5015
rect 13093 4981 13127 5015
rect 15209 4981 15243 5015
rect 17325 4981 17359 5015
rect 19441 4981 19475 5015
rect 21557 4981 21591 5015
rect 23673 4981 23707 5015
rect 25789 4981 25823 5015
rect 27905 4981 27939 5015
rect 30021 4981 30055 5015
rect 32137 4981 32171 5015
rect 34253 4981 34287 5015
rect 36369 4981 36403 5015
rect 38485 4981 38519 5015
rect 40601 4981 40635 5015
rect 42717 4981 42751 5015
rect 44833 4981 44867 5015
rect 46949 4981 46983 5015
rect 49065 4981 49099 5015
rect 51181 4981 51215 5015
rect 53297 4981 53331 5015
rect 55413 4981 55447 5015
rect 57529 4981 57563 5015
rect 59645 4981 59679 5015
rect 61761 4981 61795 5015
rect 63877 4981 63911 5015
rect 65993 4981 66027 5015
rect 68109 4981 68143 5015
rect 70225 4981 70259 5015
rect 72341 4981 72375 5015
rect 74457 4981 74491 5015
rect 76573 4981 76607 5015
rect 78689 4981 78723 5015
rect 80805 4981 80839 5015
rect 82921 4981 82955 5015
rect 85037 4981 85071 5015
rect 87153 4981 87187 5015
rect 89269 4981 89303 5015
rect 91385 4981 91419 5015
rect 93501 4981 93535 5015
rect 95617 4981 95651 5015
rect 97733 4981 97767 5015
rect 99849 4981 99883 5015
rect 101965 4981 101999 5015
rect 104081 4981 104115 5015
rect 106197 4981 106231 5015
rect 1409 4641 1443 4675
rect 3249 4641 3283 4675
rect 3525 4641 3559 4675
rect 5365 4641 5399 4675
rect 5641 4641 5675 4675
rect 7481 4641 7515 4675
rect 7757 4641 7791 4675
rect 9597 4641 9631 4675
rect 9873 4641 9907 4675
rect 11713 4641 11747 4675
rect 11989 4641 12023 4675
rect 13829 4641 13863 4675
rect 14105 4641 14139 4675
rect 15945 4641 15979 4675
rect 16221 4641 16255 4675
rect 18061 4641 18095 4675
rect 18337 4641 18371 4675
rect 20177 4641 20211 4675
rect 20453 4641 20487 4675
rect 22293 4641 22327 4675
rect 22569 4641 22603 4675
rect 24409 4641 24443 4675
rect 24685 4641 24719 4675
rect 26525 4641 26559 4675
rect 26801 4641 26835 4675
rect 28641 4641 28675 4675
rect 28917 4641 28951 4675
rect 30757 4641 30791 4675
rect 31033 4641 31067 4675
rect 32873 4641 32907 4675
rect 33149 4641 33183 4675
rect 34989 4641 35023 4675
rect 35265 4641 35299 4675
rect 37105 4641 37139 4675
rect 37381 4641 37415 4675
rect 39221 4641 39255 4675
rect 39497 4641 39531 4675
rect 41337 4641 41371 4675
rect 41613 4641 41647 4675
rect 43453 4641 43487 4675
rect 43729 4641 43763 4675
rect 45569 4641 45603 4675
rect 45845 4641 45879 4675
rect 47685 4641 47719 4675
rect 47961 4641 47995 4675
rect 49801 4641 49835 4675
rect 50077 4641 50111 4675
rect 51917 4641 51951 4675
rect 52193 4641 52227 4675
rect 54033 4641 54067 4675
rect 54309 4641 54343 4675
rect 56149 4641 56183 4675
rect 56425 4641 56459 4675
rect 58265 4641 58299 4675
rect 58541 4641 58575 4675
rect 60657 4641 60691 4675
rect 62497 4641 62531 4675
rect 62773 4641 62807 4675
rect 64613 4641 64647 4675
rect 64889 4641 64923 4675
rect 66729 4641 66763 4675
rect 67005 4641 67039 4675
rect 68845 4641 68879 4675
rect 69121 4641 69155 4675
rect 70961 4641 70995 4675
rect 71237 4641 71271 4675
rect 73077 4641 73111 4675
rect 73353 4641 73387 4675
rect 75193 4641 75227 4675
rect 75469 4641 75503 4675
rect 77585 4641 77619 4675
rect 79425 4641 79459 4675
rect 79701 4641 79735 4675
rect 81541 4641 81575 4675
rect 81817 4641 81851 4675
rect 83657 4641 83691 4675
rect 83933 4641 83967 4675
rect 85773 4641 85807 4675
rect 86049 4641 86083 4675
rect 87889 4641 87923 4675
rect 88165 4641 88199 4675
rect 90005 4641 90039 4675
rect 90281 4641 90315 4675
rect 92121 4641 92155 4675
rect 92397 4641 92431 4675
rect 94237 4641 94271 4675
rect 94513 4641 94547 4675
rect 96353 4641 96387 4675
rect 96629 4641 96663 4675
rect 98469 4641 98503 4675
rect 98745 4641 98779 4675
rect 100585 4641 100619 4675
rect 100861 4641 100895 4675
rect 102701 4641 102735 4675
rect 102977 4641 103011 4675
rect 104817 4641 104851 4675
rect 105093 4641 105127 4675
rect 1133 4573 1167 4607
rect 6745 4573 6779 4607
rect 27905 4573 27939 4607
rect 30021 4573 30055 4607
rect 38485 4573 38519 4607
rect 60381 4573 60415 4607
rect 77309 4573 77343 4607
rect 2513 4437 2547 4471
rect 4629 4437 4663 4471
rect 8861 4437 8895 4471
rect 10977 4437 11011 4471
rect 13093 4437 13127 4471
rect 15209 4437 15243 4471
rect 17325 4437 17359 4471
rect 19441 4437 19475 4471
rect 21557 4437 21591 4471
rect 23673 4437 23707 4471
rect 25789 4437 25823 4471
rect 32137 4437 32171 4471
rect 34253 4437 34287 4471
rect 36369 4437 36403 4471
rect 40601 4437 40635 4471
rect 42717 4437 42751 4471
rect 44833 4437 44867 4471
rect 46949 4437 46983 4471
rect 49065 4437 49099 4471
rect 51181 4437 51215 4471
rect 53297 4437 53331 4471
rect 55413 4437 55447 4471
rect 57529 4437 57563 4471
rect 59645 4437 59679 4471
rect 61761 4437 61795 4471
rect 63877 4437 63911 4471
rect 65993 4437 66027 4471
rect 68109 4437 68143 4471
rect 70225 4437 70259 4471
rect 72341 4437 72375 4471
rect 74457 4437 74491 4471
rect 76573 4437 76607 4471
rect 78873 4437 78907 4471
rect 80989 4437 81023 4471
rect 82921 4437 82955 4471
rect 85037 4437 85071 4471
rect 87153 4437 87187 4471
rect 89269 4437 89303 4471
rect 91385 4437 91419 4471
rect 93685 4437 93719 4471
rect 95801 4437 95835 4471
rect 97917 4437 97951 4471
rect 99849 4437 99883 4471
rect 101965 4437 101999 4471
rect 104081 4437 104115 4471
rect 106197 4437 106231 4471
rect 1133 4097 1167 4131
rect 3249 4097 3283 4131
rect 5365 4097 5399 4131
rect 7481 4097 7515 4131
rect 9597 4097 9631 4131
rect 11713 4097 11747 4131
rect 13829 4097 13863 4131
rect 15945 4097 15979 4131
rect 18061 4097 18095 4131
rect 20177 4097 20211 4131
rect 22293 4097 22327 4131
rect 24409 4097 24443 4131
rect 26525 4097 26559 4131
rect 28641 4097 28675 4131
rect 30757 4097 30791 4131
rect 32873 4097 32907 4131
rect 37105 4097 37139 4131
rect 39221 4097 39255 4131
rect 41337 4097 41371 4131
rect 43453 4097 43487 4131
rect 45569 4097 45603 4131
rect 47685 4097 47719 4131
rect 49801 4097 49835 4131
rect 51917 4097 51951 4131
rect 54033 4097 54067 4131
rect 58265 4097 58299 4131
rect 62497 4097 62531 4131
rect 64613 4097 64647 4131
rect 66729 4097 66763 4131
rect 68845 4097 68879 4131
rect 70961 4097 70995 4131
rect 73077 4097 73111 4131
rect 75193 4097 75227 4131
rect 79425 4097 79459 4131
rect 81541 4097 81575 4131
rect 83657 4097 83691 4131
rect 85773 4097 85807 4131
rect 87889 4097 87923 4131
rect 92121 4097 92155 4131
rect 94237 4097 94271 4131
rect 96353 4097 96387 4131
rect 98469 4097 98503 4131
rect 100585 4097 100619 4131
rect 102701 4097 102735 4131
rect 104817 4097 104851 4131
rect 1409 4029 1443 4063
rect 3525 4029 3559 4063
rect 5641 4029 5675 4063
rect 7757 4029 7791 4063
rect 9873 4029 9907 4063
rect 11989 4029 12023 4063
rect 14105 4029 14139 4063
rect 16221 4029 16255 4063
rect 18337 4029 18371 4063
rect 20453 4029 20487 4063
rect 22569 4029 22603 4063
rect 24685 4029 24719 4063
rect 26801 4029 26835 4063
rect 28917 4029 28951 4063
rect 31033 4029 31067 4063
rect 33149 4029 33183 4063
rect 34989 4029 35023 4063
rect 35265 4029 35299 4063
rect 37381 4029 37415 4063
rect 39497 4029 39531 4063
rect 41613 4029 41647 4063
rect 43729 4029 43763 4063
rect 45845 4029 45879 4063
rect 47961 4029 47995 4063
rect 50077 4029 50111 4063
rect 52193 4029 52227 4063
rect 54309 4029 54343 4063
rect 56149 4029 56183 4063
rect 56425 4029 56459 4063
rect 58541 4029 58575 4063
rect 60381 4029 60415 4063
rect 60657 4029 60691 4063
rect 62773 4029 62807 4063
rect 64889 4029 64923 4063
rect 67005 4029 67039 4063
rect 69121 4029 69155 4063
rect 71237 4029 71271 4063
rect 73353 4029 73387 4063
rect 75469 4029 75503 4063
rect 77309 4029 77343 4063
rect 77585 4029 77619 4063
rect 79701 4029 79735 4063
rect 81817 4029 81851 4063
rect 83933 4029 83967 4063
rect 86049 4029 86083 4063
rect 88165 4029 88199 4063
rect 90005 4029 90039 4063
rect 90281 4029 90315 4063
rect 92397 4029 92431 4063
rect 94513 4029 94547 4063
rect 96629 4029 96663 4063
rect 98745 4029 98779 4063
rect 100861 4029 100895 4063
rect 102977 4029 103011 4063
rect 105093 4029 105127 4063
rect 81081 3961 81115 3995
rect 2513 3893 2547 3927
rect 4629 3893 4663 3927
rect 6745 3893 6779 3927
rect 8861 3893 8895 3927
rect 11161 3893 11195 3927
rect 13277 3893 13311 3927
rect 15209 3893 15243 3927
rect 17325 3893 17359 3927
rect 19441 3893 19475 3927
rect 21557 3893 21591 3927
rect 23673 3893 23707 3927
rect 25789 3893 25823 3927
rect 28089 3893 28123 3927
rect 30205 3893 30239 3927
rect 32137 3893 32171 3927
rect 34253 3893 34287 3927
rect 36369 3893 36403 3927
rect 38485 3893 38519 3927
rect 40601 3893 40635 3927
rect 42717 3893 42751 3927
rect 45017 3893 45051 3927
rect 47133 3893 47167 3927
rect 49065 3893 49099 3927
rect 51181 3893 51215 3927
rect 53297 3893 53331 3927
rect 55413 3893 55447 3927
rect 57529 3893 57563 3927
rect 59645 3893 59679 3927
rect 61945 3893 61979 3927
rect 64061 3893 64095 3927
rect 65993 3893 66027 3927
rect 68109 3893 68143 3927
rect 70225 3893 70259 3927
rect 72341 3893 72375 3927
rect 74457 3893 74491 3927
rect 76757 3893 76791 3927
rect 78873 3893 78907 3927
rect 82921 3893 82955 3927
rect 85037 3893 85071 3927
rect 87153 3893 87187 3927
rect 89453 3893 89487 3927
rect 91385 3893 91419 3927
rect 93501 3893 93535 3927
rect 95801 3893 95835 3927
rect 97917 3893 97951 3927
rect 99849 3893 99883 3927
rect 101965 3893 101999 3927
rect 104081 3893 104115 3927
rect 106197 3893 106231 3927
rect 2513 3689 2547 3723
rect 10977 3689 11011 3723
rect 13093 3689 13127 3723
rect 15209 3689 15243 3723
rect 17325 3689 17359 3723
rect 27905 3689 27939 3723
rect 30021 3689 30055 3723
rect 32137 3689 32171 3723
rect 34253 3689 34287 3723
rect 44833 3689 44867 3723
rect 46949 3689 46983 3723
rect 49065 3689 49099 3723
rect 51181 3689 51215 3723
rect 63877 3689 63911 3723
rect 65993 3689 66027 3723
rect 68109 3689 68143 3723
rect 78689 3689 78723 3723
rect 80805 3689 80839 3723
rect 82921 3689 82955 3723
rect 85037 3689 85071 3723
rect 95617 3689 95651 3723
rect 99849 3689 99883 3723
rect 101965 3689 101999 3723
rect 1133 3553 1167 3587
rect 3249 3553 3283 3587
rect 5365 3553 5399 3587
rect 7481 3553 7515 3587
rect 9597 3553 9631 3587
rect 11713 3553 11747 3587
rect 13829 3553 13863 3587
rect 15945 3553 15979 3587
rect 18061 3553 18095 3587
rect 20177 3553 20211 3587
rect 22293 3553 22327 3587
rect 24409 3553 24443 3587
rect 26525 3553 26559 3587
rect 28641 3553 28675 3587
rect 30757 3553 30791 3587
rect 32873 3553 32907 3587
rect 34989 3553 35023 3587
rect 37105 3553 37139 3587
rect 39221 3553 39255 3587
rect 39497 3553 39531 3587
rect 41337 3553 41371 3587
rect 43453 3553 43487 3587
rect 45569 3553 45603 3587
rect 47685 3553 47719 3587
rect 49801 3553 49835 3587
rect 51917 3553 51951 3587
rect 54033 3553 54067 3587
rect 56149 3553 56183 3587
rect 58265 3553 58299 3587
rect 60381 3553 60415 3587
rect 62497 3553 62531 3587
rect 64613 3553 64647 3587
rect 66729 3553 66763 3587
rect 68845 3553 68879 3587
rect 70961 3553 70995 3587
rect 73077 3553 73111 3587
rect 75193 3553 75227 3587
rect 79425 3553 79459 3587
rect 81541 3553 81575 3587
rect 83657 3553 83691 3587
rect 85773 3553 85807 3587
rect 87889 3553 87923 3587
rect 90005 3553 90039 3587
rect 92121 3553 92155 3587
rect 94237 3553 94271 3587
rect 96353 3553 96387 3587
rect 98469 3553 98503 3587
rect 100585 3553 100619 3587
rect 102701 3553 102735 3587
rect 104817 3553 104851 3587
rect 1409 3485 1443 3519
rect 3525 3485 3559 3519
rect 4629 3485 4663 3519
rect 5641 3485 5675 3519
rect 6745 3485 6779 3519
rect 7757 3485 7791 3519
rect 8861 3485 8895 3519
rect 9873 3485 9907 3519
rect 11989 3485 12023 3519
rect 14105 3485 14139 3519
rect 16221 3485 16255 3519
rect 18337 3485 18371 3519
rect 19441 3485 19475 3519
rect 20453 3485 20487 3519
rect 21557 3485 21591 3519
rect 22569 3485 22603 3519
rect 23673 3485 23707 3519
rect 24685 3485 24719 3519
rect 25789 3485 25823 3519
rect 26801 3485 26835 3519
rect 28917 3485 28951 3519
rect 31033 3485 31067 3519
rect 33149 3485 33183 3519
rect 35265 3485 35299 3519
rect 36369 3485 36403 3519
rect 37381 3485 37415 3519
rect 38485 3485 38519 3519
rect 40693 3485 40727 3519
rect 41613 3485 41647 3519
rect 42717 3485 42751 3519
rect 43729 3485 43763 3519
rect 45845 3485 45879 3519
rect 47961 3485 47995 3519
rect 50077 3485 50111 3519
rect 52193 3485 52227 3519
rect 53297 3485 53331 3519
rect 54309 3485 54343 3519
rect 55413 3485 55447 3519
rect 56425 3485 56459 3519
rect 57529 3485 57563 3519
rect 58541 3485 58575 3519
rect 59645 3485 59679 3519
rect 60657 3485 60691 3519
rect 61761 3485 61795 3519
rect 62773 3485 62807 3519
rect 64889 3485 64923 3519
rect 67005 3485 67039 3519
rect 69121 3485 69155 3519
rect 70225 3485 70259 3519
rect 71237 3485 71271 3519
rect 72341 3485 72375 3519
rect 73353 3485 73387 3519
rect 74457 3485 74491 3519
rect 75469 3485 75503 3519
rect 76573 3485 76607 3519
rect 77309 3485 77343 3519
rect 77585 3485 77619 3519
rect 79701 3485 79735 3519
rect 81817 3485 81851 3519
rect 83933 3485 83967 3519
rect 86049 3485 86083 3519
rect 87153 3485 87187 3519
rect 88165 3485 88199 3519
rect 89269 3485 89303 3519
rect 90281 3485 90315 3519
rect 91385 3485 91419 3519
rect 92397 3485 92431 3519
rect 93501 3485 93535 3519
rect 94513 3485 94547 3519
rect 96629 3485 96663 3519
rect 97733 3485 97767 3519
rect 98745 3485 98779 3519
rect 100861 3485 100895 3519
rect 102977 3485 103011 3519
rect 104081 3485 104115 3519
rect 105093 3485 105127 3519
rect 106197 3485 106231 3519
rect 1225 3145 1259 3179
rect 41429 3145 41463 3179
rect 77401 3145 77435 3179
rect 87981 3145 88015 3179
rect 50721 3009 50755 3043
rect 51917 3009 51951 3043
rect 1317 2941 1351 2975
rect 3249 2941 3283 2975
rect 3433 2941 3467 2975
rect 5365 2941 5399 2975
rect 5549 2941 5583 2975
rect 7481 2941 7515 2975
rect 7665 2941 7699 2975
rect 9597 2941 9631 2975
rect 9781 2941 9815 2975
rect 11713 2941 11747 2975
rect 11897 2941 11931 2975
rect 13829 2941 13863 2975
rect 14013 2941 14047 2975
rect 15945 2941 15979 2975
rect 18061 2941 18095 2975
rect 18245 2941 18279 2975
rect 20177 2941 20211 2975
rect 20361 2941 20395 2975
rect 22293 2941 22327 2975
rect 22477 2941 22511 2975
rect 24409 2941 24443 2975
rect 24593 2941 24627 2975
rect 26525 2941 26559 2975
rect 26709 2941 26743 2975
rect 28641 2941 28675 2975
rect 28825 2941 28859 2975
rect 30757 2941 30791 2975
rect 30941 2941 30975 2975
rect 32873 2941 32907 2975
rect 34989 2941 35023 2975
rect 35173 2941 35207 2975
rect 37105 2941 37139 2975
rect 37289 2941 37323 2975
rect 39221 2941 39255 2975
rect 39405 2941 39439 2975
rect 41521 2941 41555 2975
rect 43453 2941 43487 2975
rect 43637 2941 43671 2975
rect 45569 2941 45603 2975
rect 45753 2941 45787 2975
rect 47685 2941 47719 2975
rect 47869 2941 47903 2975
rect 49801 2941 49835 2975
rect 52101 2941 52135 2975
rect 54033 2941 54067 2975
rect 54217 2941 54251 2975
rect 56149 2941 56183 2975
rect 56333 2941 56367 2975
rect 58265 2941 58299 2975
rect 58449 2941 58483 2975
rect 60381 2941 60415 2975
rect 60565 2941 60599 2975
rect 62497 2941 62531 2975
rect 62681 2941 62715 2975
rect 64613 2941 64647 2975
rect 64797 2941 64831 2975
rect 66729 2941 66763 2975
rect 68845 2941 68879 2975
rect 69029 2941 69063 2975
rect 70961 2941 70995 2975
rect 71145 2941 71179 2975
rect 73077 2941 73111 2975
rect 73261 2941 73295 2975
rect 75193 2941 75227 2975
rect 75377 2941 75411 2975
rect 77493 2941 77527 2975
rect 79425 2941 79459 2975
rect 79609 2941 79643 2975
rect 81541 2941 81575 2975
rect 81725 2941 81759 2975
rect 83657 2941 83691 2975
rect 85773 2941 85807 2975
rect 85957 2941 85991 2975
rect 88073 2941 88107 2975
rect 90005 2941 90039 2975
rect 90189 2941 90223 2975
rect 92121 2941 92155 2975
rect 92305 2941 92339 2975
rect 94237 2941 94271 2975
rect 94421 2941 94455 2975
rect 96353 2941 96387 2975
rect 96537 2941 96571 2975
rect 98469 2941 98503 2975
rect 98653 2941 98687 2975
rect 100585 2941 100619 2975
rect 100769 2941 100803 2975
rect 102701 2941 102735 2975
rect 102885 2941 102919 2975
rect 104817 2941 104851 2975
rect 105001 2941 105035 2975
rect 16129 2873 16163 2907
rect 33057 2873 33091 2907
rect 49985 2873 50019 2907
rect 50721 2873 50755 2907
rect 66913 2873 66947 2907
rect 83841 2873 83875 2907
rect 5549 2601 5583 2635
rect 20361 2601 20395 2635
rect 22477 2601 22511 2635
rect 30941 2601 30975 2635
rect 35173 2601 35207 2635
rect 41521 2601 41555 2635
rect 60565 2601 60599 2635
rect 71145 2601 71179 2635
rect 77493 2601 77527 2635
rect 96537 2601 96571 2635
rect 102885 2601 102919 2635
rect 7573 2533 7607 2567
rect 9873 2533 9907 2567
rect 11805 2533 11839 2567
rect 11989 2533 12023 2567
rect 13921 2533 13955 2567
rect 22385 2533 22419 2567
rect 24501 2533 24535 2567
rect 32965 2533 32999 2567
rect 37197 2533 37231 2567
rect 43545 2533 43579 2567
rect 45845 2533 45879 2567
rect 47777 2533 47811 2567
rect 56425 2533 56459 2567
rect 58357 2533 58391 2567
rect 58541 2533 58575 2567
rect 60473 2533 60507 2567
rect 62589 2533 62623 2567
rect 73169 2533 73203 2567
rect 79517 2533 79551 2567
rect 88165 2533 88199 2567
rect 90097 2533 90131 2567
rect 92397 2533 92431 2567
rect 94329 2533 94363 2567
rect 94513 2533 94547 2567
rect 96445 2533 96479 2567
rect 98561 2533 98595 2567
rect 102609 2533 102643 2567
rect 102793 2533 102827 2567
rect 104909 2533 104943 2567
rect 105093 2533 105127 2567
rect 1225 2465 1259 2499
rect 1409 2465 1443 2499
rect 3341 2465 3375 2499
rect 5457 2465 5491 2499
rect 9689 2465 9723 2499
rect 16037 2465 16071 2499
rect 18153 2465 18187 2499
rect 18337 2465 18371 2499
rect 20269 2465 20303 2499
rect 26617 2465 26651 2499
rect 28733 2465 28767 2499
rect 28917 2465 28951 2499
rect 30849 2465 30883 2499
rect 33149 2465 33183 2499
rect 35081 2465 35115 2499
rect 39313 2465 39347 2499
rect 41429 2465 41463 2499
rect 45661 2465 45695 2499
rect 47961 2465 47995 2499
rect 49893 2465 49927 2499
rect 52009 2465 52043 2499
rect 52193 2465 52227 2499
rect 54125 2465 54159 2499
rect 56241 2465 56275 2499
rect 64705 2465 64739 2499
rect 64889 2465 64923 2499
rect 66821 2465 66855 2499
rect 68937 2465 68971 2499
rect 69121 2465 69155 2499
rect 71053 2465 71087 2499
rect 75285 2465 75319 2499
rect 77401 2465 77435 2499
rect 79701 2465 79735 2499
rect 81633 2465 81667 2499
rect 81817 2465 81851 2499
rect 83749 2465 83783 2499
rect 85865 2465 85899 2499
rect 87981 2465 88015 2499
rect 92213 2465 92247 2499
rect 100677 2465 100711 2499
rect 7757 2397 7791 2431
rect 14105 2397 14139 2431
rect 24685 2397 24719 2431
rect 26801 2397 26835 2431
rect 37381 2397 37415 2431
rect 43729 2397 43763 2431
rect 54309 2397 54343 2431
rect 62773 2397 62807 2431
rect 73353 2397 73387 2431
rect 86049 2397 86083 2431
rect 90281 2397 90315 2431
rect 98745 2397 98779 2431
rect 16221 2329 16255 2363
rect 39497 2329 39531 2363
rect 50077 2329 50111 2363
rect 67005 2329 67039 2363
rect 83933 2329 83967 2363
rect 100861 2329 100895 2363
rect 102609 2329 102643 2363
rect 3433 2261 3467 2295
rect 75377 2261 75411 2295
rect 1133 1921 1167 1955
rect 3249 1921 3283 1955
rect 3525 1921 3559 1955
rect 5365 1921 5399 1955
rect 5641 1921 5675 1955
rect 7481 1921 7515 1955
rect 7757 1921 7791 1955
rect 9597 1921 9631 1955
rect 9873 1921 9907 1955
rect 11713 1921 11747 1955
rect 11989 1921 12023 1955
rect 13829 1921 13863 1955
rect 14105 1921 14139 1955
rect 15945 1921 15979 1955
rect 16221 1921 16255 1955
rect 18061 1921 18095 1955
rect 18337 1921 18371 1955
rect 20177 1921 20211 1955
rect 20453 1921 20487 1955
rect 22293 1921 22327 1955
rect 24409 1921 24443 1955
rect 24685 1921 24719 1955
rect 26525 1921 26559 1955
rect 26801 1921 26835 1955
rect 28641 1921 28675 1955
rect 28917 1921 28951 1955
rect 30757 1921 30791 1955
rect 31033 1921 31067 1955
rect 32873 1921 32907 1955
rect 33149 1921 33183 1955
rect 35265 1921 35299 1955
rect 37105 1921 37139 1955
rect 37381 1921 37415 1955
rect 39221 1921 39255 1955
rect 39497 1921 39531 1955
rect 41337 1921 41371 1955
rect 41613 1921 41647 1955
rect 43453 1921 43487 1955
rect 43729 1921 43763 1955
rect 45569 1921 45603 1955
rect 45845 1921 45879 1955
rect 47685 1921 47719 1955
rect 47961 1921 47995 1955
rect 49801 1921 49835 1955
rect 50077 1921 50111 1955
rect 51917 1921 51951 1955
rect 52193 1921 52227 1955
rect 54033 1921 54067 1955
rect 54309 1921 54343 1955
rect 56149 1921 56183 1955
rect 56425 1921 56459 1955
rect 58265 1921 58299 1955
rect 58541 1921 58575 1955
rect 60381 1921 60415 1955
rect 62497 1921 62531 1955
rect 62773 1921 62807 1955
rect 64613 1921 64647 1955
rect 64889 1921 64923 1955
rect 66729 1921 66763 1955
rect 67005 1921 67039 1955
rect 68845 1921 68879 1955
rect 69121 1921 69155 1955
rect 70961 1921 70995 1955
rect 71237 1921 71271 1955
rect 73077 1921 73111 1955
rect 73353 1921 73387 1955
rect 75193 1921 75227 1955
rect 75469 1921 75503 1955
rect 77585 1921 77619 1955
rect 79425 1921 79459 1955
rect 79701 1921 79735 1955
rect 81541 1921 81575 1955
rect 81817 1921 81851 1955
rect 83657 1921 83691 1955
rect 83933 1921 83967 1955
rect 85773 1921 85807 1955
rect 86049 1921 86083 1955
rect 87889 1921 87923 1955
rect 88165 1921 88199 1955
rect 90005 1921 90039 1955
rect 90281 1921 90315 1955
rect 92121 1921 92155 1955
rect 92397 1921 92431 1955
rect 94237 1921 94271 1955
rect 94513 1921 94547 1955
rect 96353 1921 96387 1955
rect 96629 1921 96663 1955
rect 98469 1921 98503 1955
rect 98745 1921 98779 1955
rect 100585 1921 100619 1955
rect 100861 1921 100895 1955
rect 102701 1921 102735 1955
rect 102977 1921 103011 1955
rect 104817 1921 104851 1955
rect 1409 1853 1443 1887
rect 22569 1853 22603 1887
rect 34989 1853 35023 1887
rect 60657 1853 60691 1887
rect 77309 1853 77343 1887
rect 105093 1853 105127 1887
rect 81081 1785 81115 1819
rect 2513 1717 2547 1751
rect 4629 1717 4663 1751
rect 6745 1717 6779 1751
rect 8861 1717 8895 1751
rect 11161 1717 11195 1751
rect 13277 1717 13311 1751
rect 15209 1717 15243 1751
rect 17325 1717 17359 1751
rect 19441 1717 19475 1751
rect 21557 1717 21591 1751
rect 23673 1717 23707 1751
rect 25789 1717 25823 1751
rect 28089 1717 28123 1751
rect 30205 1717 30239 1751
rect 32137 1717 32171 1751
rect 34253 1717 34287 1751
rect 36369 1717 36403 1751
rect 38485 1717 38519 1751
rect 40601 1717 40635 1751
rect 42717 1717 42751 1751
rect 45017 1717 45051 1751
rect 47133 1717 47167 1751
rect 49065 1717 49099 1751
rect 51181 1717 51215 1751
rect 53297 1717 53331 1751
rect 55413 1717 55447 1751
rect 57529 1717 57563 1751
rect 59645 1717 59679 1751
rect 61945 1717 61979 1751
rect 64061 1717 64095 1751
rect 65993 1717 66027 1751
rect 68109 1717 68143 1751
rect 70225 1717 70259 1751
rect 72341 1717 72375 1751
rect 74457 1717 74491 1751
rect 76573 1717 76607 1751
rect 78873 1717 78907 1751
rect 82921 1717 82955 1751
rect 85037 1717 85071 1751
rect 87153 1717 87187 1751
rect 89269 1717 89303 1751
rect 91385 1717 91419 1751
rect 93501 1717 93535 1751
rect 95801 1717 95835 1751
rect 97917 1717 97951 1751
rect 99849 1717 99883 1751
rect 101965 1717 101999 1751
rect 104081 1717 104115 1751
rect 106197 1717 106231 1751
rect 2513 1513 2547 1547
rect 8861 1513 8895 1547
rect 10977 1513 11011 1547
rect 15209 1513 15243 1547
rect 25789 1513 25823 1547
rect 27905 1513 27939 1547
rect 32137 1513 32171 1547
rect 42717 1513 42751 1547
rect 44833 1513 44867 1547
rect 49065 1513 49099 1547
rect 59645 1513 59679 1547
rect 65993 1513 66027 1547
rect 76573 1513 76607 1547
rect 78689 1513 78723 1547
rect 82921 1513 82955 1547
rect 93501 1513 93535 1547
rect 95617 1513 95651 1547
rect 99849 1513 99883 1547
rect 1133 1377 1167 1411
rect 1409 1377 1443 1411
rect 3249 1377 3283 1411
rect 3525 1377 3559 1411
rect 5365 1377 5399 1411
rect 5641 1377 5675 1411
rect 7481 1377 7515 1411
rect 7757 1377 7791 1411
rect 9597 1377 9631 1411
rect 9873 1377 9907 1411
rect 11713 1377 11747 1411
rect 11989 1377 12023 1411
rect 13829 1377 13863 1411
rect 14105 1377 14139 1411
rect 15945 1377 15979 1411
rect 16221 1377 16255 1411
rect 18061 1377 18095 1411
rect 18337 1377 18371 1411
rect 20177 1377 20211 1411
rect 20453 1377 20487 1411
rect 22293 1377 22327 1411
rect 22569 1377 22603 1411
rect 24409 1377 24443 1411
rect 24685 1377 24719 1411
rect 26525 1377 26559 1411
rect 26801 1377 26835 1411
rect 28641 1377 28675 1411
rect 28917 1377 28951 1411
rect 30757 1377 30791 1411
rect 31033 1377 31067 1411
rect 32873 1377 32907 1411
rect 33149 1377 33183 1411
rect 34989 1377 35023 1411
rect 35265 1377 35299 1411
rect 37105 1377 37139 1411
rect 37381 1377 37415 1411
rect 39221 1377 39255 1411
rect 39497 1377 39531 1411
rect 41337 1377 41371 1411
rect 41613 1377 41647 1411
rect 43453 1377 43487 1411
rect 43729 1377 43763 1411
rect 45569 1377 45603 1411
rect 45845 1377 45879 1411
rect 47685 1377 47719 1411
rect 47961 1377 47995 1411
rect 49801 1377 49835 1411
rect 50077 1377 50111 1411
rect 51917 1377 51951 1411
rect 52193 1377 52227 1411
rect 54033 1377 54067 1411
rect 54309 1377 54343 1411
rect 56149 1377 56183 1411
rect 56425 1377 56459 1411
rect 58265 1377 58299 1411
rect 58541 1377 58575 1411
rect 60381 1377 60415 1411
rect 60657 1377 60691 1411
rect 62497 1377 62531 1411
rect 62773 1377 62807 1411
rect 64613 1377 64647 1411
rect 64889 1377 64923 1411
rect 66729 1377 66763 1411
rect 67005 1377 67039 1411
rect 68845 1377 68879 1411
rect 69121 1377 69155 1411
rect 70961 1377 70995 1411
rect 71237 1377 71271 1411
rect 73077 1377 73111 1411
rect 73353 1377 73387 1411
rect 75193 1377 75227 1411
rect 75469 1377 75503 1411
rect 77309 1377 77343 1411
rect 77585 1377 77619 1411
rect 79425 1377 79459 1411
rect 79701 1377 79735 1411
rect 81541 1377 81575 1411
rect 81817 1377 81851 1411
rect 83657 1377 83691 1411
rect 83933 1377 83967 1411
rect 85773 1377 85807 1411
rect 86049 1377 86083 1411
rect 87889 1377 87923 1411
rect 88165 1377 88199 1411
rect 90005 1377 90039 1411
rect 90281 1377 90315 1411
rect 92121 1377 92155 1411
rect 92397 1377 92431 1411
rect 94237 1377 94271 1411
rect 94513 1377 94547 1411
rect 96353 1377 96387 1411
rect 96629 1377 96663 1411
rect 98469 1377 98503 1411
rect 98745 1377 98779 1411
rect 100585 1377 100619 1411
rect 100861 1377 100895 1411
rect 102701 1377 102735 1411
rect 102977 1377 103011 1411
rect 104817 1377 104851 1411
rect 105093 1377 105127 1411
rect 4629 1173 4663 1207
rect 6745 1173 6779 1207
rect 13093 1173 13127 1207
rect 17325 1173 17359 1207
rect 19441 1173 19475 1207
rect 21557 1173 21591 1207
rect 23673 1173 23707 1207
rect 30021 1173 30055 1207
rect 34253 1173 34287 1207
rect 36369 1173 36403 1207
rect 38485 1173 38519 1207
rect 40601 1173 40635 1207
rect 46949 1173 46983 1207
rect 51181 1173 51215 1207
rect 53297 1173 53331 1207
rect 55413 1173 55447 1207
rect 57529 1173 57563 1207
rect 61761 1173 61795 1207
rect 63877 1173 63911 1207
rect 68109 1173 68143 1207
rect 70225 1173 70259 1207
rect 72341 1173 72375 1207
rect 74457 1173 74491 1207
rect 80805 1173 80839 1207
rect 85037 1173 85071 1207
rect 87153 1173 87187 1207
rect 89269 1173 89303 1207
rect 91385 1173 91419 1207
rect 97733 1173 97767 1207
rect 101965 1173 101999 1207
rect 104081 1173 104115 1207
rect 106197 1173 106231 1207
<< metal1 >>
rect 1104 7642 106904 7664
rect 1104 7590 4042 7642
rect 4094 7590 4106 7642
rect 4158 7590 4170 7642
rect 4222 7590 4234 7642
rect 4286 7590 34762 7642
rect 34814 7590 34826 7642
rect 34878 7590 34890 7642
rect 34942 7590 34954 7642
rect 35006 7590 65482 7642
rect 65534 7590 65546 7642
rect 65598 7590 65610 7642
rect 65662 7590 65674 7642
rect 65726 7590 96202 7642
rect 96254 7590 96266 7642
rect 96318 7590 96330 7642
rect 96382 7590 96394 7642
rect 96446 7590 106904 7642
rect 1104 7568 106904 7590
rect 1118 7324 1124 7336
rect 1079 7296 1124 7324
rect 1118 7284 1124 7296
rect 1176 7284 1182 7336
rect 1397 7327 1455 7333
rect 1397 7324 1409 7327
rect 1228 7296 1409 7324
rect 1228 7256 1256 7296
rect 1397 7293 1409 7296
rect 1443 7293 1455 7327
rect 3234 7324 3240 7336
rect 3195 7296 3240 7324
rect 1397 7287 1455 7293
rect 3234 7284 3240 7296
rect 3292 7284 3298 7336
rect 3510 7324 3516 7336
rect 3471 7296 3516 7324
rect 3510 7284 3516 7296
rect 3568 7284 3574 7336
rect 5258 7284 5264 7336
rect 5316 7324 5322 7336
rect 5353 7327 5411 7333
rect 5353 7324 5365 7327
rect 5316 7296 5365 7324
rect 5316 7284 5322 7296
rect 5353 7293 5365 7296
rect 5399 7293 5411 7327
rect 5626 7324 5632 7336
rect 5587 7296 5632 7324
rect 5353 7287 5411 7293
rect 5626 7284 5632 7296
rect 5684 7284 5690 7336
rect 7374 7284 7380 7336
rect 7432 7324 7438 7336
rect 7469 7327 7527 7333
rect 7469 7324 7481 7327
rect 7432 7296 7481 7324
rect 7432 7284 7438 7296
rect 7469 7293 7481 7296
rect 7515 7293 7527 7327
rect 7742 7324 7748 7336
rect 7703 7296 7748 7324
rect 7469 7287 7527 7293
rect 7742 7284 7748 7296
rect 7800 7284 7806 7336
rect 9582 7324 9588 7336
rect 9543 7296 9588 7324
rect 9582 7284 9588 7296
rect 9640 7284 9646 7336
rect 9858 7324 9864 7336
rect 9819 7296 9864 7324
rect 9858 7284 9864 7296
rect 9916 7284 9922 7336
rect 11698 7324 11704 7336
rect 11659 7296 11704 7324
rect 11698 7284 11704 7296
rect 11756 7284 11762 7336
rect 11974 7324 11980 7336
rect 11935 7296 11980 7324
rect 11974 7284 11980 7296
rect 12032 7284 12038 7336
rect 13814 7324 13820 7336
rect 13775 7296 13820 7324
rect 13814 7284 13820 7296
rect 13872 7284 13878 7336
rect 14090 7324 14096 7336
rect 14051 7296 14096 7324
rect 14090 7284 14096 7296
rect 14148 7284 14154 7336
rect 15930 7324 15936 7336
rect 15891 7296 15936 7324
rect 15930 7284 15936 7296
rect 15988 7284 15994 7336
rect 16206 7324 16212 7336
rect 16167 7296 16212 7324
rect 16206 7284 16212 7296
rect 16264 7284 16270 7336
rect 18046 7324 18052 7336
rect 18007 7296 18052 7324
rect 18046 7284 18052 7296
rect 18104 7284 18110 7336
rect 18322 7324 18328 7336
rect 18283 7296 18328 7324
rect 18322 7284 18328 7296
rect 18380 7284 18386 7336
rect 20070 7284 20076 7336
rect 20128 7324 20134 7336
rect 20165 7327 20223 7333
rect 20165 7324 20177 7327
rect 20128 7296 20177 7324
rect 20128 7284 20134 7296
rect 20165 7293 20177 7296
rect 20211 7293 20223 7327
rect 20438 7324 20444 7336
rect 20399 7296 20444 7324
rect 20165 7287 20223 7293
rect 20438 7284 20444 7296
rect 20496 7284 20502 7336
rect 22186 7284 22192 7336
rect 22244 7324 22250 7336
rect 22281 7327 22339 7333
rect 22281 7324 22293 7327
rect 22244 7296 22293 7324
rect 22244 7284 22250 7296
rect 22281 7293 22293 7296
rect 22327 7293 22339 7327
rect 22554 7324 22560 7336
rect 22515 7296 22560 7324
rect 22281 7287 22339 7293
rect 22554 7284 22560 7296
rect 22612 7284 22618 7336
rect 24394 7324 24400 7336
rect 24355 7296 24400 7324
rect 24394 7284 24400 7296
rect 24452 7284 24458 7336
rect 24670 7324 24676 7336
rect 24631 7296 24676 7324
rect 24670 7284 24676 7296
rect 24728 7284 24734 7336
rect 26510 7324 26516 7336
rect 26471 7296 26516 7324
rect 26510 7284 26516 7296
rect 26568 7284 26574 7336
rect 26786 7324 26792 7336
rect 26747 7296 26792 7324
rect 26786 7284 26792 7296
rect 26844 7284 26850 7336
rect 28626 7324 28632 7336
rect 28587 7296 28632 7324
rect 28626 7284 28632 7296
rect 28684 7284 28690 7336
rect 28902 7324 28908 7336
rect 28863 7296 28908 7324
rect 28902 7284 28908 7296
rect 28960 7284 28966 7336
rect 30742 7324 30748 7336
rect 30703 7296 30748 7324
rect 30742 7284 30748 7296
rect 30800 7284 30806 7336
rect 31018 7324 31024 7336
rect 30979 7296 31024 7324
rect 31018 7284 31024 7296
rect 31076 7284 31082 7336
rect 32858 7324 32864 7336
rect 32819 7296 32864 7324
rect 32858 7284 32864 7296
rect 32916 7284 32922 7336
rect 33134 7324 33140 7336
rect 33095 7296 33140 7324
rect 33134 7284 33140 7296
rect 33192 7284 33198 7336
rect 34977 7327 35035 7333
rect 34977 7293 34989 7327
rect 35023 7324 35035 7327
rect 35066 7324 35072 7336
rect 35023 7296 35072 7324
rect 35023 7293 35035 7296
rect 34977 7287 35035 7293
rect 35066 7284 35072 7296
rect 35124 7284 35130 7336
rect 35250 7324 35256 7336
rect 35211 7296 35256 7324
rect 35250 7284 35256 7296
rect 35308 7284 35314 7336
rect 37090 7324 37096 7336
rect 37051 7296 37096 7324
rect 37090 7284 37096 7296
rect 37148 7284 37154 7336
rect 37366 7324 37372 7336
rect 37327 7296 37372 7324
rect 37366 7284 37372 7296
rect 37424 7284 37430 7336
rect 39206 7324 39212 7336
rect 39167 7296 39212 7324
rect 39206 7284 39212 7296
rect 39264 7284 39270 7336
rect 39482 7324 39488 7336
rect 39443 7296 39488 7324
rect 39482 7284 39488 7296
rect 39540 7284 39546 7336
rect 41230 7284 41236 7336
rect 41288 7324 41294 7336
rect 41325 7327 41383 7333
rect 41325 7324 41337 7327
rect 41288 7296 41337 7324
rect 41288 7284 41294 7296
rect 41325 7293 41337 7296
rect 41371 7293 41383 7327
rect 41598 7324 41604 7336
rect 41559 7296 41604 7324
rect 41325 7287 41383 7293
rect 41598 7284 41604 7296
rect 41656 7284 41662 7336
rect 43438 7324 43444 7336
rect 43399 7296 43444 7324
rect 43438 7284 43444 7296
rect 43496 7284 43502 7336
rect 43714 7324 43720 7336
rect 43675 7296 43720 7324
rect 43714 7284 43720 7296
rect 43772 7284 43778 7336
rect 45554 7324 45560 7336
rect 45515 7296 45560 7324
rect 45554 7284 45560 7296
rect 45612 7284 45618 7336
rect 45830 7324 45836 7336
rect 45791 7296 45836 7324
rect 45830 7284 45836 7296
rect 45888 7284 45894 7336
rect 47670 7324 47676 7336
rect 47631 7296 47676 7324
rect 47670 7284 47676 7296
rect 47728 7284 47734 7336
rect 47946 7324 47952 7336
rect 47907 7296 47952 7324
rect 47946 7284 47952 7296
rect 48004 7284 48010 7336
rect 49786 7324 49792 7336
rect 49747 7296 49792 7324
rect 49786 7284 49792 7296
rect 49844 7284 49850 7336
rect 50065 7327 50123 7333
rect 50065 7293 50077 7327
rect 50111 7324 50123 7327
rect 51166 7324 51172 7336
rect 50111 7296 51172 7324
rect 50111 7293 50123 7296
rect 50065 7287 50123 7293
rect 51166 7284 51172 7296
rect 51224 7284 51230 7336
rect 51902 7324 51908 7336
rect 51863 7296 51908 7324
rect 51902 7284 51908 7296
rect 51960 7284 51966 7336
rect 52178 7324 52184 7336
rect 52139 7296 52184 7324
rect 52178 7284 52184 7296
rect 52236 7284 52242 7336
rect 54018 7324 54024 7336
rect 53979 7296 54024 7324
rect 54018 7284 54024 7296
rect 54076 7284 54082 7336
rect 54294 7324 54300 7336
rect 54255 7296 54300 7324
rect 54294 7284 54300 7296
rect 54352 7284 54358 7336
rect 56042 7284 56048 7336
rect 56100 7324 56106 7336
rect 56137 7327 56195 7333
rect 56137 7324 56149 7327
rect 56100 7296 56149 7324
rect 56100 7284 56106 7296
rect 56137 7293 56149 7296
rect 56183 7293 56195 7327
rect 56410 7324 56416 7336
rect 56371 7296 56416 7324
rect 56137 7287 56195 7293
rect 56410 7284 56416 7296
rect 56468 7284 56474 7336
rect 58158 7284 58164 7336
rect 58216 7324 58222 7336
rect 58253 7327 58311 7333
rect 58253 7324 58265 7327
rect 58216 7296 58265 7324
rect 58216 7284 58222 7296
rect 58253 7293 58265 7296
rect 58299 7293 58311 7327
rect 58526 7324 58532 7336
rect 58487 7296 58532 7324
rect 58253 7287 58311 7293
rect 58526 7284 58532 7296
rect 58584 7284 58590 7336
rect 60366 7284 60372 7336
rect 60424 7324 60430 7336
rect 60642 7324 60648 7336
rect 60424 7296 60469 7324
rect 60603 7296 60648 7324
rect 60424 7284 60430 7296
rect 60642 7284 60648 7296
rect 60700 7284 60706 7336
rect 62482 7324 62488 7336
rect 62443 7296 62488 7324
rect 62482 7284 62488 7296
rect 62540 7284 62546 7336
rect 62758 7324 62764 7336
rect 62719 7296 62764 7324
rect 62758 7284 62764 7296
rect 62816 7284 62822 7336
rect 64598 7324 64604 7336
rect 64559 7296 64604 7324
rect 64598 7284 64604 7296
rect 64656 7284 64662 7336
rect 64874 7324 64880 7336
rect 64835 7296 64880 7324
rect 64874 7284 64880 7296
rect 64932 7284 64938 7336
rect 66714 7324 66720 7336
rect 66675 7296 66720 7324
rect 66714 7284 66720 7296
rect 66772 7284 66778 7336
rect 66990 7324 66996 7336
rect 66951 7296 66996 7324
rect 66990 7284 66996 7296
rect 67048 7284 67054 7336
rect 68830 7324 68836 7336
rect 68791 7296 68836 7324
rect 68830 7284 68836 7296
rect 68888 7284 68894 7336
rect 69106 7324 69112 7336
rect 69067 7296 69112 7324
rect 69106 7284 69112 7296
rect 69164 7284 69170 7336
rect 70854 7284 70860 7336
rect 70912 7324 70918 7336
rect 70949 7327 71007 7333
rect 70949 7324 70961 7327
rect 70912 7296 70961 7324
rect 70912 7284 70918 7296
rect 70949 7293 70961 7296
rect 70995 7293 71007 7327
rect 71222 7324 71228 7336
rect 71183 7296 71228 7324
rect 70949 7287 71007 7293
rect 71222 7284 71228 7296
rect 71280 7284 71286 7336
rect 72970 7284 72976 7336
rect 73028 7324 73034 7336
rect 73065 7327 73123 7333
rect 73065 7324 73077 7327
rect 73028 7296 73077 7324
rect 73028 7284 73034 7296
rect 73065 7293 73077 7296
rect 73111 7293 73123 7327
rect 73338 7324 73344 7336
rect 73299 7296 73344 7324
rect 73065 7287 73123 7293
rect 73338 7284 73344 7296
rect 73396 7284 73402 7336
rect 75086 7284 75092 7336
rect 75144 7324 75150 7336
rect 75181 7327 75239 7333
rect 75181 7324 75193 7327
rect 75144 7296 75193 7324
rect 75144 7284 75150 7296
rect 75181 7293 75193 7296
rect 75227 7293 75239 7327
rect 75454 7324 75460 7336
rect 75415 7296 75460 7324
rect 75181 7287 75239 7293
rect 75454 7284 75460 7296
rect 75512 7284 75518 7336
rect 77202 7284 77208 7336
rect 77260 7324 77266 7336
rect 77297 7327 77355 7333
rect 77297 7324 77309 7327
rect 77260 7296 77309 7324
rect 77260 7284 77266 7296
rect 77297 7293 77309 7296
rect 77343 7293 77355 7327
rect 77570 7324 77576 7336
rect 77531 7296 77576 7324
rect 77297 7287 77355 7293
rect 77570 7284 77576 7296
rect 77628 7284 77634 7336
rect 79318 7284 79324 7336
rect 79376 7324 79382 7336
rect 79413 7327 79471 7333
rect 79413 7324 79425 7327
rect 79376 7296 79425 7324
rect 79376 7284 79382 7296
rect 79413 7293 79425 7296
rect 79459 7293 79471 7327
rect 79686 7324 79692 7336
rect 79647 7296 79692 7324
rect 79413 7287 79471 7293
rect 79686 7284 79692 7296
rect 79744 7284 79750 7336
rect 81434 7284 81440 7336
rect 81492 7324 81498 7336
rect 81529 7327 81587 7333
rect 81529 7324 81541 7327
rect 81492 7296 81541 7324
rect 81492 7284 81498 7296
rect 81529 7293 81541 7296
rect 81575 7293 81587 7327
rect 81802 7324 81808 7336
rect 81763 7296 81808 7324
rect 81529 7287 81587 7293
rect 81802 7284 81808 7296
rect 81860 7284 81866 7336
rect 83550 7284 83556 7336
rect 83608 7324 83614 7336
rect 83645 7327 83703 7333
rect 83645 7324 83657 7327
rect 83608 7296 83657 7324
rect 83608 7284 83614 7296
rect 83645 7293 83657 7296
rect 83691 7293 83703 7327
rect 83918 7324 83924 7336
rect 83879 7296 83924 7324
rect 83645 7287 83703 7293
rect 83918 7284 83924 7296
rect 83976 7284 83982 7336
rect 85666 7284 85672 7336
rect 85724 7324 85730 7336
rect 85761 7327 85819 7333
rect 85761 7324 85773 7327
rect 85724 7296 85773 7324
rect 85724 7284 85730 7296
rect 85761 7293 85773 7296
rect 85807 7293 85819 7327
rect 86034 7324 86040 7336
rect 85995 7296 86040 7324
rect 85761 7287 85819 7293
rect 86034 7284 86040 7296
rect 86092 7284 86098 7336
rect 87782 7284 87788 7336
rect 87840 7324 87846 7336
rect 87877 7327 87935 7333
rect 87877 7324 87889 7327
rect 87840 7296 87889 7324
rect 87840 7284 87846 7296
rect 87877 7293 87889 7296
rect 87923 7293 87935 7327
rect 88150 7324 88156 7336
rect 88111 7296 88156 7324
rect 87877 7287 87935 7293
rect 88150 7284 88156 7296
rect 88208 7284 88214 7336
rect 89898 7284 89904 7336
rect 89956 7324 89962 7336
rect 89993 7327 90051 7333
rect 89993 7324 90005 7327
rect 89956 7296 90005 7324
rect 89956 7284 89962 7296
rect 89993 7293 90005 7296
rect 90039 7293 90051 7327
rect 90266 7324 90272 7336
rect 90227 7296 90272 7324
rect 89993 7287 90051 7293
rect 90266 7284 90272 7296
rect 90324 7284 90330 7336
rect 92014 7284 92020 7336
rect 92072 7324 92078 7336
rect 92109 7327 92167 7333
rect 92109 7324 92121 7327
rect 92072 7296 92121 7324
rect 92072 7284 92078 7296
rect 92109 7293 92121 7296
rect 92155 7293 92167 7327
rect 92382 7324 92388 7336
rect 92343 7296 92388 7324
rect 92109 7287 92167 7293
rect 92382 7284 92388 7296
rect 92440 7284 92446 7336
rect 94222 7324 94228 7336
rect 94183 7296 94228 7324
rect 94222 7284 94228 7296
rect 94280 7284 94286 7336
rect 94498 7324 94504 7336
rect 94459 7296 94504 7324
rect 94498 7284 94504 7296
rect 94556 7284 94562 7336
rect 96062 7284 96068 7336
rect 96120 7324 96126 7336
rect 96341 7327 96399 7333
rect 96341 7324 96353 7327
rect 96120 7296 96353 7324
rect 96120 7284 96126 7296
rect 96341 7293 96353 7296
rect 96387 7293 96399 7327
rect 96614 7324 96620 7336
rect 96575 7296 96620 7324
rect 96341 7287 96399 7293
rect 96614 7284 96620 7296
rect 96672 7284 96678 7336
rect 98362 7284 98368 7336
rect 98420 7324 98426 7336
rect 98457 7327 98515 7333
rect 98457 7324 98469 7327
rect 98420 7296 98469 7324
rect 98420 7284 98426 7296
rect 98457 7293 98469 7296
rect 98503 7293 98515 7327
rect 98730 7324 98736 7336
rect 98691 7296 98736 7324
rect 98457 7287 98515 7293
rect 98730 7284 98736 7296
rect 98788 7284 98794 7336
rect 100478 7284 100484 7336
rect 100536 7324 100542 7336
rect 100573 7327 100631 7333
rect 100573 7324 100585 7327
rect 100536 7296 100585 7324
rect 100536 7284 100542 7296
rect 100573 7293 100585 7296
rect 100619 7293 100631 7327
rect 100846 7324 100852 7336
rect 100807 7296 100852 7324
rect 100573 7287 100631 7293
rect 100846 7284 100852 7296
rect 100904 7284 100910 7336
rect 102686 7324 102692 7336
rect 102647 7296 102692 7324
rect 102686 7284 102692 7296
rect 102744 7284 102750 7336
rect 102962 7324 102968 7336
rect 102923 7296 102968 7324
rect 102962 7284 102968 7296
rect 103020 7284 103026 7336
rect 104802 7324 104808 7336
rect 104763 7296 104808 7324
rect 104802 7284 104808 7296
rect 104860 7284 104866 7336
rect 105078 7324 105084 7336
rect 105039 7296 105084 7324
rect 105078 7284 105084 7296
rect 105136 7284 105142 7336
rect 11238 7256 11244 7268
rect 1044 7228 1256 7256
rect 11199 7228 11244 7256
rect 1044 6984 1072 7228
rect 11238 7216 11244 7228
rect 11296 7216 11302 7268
rect 13354 7256 13360 7268
rect 13315 7228 13360 7256
rect 13354 7216 13360 7228
rect 13412 7216 13418 7268
rect 23934 7256 23940 7268
rect 23895 7228 23940 7256
rect 23934 7216 23940 7228
rect 23992 7216 23998 7268
rect 30282 7256 30288 7268
rect 30243 7228 30288 7256
rect 30282 7216 30288 7228
rect 30340 7216 30346 7268
rect 47210 7256 47216 7268
rect 47171 7228 47216 7256
rect 47210 7216 47216 7228
rect 47268 7216 47274 7268
rect 64138 7256 64144 7268
rect 64099 7228 64144 7256
rect 64138 7216 64144 7228
rect 64196 7216 64202 7268
rect 78950 7256 78956 7268
rect 78911 7228 78956 7256
rect 78950 7216 78956 7228
rect 79008 7216 79014 7268
rect 81069 7259 81127 7265
rect 81069 7225 81081 7259
rect 81115 7256 81127 7259
rect 81342 7256 81348 7268
rect 81115 7228 81348 7256
rect 81115 7225 81127 7228
rect 81069 7219 81127 7225
rect 81342 7216 81348 7228
rect 81400 7216 81406 7268
rect 95878 7256 95884 7268
rect 95839 7228 95884 7256
rect 95878 7216 95884 7228
rect 95936 7216 95942 7268
rect 97997 7259 98055 7265
rect 97997 7225 98009 7259
rect 98043 7256 98055 7259
rect 98086 7256 98092 7268
rect 98043 7228 98092 7256
rect 98043 7225 98055 7228
rect 97997 7219 98055 7225
rect 98086 7216 98092 7228
rect 98144 7216 98150 7268
rect 2501 7191 2559 7197
rect 2501 7157 2513 7191
rect 2547 7188 2559 7191
rect 2590 7188 2596 7200
rect 2547 7160 2596 7188
rect 2547 7157 2559 7160
rect 2501 7151 2559 7157
rect 2590 7148 2596 7160
rect 2648 7148 2654 7200
rect 4522 7148 4528 7200
rect 4580 7188 4586 7200
rect 4617 7191 4675 7197
rect 4617 7188 4629 7191
rect 4580 7160 4629 7188
rect 4580 7148 4586 7160
rect 4617 7157 4629 7160
rect 4663 7157 4675 7191
rect 4617 7151 4675 7157
rect 6638 7148 6644 7200
rect 6696 7188 6702 7200
rect 6733 7191 6791 7197
rect 6733 7188 6745 7191
rect 6696 7160 6745 7188
rect 6696 7148 6702 7160
rect 6733 7157 6745 7160
rect 6779 7157 6791 7191
rect 6733 7151 6791 7157
rect 8938 7148 8944 7200
rect 8996 7188 9002 7200
rect 9033 7191 9091 7197
rect 9033 7188 9045 7191
rect 8996 7160 9045 7188
rect 8996 7148 9002 7160
rect 9033 7157 9045 7160
rect 9079 7157 9091 7191
rect 9033 7151 9091 7157
rect 15102 7148 15108 7200
rect 15160 7188 15166 7200
rect 15197 7191 15255 7197
rect 15197 7188 15209 7191
rect 15160 7160 15209 7188
rect 15160 7148 15166 7160
rect 15197 7157 15209 7160
rect 15243 7157 15255 7191
rect 15197 7151 15255 7157
rect 17218 7148 17224 7200
rect 17276 7188 17282 7200
rect 17313 7191 17371 7197
rect 17313 7188 17325 7191
rect 17276 7160 17325 7188
rect 17276 7148 17282 7160
rect 17313 7157 17325 7160
rect 17359 7157 17371 7191
rect 17313 7151 17371 7157
rect 19242 7148 19248 7200
rect 19300 7188 19306 7200
rect 19429 7191 19487 7197
rect 19429 7188 19441 7191
rect 19300 7160 19441 7188
rect 19300 7148 19306 7160
rect 19429 7157 19441 7160
rect 19475 7157 19487 7191
rect 19429 7151 19487 7157
rect 21450 7148 21456 7200
rect 21508 7188 21514 7200
rect 21545 7191 21603 7197
rect 21545 7188 21557 7191
rect 21508 7160 21557 7188
rect 21508 7148 21514 7160
rect 21545 7157 21557 7160
rect 21591 7157 21603 7191
rect 21545 7151 21603 7157
rect 25866 7148 25872 7200
rect 25924 7188 25930 7200
rect 25961 7191 26019 7197
rect 25961 7188 25973 7191
rect 25924 7160 25973 7188
rect 25924 7148 25930 7160
rect 25961 7157 25973 7160
rect 26007 7157 26019 7191
rect 25961 7151 26019 7157
rect 27982 7148 27988 7200
rect 28040 7188 28046 7200
rect 28077 7191 28135 7197
rect 28077 7188 28089 7191
rect 28040 7160 28089 7188
rect 28040 7148 28046 7160
rect 28077 7157 28089 7160
rect 28123 7157 28135 7191
rect 28077 7151 28135 7157
rect 32030 7148 32036 7200
rect 32088 7188 32094 7200
rect 32125 7191 32183 7197
rect 32125 7188 32137 7191
rect 32088 7160 32137 7188
rect 32088 7148 32094 7160
rect 32125 7157 32137 7160
rect 32171 7157 32183 7191
rect 32125 7151 32183 7157
rect 34146 7148 34152 7200
rect 34204 7188 34210 7200
rect 34241 7191 34299 7197
rect 34241 7188 34253 7191
rect 34204 7160 34253 7188
rect 34204 7148 34210 7160
rect 34241 7157 34253 7160
rect 34287 7157 34299 7191
rect 34241 7151 34299 7157
rect 36170 7148 36176 7200
rect 36228 7188 36234 7200
rect 36357 7191 36415 7197
rect 36357 7188 36369 7191
rect 36228 7160 36369 7188
rect 36228 7148 36234 7160
rect 36357 7157 36369 7160
rect 36403 7157 36415 7191
rect 36357 7151 36415 7157
rect 38378 7148 38384 7200
rect 38436 7188 38442 7200
rect 38473 7191 38531 7197
rect 38473 7188 38485 7191
rect 38436 7160 38485 7188
rect 38436 7148 38442 7160
rect 38473 7157 38485 7160
rect 38519 7157 38531 7191
rect 38473 7151 38531 7157
rect 40494 7148 40500 7200
rect 40552 7188 40558 7200
rect 40589 7191 40647 7197
rect 40589 7188 40601 7191
rect 40552 7160 40601 7188
rect 40552 7148 40558 7160
rect 40589 7157 40601 7160
rect 40635 7157 40647 7191
rect 42886 7188 42892 7200
rect 42847 7160 42892 7188
rect 40589 7151 40647 7157
rect 42886 7148 42892 7160
rect 42944 7148 42950 7200
rect 44910 7148 44916 7200
rect 44968 7188 44974 7200
rect 45005 7191 45063 7197
rect 45005 7188 45017 7191
rect 44968 7160 45017 7188
rect 44968 7148 44974 7160
rect 45005 7157 45017 7160
rect 45051 7157 45063 7191
rect 45005 7151 45063 7157
rect 48958 7148 48964 7200
rect 49016 7188 49022 7200
rect 49053 7191 49111 7197
rect 49053 7188 49065 7191
rect 49016 7160 49065 7188
rect 49016 7148 49022 7160
rect 49053 7157 49065 7160
rect 49099 7157 49111 7191
rect 49053 7151 49111 7157
rect 51074 7148 51080 7200
rect 51132 7188 51138 7200
rect 51169 7191 51227 7197
rect 51169 7188 51181 7191
rect 51132 7160 51181 7188
rect 51132 7148 51138 7160
rect 51169 7157 51181 7160
rect 51215 7157 51227 7191
rect 53282 7188 53288 7200
rect 53243 7160 53288 7188
rect 51169 7151 51227 7157
rect 53282 7148 53288 7160
rect 53340 7148 53346 7200
rect 55306 7148 55312 7200
rect 55364 7188 55370 7200
rect 55401 7191 55459 7197
rect 55401 7188 55413 7191
rect 55364 7160 55413 7188
rect 55364 7148 55370 7160
rect 55401 7157 55413 7160
rect 55447 7157 55459 7191
rect 55401 7151 55459 7157
rect 57422 7148 57428 7200
rect 57480 7188 57486 7200
rect 57517 7191 57575 7197
rect 57517 7188 57529 7191
rect 57480 7160 57529 7188
rect 57480 7148 57486 7160
rect 57517 7157 57529 7160
rect 57563 7157 57575 7191
rect 57517 7151 57575 7157
rect 59722 7148 59728 7200
rect 59780 7188 59786 7200
rect 59817 7191 59875 7197
rect 59817 7188 59829 7191
rect 59780 7160 59829 7188
rect 59780 7148 59786 7160
rect 59817 7157 59829 7160
rect 59863 7157 59875 7191
rect 59817 7151 59875 7157
rect 61838 7148 61844 7200
rect 61896 7188 61902 7200
rect 61933 7191 61991 7197
rect 61933 7188 61945 7191
rect 61896 7160 61945 7188
rect 61896 7148 61902 7160
rect 61933 7157 61945 7160
rect 61979 7157 61991 7191
rect 61933 7151 61991 7157
rect 65886 7148 65892 7200
rect 65944 7188 65950 7200
rect 65981 7191 66039 7197
rect 65981 7188 65993 7191
rect 65944 7160 65993 7188
rect 65944 7148 65950 7160
rect 65981 7157 65993 7160
rect 66027 7157 66039 7191
rect 65981 7151 66039 7157
rect 68002 7148 68008 7200
rect 68060 7188 68066 7200
rect 68097 7191 68155 7197
rect 68097 7188 68109 7191
rect 68060 7160 68109 7188
rect 68060 7148 68066 7160
rect 68097 7157 68109 7160
rect 68143 7157 68155 7191
rect 70210 7188 70216 7200
rect 70171 7160 70216 7188
rect 68097 7151 68155 7157
rect 70210 7148 70216 7160
rect 70268 7148 70274 7200
rect 72234 7148 72240 7200
rect 72292 7188 72298 7200
rect 72329 7191 72387 7197
rect 72329 7188 72341 7191
rect 72292 7160 72341 7188
rect 72292 7148 72298 7160
rect 72329 7157 72341 7160
rect 72375 7157 72387 7191
rect 72329 7151 72387 7157
rect 74350 7148 74356 7200
rect 74408 7188 74414 7200
rect 74445 7191 74503 7197
rect 74445 7188 74457 7191
rect 74408 7160 74457 7188
rect 74408 7148 74414 7160
rect 74445 7157 74457 7160
rect 74491 7157 74503 7191
rect 74445 7151 74503 7157
rect 76650 7148 76656 7200
rect 76708 7188 76714 7200
rect 76745 7191 76803 7197
rect 76745 7188 76757 7191
rect 76708 7160 76757 7188
rect 76708 7148 76714 7160
rect 76745 7157 76757 7160
rect 76791 7157 76803 7191
rect 76745 7151 76803 7157
rect 82814 7148 82820 7200
rect 82872 7188 82878 7200
rect 82909 7191 82967 7197
rect 82909 7188 82921 7191
rect 82872 7160 82921 7188
rect 82872 7148 82878 7160
rect 82909 7157 82921 7160
rect 82955 7157 82967 7191
rect 82909 7151 82967 7157
rect 85114 7148 85120 7200
rect 85172 7188 85178 7200
rect 85209 7191 85267 7197
rect 85209 7188 85221 7191
rect 85172 7160 85221 7188
rect 85172 7148 85178 7160
rect 85209 7157 85221 7160
rect 85255 7157 85267 7191
rect 87138 7188 87144 7200
rect 87099 7160 87144 7188
rect 85209 7151 85267 7157
rect 87138 7148 87144 7160
rect 87196 7148 87202 7200
rect 89162 7148 89168 7200
rect 89220 7188 89226 7200
rect 89257 7191 89315 7197
rect 89257 7188 89269 7191
rect 89220 7160 89269 7188
rect 89220 7148 89226 7160
rect 89257 7157 89269 7160
rect 89303 7157 89315 7191
rect 89257 7151 89315 7157
rect 91373 7191 91431 7197
rect 91373 7157 91385 7191
rect 91419 7188 91431 7191
rect 91462 7188 91468 7200
rect 91419 7160 91468 7188
rect 91419 7157 91431 7160
rect 91373 7151 91431 7157
rect 91462 7148 91468 7160
rect 91520 7148 91526 7200
rect 93578 7148 93584 7200
rect 93636 7188 93642 7200
rect 93673 7191 93731 7197
rect 93673 7188 93685 7191
rect 93636 7160 93685 7188
rect 93636 7148 93642 7160
rect 93673 7157 93685 7160
rect 93719 7157 93731 7191
rect 93673 7151 93731 7157
rect 99742 7148 99748 7200
rect 99800 7188 99806 7200
rect 99837 7191 99895 7197
rect 99837 7188 99849 7191
rect 99800 7160 99849 7188
rect 99800 7148 99806 7160
rect 99837 7157 99849 7160
rect 99883 7157 99895 7191
rect 99837 7151 99895 7157
rect 101858 7148 101864 7200
rect 101916 7188 101922 7200
rect 101953 7191 102011 7197
rect 101953 7188 101965 7191
rect 101916 7160 101965 7188
rect 101916 7148 101922 7160
rect 101953 7157 101965 7160
rect 101999 7157 102011 7191
rect 101953 7151 102011 7157
rect 103882 7148 103888 7200
rect 103940 7188 103946 7200
rect 104069 7191 104127 7197
rect 104069 7188 104081 7191
rect 103940 7160 104081 7188
rect 103940 7148 103946 7160
rect 104069 7157 104081 7160
rect 104115 7157 104127 7191
rect 106182 7188 106188 7200
rect 106143 7160 106188 7188
rect 104069 7151 104127 7157
rect 106182 7148 106188 7160
rect 106240 7148 106246 7200
rect 1104 7098 106904 7120
rect 1104 7046 19402 7098
rect 19454 7046 19466 7098
rect 19518 7046 19530 7098
rect 19582 7046 19594 7098
rect 19646 7046 50122 7098
rect 50174 7046 50186 7098
rect 50238 7046 50250 7098
rect 50302 7046 50314 7098
rect 50366 7046 80842 7098
rect 80894 7046 80906 7098
rect 80958 7046 80970 7098
rect 81022 7046 81034 7098
rect 81086 7046 106904 7098
rect 1104 7024 106904 7046
rect 2501 6987 2559 6993
rect 2501 6984 2513 6987
rect 1044 6956 2513 6984
rect 2501 6953 2513 6956
rect 2547 6953 2559 6987
rect 2501 6947 2559 6953
rect 3510 6944 3516 6996
rect 3568 6984 3574 6996
rect 4617 6987 4675 6993
rect 4617 6984 4629 6987
rect 3568 6956 4629 6984
rect 3568 6944 3574 6956
rect 4617 6953 4629 6956
rect 4663 6953 4675 6987
rect 4617 6947 4675 6953
rect 5626 6944 5632 6996
rect 5684 6984 5690 6996
rect 6733 6987 6791 6993
rect 6733 6984 6745 6987
rect 5684 6956 6745 6984
rect 5684 6944 5690 6956
rect 6733 6953 6745 6956
rect 6779 6953 6791 6987
rect 6733 6947 6791 6953
rect 7742 6944 7748 6996
rect 7800 6984 7806 6996
rect 8849 6987 8907 6993
rect 8849 6984 8861 6987
rect 7800 6956 8861 6984
rect 7800 6944 7806 6956
rect 8849 6953 8861 6956
rect 8895 6953 8907 6987
rect 8849 6947 8907 6953
rect 9858 6944 9864 6996
rect 9916 6984 9922 6996
rect 10965 6987 11023 6993
rect 10965 6984 10977 6987
rect 9916 6956 10977 6984
rect 9916 6944 9922 6956
rect 10965 6953 10977 6956
rect 11011 6953 11023 6987
rect 10965 6947 11023 6953
rect 11974 6944 11980 6996
rect 12032 6984 12038 6996
rect 13081 6987 13139 6993
rect 13081 6984 13093 6987
rect 12032 6956 13093 6984
rect 12032 6944 12038 6956
rect 13081 6953 13093 6956
rect 13127 6953 13139 6987
rect 13081 6947 13139 6953
rect 14090 6944 14096 6996
rect 14148 6984 14154 6996
rect 15197 6987 15255 6993
rect 15197 6984 15209 6987
rect 14148 6956 15209 6984
rect 14148 6944 14154 6956
rect 15197 6953 15209 6956
rect 15243 6953 15255 6987
rect 15197 6947 15255 6953
rect 16206 6944 16212 6996
rect 16264 6984 16270 6996
rect 17313 6987 17371 6993
rect 17313 6984 17325 6987
rect 16264 6956 17325 6984
rect 16264 6944 16270 6956
rect 17313 6953 17325 6956
rect 17359 6953 17371 6987
rect 17313 6947 17371 6953
rect 18322 6944 18328 6996
rect 18380 6984 18386 6996
rect 19429 6987 19487 6993
rect 19429 6984 19441 6987
rect 18380 6956 19441 6984
rect 18380 6944 18386 6956
rect 19429 6953 19441 6956
rect 19475 6953 19487 6987
rect 19429 6947 19487 6953
rect 20438 6944 20444 6996
rect 20496 6984 20502 6996
rect 21545 6987 21603 6993
rect 21545 6984 21557 6987
rect 20496 6956 21557 6984
rect 20496 6944 20502 6956
rect 21545 6953 21557 6956
rect 21591 6953 21603 6987
rect 21545 6947 21603 6953
rect 22554 6944 22560 6996
rect 22612 6984 22618 6996
rect 23661 6987 23719 6993
rect 23661 6984 23673 6987
rect 22612 6956 23673 6984
rect 22612 6944 22618 6956
rect 23661 6953 23673 6956
rect 23707 6953 23719 6987
rect 23661 6947 23719 6953
rect 24670 6944 24676 6996
rect 24728 6984 24734 6996
rect 25777 6987 25835 6993
rect 25777 6984 25789 6987
rect 24728 6956 25789 6984
rect 24728 6944 24734 6956
rect 25777 6953 25789 6956
rect 25823 6953 25835 6987
rect 25777 6947 25835 6953
rect 26786 6944 26792 6996
rect 26844 6984 26850 6996
rect 27893 6987 27951 6993
rect 27893 6984 27905 6987
rect 26844 6956 27905 6984
rect 26844 6944 26850 6956
rect 27893 6953 27905 6956
rect 27939 6953 27951 6987
rect 27893 6947 27951 6953
rect 28902 6944 28908 6996
rect 28960 6984 28966 6996
rect 30009 6987 30067 6993
rect 30009 6984 30021 6987
rect 28960 6956 30021 6984
rect 28960 6944 28966 6956
rect 30009 6953 30021 6956
rect 30055 6953 30067 6987
rect 30009 6947 30067 6953
rect 31018 6944 31024 6996
rect 31076 6984 31082 6996
rect 32125 6987 32183 6993
rect 32125 6984 32137 6987
rect 31076 6956 32137 6984
rect 31076 6944 31082 6956
rect 32125 6953 32137 6956
rect 32171 6953 32183 6987
rect 32125 6947 32183 6953
rect 33134 6944 33140 6996
rect 33192 6984 33198 6996
rect 34241 6987 34299 6993
rect 34241 6984 34253 6987
rect 33192 6956 34253 6984
rect 33192 6944 33198 6956
rect 34241 6953 34253 6956
rect 34287 6953 34299 6987
rect 34241 6947 34299 6953
rect 35250 6944 35256 6996
rect 35308 6984 35314 6996
rect 36357 6987 36415 6993
rect 36357 6984 36369 6987
rect 35308 6956 36369 6984
rect 35308 6944 35314 6956
rect 36357 6953 36369 6956
rect 36403 6953 36415 6987
rect 36357 6947 36415 6953
rect 37366 6944 37372 6996
rect 37424 6984 37430 6996
rect 38473 6987 38531 6993
rect 38473 6984 38485 6987
rect 37424 6956 38485 6984
rect 37424 6944 37430 6956
rect 38473 6953 38485 6956
rect 38519 6953 38531 6987
rect 38473 6947 38531 6953
rect 39482 6944 39488 6996
rect 39540 6984 39546 6996
rect 40589 6987 40647 6993
rect 40589 6984 40601 6987
rect 39540 6956 40601 6984
rect 39540 6944 39546 6956
rect 40589 6953 40601 6956
rect 40635 6953 40647 6987
rect 40589 6947 40647 6953
rect 41598 6944 41604 6996
rect 41656 6984 41662 6996
rect 42705 6987 42763 6993
rect 42705 6984 42717 6987
rect 41656 6956 42717 6984
rect 41656 6944 41662 6956
rect 42705 6953 42717 6956
rect 42751 6953 42763 6987
rect 42705 6947 42763 6953
rect 43714 6944 43720 6996
rect 43772 6984 43778 6996
rect 44821 6987 44879 6993
rect 44821 6984 44833 6987
rect 43772 6956 44833 6984
rect 43772 6944 43778 6956
rect 44821 6953 44833 6956
rect 44867 6953 44879 6987
rect 44821 6947 44879 6953
rect 45830 6944 45836 6996
rect 45888 6984 45894 6996
rect 46937 6987 46995 6993
rect 46937 6984 46949 6987
rect 45888 6956 46949 6984
rect 45888 6944 45894 6956
rect 46937 6953 46949 6956
rect 46983 6953 46995 6987
rect 46937 6947 46995 6953
rect 47946 6944 47952 6996
rect 48004 6984 48010 6996
rect 49053 6987 49111 6993
rect 49053 6984 49065 6987
rect 48004 6956 49065 6984
rect 48004 6944 48010 6956
rect 49053 6953 49065 6956
rect 49099 6953 49111 6987
rect 51166 6984 51172 6996
rect 51127 6956 51172 6984
rect 49053 6947 49111 6953
rect 51166 6944 51172 6956
rect 51224 6944 51230 6996
rect 52178 6944 52184 6996
rect 52236 6984 52242 6996
rect 53285 6987 53343 6993
rect 53285 6984 53297 6987
rect 52236 6956 53297 6984
rect 52236 6944 52242 6956
rect 53285 6953 53297 6956
rect 53331 6953 53343 6987
rect 53285 6947 53343 6953
rect 54294 6944 54300 6996
rect 54352 6984 54358 6996
rect 55401 6987 55459 6993
rect 55401 6984 55413 6987
rect 54352 6956 55413 6984
rect 54352 6944 54358 6956
rect 55401 6953 55413 6956
rect 55447 6953 55459 6987
rect 55401 6947 55459 6953
rect 56410 6944 56416 6996
rect 56468 6984 56474 6996
rect 57517 6987 57575 6993
rect 57517 6984 57529 6987
rect 56468 6956 57529 6984
rect 56468 6944 56474 6956
rect 57517 6953 57529 6956
rect 57563 6953 57575 6987
rect 57517 6947 57575 6953
rect 58526 6944 58532 6996
rect 58584 6984 58590 6996
rect 59633 6987 59691 6993
rect 59633 6984 59645 6987
rect 58584 6956 59645 6984
rect 58584 6944 58590 6956
rect 59633 6953 59645 6956
rect 59679 6953 59691 6987
rect 59633 6947 59691 6953
rect 60642 6944 60648 6996
rect 60700 6984 60706 6996
rect 61749 6987 61807 6993
rect 61749 6984 61761 6987
rect 60700 6956 61761 6984
rect 60700 6944 60706 6956
rect 61749 6953 61761 6956
rect 61795 6953 61807 6987
rect 61749 6947 61807 6953
rect 62758 6944 62764 6996
rect 62816 6984 62822 6996
rect 63865 6987 63923 6993
rect 63865 6984 63877 6987
rect 62816 6956 63877 6984
rect 62816 6944 62822 6956
rect 63865 6953 63877 6956
rect 63911 6953 63923 6987
rect 63865 6947 63923 6953
rect 64874 6944 64880 6996
rect 64932 6984 64938 6996
rect 65981 6987 66039 6993
rect 65981 6984 65993 6987
rect 64932 6956 65993 6984
rect 64932 6944 64938 6956
rect 65981 6953 65993 6956
rect 66027 6953 66039 6987
rect 65981 6947 66039 6953
rect 66990 6944 66996 6996
rect 67048 6984 67054 6996
rect 68097 6987 68155 6993
rect 68097 6984 68109 6987
rect 67048 6956 68109 6984
rect 67048 6944 67054 6956
rect 68097 6953 68109 6956
rect 68143 6953 68155 6987
rect 68097 6947 68155 6953
rect 69106 6944 69112 6996
rect 69164 6984 69170 6996
rect 70213 6987 70271 6993
rect 70213 6984 70225 6987
rect 69164 6956 70225 6984
rect 69164 6944 69170 6956
rect 70213 6953 70225 6956
rect 70259 6953 70271 6987
rect 70213 6947 70271 6953
rect 71222 6944 71228 6996
rect 71280 6984 71286 6996
rect 72329 6987 72387 6993
rect 72329 6984 72341 6987
rect 71280 6956 72341 6984
rect 71280 6944 71286 6956
rect 72329 6953 72341 6956
rect 72375 6953 72387 6987
rect 72329 6947 72387 6953
rect 73338 6944 73344 6996
rect 73396 6984 73402 6996
rect 74445 6987 74503 6993
rect 74445 6984 74457 6987
rect 73396 6956 74457 6984
rect 73396 6944 73402 6956
rect 74445 6953 74457 6956
rect 74491 6953 74503 6987
rect 74445 6947 74503 6953
rect 75454 6944 75460 6996
rect 75512 6984 75518 6996
rect 76561 6987 76619 6993
rect 76561 6984 76573 6987
rect 75512 6956 76573 6984
rect 75512 6944 75518 6956
rect 76561 6953 76573 6956
rect 76607 6953 76619 6987
rect 76561 6947 76619 6953
rect 77570 6944 77576 6996
rect 77628 6984 77634 6996
rect 78677 6987 78735 6993
rect 78677 6984 78689 6987
rect 77628 6956 78689 6984
rect 77628 6944 77634 6956
rect 78677 6953 78689 6956
rect 78723 6953 78735 6987
rect 78677 6947 78735 6953
rect 79686 6944 79692 6996
rect 79744 6984 79750 6996
rect 80793 6987 80851 6993
rect 80793 6984 80805 6987
rect 79744 6956 80805 6984
rect 79744 6944 79750 6956
rect 80793 6953 80805 6956
rect 80839 6953 80851 6987
rect 80793 6947 80851 6953
rect 81802 6944 81808 6996
rect 81860 6984 81866 6996
rect 82909 6987 82967 6993
rect 82909 6984 82921 6987
rect 81860 6956 82921 6984
rect 81860 6944 81866 6956
rect 82909 6953 82921 6956
rect 82955 6953 82967 6987
rect 82909 6947 82967 6953
rect 83918 6944 83924 6996
rect 83976 6984 83982 6996
rect 85025 6987 85083 6993
rect 85025 6984 85037 6987
rect 83976 6956 85037 6984
rect 83976 6944 83982 6956
rect 85025 6953 85037 6956
rect 85071 6953 85083 6987
rect 85025 6947 85083 6953
rect 86034 6944 86040 6996
rect 86092 6984 86098 6996
rect 87141 6987 87199 6993
rect 87141 6984 87153 6987
rect 86092 6956 87153 6984
rect 86092 6944 86098 6956
rect 87141 6953 87153 6956
rect 87187 6953 87199 6987
rect 87141 6947 87199 6953
rect 88150 6944 88156 6996
rect 88208 6984 88214 6996
rect 89257 6987 89315 6993
rect 89257 6984 89269 6987
rect 88208 6956 89269 6984
rect 88208 6944 88214 6956
rect 89257 6953 89269 6956
rect 89303 6953 89315 6987
rect 89257 6947 89315 6953
rect 90266 6944 90272 6996
rect 90324 6984 90330 6996
rect 91373 6987 91431 6993
rect 91373 6984 91385 6987
rect 90324 6956 91385 6984
rect 90324 6944 90330 6956
rect 91373 6953 91385 6956
rect 91419 6953 91431 6987
rect 91373 6947 91431 6953
rect 92382 6944 92388 6996
rect 92440 6984 92446 6996
rect 93489 6987 93547 6993
rect 93489 6984 93501 6987
rect 92440 6956 93501 6984
rect 92440 6944 92446 6956
rect 93489 6953 93501 6956
rect 93535 6953 93547 6987
rect 93489 6947 93547 6953
rect 94498 6944 94504 6996
rect 94556 6984 94562 6996
rect 95605 6987 95663 6993
rect 95605 6984 95617 6987
rect 94556 6956 95617 6984
rect 94556 6944 94562 6956
rect 95605 6953 95617 6956
rect 95651 6953 95663 6987
rect 95605 6947 95663 6953
rect 96614 6944 96620 6996
rect 96672 6984 96678 6996
rect 97721 6987 97779 6993
rect 97721 6984 97733 6987
rect 96672 6956 97733 6984
rect 96672 6944 96678 6956
rect 97721 6953 97733 6956
rect 97767 6953 97779 6987
rect 97721 6947 97779 6953
rect 98730 6944 98736 6996
rect 98788 6984 98794 6996
rect 99837 6987 99895 6993
rect 99837 6984 99849 6987
rect 98788 6956 99849 6984
rect 98788 6944 98794 6956
rect 99837 6953 99849 6956
rect 99883 6953 99895 6987
rect 99837 6947 99895 6953
rect 100846 6944 100852 6996
rect 100904 6984 100910 6996
rect 101953 6987 102011 6993
rect 101953 6984 101965 6987
rect 100904 6956 101965 6984
rect 100904 6944 100910 6956
rect 101953 6953 101965 6956
rect 101999 6953 102011 6987
rect 101953 6947 102011 6953
rect 102962 6944 102968 6996
rect 103020 6984 103026 6996
rect 104069 6987 104127 6993
rect 104069 6984 104081 6987
rect 103020 6956 104081 6984
rect 103020 6944 103026 6956
rect 104069 6953 104081 6956
rect 104115 6953 104127 6987
rect 104069 6947 104127 6953
rect 105078 6944 105084 6996
rect 105136 6984 105142 6996
rect 106185 6987 106243 6993
rect 106185 6984 106197 6987
rect 105136 6956 106197 6984
rect 105136 6944 105142 6956
rect 106185 6953 106197 6956
rect 106231 6953 106243 6987
rect 106185 6947 106243 6953
rect 1118 6848 1124 6860
rect 1079 6820 1124 6848
rect 1118 6808 1124 6820
rect 1176 6808 1182 6860
rect 3234 6848 3240 6860
rect 3195 6820 3240 6848
rect 3234 6808 3240 6820
rect 3292 6808 3298 6860
rect 5258 6808 5264 6860
rect 5316 6848 5322 6860
rect 5353 6851 5411 6857
rect 5353 6848 5365 6851
rect 5316 6820 5365 6848
rect 5316 6808 5322 6820
rect 5353 6817 5365 6820
rect 5399 6817 5411 6851
rect 5353 6811 5411 6817
rect 7374 6808 7380 6860
rect 7432 6848 7438 6860
rect 7469 6851 7527 6857
rect 7469 6848 7481 6851
rect 7432 6820 7481 6848
rect 7432 6808 7438 6820
rect 7469 6817 7481 6820
rect 7515 6817 7527 6851
rect 9582 6848 9588 6860
rect 9543 6820 9588 6848
rect 7469 6811 7527 6817
rect 9582 6808 9588 6820
rect 9640 6808 9646 6860
rect 11698 6848 11704 6860
rect 11659 6820 11704 6848
rect 11698 6808 11704 6820
rect 11756 6808 11762 6860
rect 13814 6848 13820 6860
rect 13775 6820 13820 6848
rect 13814 6808 13820 6820
rect 13872 6808 13878 6860
rect 15930 6848 15936 6860
rect 15891 6820 15936 6848
rect 15930 6808 15936 6820
rect 15988 6808 15994 6860
rect 18046 6848 18052 6860
rect 18007 6820 18052 6848
rect 18046 6808 18052 6820
rect 18104 6808 18110 6860
rect 20070 6808 20076 6860
rect 20128 6848 20134 6860
rect 20165 6851 20223 6857
rect 20165 6848 20177 6851
rect 20128 6820 20177 6848
rect 20128 6808 20134 6820
rect 20165 6817 20177 6820
rect 20211 6817 20223 6851
rect 20165 6811 20223 6817
rect 22186 6808 22192 6860
rect 22244 6848 22250 6860
rect 22281 6851 22339 6857
rect 22281 6848 22293 6851
rect 22244 6820 22293 6848
rect 22244 6808 22250 6820
rect 22281 6817 22293 6820
rect 22327 6817 22339 6851
rect 24394 6848 24400 6860
rect 24355 6820 24400 6848
rect 22281 6811 22339 6817
rect 24394 6808 24400 6820
rect 24452 6808 24458 6860
rect 26510 6848 26516 6860
rect 26471 6820 26516 6848
rect 26510 6808 26516 6820
rect 26568 6808 26574 6860
rect 28626 6848 28632 6860
rect 28587 6820 28632 6848
rect 28626 6808 28632 6820
rect 28684 6808 28690 6860
rect 30742 6848 30748 6860
rect 30703 6820 30748 6848
rect 30742 6808 30748 6820
rect 30800 6808 30806 6860
rect 32858 6848 32864 6860
rect 32819 6820 32864 6848
rect 32858 6808 32864 6820
rect 32916 6808 32922 6860
rect 34977 6851 35035 6857
rect 34977 6817 34989 6851
rect 35023 6848 35035 6851
rect 35066 6848 35072 6860
rect 35023 6820 35072 6848
rect 35023 6817 35035 6820
rect 34977 6811 35035 6817
rect 35066 6808 35072 6820
rect 35124 6808 35130 6860
rect 37090 6848 37096 6860
rect 37051 6820 37096 6848
rect 37090 6808 37096 6820
rect 37148 6808 37154 6860
rect 39206 6848 39212 6860
rect 39167 6820 39212 6848
rect 39206 6808 39212 6820
rect 39264 6808 39270 6860
rect 41230 6808 41236 6860
rect 41288 6848 41294 6860
rect 41325 6851 41383 6857
rect 41325 6848 41337 6851
rect 41288 6820 41337 6848
rect 41288 6808 41294 6820
rect 41325 6817 41337 6820
rect 41371 6817 41383 6851
rect 43438 6848 43444 6860
rect 43399 6820 43444 6848
rect 41325 6811 41383 6817
rect 43438 6808 43444 6820
rect 43496 6808 43502 6860
rect 45554 6848 45560 6860
rect 45515 6820 45560 6848
rect 45554 6808 45560 6820
rect 45612 6808 45618 6860
rect 47670 6848 47676 6860
rect 47631 6820 47676 6848
rect 47670 6808 47676 6820
rect 47728 6808 47734 6860
rect 49786 6848 49792 6860
rect 49747 6820 49792 6848
rect 49786 6808 49792 6820
rect 49844 6808 49850 6860
rect 51902 6848 51908 6860
rect 51863 6820 51908 6848
rect 51902 6808 51908 6820
rect 51960 6808 51966 6860
rect 54018 6848 54024 6860
rect 53979 6820 54024 6848
rect 54018 6808 54024 6820
rect 54076 6808 54082 6860
rect 56042 6808 56048 6860
rect 56100 6848 56106 6860
rect 56137 6851 56195 6857
rect 56137 6848 56149 6851
rect 56100 6820 56149 6848
rect 56100 6808 56106 6820
rect 56137 6817 56149 6820
rect 56183 6817 56195 6851
rect 56137 6811 56195 6817
rect 58158 6808 58164 6860
rect 58216 6848 58222 6860
rect 58253 6851 58311 6857
rect 58253 6848 58265 6851
rect 58216 6820 58265 6848
rect 58216 6808 58222 6820
rect 58253 6817 58265 6820
rect 58299 6817 58311 6851
rect 62482 6848 62488 6860
rect 62443 6820 62488 6848
rect 58253 6811 58311 6817
rect 62482 6808 62488 6820
rect 62540 6808 62546 6860
rect 64598 6848 64604 6860
rect 64559 6820 64604 6848
rect 64598 6808 64604 6820
rect 64656 6808 64662 6860
rect 66714 6848 66720 6860
rect 66675 6820 66720 6848
rect 66714 6808 66720 6820
rect 66772 6808 66778 6860
rect 68830 6848 68836 6860
rect 68791 6820 68836 6848
rect 68830 6808 68836 6820
rect 68888 6808 68894 6860
rect 70854 6808 70860 6860
rect 70912 6848 70918 6860
rect 70949 6851 71007 6857
rect 70949 6848 70961 6851
rect 70912 6820 70961 6848
rect 70912 6808 70918 6820
rect 70949 6817 70961 6820
rect 70995 6817 71007 6851
rect 70949 6811 71007 6817
rect 72970 6808 72976 6860
rect 73028 6848 73034 6860
rect 73065 6851 73123 6857
rect 73065 6848 73077 6851
rect 73028 6820 73077 6848
rect 73028 6808 73034 6820
rect 73065 6817 73077 6820
rect 73111 6817 73123 6851
rect 73065 6811 73123 6817
rect 75086 6808 75092 6860
rect 75144 6848 75150 6860
rect 75181 6851 75239 6857
rect 75181 6848 75193 6851
rect 75144 6820 75193 6848
rect 75144 6808 75150 6820
rect 75181 6817 75193 6820
rect 75227 6817 75239 6851
rect 75181 6811 75239 6817
rect 79318 6808 79324 6860
rect 79376 6848 79382 6860
rect 79413 6851 79471 6857
rect 79413 6848 79425 6851
rect 79376 6820 79425 6848
rect 79376 6808 79382 6820
rect 79413 6817 79425 6820
rect 79459 6817 79471 6851
rect 79413 6811 79471 6817
rect 81434 6808 81440 6860
rect 81492 6848 81498 6860
rect 81529 6851 81587 6857
rect 81529 6848 81541 6851
rect 81492 6820 81541 6848
rect 81492 6808 81498 6820
rect 81529 6817 81541 6820
rect 81575 6817 81587 6851
rect 81529 6811 81587 6817
rect 83550 6808 83556 6860
rect 83608 6848 83614 6860
rect 83645 6851 83703 6857
rect 83645 6848 83657 6851
rect 83608 6820 83657 6848
rect 83608 6808 83614 6820
rect 83645 6817 83657 6820
rect 83691 6817 83703 6851
rect 83645 6811 83703 6817
rect 85666 6808 85672 6860
rect 85724 6848 85730 6860
rect 85761 6851 85819 6857
rect 85761 6848 85773 6851
rect 85724 6820 85773 6848
rect 85724 6808 85730 6820
rect 85761 6817 85773 6820
rect 85807 6817 85819 6851
rect 85761 6811 85819 6817
rect 87782 6808 87788 6860
rect 87840 6848 87846 6860
rect 87877 6851 87935 6857
rect 87877 6848 87889 6851
rect 87840 6820 87889 6848
rect 87840 6808 87846 6820
rect 87877 6817 87889 6820
rect 87923 6817 87935 6851
rect 87877 6811 87935 6817
rect 89898 6808 89904 6860
rect 89956 6848 89962 6860
rect 89993 6851 90051 6857
rect 89993 6848 90005 6851
rect 89956 6820 90005 6848
rect 89956 6808 89962 6820
rect 89993 6817 90005 6820
rect 90039 6817 90051 6851
rect 89993 6811 90051 6817
rect 92014 6808 92020 6860
rect 92072 6848 92078 6860
rect 92109 6851 92167 6857
rect 92109 6848 92121 6851
rect 92072 6820 92121 6848
rect 92072 6808 92078 6820
rect 92109 6817 92121 6820
rect 92155 6817 92167 6851
rect 94222 6848 94228 6860
rect 94183 6820 94228 6848
rect 92109 6811 92167 6817
rect 94222 6808 94228 6820
rect 94280 6808 94286 6860
rect 96062 6808 96068 6860
rect 96120 6848 96126 6860
rect 96341 6851 96399 6857
rect 96341 6848 96353 6851
rect 96120 6820 96353 6848
rect 96120 6808 96126 6820
rect 96341 6817 96353 6820
rect 96387 6817 96399 6851
rect 96341 6811 96399 6817
rect 98362 6808 98368 6860
rect 98420 6848 98426 6860
rect 98457 6851 98515 6857
rect 98457 6848 98469 6851
rect 98420 6820 98469 6848
rect 98420 6808 98426 6820
rect 98457 6817 98469 6820
rect 98503 6817 98515 6851
rect 98457 6811 98515 6817
rect 100478 6808 100484 6860
rect 100536 6848 100542 6860
rect 100573 6851 100631 6857
rect 100573 6848 100585 6851
rect 100536 6820 100585 6848
rect 100536 6808 100542 6820
rect 100573 6817 100585 6820
rect 100619 6817 100631 6851
rect 102686 6848 102692 6860
rect 102647 6820 102692 6848
rect 100573 6811 100631 6817
rect 102686 6808 102692 6820
rect 102744 6808 102750 6860
rect 104802 6848 104808 6860
rect 104763 6820 104808 6848
rect 104802 6808 104808 6820
rect 104860 6808 104866 6860
rect 1397 6783 1455 6789
rect 1397 6749 1409 6783
rect 1443 6780 1455 6783
rect 2130 6780 2136 6792
rect 1443 6752 2136 6780
rect 1443 6749 1455 6752
rect 1397 6743 1455 6749
rect 2130 6740 2136 6752
rect 2188 6740 2194 6792
rect 3510 6780 3516 6792
rect 3471 6752 3516 6780
rect 3510 6740 3516 6752
rect 3568 6740 3574 6792
rect 5626 6780 5632 6792
rect 5587 6752 5632 6780
rect 5626 6740 5632 6752
rect 5684 6740 5690 6792
rect 7742 6780 7748 6792
rect 7703 6752 7748 6780
rect 7742 6740 7748 6752
rect 7800 6740 7806 6792
rect 9858 6780 9864 6792
rect 9819 6752 9864 6780
rect 9858 6740 9864 6752
rect 9916 6740 9922 6792
rect 11974 6780 11980 6792
rect 11935 6752 11980 6780
rect 11974 6740 11980 6752
rect 12032 6740 12038 6792
rect 14090 6780 14096 6792
rect 14051 6752 14096 6780
rect 14090 6740 14096 6752
rect 14148 6740 14154 6792
rect 16206 6780 16212 6792
rect 16167 6752 16212 6780
rect 16206 6740 16212 6752
rect 16264 6740 16270 6792
rect 18322 6780 18328 6792
rect 18283 6752 18328 6780
rect 18322 6740 18328 6752
rect 18380 6740 18386 6792
rect 20438 6780 20444 6792
rect 20399 6752 20444 6780
rect 20438 6740 20444 6752
rect 20496 6740 20502 6792
rect 22554 6780 22560 6792
rect 22515 6752 22560 6780
rect 22554 6740 22560 6752
rect 22612 6740 22618 6792
rect 24670 6780 24676 6792
rect 24631 6752 24676 6780
rect 24670 6740 24676 6752
rect 24728 6740 24734 6792
rect 26786 6780 26792 6792
rect 26747 6752 26792 6780
rect 26786 6740 26792 6752
rect 26844 6740 26850 6792
rect 28902 6780 28908 6792
rect 28863 6752 28908 6780
rect 28902 6740 28908 6752
rect 28960 6740 28966 6792
rect 31018 6780 31024 6792
rect 30979 6752 31024 6780
rect 31018 6740 31024 6752
rect 31076 6740 31082 6792
rect 33134 6780 33140 6792
rect 33095 6752 33140 6780
rect 33134 6740 33140 6752
rect 33192 6740 33198 6792
rect 35250 6780 35256 6792
rect 35211 6752 35256 6780
rect 35250 6740 35256 6752
rect 35308 6740 35314 6792
rect 37366 6780 37372 6792
rect 37327 6752 37372 6780
rect 37366 6740 37372 6752
rect 37424 6740 37430 6792
rect 39390 6740 39396 6792
rect 39448 6780 39454 6792
rect 39485 6783 39543 6789
rect 39485 6780 39497 6783
rect 39448 6752 39497 6780
rect 39448 6740 39454 6752
rect 39485 6749 39497 6752
rect 39531 6749 39543 6783
rect 41598 6780 41604 6792
rect 41559 6752 41604 6780
rect 39485 6743 39543 6749
rect 41598 6740 41604 6752
rect 41656 6740 41662 6792
rect 43714 6780 43720 6792
rect 43675 6752 43720 6780
rect 43714 6740 43720 6752
rect 43772 6740 43778 6792
rect 45830 6780 45836 6792
rect 45791 6752 45836 6780
rect 45830 6740 45836 6752
rect 45888 6740 45894 6792
rect 47946 6780 47952 6792
rect 47907 6752 47952 6780
rect 47946 6740 47952 6752
rect 48004 6740 48010 6792
rect 50062 6740 50068 6792
rect 50120 6780 50126 6792
rect 52178 6780 52184 6792
rect 50120 6752 50165 6780
rect 52139 6752 52184 6780
rect 50120 6740 50126 6752
rect 52178 6740 52184 6752
rect 52236 6740 52242 6792
rect 54294 6780 54300 6792
rect 54255 6752 54300 6780
rect 54294 6740 54300 6752
rect 54352 6740 54358 6792
rect 56410 6780 56416 6792
rect 56371 6752 56416 6780
rect 56410 6740 56416 6752
rect 56468 6740 56474 6792
rect 58526 6780 58532 6792
rect 58487 6752 58532 6780
rect 58526 6740 58532 6752
rect 58584 6740 58590 6792
rect 60366 6740 60372 6792
rect 60424 6780 60430 6792
rect 60642 6780 60648 6792
rect 60424 6752 60469 6780
rect 60603 6752 60648 6780
rect 60424 6740 60430 6752
rect 60642 6740 60648 6752
rect 60700 6740 60706 6792
rect 62758 6780 62764 6792
rect 62719 6752 62764 6780
rect 62758 6740 62764 6752
rect 62816 6740 62822 6792
rect 64874 6780 64880 6792
rect 64835 6752 64880 6780
rect 64874 6740 64880 6752
rect 64932 6740 64938 6792
rect 66990 6780 66996 6792
rect 66951 6752 66996 6780
rect 66990 6740 66996 6752
rect 67048 6740 67054 6792
rect 69106 6780 69112 6792
rect 69067 6752 69112 6780
rect 69106 6740 69112 6752
rect 69164 6740 69170 6792
rect 71222 6780 71228 6792
rect 71183 6752 71228 6780
rect 71222 6740 71228 6752
rect 71280 6740 71286 6792
rect 73338 6780 73344 6792
rect 73299 6752 73344 6780
rect 73338 6740 73344 6752
rect 73396 6740 73402 6792
rect 75362 6740 75368 6792
rect 75420 6780 75426 6792
rect 75457 6783 75515 6789
rect 75457 6780 75469 6783
rect 75420 6752 75469 6780
rect 75420 6740 75426 6752
rect 75457 6749 75469 6752
rect 75503 6749 75515 6783
rect 77294 6780 77300 6792
rect 77255 6752 77300 6780
rect 75457 6743 75515 6749
rect 77294 6740 77300 6752
rect 77352 6740 77358 6792
rect 77570 6780 77576 6792
rect 77531 6752 77576 6780
rect 77570 6740 77576 6752
rect 77628 6740 77634 6792
rect 79686 6780 79692 6792
rect 79647 6752 79692 6780
rect 79686 6740 79692 6752
rect 79744 6740 79750 6792
rect 81802 6780 81808 6792
rect 81763 6752 81808 6780
rect 81802 6740 81808 6752
rect 81860 6740 81866 6792
rect 83918 6780 83924 6792
rect 83879 6752 83924 6780
rect 83918 6740 83924 6752
rect 83976 6740 83982 6792
rect 85942 6740 85948 6792
rect 86000 6780 86006 6792
rect 86037 6783 86095 6789
rect 86037 6780 86049 6783
rect 86000 6752 86049 6780
rect 86000 6740 86006 6752
rect 86037 6749 86049 6752
rect 86083 6749 86095 6783
rect 88150 6780 88156 6792
rect 88111 6752 88156 6780
rect 86037 6743 86095 6749
rect 88150 6740 88156 6752
rect 88208 6740 88214 6792
rect 90266 6780 90272 6792
rect 90227 6752 90272 6780
rect 90266 6740 90272 6752
rect 90324 6740 90330 6792
rect 92382 6780 92388 6792
rect 92343 6752 92388 6780
rect 92382 6740 92388 6752
rect 92440 6740 92446 6792
rect 94498 6780 94504 6792
rect 94459 6752 94504 6780
rect 94498 6740 94504 6752
rect 94556 6740 94562 6792
rect 96614 6780 96620 6792
rect 96575 6752 96620 6780
rect 96614 6740 96620 6752
rect 96672 6740 96678 6792
rect 98730 6780 98736 6792
rect 98691 6752 98736 6780
rect 98730 6740 98736 6752
rect 98788 6740 98794 6792
rect 100846 6780 100852 6792
rect 100807 6752 100852 6780
rect 100846 6740 100852 6752
rect 100904 6740 100910 6792
rect 102962 6780 102968 6792
rect 102923 6752 102968 6780
rect 102962 6740 102968 6752
rect 103020 6740 103026 6792
rect 105078 6780 105084 6792
rect 105039 6752 105084 6780
rect 105078 6740 105084 6752
rect 105136 6740 105142 6792
rect 1104 6554 106904 6576
rect 1104 6502 4042 6554
rect 4094 6502 4106 6554
rect 4158 6502 4170 6554
rect 4222 6502 4234 6554
rect 4286 6502 34762 6554
rect 34814 6502 34826 6554
rect 34878 6502 34890 6554
rect 34942 6502 34954 6554
rect 35006 6502 65482 6554
rect 65534 6502 65546 6554
rect 65598 6502 65610 6554
rect 65662 6502 65674 6554
rect 65726 6502 96202 6554
rect 96254 6502 96266 6554
rect 96318 6502 96330 6554
rect 96382 6502 96394 6554
rect 96446 6502 106904 6554
rect 1104 6480 106904 6502
rect 2130 6332 2136 6384
rect 2188 6372 2194 6384
rect 3237 6375 3295 6381
rect 3237 6372 3249 6375
rect 2188 6344 3249 6372
rect 2188 6332 2194 6344
rect 3237 6341 3249 6344
rect 3283 6341 3295 6375
rect 3237 6335 3295 6341
rect 3421 6239 3479 6245
rect 3421 6205 3433 6239
rect 3467 6236 3479 6239
rect 3510 6236 3516 6248
rect 3467 6208 3516 6236
rect 3467 6205 3479 6208
rect 3421 6199 3479 6205
rect 3510 6196 3516 6208
rect 3568 6196 3574 6248
rect 5537 6239 5595 6245
rect 5537 6205 5549 6239
rect 5583 6236 5595 6239
rect 5626 6236 5632 6248
rect 5583 6208 5632 6236
rect 5583 6205 5595 6208
rect 5537 6199 5595 6205
rect 5626 6196 5632 6208
rect 5684 6236 5690 6248
rect 7469 6239 7527 6245
rect 7469 6236 7481 6239
rect 5684 6208 7481 6236
rect 5684 6196 5690 6208
rect 7469 6205 7481 6208
rect 7515 6205 7527 6239
rect 7469 6199 7527 6205
rect 7653 6239 7711 6245
rect 7653 6205 7665 6239
rect 7699 6236 7711 6239
rect 7742 6236 7748 6248
rect 7699 6208 7748 6236
rect 7699 6205 7711 6208
rect 7653 6199 7711 6205
rect 7742 6196 7748 6208
rect 7800 6236 7806 6248
rect 9585 6239 9643 6245
rect 9585 6236 9597 6239
rect 7800 6208 9597 6236
rect 7800 6196 7806 6208
rect 9585 6205 9597 6208
rect 9631 6205 9643 6239
rect 9585 6199 9643 6205
rect 9769 6239 9827 6245
rect 9769 6205 9781 6239
rect 9815 6236 9827 6239
rect 9858 6236 9864 6248
rect 9815 6208 9864 6236
rect 9815 6205 9827 6208
rect 9769 6199 9827 6205
rect 9858 6196 9864 6208
rect 9916 6236 9922 6248
rect 11701 6239 11759 6245
rect 11701 6236 11713 6239
rect 9916 6208 11713 6236
rect 9916 6196 9922 6208
rect 11701 6205 11713 6208
rect 11747 6205 11759 6239
rect 11701 6199 11759 6205
rect 11885 6239 11943 6245
rect 11885 6205 11897 6239
rect 11931 6236 11943 6239
rect 11974 6236 11980 6248
rect 11931 6208 11980 6236
rect 11931 6205 11943 6208
rect 11885 6199 11943 6205
rect 11974 6196 11980 6208
rect 12032 6236 12038 6248
rect 13817 6239 13875 6245
rect 13817 6236 13829 6239
rect 12032 6208 13829 6236
rect 12032 6196 12038 6208
rect 13817 6205 13829 6208
rect 13863 6205 13875 6239
rect 13817 6199 13875 6205
rect 14001 6239 14059 6245
rect 14001 6205 14013 6239
rect 14047 6236 14059 6239
rect 14090 6236 14096 6248
rect 14047 6208 14096 6236
rect 14047 6205 14059 6208
rect 14001 6199 14059 6205
rect 14090 6196 14096 6208
rect 14148 6236 14154 6248
rect 15933 6239 15991 6245
rect 15933 6236 15945 6239
rect 14148 6208 15945 6236
rect 14148 6196 14154 6208
rect 15933 6205 15945 6208
rect 15979 6205 15991 6239
rect 15933 6199 15991 6205
rect 16117 6239 16175 6245
rect 16117 6205 16129 6239
rect 16163 6236 16175 6239
rect 16206 6236 16212 6248
rect 16163 6208 16212 6236
rect 16163 6205 16175 6208
rect 16117 6199 16175 6205
rect 16206 6196 16212 6208
rect 16264 6236 16270 6248
rect 18049 6239 18107 6245
rect 18049 6236 18061 6239
rect 16264 6208 18061 6236
rect 16264 6196 16270 6208
rect 18049 6205 18061 6208
rect 18095 6205 18107 6239
rect 18049 6199 18107 6205
rect 18233 6239 18291 6245
rect 18233 6205 18245 6239
rect 18279 6236 18291 6239
rect 18322 6236 18328 6248
rect 18279 6208 18328 6236
rect 18279 6205 18291 6208
rect 18233 6199 18291 6205
rect 18322 6196 18328 6208
rect 18380 6236 18386 6248
rect 20165 6239 20223 6245
rect 20165 6236 20177 6239
rect 18380 6208 20177 6236
rect 18380 6196 18386 6208
rect 20165 6205 20177 6208
rect 20211 6205 20223 6239
rect 20165 6199 20223 6205
rect 20349 6239 20407 6245
rect 20349 6205 20361 6239
rect 20395 6236 20407 6239
rect 20438 6236 20444 6248
rect 20395 6208 20444 6236
rect 20395 6205 20407 6208
rect 20349 6199 20407 6205
rect 20438 6196 20444 6208
rect 20496 6236 20502 6248
rect 22281 6239 22339 6245
rect 22281 6236 22293 6239
rect 20496 6208 22293 6236
rect 20496 6196 20502 6208
rect 22281 6205 22293 6208
rect 22327 6205 22339 6239
rect 22281 6199 22339 6205
rect 22465 6239 22523 6245
rect 22465 6205 22477 6239
rect 22511 6236 22523 6239
rect 22554 6236 22560 6248
rect 22511 6208 22560 6236
rect 22511 6205 22523 6208
rect 22465 6199 22523 6205
rect 22554 6196 22560 6208
rect 22612 6236 22618 6248
rect 24397 6239 24455 6245
rect 24397 6236 24409 6239
rect 22612 6208 24409 6236
rect 22612 6196 22618 6208
rect 24397 6205 24409 6208
rect 24443 6205 24455 6239
rect 24397 6199 24455 6205
rect 24581 6239 24639 6245
rect 24581 6205 24593 6239
rect 24627 6236 24639 6239
rect 24670 6236 24676 6248
rect 24627 6208 24676 6236
rect 24627 6205 24639 6208
rect 24581 6199 24639 6205
rect 24670 6196 24676 6208
rect 24728 6236 24734 6248
rect 26513 6239 26571 6245
rect 26513 6236 26525 6239
rect 24728 6208 26525 6236
rect 24728 6196 24734 6208
rect 26513 6205 26525 6208
rect 26559 6205 26571 6239
rect 26513 6199 26571 6205
rect 26697 6239 26755 6245
rect 26697 6205 26709 6239
rect 26743 6236 26755 6239
rect 26786 6236 26792 6248
rect 26743 6208 26792 6236
rect 26743 6205 26755 6208
rect 26697 6199 26755 6205
rect 26786 6196 26792 6208
rect 26844 6236 26850 6248
rect 28629 6239 28687 6245
rect 28629 6236 28641 6239
rect 26844 6208 28641 6236
rect 26844 6196 26850 6208
rect 28629 6205 28641 6208
rect 28675 6205 28687 6239
rect 28629 6199 28687 6205
rect 28813 6239 28871 6245
rect 28813 6205 28825 6239
rect 28859 6236 28871 6239
rect 28902 6236 28908 6248
rect 28859 6208 28908 6236
rect 28859 6205 28871 6208
rect 28813 6199 28871 6205
rect 28902 6196 28908 6208
rect 28960 6236 28966 6248
rect 30745 6239 30803 6245
rect 30745 6236 30757 6239
rect 28960 6208 30757 6236
rect 28960 6196 28966 6208
rect 30745 6205 30757 6208
rect 30791 6205 30803 6239
rect 30745 6199 30803 6205
rect 30929 6239 30987 6245
rect 30929 6205 30941 6239
rect 30975 6236 30987 6239
rect 31018 6236 31024 6248
rect 30975 6208 31024 6236
rect 30975 6205 30987 6208
rect 30929 6199 30987 6205
rect 31018 6196 31024 6208
rect 31076 6236 31082 6248
rect 32861 6239 32919 6245
rect 32861 6236 32873 6239
rect 31076 6208 32873 6236
rect 31076 6196 31082 6208
rect 32861 6205 32873 6208
rect 32907 6205 32919 6239
rect 32861 6199 32919 6205
rect 33045 6239 33103 6245
rect 33045 6205 33057 6239
rect 33091 6236 33103 6239
rect 33134 6236 33140 6248
rect 33091 6208 33140 6236
rect 33091 6205 33103 6208
rect 33045 6199 33103 6205
rect 33134 6196 33140 6208
rect 33192 6236 33198 6248
rect 34977 6239 35035 6245
rect 34977 6236 34989 6239
rect 33192 6208 34989 6236
rect 33192 6196 33198 6208
rect 34977 6205 34989 6208
rect 35023 6205 35035 6239
rect 34977 6199 35035 6205
rect 35161 6239 35219 6245
rect 35161 6205 35173 6239
rect 35207 6236 35219 6239
rect 35250 6236 35256 6248
rect 35207 6208 35256 6236
rect 35207 6205 35219 6208
rect 35161 6199 35219 6205
rect 35250 6196 35256 6208
rect 35308 6236 35314 6248
rect 37093 6239 37151 6245
rect 37093 6236 37105 6239
rect 35308 6208 37105 6236
rect 35308 6196 35314 6208
rect 37093 6205 37105 6208
rect 37139 6205 37151 6239
rect 37093 6199 37151 6205
rect 37277 6239 37335 6245
rect 37277 6205 37289 6239
rect 37323 6236 37335 6239
rect 37366 6236 37372 6248
rect 37323 6208 37372 6236
rect 37323 6205 37335 6208
rect 37277 6199 37335 6205
rect 37366 6196 37372 6208
rect 37424 6236 37430 6248
rect 39209 6239 39267 6245
rect 39209 6236 39221 6239
rect 37424 6208 39221 6236
rect 37424 6196 37430 6208
rect 39209 6205 39221 6208
rect 39255 6205 39267 6239
rect 39209 6199 39267 6205
rect 41509 6239 41567 6245
rect 41509 6205 41521 6239
rect 41555 6236 41567 6239
rect 41598 6236 41604 6248
rect 41555 6208 41604 6236
rect 41555 6205 41567 6208
rect 41509 6199 41567 6205
rect 41598 6196 41604 6208
rect 41656 6236 41662 6248
rect 43441 6239 43499 6245
rect 43441 6236 43453 6239
rect 41656 6208 43453 6236
rect 41656 6196 41662 6208
rect 43441 6205 43453 6208
rect 43487 6205 43499 6239
rect 43441 6199 43499 6205
rect 43625 6239 43683 6245
rect 43625 6205 43637 6239
rect 43671 6236 43683 6239
rect 43714 6236 43720 6248
rect 43671 6208 43720 6236
rect 43671 6205 43683 6208
rect 43625 6199 43683 6205
rect 43714 6196 43720 6208
rect 43772 6236 43778 6248
rect 45557 6239 45615 6245
rect 45557 6236 45569 6239
rect 43772 6208 45569 6236
rect 43772 6196 43778 6208
rect 45557 6205 45569 6208
rect 45603 6205 45615 6239
rect 45557 6199 45615 6205
rect 45741 6239 45799 6245
rect 45741 6205 45753 6239
rect 45787 6236 45799 6239
rect 45830 6236 45836 6248
rect 45787 6208 45836 6236
rect 45787 6205 45799 6208
rect 45741 6199 45799 6205
rect 45830 6196 45836 6208
rect 45888 6236 45894 6248
rect 47673 6239 47731 6245
rect 47673 6236 47685 6239
rect 45888 6208 47685 6236
rect 45888 6196 45894 6208
rect 47673 6205 47685 6208
rect 47719 6205 47731 6239
rect 47673 6199 47731 6205
rect 47857 6239 47915 6245
rect 47857 6205 47869 6239
rect 47903 6236 47915 6239
rect 47946 6236 47952 6248
rect 47903 6208 47952 6236
rect 47903 6205 47915 6208
rect 47857 6199 47915 6205
rect 47946 6196 47952 6208
rect 48004 6236 48010 6248
rect 49789 6239 49847 6245
rect 49789 6236 49801 6239
rect 48004 6208 49801 6236
rect 48004 6196 48010 6208
rect 49789 6205 49801 6208
rect 49835 6205 49847 6239
rect 49789 6199 49847 6205
rect 49973 6239 50031 6245
rect 49973 6205 49985 6239
rect 50019 6205 50031 6239
rect 49973 6199 50031 6205
rect 52089 6239 52147 6245
rect 52089 6205 52101 6239
rect 52135 6236 52147 6239
rect 52178 6236 52184 6248
rect 52135 6208 52184 6236
rect 52135 6205 52147 6208
rect 52089 6199 52147 6205
rect 3528 6168 3556 6196
rect 5353 6171 5411 6177
rect 5353 6168 5365 6171
rect 3528 6140 5365 6168
rect 5353 6137 5365 6140
rect 5399 6137 5411 6171
rect 39390 6168 39396 6180
rect 39351 6140 39396 6168
rect 5353 6131 5411 6137
rect 39390 6128 39396 6140
rect 39448 6168 39454 6180
rect 41325 6171 41383 6177
rect 41325 6168 41337 6171
rect 39448 6140 41337 6168
rect 39448 6128 39454 6140
rect 41325 6137 41337 6140
rect 41371 6137 41383 6171
rect 41325 6131 41383 6137
rect 49988 6168 50016 6199
rect 52178 6196 52184 6208
rect 52236 6236 52242 6248
rect 54021 6239 54079 6245
rect 54021 6236 54033 6239
rect 52236 6208 54033 6236
rect 52236 6196 52242 6208
rect 54021 6205 54033 6208
rect 54067 6205 54079 6239
rect 54021 6199 54079 6205
rect 54205 6239 54263 6245
rect 54205 6205 54217 6239
rect 54251 6236 54263 6239
rect 54294 6236 54300 6248
rect 54251 6208 54300 6236
rect 54251 6205 54263 6208
rect 54205 6199 54263 6205
rect 54294 6196 54300 6208
rect 54352 6236 54358 6248
rect 56137 6239 56195 6245
rect 56137 6236 56149 6239
rect 54352 6208 56149 6236
rect 54352 6196 54358 6208
rect 56137 6205 56149 6208
rect 56183 6205 56195 6239
rect 56137 6199 56195 6205
rect 56321 6239 56379 6245
rect 56321 6205 56333 6239
rect 56367 6236 56379 6239
rect 56410 6236 56416 6248
rect 56367 6208 56416 6236
rect 56367 6205 56379 6208
rect 56321 6199 56379 6205
rect 56410 6196 56416 6208
rect 56468 6236 56474 6248
rect 58253 6239 58311 6245
rect 58253 6236 58265 6239
rect 56468 6208 58265 6236
rect 56468 6196 56474 6208
rect 58253 6205 58265 6208
rect 58299 6205 58311 6239
rect 58253 6199 58311 6205
rect 58437 6239 58495 6245
rect 58437 6205 58449 6239
rect 58483 6236 58495 6239
rect 58526 6236 58532 6248
rect 58483 6208 58532 6236
rect 58483 6205 58495 6208
rect 58437 6199 58495 6205
rect 58526 6196 58532 6208
rect 58584 6236 58590 6248
rect 60369 6239 60427 6245
rect 60369 6236 60381 6239
rect 58584 6208 60381 6236
rect 58584 6196 58590 6208
rect 60369 6205 60381 6208
rect 60415 6205 60427 6239
rect 60369 6199 60427 6205
rect 60553 6239 60611 6245
rect 60553 6205 60565 6239
rect 60599 6236 60611 6239
rect 60642 6236 60648 6248
rect 60599 6208 60648 6236
rect 60599 6205 60611 6208
rect 60553 6199 60611 6205
rect 60642 6196 60648 6208
rect 60700 6236 60706 6248
rect 62485 6239 62543 6245
rect 62485 6236 62497 6239
rect 60700 6208 62497 6236
rect 60700 6196 60706 6208
rect 62485 6205 62497 6208
rect 62531 6205 62543 6239
rect 62485 6199 62543 6205
rect 62669 6239 62727 6245
rect 62669 6205 62681 6239
rect 62715 6236 62727 6239
rect 62758 6236 62764 6248
rect 62715 6208 62764 6236
rect 62715 6205 62727 6208
rect 62669 6199 62727 6205
rect 62758 6196 62764 6208
rect 62816 6236 62822 6248
rect 64601 6239 64659 6245
rect 64601 6236 64613 6239
rect 62816 6208 64613 6236
rect 62816 6196 62822 6208
rect 64601 6205 64613 6208
rect 64647 6205 64659 6239
rect 64601 6199 64659 6205
rect 64785 6239 64843 6245
rect 64785 6205 64797 6239
rect 64831 6236 64843 6239
rect 64874 6236 64880 6248
rect 64831 6208 64880 6236
rect 64831 6205 64843 6208
rect 64785 6199 64843 6205
rect 64874 6196 64880 6208
rect 64932 6236 64938 6248
rect 66717 6239 66775 6245
rect 66717 6236 66729 6239
rect 64932 6208 66729 6236
rect 64932 6196 64938 6208
rect 66717 6205 66729 6208
rect 66763 6205 66775 6239
rect 66717 6199 66775 6205
rect 66901 6239 66959 6245
rect 66901 6205 66913 6239
rect 66947 6236 66959 6239
rect 66990 6236 66996 6248
rect 66947 6208 66996 6236
rect 66947 6205 66959 6208
rect 66901 6199 66959 6205
rect 66990 6196 66996 6208
rect 67048 6236 67054 6248
rect 68833 6239 68891 6245
rect 68833 6236 68845 6239
rect 67048 6208 68845 6236
rect 67048 6196 67054 6208
rect 68833 6205 68845 6208
rect 68879 6205 68891 6239
rect 68833 6199 68891 6205
rect 69017 6239 69075 6245
rect 69017 6205 69029 6239
rect 69063 6236 69075 6239
rect 69106 6236 69112 6248
rect 69063 6208 69112 6236
rect 69063 6205 69075 6208
rect 69017 6199 69075 6205
rect 69106 6196 69112 6208
rect 69164 6236 69170 6248
rect 70949 6239 71007 6245
rect 70949 6236 70961 6239
rect 69164 6208 70961 6236
rect 69164 6196 69170 6208
rect 70949 6205 70961 6208
rect 70995 6205 71007 6239
rect 70949 6199 71007 6205
rect 71133 6239 71191 6245
rect 71133 6205 71145 6239
rect 71179 6236 71191 6239
rect 71222 6236 71228 6248
rect 71179 6208 71228 6236
rect 71179 6205 71191 6208
rect 71133 6199 71191 6205
rect 71222 6196 71228 6208
rect 71280 6236 71286 6248
rect 73065 6239 73123 6245
rect 73065 6236 73077 6239
rect 71280 6208 73077 6236
rect 71280 6196 71286 6208
rect 73065 6205 73077 6208
rect 73111 6205 73123 6239
rect 73065 6199 73123 6205
rect 73249 6239 73307 6245
rect 73249 6205 73261 6239
rect 73295 6236 73307 6239
rect 73338 6236 73344 6248
rect 73295 6208 73344 6236
rect 73295 6205 73307 6208
rect 73249 6199 73307 6205
rect 73338 6196 73344 6208
rect 73396 6236 73402 6248
rect 75181 6239 75239 6245
rect 75181 6236 75193 6239
rect 73396 6208 75193 6236
rect 73396 6196 73402 6208
rect 75181 6205 75193 6208
rect 75227 6205 75239 6239
rect 75181 6199 75239 6205
rect 77481 6239 77539 6245
rect 77481 6205 77493 6239
rect 77527 6236 77539 6239
rect 77570 6236 77576 6248
rect 77527 6208 77576 6236
rect 77527 6205 77539 6208
rect 77481 6199 77539 6205
rect 77570 6196 77576 6208
rect 77628 6236 77634 6248
rect 79413 6239 79471 6245
rect 79413 6236 79425 6239
rect 77628 6208 79425 6236
rect 77628 6196 77634 6208
rect 79413 6205 79425 6208
rect 79459 6205 79471 6239
rect 79413 6199 79471 6205
rect 79597 6239 79655 6245
rect 79597 6205 79609 6239
rect 79643 6236 79655 6239
rect 79686 6236 79692 6248
rect 79643 6208 79692 6236
rect 79643 6205 79655 6208
rect 79597 6199 79655 6205
rect 79686 6196 79692 6208
rect 79744 6236 79750 6248
rect 81529 6239 81587 6245
rect 81529 6236 81541 6239
rect 79744 6208 81541 6236
rect 79744 6196 79750 6208
rect 81529 6205 81541 6208
rect 81575 6205 81587 6239
rect 81529 6199 81587 6205
rect 81713 6239 81771 6245
rect 81713 6205 81725 6239
rect 81759 6236 81771 6239
rect 81802 6236 81808 6248
rect 81759 6208 81808 6236
rect 81759 6205 81771 6208
rect 81713 6199 81771 6205
rect 81802 6196 81808 6208
rect 81860 6236 81866 6248
rect 83645 6239 83703 6245
rect 83645 6236 83657 6239
rect 81860 6208 83657 6236
rect 81860 6196 81866 6208
rect 83645 6205 83657 6208
rect 83691 6205 83703 6239
rect 83645 6199 83703 6205
rect 83829 6239 83887 6245
rect 83829 6205 83841 6239
rect 83875 6236 83887 6239
rect 83918 6236 83924 6248
rect 83875 6208 83924 6236
rect 83875 6205 83887 6208
rect 83829 6199 83887 6205
rect 83918 6196 83924 6208
rect 83976 6236 83982 6248
rect 85761 6239 85819 6245
rect 85761 6236 85773 6239
rect 83976 6208 85773 6236
rect 83976 6196 83982 6208
rect 85761 6205 85773 6208
rect 85807 6205 85819 6239
rect 85761 6199 85819 6205
rect 88061 6239 88119 6245
rect 88061 6205 88073 6239
rect 88107 6236 88119 6239
rect 88150 6236 88156 6248
rect 88107 6208 88156 6236
rect 88107 6205 88119 6208
rect 88061 6199 88119 6205
rect 88150 6196 88156 6208
rect 88208 6236 88214 6248
rect 89993 6239 90051 6245
rect 89993 6236 90005 6239
rect 88208 6208 90005 6236
rect 88208 6196 88214 6208
rect 89993 6205 90005 6208
rect 90039 6205 90051 6239
rect 89993 6199 90051 6205
rect 90177 6239 90235 6245
rect 90177 6205 90189 6239
rect 90223 6236 90235 6239
rect 90266 6236 90272 6248
rect 90223 6208 90272 6236
rect 90223 6205 90235 6208
rect 90177 6199 90235 6205
rect 90266 6196 90272 6208
rect 90324 6236 90330 6248
rect 92109 6239 92167 6245
rect 92109 6236 92121 6239
rect 90324 6208 92121 6236
rect 90324 6196 90330 6208
rect 92109 6205 92121 6208
rect 92155 6205 92167 6239
rect 92109 6199 92167 6205
rect 92293 6239 92351 6245
rect 92293 6205 92305 6239
rect 92339 6236 92351 6239
rect 92382 6236 92388 6248
rect 92339 6208 92388 6236
rect 92339 6205 92351 6208
rect 92293 6199 92351 6205
rect 92382 6196 92388 6208
rect 92440 6236 92446 6248
rect 94225 6239 94283 6245
rect 94225 6236 94237 6239
rect 92440 6208 94237 6236
rect 92440 6196 92446 6208
rect 94225 6205 94237 6208
rect 94271 6205 94283 6239
rect 94225 6199 94283 6205
rect 94409 6239 94467 6245
rect 94409 6205 94421 6239
rect 94455 6236 94467 6239
rect 94498 6236 94504 6248
rect 94455 6208 94504 6236
rect 94455 6205 94467 6208
rect 94409 6199 94467 6205
rect 94498 6196 94504 6208
rect 94556 6236 94562 6248
rect 96341 6239 96399 6245
rect 96341 6236 96353 6239
rect 94556 6208 96353 6236
rect 94556 6196 94562 6208
rect 96341 6205 96353 6208
rect 96387 6205 96399 6239
rect 96341 6199 96399 6205
rect 96525 6239 96583 6245
rect 96525 6205 96537 6239
rect 96571 6236 96583 6239
rect 96614 6236 96620 6248
rect 96571 6208 96620 6236
rect 96571 6205 96583 6208
rect 96525 6199 96583 6205
rect 96614 6196 96620 6208
rect 96672 6236 96678 6248
rect 98457 6239 98515 6245
rect 98457 6236 98469 6239
rect 96672 6208 98469 6236
rect 96672 6196 96678 6208
rect 98457 6205 98469 6208
rect 98503 6205 98515 6239
rect 98457 6199 98515 6205
rect 98641 6239 98699 6245
rect 98641 6205 98653 6239
rect 98687 6236 98699 6239
rect 98730 6236 98736 6248
rect 98687 6208 98736 6236
rect 98687 6205 98699 6208
rect 98641 6199 98699 6205
rect 98730 6196 98736 6208
rect 98788 6236 98794 6248
rect 100573 6239 100631 6245
rect 100573 6236 100585 6239
rect 98788 6208 100585 6236
rect 98788 6196 98794 6208
rect 100573 6205 100585 6208
rect 100619 6205 100631 6239
rect 100573 6199 100631 6205
rect 100757 6239 100815 6245
rect 100757 6205 100769 6239
rect 100803 6236 100815 6239
rect 100846 6236 100852 6248
rect 100803 6208 100852 6236
rect 100803 6205 100815 6208
rect 100757 6199 100815 6205
rect 100846 6196 100852 6208
rect 100904 6236 100910 6248
rect 102689 6239 102747 6245
rect 102689 6236 102701 6239
rect 100904 6208 102701 6236
rect 100904 6196 100910 6208
rect 102689 6205 102701 6208
rect 102735 6205 102747 6239
rect 102689 6199 102747 6205
rect 102873 6239 102931 6245
rect 102873 6205 102885 6239
rect 102919 6236 102931 6239
rect 102962 6236 102968 6248
rect 102919 6208 102968 6236
rect 102919 6205 102931 6208
rect 102873 6199 102931 6205
rect 102962 6196 102968 6208
rect 103020 6236 103026 6248
rect 104805 6239 104863 6245
rect 104805 6236 104817 6239
rect 103020 6208 104817 6236
rect 103020 6196 103026 6208
rect 104805 6205 104817 6208
rect 104851 6205 104863 6239
rect 104805 6199 104863 6205
rect 104989 6239 105047 6245
rect 104989 6205 105001 6239
rect 105035 6236 105047 6239
rect 105078 6236 105084 6248
rect 105035 6208 105084 6236
rect 105035 6205 105047 6208
rect 104989 6199 105047 6205
rect 105078 6196 105084 6208
rect 105136 6196 105142 6248
rect 50062 6168 50068 6180
rect 49988 6140 50068 6168
rect 49988 6100 50016 6140
rect 50062 6128 50068 6140
rect 50120 6128 50126 6180
rect 75362 6168 75368 6180
rect 75323 6140 75368 6168
rect 75362 6128 75368 6140
rect 75420 6168 75426 6180
rect 77297 6171 77355 6177
rect 77297 6168 77309 6171
rect 75420 6140 77309 6168
rect 75420 6128 75426 6140
rect 77297 6137 77309 6140
rect 77343 6137 77355 6171
rect 85942 6168 85948 6180
rect 85903 6140 85948 6168
rect 77297 6131 77355 6137
rect 85942 6128 85948 6140
rect 86000 6168 86006 6180
rect 87877 6171 87935 6177
rect 87877 6168 87889 6171
rect 86000 6140 87889 6168
rect 86000 6128 86006 6140
rect 87877 6137 87889 6140
rect 87923 6137 87935 6171
rect 87877 6131 87935 6137
rect 51997 6103 52055 6109
rect 51997 6100 52009 6103
rect 49988 6072 52009 6100
rect 51997 6069 52009 6072
rect 52043 6069 52055 6103
rect 51997 6063 52055 6069
rect 1104 6010 106904 6032
rect 1104 5958 19402 6010
rect 19454 5958 19466 6010
rect 19518 5958 19530 6010
rect 19582 5958 19594 6010
rect 19646 5958 50122 6010
rect 50174 5958 50186 6010
rect 50238 5958 50250 6010
rect 50302 5958 50314 6010
rect 50366 5958 80842 6010
rect 80894 5958 80906 6010
rect 80958 5958 80970 6010
rect 81022 5958 81034 6010
rect 81086 5958 106904 6010
rect 1104 5936 106904 5958
rect 20349 5899 20407 5905
rect 20349 5865 20361 5899
rect 20395 5896 20407 5899
rect 22465 5899 22523 5905
rect 20395 5868 22416 5896
rect 20395 5865 20407 5868
rect 20349 5859 20407 5865
rect 22388 5840 22416 5868
rect 22465 5865 22477 5899
rect 22511 5865 22523 5899
rect 22465 5859 22523 5865
rect 30929 5899 30987 5905
rect 30929 5865 30941 5899
rect 30975 5865 30987 5899
rect 30929 5859 30987 5865
rect 35161 5899 35219 5905
rect 35161 5865 35173 5899
rect 35207 5896 35219 5899
rect 41509 5899 41567 5905
rect 35207 5868 37228 5896
rect 35207 5865 35219 5868
rect 35161 5859 35219 5865
rect 9861 5831 9919 5837
rect 9861 5797 9873 5831
rect 9907 5828 9919 5831
rect 11793 5831 11851 5837
rect 11793 5828 11805 5831
rect 9907 5800 11805 5828
rect 9907 5797 9919 5800
rect 9861 5791 9919 5797
rect 11793 5797 11805 5800
rect 11839 5828 11851 5831
rect 11882 5828 11888 5840
rect 11839 5800 11888 5828
rect 11839 5797 11851 5800
rect 11793 5791 11851 5797
rect 11882 5788 11888 5800
rect 11940 5788 11946 5840
rect 11977 5831 12035 5837
rect 11977 5797 11989 5831
rect 12023 5828 12035 5831
rect 13909 5831 13967 5837
rect 13909 5828 13921 5831
rect 12023 5800 13921 5828
rect 12023 5797 12035 5800
rect 11977 5791 12035 5797
rect 13909 5797 13921 5800
rect 13955 5828 13967 5831
rect 14090 5828 14096 5840
rect 13955 5800 14096 5828
rect 13955 5797 13967 5800
rect 13909 5791 13967 5797
rect 14090 5788 14096 5800
rect 14148 5788 14154 5840
rect 22370 5828 22376 5840
rect 22331 5800 22376 5828
rect 22370 5788 22376 5800
rect 22428 5788 22434 5840
rect 22480 5828 22508 5859
rect 24489 5831 24547 5837
rect 24489 5828 24501 5831
rect 22480 5800 24501 5828
rect 24489 5797 24501 5800
rect 24535 5828 24547 5831
rect 24670 5828 24676 5840
rect 24535 5800 24676 5828
rect 24535 5797 24547 5800
rect 24489 5791 24547 5797
rect 24670 5788 24676 5800
rect 24728 5788 24734 5840
rect 30944 5828 30972 5859
rect 32953 5831 33011 5837
rect 32953 5828 32965 5831
rect 30944 5800 32965 5828
rect 32953 5797 32965 5800
rect 32999 5828 33011 5831
rect 33042 5828 33048 5840
rect 32999 5800 33048 5828
rect 32999 5797 33011 5800
rect 32953 5791 33011 5797
rect 33042 5788 33048 5800
rect 33100 5788 33106 5840
rect 37200 5837 37228 5868
rect 41509 5865 41521 5899
rect 41555 5865 41567 5899
rect 41509 5859 41567 5865
rect 60553 5899 60611 5905
rect 60553 5865 60565 5899
rect 60599 5865 60611 5899
rect 60553 5859 60611 5865
rect 71133 5899 71191 5905
rect 71133 5865 71145 5899
rect 71179 5896 71191 5899
rect 77481 5899 77539 5905
rect 71179 5868 73200 5896
rect 71179 5865 71191 5868
rect 71133 5859 71191 5865
rect 37185 5831 37243 5837
rect 37185 5797 37197 5831
rect 37231 5828 37243 5831
rect 37366 5828 37372 5840
rect 37231 5800 37372 5828
rect 37231 5797 37243 5800
rect 37185 5791 37243 5797
rect 37366 5788 37372 5800
rect 37424 5788 37430 5840
rect 41233 5831 41291 5837
rect 41233 5797 41245 5831
rect 41279 5828 41291 5831
rect 41417 5831 41475 5837
rect 41417 5828 41429 5831
rect 41279 5800 41429 5828
rect 41279 5797 41291 5800
rect 41233 5791 41291 5797
rect 41417 5797 41429 5800
rect 41463 5797 41475 5831
rect 41524 5828 41552 5859
rect 43533 5831 43591 5837
rect 43533 5828 43545 5831
rect 41524 5800 43545 5828
rect 41417 5791 41475 5797
rect 43533 5797 43545 5800
rect 43579 5828 43591 5831
rect 43714 5828 43720 5840
rect 43579 5800 43720 5828
rect 43579 5797 43591 5800
rect 43533 5791 43591 5797
rect 43714 5788 43720 5800
rect 43772 5788 43778 5840
rect 45833 5831 45891 5837
rect 45833 5797 45845 5831
rect 45879 5828 45891 5831
rect 47765 5831 47823 5837
rect 47765 5828 47777 5831
rect 45879 5800 47777 5828
rect 45879 5797 45891 5800
rect 45833 5791 45891 5797
rect 47765 5797 47777 5800
rect 47811 5828 47823 5831
rect 47854 5828 47860 5840
rect 47811 5800 47860 5828
rect 47811 5797 47823 5800
rect 47765 5791 47823 5797
rect 47854 5788 47860 5800
rect 47912 5788 47918 5840
rect 56413 5831 56471 5837
rect 56413 5797 56425 5831
rect 56459 5828 56471 5831
rect 58345 5831 58403 5837
rect 58345 5828 58357 5831
rect 56459 5800 58357 5828
rect 56459 5797 56471 5800
rect 56413 5791 56471 5797
rect 58345 5797 58357 5800
rect 58391 5828 58403 5831
rect 58434 5828 58440 5840
rect 58391 5800 58440 5828
rect 58391 5797 58403 5800
rect 58345 5791 58403 5797
rect 58434 5788 58440 5800
rect 58492 5788 58498 5840
rect 58529 5831 58587 5837
rect 58529 5797 58541 5831
rect 58575 5828 58587 5831
rect 60458 5828 60464 5840
rect 58575 5800 60464 5828
rect 58575 5797 58587 5800
rect 58529 5791 58587 5797
rect 60458 5788 60464 5800
rect 60516 5788 60522 5840
rect 60568 5828 60596 5859
rect 62577 5831 62635 5837
rect 62577 5828 62589 5831
rect 60568 5800 62589 5828
rect 62577 5797 62589 5800
rect 62623 5828 62635 5831
rect 62758 5828 62764 5840
rect 62623 5800 62764 5828
rect 62623 5797 62635 5800
rect 62577 5791 62635 5797
rect 62758 5788 62764 5800
rect 62816 5788 62822 5840
rect 73172 5837 73200 5868
rect 77481 5865 77493 5899
rect 77527 5865 77539 5899
rect 77481 5859 77539 5865
rect 81713 5899 81771 5905
rect 81713 5865 81725 5899
rect 81759 5865 81771 5899
rect 81713 5859 81771 5865
rect 102873 5899 102931 5905
rect 102873 5865 102885 5899
rect 102919 5896 102931 5899
rect 102919 5868 104940 5896
rect 102919 5865 102931 5868
rect 102873 5859 102931 5865
rect 73157 5831 73215 5837
rect 73157 5797 73169 5831
rect 73203 5828 73215 5831
rect 73338 5828 73344 5840
rect 73203 5800 73344 5828
rect 73203 5797 73215 5800
rect 73157 5791 73215 5797
rect 73338 5788 73344 5800
rect 73396 5788 73402 5840
rect 77389 5831 77447 5837
rect 77389 5797 77401 5831
rect 77435 5797 77447 5831
rect 77496 5828 77524 5859
rect 79505 5831 79563 5837
rect 79505 5828 79517 5831
rect 77496 5800 79517 5828
rect 77389 5791 77447 5797
rect 79505 5797 79517 5800
rect 79551 5828 79563 5831
rect 79594 5828 79600 5840
rect 79551 5800 79600 5828
rect 79551 5797 79563 5800
rect 79505 5791 79563 5797
rect 1213 5763 1271 5769
rect 1213 5729 1225 5763
rect 1259 5760 1271 5763
rect 1302 5760 1308 5772
rect 1259 5732 1308 5760
rect 1259 5729 1271 5732
rect 1213 5723 1271 5729
rect 1302 5720 1308 5732
rect 1360 5720 1366 5772
rect 1397 5763 1455 5769
rect 1397 5729 1409 5763
rect 1443 5760 1455 5763
rect 3329 5763 3387 5769
rect 3329 5760 3341 5763
rect 1443 5732 3341 5760
rect 1443 5729 1455 5732
rect 1397 5723 1455 5729
rect 3329 5729 3341 5732
rect 3375 5760 3387 5763
rect 3510 5760 3516 5772
rect 3375 5732 3516 5760
rect 3375 5729 3387 5732
rect 3329 5723 3387 5729
rect 3510 5720 3516 5732
rect 3568 5720 3574 5772
rect 5445 5763 5503 5769
rect 5445 5729 5457 5763
rect 5491 5729 5503 5763
rect 5445 5723 5503 5729
rect 5629 5763 5687 5769
rect 5629 5729 5641 5763
rect 5675 5760 5687 5763
rect 7561 5763 7619 5769
rect 7561 5760 7573 5763
rect 5675 5732 7573 5760
rect 5675 5729 5687 5732
rect 5629 5723 5687 5729
rect 7561 5729 7573 5732
rect 7607 5760 7619 5763
rect 7650 5760 7656 5772
rect 7607 5732 7656 5760
rect 7607 5729 7619 5732
rect 7561 5723 7619 5729
rect 5460 5624 5488 5723
rect 7650 5720 7656 5732
rect 7708 5720 7714 5772
rect 9677 5763 9735 5769
rect 9677 5729 9689 5763
rect 9723 5729 9735 5763
rect 16025 5763 16083 5769
rect 16025 5760 16037 5763
rect 9677 5723 9735 5729
rect 14108 5732 16037 5760
rect 7745 5695 7803 5701
rect 7745 5661 7757 5695
rect 7791 5692 7803 5695
rect 9692 5692 9720 5723
rect 9858 5692 9864 5704
rect 7791 5664 9864 5692
rect 7791 5661 7803 5664
rect 7745 5655 7803 5661
rect 9858 5652 9864 5664
rect 9916 5652 9922 5704
rect 14108 5701 14136 5732
rect 16025 5729 16037 5732
rect 16071 5760 16083 5763
rect 16206 5760 16212 5772
rect 16071 5732 16212 5760
rect 16071 5729 16083 5732
rect 16025 5723 16083 5729
rect 16206 5720 16212 5732
rect 16264 5720 16270 5772
rect 18141 5763 18199 5769
rect 18141 5729 18153 5763
rect 18187 5729 18199 5763
rect 18141 5723 18199 5729
rect 18325 5763 18383 5769
rect 18325 5729 18337 5763
rect 18371 5760 18383 5763
rect 20257 5763 20315 5769
rect 20257 5760 20269 5763
rect 18371 5732 20269 5760
rect 18371 5729 18383 5732
rect 18325 5723 18383 5729
rect 20257 5729 20269 5732
rect 20303 5760 20315 5763
rect 20438 5760 20444 5772
rect 20303 5732 20444 5760
rect 20303 5729 20315 5732
rect 20257 5723 20315 5729
rect 14093 5695 14151 5701
rect 14093 5661 14105 5695
rect 14139 5661 14151 5695
rect 14093 5655 14151 5661
rect 5626 5624 5632 5636
rect 5460 5596 5632 5624
rect 3421 5559 3479 5565
rect 3421 5525 3433 5559
rect 3467 5556 3479 5559
rect 5460 5556 5488 5596
rect 5626 5584 5632 5596
rect 5684 5584 5690 5636
rect 16209 5627 16267 5633
rect 16209 5593 16221 5627
rect 16255 5624 16267 5627
rect 18156 5624 18184 5723
rect 20438 5720 20444 5732
rect 20496 5720 20502 5772
rect 26605 5763 26663 5769
rect 26605 5729 26617 5763
rect 26651 5729 26663 5763
rect 26605 5723 26663 5729
rect 28721 5763 28779 5769
rect 28721 5729 28733 5763
rect 28767 5729 28779 5763
rect 28721 5723 28779 5729
rect 28905 5763 28963 5769
rect 28905 5729 28917 5763
rect 28951 5760 28963 5763
rect 30837 5763 30895 5769
rect 30837 5760 30849 5763
rect 28951 5732 30849 5760
rect 28951 5729 28963 5732
rect 28905 5723 28963 5729
rect 30837 5729 30849 5732
rect 30883 5760 30895 5763
rect 31018 5760 31024 5772
rect 30883 5732 31024 5760
rect 30883 5729 30895 5732
rect 30837 5723 30895 5729
rect 24673 5695 24731 5701
rect 24673 5661 24685 5695
rect 24719 5692 24731 5695
rect 26620 5692 26648 5723
rect 26694 5692 26700 5704
rect 24719 5664 26700 5692
rect 24719 5661 24731 5664
rect 24673 5655 24731 5661
rect 26694 5652 26700 5664
rect 26752 5652 26758 5704
rect 26789 5695 26847 5701
rect 26789 5661 26801 5695
rect 26835 5692 26847 5695
rect 28736 5692 28764 5723
rect 31018 5720 31024 5732
rect 31076 5720 31082 5772
rect 33137 5763 33195 5769
rect 33137 5729 33149 5763
rect 33183 5760 33195 5763
rect 35069 5763 35127 5769
rect 35069 5760 35081 5763
rect 33183 5732 35081 5760
rect 33183 5729 33195 5732
rect 33137 5723 33195 5729
rect 35069 5729 35081 5732
rect 35115 5760 35127 5763
rect 35250 5760 35256 5772
rect 35115 5732 35256 5760
rect 35115 5729 35127 5732
rect 35069 5723 35127 5729
rect 35250 5720 35256 5732
rect 35308 5720 35314 5772
rect 39301 5763 39359 5769
rect 39301 5729 39313 5763
rect 39347 5729 39359 5763
rect 39301 5723 39359 5729
rect 45649 5763 45707 5769
rect 45649 5729 45661 5763
rect 45695 5729 45707 5763
rect 45649 5723 45707 5729
rect 47949 5763 48007 5769
rect 47949 5729 47961 5763
rect 47995 5760 48007 5763
rect 49881 5763 49939 5769
rect 49881 5760 49893 5763
rect 47995 5732 49893 5760
rect 47995 5729 48007 5732
rect 47949 5723 48007 5729
rect 49881 5729 49893 5732
rect 49927 5760 49939 5763
rect 50062 5760 50068 5772
rect 49927 5732 50068 5760
rect 49927 5729 49939 5732
rect 49881 5723 49939 5729
rect 28810 5692 28816 5704
rect 26835 5664 28816 5692
rect 26835 5661 26847 5664
rect 26789 5655 26847 5661
rect 28810 5652 28816 5664
rect 28868 5652 28874 5704
rect 37369 5695 37427 5701
rect 37369 5661 37381 5695
rect 37415 5692 37427 5695
rect 39316 5692 39344 5723
rect 39482 5692 39488 5704
rect 37415 5664 39488 5692
rect 37415 5661 37427 5664
rect 37369 5655 37427 5661
rect 39482 5652 39488 5664
rect 39540 5652 39546 5704
rect 43717 5695 43775 5701
rect 43717 5661 43729 5695
rect 43763 5692 43775 5695
rect 45664 5692 45692 5723
rect 50062 5720 50068 5732
rect 50120 5720 50126 5772
rect 51997 5763 52055 5769
rect 51997 5729 52009 5763
rect 52043 5729 52055 5763
rect 51997 5723 52055 5729
rect 52181 5763 52239 5769
rect 52181 5729 52193 5763
rect 52227 5760 52239 5763
rect 54113 5763 54171 5769
rect 54113 5760 54125 5763
rect 52227 5732 54125 5760
rect 52227 5729 52239 5732
rect 52181 5723 52239 5729
rect 54113 5729 54125 5732
rect 54159 5760 54171 5763
rect 54202 5760 54208 5772
rect 54159 5732 54208 5760
rect 54159 5729 54171 5732
rect 54113 5723 54171 5729
rect 45830 5692 45836 5704
rect 43763 5664 45836 5692
rect 43763 5661 43775 5664
rect 43717 5655 43775 5661
rect 45830 5652 45836 5664
rect 45888 5652 45894 5704
rect 18322 5624 18328 5636
rect 16255 5596 18328 5624
rect 16255 5593 16267 5596
rect 16209 5587 16267 5593
rect 18322 5584 18328 5596
rect 18380 5584 18386 5636
rect 50065 5627 50123 5633
rect 50065 5593 50077 5627
rect 50111 5624 50123 5627
rect 52012 5624 52040 5723
rect 54202 5720 54208 5732
rect 54260 5720 54266 5772
rect 56229 5763 56287 5769
rect 56229 5729 56241 5763
rect 56275 5729 56287 5763
rect 64693 5763 64751 5769
rect 64693 5760 64705 5763
rect 56229 5723 56287 5729
rect 62776 5732 64705 5760
rect 54297 5695 54355 5701
rect 54297 5661 54309 5695
rect 54343 5692 54355 5695
rect 56244 5692 56272 5723
rect 56410 5692 56416 5704
rect 54343 5664 56416 5692
rect 54343 5661 54355 5664
rect 54297 5655 54355 5661
rect 56410 5652 56416 5664
rect 56468 5652 56474 5704
rect 62776 5701 62804 5732
rect 64693 5729 64705 5732
rect 64739 5760 64751 5763
rect 64782 5760 64788 5772
rect 64739 5732 64788 5760
rect 64739 5729 64751 5732
rect 64693 5723 64751 5729
rect 64782 5720 64788 5732
rect 64840 5720 64846 5772
rect 64877 5763 64935 5769
rect 64877 5729 64889 5763
rect 64923 5760 64935 5763
rect 66809 5763 66867 5769
rect 66809 5760 66821 5763
rect 64923 5732 66821 5760
rect 64923 5729 64935 5732
rect 64877 5723 64935 5729
rect 66809 5729 66821 5732
rect 66855 5760 66867 5763
rect 66990 5760 66996 5772
rect 66855 5732 66996 5760
rect 66855 5729 66867 5732
rect 66809 5723 66867 5729
rect 66990 5720 66996 5732
rect 67048 5720 67054 5772
rect 68925 5763 68983 5769
rect 68925 5729 68937 5763
rect 68971 5729 68983 5763
rect 68925 5723 68983 5729
rect 69109 5763 69167 5769
rect 69109 5729 69121 5763
rect 69155 5760 69167 5763
rect 71041 5763 71099 5769
rect 71041 5760 71053 5763
rect 69155 5732 71053 5760
rect 69155 5729 69167 5732
rect 69109 5723 69167 5729
rect 71041 5729 71053 5732
rect 71087 5760 71099 5763
rect 71222 5760 71228 5772
rect 71087 5732 71228 5760
rect 71087 5729 71099 5732
rect 71041 5723 71099 5729
rect 62761 5695 62819 5701
rect 62761 5661 62773 5695
rect 62807 5661 62819 5695
rect 62761 5655 62819 5661
rect 52178 5624 52184 5636
rect 50111 5596 52184 5624
rect 50111 5593 50123 5596
rect 50065 5587 50123 5593
rect 52178 5584 52184 5596
rect 52236 5584 52242 5636
rect 66993 5627 67051 5633
rect 66993 5593 67005 5627
rect 67039 5624 67051 5627
rect 68940 5624 68968 5723
rect 71222 5720 71228 5732
rect 71280 5720 71286 5772
rect 75273 5763 75331 5769
rect 75273 5729 75285 5763
rect 75319 5729 75331 5763
rect 75273 5723 75331 5729
rect 73341 5695 73399 5701
rect 73341 5661 73353 5695
rect 73387 5692 73399 5695
rect 75288 5692 75316 5723
rect 75454 5692 75460 5704
rect 73387 5664 75460 5692
rect 73387 5661 73399 5664
rect 73341 5655 73399 5661
rect 75454 5652 75460 5664
rect 75512 5652 75518 5704
rect 69106 5624 69112 5636
rect 67039 5596 69112 5624
rect 67039 5593 67051 5596
rect 66993 5587 67051 5593
rect 69106 5584 69112 5596
rect 69164 5584 69170 5636
rect 3467 5528 5488 5556
rect 39393 5559 39451 5565
rect 3467 5525 3479 5528
rect 3421 5519 3479 5525
rect 39393 5525 39405 5559
rect 39439 5556 39451 5559
rect 41233 5559 41291 5565
rect 41233 5556 41245 5559
rect 39439 5528 41245 5556
rect 39439 5525 39451 5528
rect 39393 5519 39451 5525
rect 41233 5525 41245 5528
rect 41279 5556 41291 5559
rect 41598 5556 41604 5568
rect 41279 5528 41604 5556
rect 41279 5525 41291 5528
rect 41233 5519 41291 5525
rect 41598 5516 41604 5528
rect 41656 5516 41662 5568
rect 75365 5559 75423 5565
rect 75365 5525 75377 5559
rect 75411 5556 75423 5559
rect 77404 5556 77432 5791
rect 79594 5788 79600 5800
rect 79652 5788 79658 5840
rect 81728 5828 81756 5859
rect 83737 5831 83795 5837
rect 83737 5828 83749 5831
rect 81728 5800 83749 5828
rect 83737 5797 83749 5800
rect 83783 5828 83795 5831
rect 83918 5828 83924 5840
rect 83783 5800 83924 5828
rect 83783 5797 83795 5800
rect 83737 5791 83795 5797
rect 83918 5788 83924 5800
rect 83976 5788 83982 5840
rect 87785 5831 87843 5837
rect 87785 5797 87797 5831
rect 87831 5828 87843 5831
rect 87969 5831 88027 5837
rect 87969 5828 87981 5831
rect 87831 5800 87981 5828
rect 87831 5797 87843 5800
rect 87785 5791 87843 5797
rect 87969 5797 87981 5800
rect 88015 5797 88027 5831
rect 87969 5791 88027 5797
rect 88153 5831 88211 5837
rect 88153 5797 88165 5831
rect 88199 5828 88211 5831
rect 90085 5831 90143 5837
rect 90085 5828 90097 5831
rect 88199 5800 90097 5828
rect 88199 5797 88211 5800
rect 88153 5791 88211 5797
rect 90085 5797 90097 5800
rect 90131 5828 90143 5831
rect 90266 5828 90272 5840
rect 90131 5800 90272 5828
rect 90131 5797 90143 5800
rect 90085 5791 90143 5797
rect 90266 5788 90272 5800
rect 90324 5788 90330 5840
rect 92385 5831 92443 5837
rect 92385 5797 92397 5831
rect 92431 5828 92443 5831
rect 94317 5831 94375 5837
rect 94317 5828 94329 5831
rect 92431 5800 94329 5828
rect 92431 5797 92443 5800
rect 92385 5791 92443 5797
rect 94317 5797 94329 5800
rect 94363 5828 94375 5831
rect 94406 5828 94412 5840
rect 94363 5800 94412 5828
rect 94363 5797 94375 5800
rect 94317 5791 94375 5797
rect 94406 5788 94412 5800
rect 94464 5788 94470 5840
rect 94501 5831 94559 5837
rect 94501 5797 94513 5831
rect 94547 5828 94559 5831
rect 96430 5828 96436 5840
rect 94547 5800 96436 5828
rect 94547 5797 94559 5800
rect 94501 5791 94559 5797
rect 96430 5788 96436 5800
rect 96488 5828 96494 5840
rect 104912 5837 104940 5868
rect 104897 5831 104955 5837
rect 96488 5800 96533 5828
rect 96488 5788 96494 5800
rect 104897 5797 104909 5831
rect 104943 5797 104955 5831
rect 105078 5828 105084 5840
rect 105039 5800 105084 5828
rect 104897 5791 104955 5797
rect 79689 5763 79747 5769
rect 79689 5729 79701 5763
rect 79735 5760 79747 5763
rect 81621 5763 81679 5769
rect 81621 5760 81633 5763
rect 79735 5732 81633 5760
rect 79735 5729 79747 5732
rect 79689 5723 79747 5729
rect 81621 5729 81633 5732
rect 81667 5760 81679 5763
rect 81802 5760 81808 5772
rect 81667 5732 81808 5760
rect 81667 5729 81679 5732
rect 81621 5723 81679 5729
rect 81802 5720 81808 5732
rect 81860 5720 81866 5772
rect 85853 5763 85911 5769
rect 85853 5760 85865 5763
rect 83936 5732 85865 5760
rect 83936 5701 83964 5732
rect 85853 5729 85865 5732
rect 85899 5760 85911 5763
rect 86034 5760 86040 5772
rect 85899 5732 86040 5760
rect 85899 5729 85911 5732
rect 85853 5723 85911 5729
rect 86034 5720 86040 5732
rect 86092 5720 86098 5772
rect 92201 5763 92259 5769
rect 92201 5729 92213 5763
rect 92247 5729 92259 5763
rect 92201 5723 92259 5729
rect 96617 5763 96675 5769
rect 96617 5729 96629 5763
rect 96663 5760 96675 5763
rect 98549 5763 98607 5769
rect 98549 5760 98561 5763
rect 96663 5732 98561 5760
rect 96663 5729 96675 5732
rect 96617 5723 96675 5729
rect 98549 5729 98561 5732
rect 98595 5760 98607 5763
rect 98638 5760 98644 5772
rect 98595 5732 98644 5760
rect 98595 5729 98607 5732
rect 98549 5723 98607 5729
rect 83921 5695 83979 5701
rect 83921 5661 83933 5695
rect 83967 5661 83979 5695
rect 83921 5655 83979 5661
rect 90269 5695 90327 5701
rect 90269 5661 90281 5695
rect 90315 5692 90327 5695
rect 92216 5692 92244 5723
rect 98638 5720 98644 5732
rect 98696 5720 98702 5772
rect 100665 5763 100723 5769
rect 100665 5760 100677 5763
rect 98748 5732 100677 5760
rect 92382 5692 92388 5704
rect 90315 5664 92388 5692
rect 90315 5661 90327 5664
rect 90269 5655 90327 5661
rect 92382 5652 92388 5664
rect 92440 5652 92446 5704
rect 98748 5701 98776 5732
rect 100665 5729 100677 5732
rect 100711 5760 100723 5763
rect 100754 5760 100760 5772
rect 100711 5732 100760 5760
rect 100711 5729 100723 5732
rect 100665 5723 100723 5729
rect 100754 5720 100760 5732
rect 100812 5720 100818 5772
rect 100849 5763 100907 5769
rect 100849 5729 100861 5763
rect 100895 5760 100907 5763
rect 102781 5763 102839 5769
rect 102781 5760 102793 5763
rect 100895 5732 102793 5760
rect 100895 5729 100907 5732
rect 100849 5723 100907 5729
rect 102781 5729 102793 5732
rect 102827 5760 102839 5763
rect 102962 5760 102968 5772
rect 102827 5732 102968 5760
rect 102827 5729 102839 5732
rect 102781 5723 102839 5729
rect 102962 5720 102968 5732
rect 103020 5720 103026 5772
rect 104912 5760 104940 5791
rect 105078 5788 105084 5800
rect 105136 5788 105142 5840
rect 104986 5760 104992 5772
rect 104912 5732 104992 5760
rect 104986 5720 104992 5732
rect 105044 5720 105050 5772
rect 98733 5695 98791 5701
rect 98733 5661 98745 5695
rect 98779 5661 98791 5695
rect 98733 5655 98791 5661
rect 77570 5556 77576 5568
rect 75411 5528 77576 5556
rect 75411 5525 75423 5528
rect 75365 5519 75423 5525
rect 77570 5516 77576 5528
rect 77628 5516 77634 5568
rect 85945 5559 86003 5565
rect 85945 5525 85957 5559
rect 85991 5556 86003 5559
rect 87785 5559 87843 5565
rect 87785 5556 87797 5559
rect 85991 5528 87797 5556
rect 85991 5525 86003 5528
rect 85945 5519 86003 5525
rect 87785 5525 87797 5528
rect 87831 5556 87843 5559
rect 88150 5556 88156 5568
rect 87831 5528 88156 5556
rect 87831 5525 87843 5528
rect 87785 5519 87843 5525
rect 88150 5516 88156 5528
rect 88208 5516 88214 5568
rect 1104 5466 106904 5488
rect 1104 5414 4042 5466
rect 4094 5414 4106 5466
rect 4158 5414 4170 5466
rect 4222 5414 4234 5466
rect 4286 5414 34762 5466
rect 34814 5414 34826 5466
rect 34878 5414 34890 5466
rect 34942 5414 34954 5466
rect 35006 5414 65482 5466
rect 65534 5414 65546 5466
rect 65598 5414 65610 5466
rect 65662 5414 65674 5466
rect 65726 5414 96202 5466
rect 96254 5414 96266 5466
rect 96318 5414 96330 5466
rect 96382 5414 96394 5466
rect 96446 5414 106904 5466
rect 1104 5392 106904 5414
rect 1118 5216 1124 5228
rect 1079 5188 1124 5216
rect 1118 5176 1124 5188
rect 1176 5176 1182 5228
rect 1302 5176 1308 5228
rect 1360 5216 1366 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 1360 5188 1409 5216
rect 1360 5176 1366 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 3234 5216 3240 5228
rect 3195 5188 3240 5216
rect 1397 5179 1455 5185
rect 3234 5176 3240 5188
rect 3292 5176 3298 5228
rect 3510 5216 3516 5228
rect 3471 5188 3516 5216
rect 3510 5176 3516 5188
rect 3568 5176 3574 5228
rect 5258 5176 5264 5228
rect 5316 5216 5322 5228
rect 5353 5219 5411 5225
rect 5353 5216 5365 5219
rect 5316 5188 5365 5216
rect 5316 5176 5322 5188
rect 5353 5185 5365 5188
rect 5399 5185 5411 5219
rect 5626 5216 5632 5228
rect 5587 5188 5632 5216
rect 5353 5179 5411 5185
rect 5626 5176 5632 5188
rect 5684 5176 5690 5228
rect 7374 5176 7380 5228
rect 7432 5216 7438 5228
rect 7469 5219 7527 5225
rect 7469 5216 7481 5219
rect 7432 5188 7481 5216
rect 7432 5176 7438 5188
rect 7469 5185 7481 5188
rect 7515 5185 7527 5219
rect 7469 5179 7527 5185
rect 7650 5176 7656 5228
rect 7708 5216 7714 5228
rect 7745 5219 7803 5225
rect 7745 5216 7757 5219
rect 7708 5188 7757 5216
rect 7708 5176 7714 5188
rect 7745 5185 7757 5188
rect 7791 5185 7803 5219
rect 9582 5216 9588 5228
rect 9543 5188 9588 5216
rect 7745 5179 7803 5185
rect 9582 5176 9588 5188
rect 9640 5176 9646 5228
rect 9858 5216 9864 5228
rect 9819 5188 9864 5216
rect 9858 5176 9864 5188
rect 9916 5176 9922 5228
rect 11698 5216 11704 5228
rect 11659 5188 11704 5216
rect 11698 5176 11704 5188
rect 11756 5176 11762 5228
rect 11882 5176 11888 5228
rect 11940 5216 11946 5228
rect 11977 5219 12035 5225
rect 11977 5216 11989 5219
rect 11940 5188 11989 5216
rect 11940 5176 11946 5188
rect 11977 5185 11989 5188
rect 12023 5185 12035 5219
rect 13814 5216 13820 5228
rect 13775 5188 13820 5216
rect 11977 5179 12035 5185
rect 13814 5176 13820 5188
rect 13872 5176 13878 5228
rect 14090 5216 14096 5228
rect 14051 5188 14096 5216
rect 14090 5176 14096 5188
rect 14148 5176 14154 5228
rect 15930 5216 15936 5228
rect 15891 5188 15936 5216
rect 15930 5176 15936 5188
rect 15988 5176 15994 5228
rect 16206 5216 16212 5228
rect 16167 5188 16212 5216
rect 16206 5176 16212 5188
rect 16264 5176 16270 5228
rect 18046 5216 18052 5228
rect 18007 5188 18052 5216
rect 18046 5176 18052 5188
rect 18104 5176 18110 5228
rect 18322 5216 18328 5228
rect 18283 5188 18328 5216
rect 18322 5176 18328 5188
rect 18380 5176 18386 5228
rect 20070 5176 20076 5228
rect 20128 5216 20134 5228
rect 20165 5219 20223 5225
rect 20165 5216 20177 5219
rect 20128 5188 20177 5216
rect 20128 5176 20134 5188
rect 20165 5185 20177 5188
rect 20211 5185 20223 5219
rect 20438 5216 20444 5228
rect 20399 5188 20444 5216
rect 20165 5179 20223 5185
rect 20438 5176 20444 5188
rect 20496 5176 20502 5228
rect 22186 5176 22192 5228
rect 22244 5216 22250 5228
rect 22281 5219 22339 5225
rect 22281 5216 22293 5219
rect 22244 5188 22293 5216
rect 22244 5176 22250 5188
rect 22281 5185 22293 5188
rect 22327 5185 22339 5219
rect 22281 5179 22339 5185
rect 22462 5176 22468 5228
rect 22520 5216 22526 5228
rect 22557 5219 22615 5225
rect 22557 5216 22569 5219
rect 22520 5188 22569 5216
rect 22520 5176 22526 5188
rect 22557 5185 22569 5188
rect 22603 5185 22615 5219
rect 22557 5179 22615 5185
rect 23750 5176 23756 5228
rect 23808 5216 23814 5228
rect 23934 5216 23940 5228
rect 23808 5188 23940 5216
rect 23808 5176 23814 5188
rect 23934 5176 23940 5188
rect 23992 5176 23998 5228
rect 24394 5216 24400 5228
rect 24355 5188 24400 5216
rect 24394 5176 24400 5188
rect 24452 5176 24458 5228
rect 24670 5216 24676 5228
rect 24631 5188 24676 5216
rect 24670 5176 24676 5188
rect 24728 5176 24734 5228
rect 26510 5216 26516 5228
rect 26471 5188 26516 5216
rect 26510 5176 26516 5188
rect 26568 5176 26574 5228
rect 26694 5176 26700 5228
rect 26752 5216 26758 5228
rect 26789 5219 26847 5225
rect 26789 5216 26801 5219
rect 26752 5188 26801 5216
rect 26752 5176 26758 5188
rect 26789 5185 26801 5188
rect 26835 5185 26847 5219
rect 28626 5216 28632 5228
rect 28587 5188 28632 5216
rect 26789 5179 26847 5185
rect 28626 5176 28632 5188
rect 28684 5176 28690 5228
rect 28810 5176 28816 5228
rect 28868 5216 28874 5228
rect 28905 5219 28963 5225
rect 28905 5216 28917 5219
rect 28868 5188 28917 5216
rect 28868 5176 28874 5188
rect 28905 5185 28917 5188
rect 28951 5185 28963 5219
rect 30742 5216 30748 5228
rect 30703 5188 30748 5216
rect 28905 5179 28963 5185
rect 30742 5176 30748 5188
rect 30800 5176 30806 5228
rect 31018 5216 31024 5228
rect 30979 5188 31024 5216
rect 31018 5176 31024 5188
rect 31076 5176 31082 5228
rect 32858 5216 32864 5228
rect 32819 5188 32864 5216
rect 32858 5176 32864 5188
rect 32916 5176 32922 5228
rect 33042 5176 33048 5228
rect 33100 5216 33106 5228
rect 33137 5219 33195 5225
rect 33137 5216 33149 5219
rect 33100 5188 33149 5216
rect 33100 5176 33106 5188
rect 33137 5185 33149 5188
rect 33183 5185 33195 5219
rect 35250 5216 35256 5228
rect 35211 5188 35256 5216
rect 33137 5179 33195 5185
rect 35250 5176 35256 5188
rect 35308 5176 35314 5228
rect 37090 5216 37096 5228
rect 37051 5188 37096 5216
rect 37090 5176 37096 5188
rect 37148 5176 37154 5228
rect 37366 5216 37372 5228
rect 37327 5188 37372 5216
rect 37366 5176 37372 5188
rect 37424 5176 37430 5228
rect 39206 5216 39212 5228
rect 39167 5188 39212 5216
rect 39206 5176 39212 5188
rect 39264 5176 39270 5228
rect 39482 5216 39488 5228
rect 39443 5188 39488 5216
rect 39482 5176 39488 5188
rect 39540 5176 39546 5228
rect 41230 5176 41236 5228
rect 41288 5216 41294 5228
rect 41325 5219 41383 5225
rect 41325 5216 41337 5219
rect 41288 5188 41337 5216
rect 41288 5176 41294 5188
rect 41325 5185 41337 5188
rect 41371 5185 41383 5219
rect 41598 5216 41604 5228
rect 41559 5188 41604 5216
rect 41325 5179 41383 5185
rect 41598 5176 41604 5188
rect 41656 5176 41662 5228
rect 43438 5216 43444 5228
rect 43399 5188 43444 5216
rect 43438 5176 43444 5188
rect 43496 5176 43502 5228
rect 43714 5216 43720 5228
rect 43675 5188 43720 5216
rect 43714 5176 43720 5188
rect 43772 5176 43778 5228
rect 45554 5216 45560 5228
rect 45515 5188 45560 5216
rect 45554 5176 45560 5188
rect 45612 5176 45618 5228
rect 45830 5216 45836 5228
rect 45791 5188 45836 5216
rect 45830 5176 45836 5188
rect 45888 5176 45894 5228
rect 47670 5216 47676 5228
rect 47631 5188 47676 5216
rect 47670 5176 47676 5188
rect 47728 5176 47734 5228
rect 47854 5176 47860 5228
rect 47912 5216 47918 5228
rect 47949 5219 48007 5225
rect 47949 5216 47961 5219
rect 47912 5188 47961 5216
rect 47912 5176 47918 5188
rect 47949 5185 47961 5188
rect 47995 5185 48007 5219
rect 49786 5216 49792 5228
rect 49747 5188 49792 5216
rect 47949 5179 48007 5185
rect 49786 5176 49792 5188
rect 49844 5176 49850 5228
rect 50062 5176 50068 5228
rect 50120 5216 50126 5228
rect 51902 5216 51908 5228
rect 50120 5188 50165 5216
rect 51863 5188 51908 5216
rect 50120 5176 50126 5188
rect 51902 5176 51908 5188
rect 51960 5176 51966 5228
rect 52178 5216 52184 5228
rect 52139 5188 52184 5216
rect 52178 5176 52184 5188
rect 52236 5176 52242 5228
rect 54018 5216 54024 5228
rect 53979 5188 54024 5216
rect 54018 5176 54024 5188
rect 54076 5176 54082 5228
rect 54202 5176 54208 5228
rect 54260 5216 54266 5228
rect 54297 5219 54355 5225
rect 54297 5216 54309 5219
rect 54260 5188 54309 5216
rect 54260 5176 54266 5188
rect 54297 5185 54309 5188
rect 54343 5185 54355 5219
rect 54297 5179 54355 5185
rect 56042 5176 56048 5228
rect 56100 5216 56106 5228
rect 56137 5219 56195 5225
rect 56137 5216 56149 5219
rect 56100 5188 56149 5216
rect 56100 5176 56106 5188
rect 56137 5185 56149 5188
rect 56183 5185 56195 5219
rect 56410 5216 56416 5228
rect 56371 5188 56416 5216
rect 56137 5179 56195 5185
rect 56410 5176 56416 5188
rect 56468 5176 56474 5228
rect 58158 5176 58164 5228
rect 58216 5216 58222 5228
rect 58253 5219 58311 5225
rect 58253 5216 58265 5219
rect 58216 5188 58265 5216
rect 58216 5176 58222 5188
rect 58253 5185 58265 5188
rect 58299 5185 58311 5219
rect 58253 5179 58311 5185
rect 58434 5176 58440 5228
rect 58492 5216 58498 5228
rect 58529 5219 58587 5225
rect 58529 5216 58541 5219
rect 58492 5188 58541 5216
rect 58492 5176 58498 5188
rect 58529 5185 58541 5188
rect 58575 5185 58587 5219
rect 58529 5179 58587 5185
rect 60550 5176 60556 5228
rect 60608 5216 60614 5228
rect 60645 5219 60703 5225
rect 60645 5216 60657 5219
rect 60608 5188 60657 5216
rect 60608 5176 60614 5188
rect 60645 5185 60657 5188
rect 60691 5185 60703 5219
rect 62482 5216 62488 5228
rect 62443 5188 62488 5216
rect 60645 5179 60703 5185
rect 62482 5176 62488 5188
rect 62540 5176 62546 5228
rect 62758 5216 62764 5228
rect 62719 5188 62764 5216
rect 62758 5176 62764 5188
rect 62816 5176 62822 5228
rect 64598 5216 64604 5228
rect 64559 5188 64604 5216
rect 64598 5176 64604 5188
rect 64656 5176 64662 5228
rect 64782 5176 64788 5228
rect 64840 5216 64846 5228
rect 64877 5219 64935 5225
rect 64877 5216 64889 5219
rect 64840 5188 64889 5216
rect 64840 5176 64846 5188
rect 64877 5185 64889 5188
rect 64923 5185 64935 5219
rect 66714 5216 66720 5228
rect 66675 5188 66720 5216
rect 64877 5179 64935 5185
rect 66714 5176 66720 5188
rect 66772 5176 66778 5228
rect 66990 5216 66996 5228
rect 66951 5188 66996 5216
rect 66990 5176 66996 5188
rect 67048 5176 67054 5228
rect 68830 5216 68836 5228
rect 68791 5188 68836 5216
rect 68830 5176 68836 5188
rect 68888 5176 68894 5228
rect 69106 5216 69112 5228
rect 69067 5188 69112 5216
rect 69106 5176 69112 5188
rect 69164 5176 69170 5228
rect 70854 5176 70860 5228
rect 70912 5216 70918 5228
rect 70949 5219 71007 5225
rect 70949 5216 70961 5219
rect 70912 5188 70961 5216
rect 70912 5176 70918 5188
rect 70949 5185 70961 5188
rect 70995 5185 71007 5219
rect 71222 5216 71228 5228
rect 71183 5188 71228 5216
rect 70949 5179 71007 5185
rect 71222 5176 71228 5188
rect 71280 5176 71286 5228
rect 72970 5176 72976 5228
rect 73028 5216 73034 5228
rect 73065 5219 73123 5225
rect 73065 5216 73077 5219
rect 73028 5188 73077 5216
rect 73028 5176 73034 5188
rect 73065 5185 73077 5188
rect 73111 5185 73123 5219
rect 73338 5216 73344 5228
rect 73299 5188 73344 5216
rect 73065 5179 73123 5185
rect 73338 5176 73344 5188
rect 73396 5176 73402 5228
rect 75086 5176 75092 5228
rect 75144 5216 75150 5228
rect 75181 5219 75239 5225
rect 75181 5216 75193 5219
rect 75144 5188 75193 5216
rect 75144 5176 75150 5188
rect 75181 5185 75193 5188
rect 75227 5185 75239 5219
rect 75454 5216 75460 5228
rect 75415 5188 75460 5216
rect 75181 5179 75239 5185
rect 75454 5176 75460 5188
rect 75512 5176 75518 5228
rect 77570 5216 77576 5228
rect 77531 5188 77576 5216
rect 77570 5176 77576 5188
rect 77628 5176 77634 5228
rect 79318 5176 79324 5228
rect 79376 5216 79382 5228
rect 79413 5219 79471 5225
rect 79413 5216 79425 5219
rect 79376 5188 79425 5216
rect 79376 5176 79382 5188
rect 79413 5185 79425 5188
rect 79459 5185 79471 5219
rect 79413 5179 79471 5185
rect 79594 5176 79600 5228
rect 79652 5216 79658 5228
rect 79689 5219 79747 5225
rect 79689 5216 79701 5219
rect 79652 5188 79701 5216
rect 79652 5176 79658 5188
rect 79689 5185 79701 5188
rect 79735 5185 79747 5219
rect 79689 5179 79747 5185
rect 81434 5176 81440 5228
rect 81492 5216 81498 5228
rect 81529 5219 81587 5225
rect 81529 5216 81541 5219
rect 81492 5188 81541 5216
rect 81492 5176 81498 5188
rect 81529 5185 81541 5188
rect 81575 5185 81587 5219
rect 81802 5216 81808 5228
rect 81763 5188 81808 5216
rect 81529 5179 81587 5185
rect 81802 5176 81808 5188
rect 81860 5176 81866 5228
rect 83550 5176 83556 5228
rect 83608 5216 83614 5228
rect 83645 5219 83703 5225
rect 83645 5216 83657 5219
rect 83608 5188 83657 5216
rect 83608 5176 83614 5188
rect 83645 5185 83657 5188
rect 83691 5185 83703 5219
rect 83918 5216 83924 5228
rect 83879 5188 83924 5216
rect 83645 5179 83703 5185
rect 83918 5176 83924 5188
rect 83976 5176 83982 5228
rect 85666 5176 85672 5228
rect 85724 5216 85730 5228
rect 85761 5219 85819 5225
rect 85761 5216 85773 5219
rect 85724 5188 85773 5216
rect 85724 5176 85730 5188
rect 85761 5185 85773 5188
rect 85807 5185 85819 5219
rect 86034 5216 86040 5228
rect 85995 5188 86040 5216
rect 85761 5179 85819 5185
rect 86034 5176 86040 5188
rect 86092 5176 86098 5228
rect 87782 5176 87788 5228
rect 87840 5216 87846 5228
rect 87877 5219 87935 5225
rect 87877 5216 87889 5219
rect 87840 5188 87889 5216
rect 87840 5176 87846 5188
rect 87877 5185 87889 5188
rect 87923 5185 87935 5219
rect 88150 5216 88156 5228
rect 88111 5188 88156 5216
rect 87877 5179 87935 5185
rect 88150 5176 88156 5188
rect 88208 5176 88214 5228
rect 89898 5176 89904 5228
rect 89956 5216 89962 5228
rect 89993 5219 90051 5225
rect 89993 5216 90005 5219
rect 89956 5188 90005 5216
rect 89956 5176 89962 5188
rect 89993 5185 90005 5188
rect 90039 5185 90051 5219
rect 90266 5216 90272 5228
rect 90227 5188 90272 5216
rect 89993 5179 90051 5185
rect 90266 5176 90272 5188
rect 90324 5176 90330 5228
rect 92014 5176 92020 5228
rect 92072 5216 92078 5228
rect 92109 5219 92167 5225
rect 92109 5216 92121 5219
rect 92072 5188 92121 5216
rect 92072 5176 92078 5188
rect 92109 5185 92121 5188
rect 92155 5185 92167 5219
rect 92382 5216 92388 5228
rect 92343 5188 92388 5216
rect 92109 5179 92167 5185
rect 92382 5176 92388 5188
rect 92440 5176 92446 5228
rect 94222 5216 94228 5228
rect 94183 5188 94228 5216
rect 94222 5176 94228 5188
rect 94280 5176 94286 5228
rect 94406 5176 94412 5228
rect 94464 5216 94470 5228
rect 94501 5219 94559 5225
rect 94501 5216 94513 5219
rect 94464 5188 94513 5216
rect 94464 5176 94470 5188
rect 94501 5185 94513 5188
rect 94547 5185 94559 5219
rect 94501 5179 94559 5185
rect 96062 5176 96068 5228
rect 96120 5216 96126 5228
rect 96341 5219 96399 5225
rect 96341 5216 96353 5219
rect 96120 5188 96353 5216
rect 96120 5176 96126 5188
rect 96341 5185 96353 5188
rect 96387 5185 96399 5219
rect 96341 5179 96399 5185
rect 96522 5176 96528 5228
rect 96580 5216 96586 5228
rect 96617 5219 96675 5225
rect 96617 5216 96629 5219
rect 96580 5188 96629 5216
rect 96580 5176 96586 5188
rect 96617 5185 96629 5188
rect 96663 5185 96675 5219
rect 96617 5179 96675 5185
rect 98362 5176 98368 5228
rect 98420 5216 98426 5228
rect 98457 5219 98515 5225
rect 98457 5216 98469 5219
rect 98420 5188 98469 5216
rect 98420 5176 98426 5188
rect 98457 5185 98469 5188
rect 98503 5185 98515 5219
rect 98457 5179 98515 5185
rect 98638 5176 98644 5228
rect 98696 5216 98702 5228
rect 98733 5219 98791 5225
rect 98733 5216 98745 5219
rect 98696 5188 98745 5216
rect 98696 5176 98702 5188
rect 98733 5185 98745 5188
rect 98779 5185 98791 5219
rect 98733 5179 98791 5185
rect 100478 5176 100484 5228
rect 100536 5216 100542 5228
rect 100573 5219 100631 5225
rect 100573 5216 100585 5219
rect 100536 5188 100585 5216
rect 100536 5176 100542 5188
rect 100573 5185 100585 5188
rect 100619 5185 100631 5219
rect 100573 5179 100631 5185
rect 100754 5176 100760 5228
rect 100812 5216 100818 5228
rect 100849 5219 100907 5225
rect 100849 5216 100861 5219
rect 100812 5188 100861 5216
rect 100812 5176 100818 5188
rect 100849 5185 100861 5188
rect 100895 5185 100907 5219
rect 102686 5216 102692 5228
rect 102647 5188 102692 5216
rect 100849 5179 100907 5185
rect 102686 5176 102692 5188
rect 102744 5176 102750 5228
rect 102962 5216 102968 5228
rect 102923 5188 102968 5216
rect 102962 5176 102968 5188
rect 103020 5176 103026 5228
rect 104802 5216 104808 5228
rect 104763 5188 104808 5216
rect 104802 5176 104808 5188
rect 104860 5176 104866 5228
rect 104986 5176 104992 5228
rect 105044 5216 105050 5228
rect 105081 5219 105139 5225
rect 105081 5216 105093 5219
rect 105044 5188 105093 5216
rect 105044 5176 105050 5188
rect 105081 5185 105093 5188
rect 105127 5185 105139 5219
rect 105081 5179 105139 5185
rect 34977 5151 35035 5157
rect 34977 5117 34989 5151
rect 35023 5148 35035 5151
rect 35066 5148 35072 5160
rect 35023 5120 35072 5148
rect 35023 5117 35035 5120
rect 34977 5111 35035 5117
rect 35066 5108 35072 5120
rect 35124 5108 35130 5160
rect 60366 5108 60372 5160
rect 60424 5148 60430 5160
rect 60424 5120 60469 5148
rect 60424 5108 60430 5120
rect 77294 5108 77300 5160
rect 77352 5148 77358 5160
rect 77352 5120 77397 5148
rect 77352 5108 77358 5120
rect 2501 5015 2559 5021
rect 2501 5012 2513 5015
rect 1044 4984 2513 5012
rect 1044 4672 1072 4984
rect 2501 4981 2513 4984
rect 2547 4981 2559 5015
rect 2501 4975 2559 4981
rect 3510 4972 3516 5024
rect 3568 5012 3574 5024
rect 4617 5015 4675 5021
rect 4617 5012 4629 5015
rect 3568 4984 4629 5012
rect 3568 4972 3574 4984
rect 4617 4981 4629 4984
rect 4663 4981 4675 5015
rect 4617 4975 4675 4981
rect 5626 4972 5632 5024
rect 5684 5012 5690 5024
rect 6733 5015 6791 5021
rect 6733 5012 6745 5015
rect 5684 4984 6745 5012
rect 5684 4972 5690 4984
rect 6733 4981 6745 4984
rect 6779 4981 6791 5015
rect 6733 4975 6791 4981
rect 7742 4972 7748 5024
rect 7800 5012 7806 5024
rect 8849 5015 8907 5021
rect 8849 5012 8861 5015
rect 7800 4984 8861 5012
rect 7800 4972 7806 4984
rect 8849 4981 8861 4984
rect 8895 4981 8907 5015
rect 8849 4975 8907 4981
rect 9858 4972 9864 5024
rect 9916 5012 9922 5024
rect 10965 5015 11023 5021
rect 10965 5012 10977 5015
rect 9916 4984 10977 5012
rect 9916 4972 9922 4984
rect 10965 4981 10977 4984
rect 11011 4981 11023 5015
rect 10965 4975 11023 4981
rect 11974 4972 11980 5024
rect 12032 5012 12038 5024
rect 13081 5015 13139 5021
rect 13081 5012 13093 5015
rect 12032 4984 13093 5012
rect 12032 4972 12038 4984
rect 13081 4981 13093 4984
rect 13127 4981 13139 5015
rect 13081 4975 13139 4981
rect 14090 4972 14096 5024
rect 14148 5012 14154 5024
rect 15197 5015 15255 5021
rect 15197 5012 15209 5015
rect 14148 4984 15209 5012
rect 14148 4972 14154 4984
rect 15197 4981 15209 4984
rect 15243 4981 15255 5015
rect 15197 4975 15255 4981
rect 16206 4972 16212 5024
rect 16264 5012 16270 5024
rect 17313 5015 17371 5021
rect 17313 5012 17325 5015
rect 16264 4984 17325 5012
rect 16264 4972 16270 4984
rect 17313 4981 17325 4984
rect 17359 4981 17371 5015
rect 17313 4975 17371 4981
rect 18322 4972 18328 5024
rect 18380 5012 18386 5024
rect 19429 5015 19487 5021
rect 19429 5012 19441 5015
rect 18380 4984 19441 5012
rect 18380 4972 18386 4984
rect 19429 4981 19441 4984
rect 19475 4981 19487 5015
rect 19429 4975 19487 4981
rect 20438 4972 20444 5024
rect 20496 5012 20502 5024
rect 21545 5015 21603 5021
rect 21545 5012 21557 5015
rect 20496 4984 21557 5012
rect 20496 4972 20502 4984
rect 21545 4981 21557 4984
rect 21591 4981 21603 5015
rect 21545 4975 21603 4981
rect 22554 4972 22560 5024
rect 22612 5012 22618 5024
rect 23661 5015 23719 5021
rect 23661 5012 23673 5015
rect 22612 4984 23673 5012
rect 22612 4972 22618 4984
rect 23661 4981 23673 4984
rect 23707 4981 23719 5015
rect 23661 4975 23719 4981
rect 24670 4972 24676 5024
rect 24728 5012 24734 5024
rect 25777 5015 25835 5021
rect 25777 5012 25789 5015
rect 24728 4984 25789 5012
rect 24728 4972 24734 4984
rect 25777 4981 25789 4984
rect 25823 4981 25835 5015
rect 25777 4975 25835 4981
rect 26786 4972 26792 5024
rect 26844 5012 26850 5024
rect 27893 5015 27951 5021
rect 27893 5012 27905 5015
rect 26844 4984 27905 5012
rect 26844 4972 26850 4984
rect 27893 4981 27905 4984
rect 27939 4981 27951 5015
rect 27893 4975 27951 4981
rect 28902 4972 28908 5024
rect 28960 5012 28966 5024
rect 30009 5015 30067 5021
rect 30009 5012 30021 5015
rect 28960 4984 30021 5012
rect 28960 4972 28966 4984
rect 30009 4981 30021 4984
rect 30055 4981 30067 5015
rect 30009 4975 30067 4981
rect 31018 4972 31024 5024
rect 31076 5012 31082 5024
rect 32125 5015 32183 5021
rect 32125 5012 32137 5015
rect 31076 4984 32137 5012
rect 31076 4972 31082 4984
rect 32125 4981 32137 4984
rect 32171 4981 32183 5015
rect 32125 4975 32183 4981
rect 33134 4972 33140 5024
rect 33192 5012 33198 5024
rect 34241 5015 34299 5021
rect 34241 5012 34253 5015
rect 33192 4984 34253 5012
rect 33192 4972 33198 4984
rect 34241 4981 34253 4984
rect 34287 4981 34299 5015
rect 34241 4975 34299 4981
rect 35250 4972 35256 5024
rect 35308 5012 35314 5024
rect 36357 5015 36415 5021
rect 36357 5012 36369 5015
rect 35308 4984 36369 5012
rect 35308 4972 35314 4984
rect 36357 4981 36369 4984
rect 36403 4981 36415 5015
rect 36357 4975 36415 4981
rect 37366 4972 37372 5024
rect 37424 5012 37430 5024
rect 38473 5015 38531 5021
rect 38473 5012 38485 5015
rect 37424 4984 38485 5012
rect 37424 4972 37430 4984
rect 38473 4981 38485 4984
rect 38519 4981 38531 5015
rect 38473 4975 38531 4981
rect 39482 4972 39488 5024
rect 39540 5012 39546 5024
rect 40589 5015 40647 5021
rect 40589 5012 40601 5015
rect 39540 4984 40601 5012
rect 39540 4972 39546 4984
rect 40589 4981 40601 4984
rect 40635 4981 40647 5015
rect 40589 4975 40647 4981
rect 41598 4972 41604 5024
rect 41656 5012 41662 5024
rect 42705 5015 42763 5021
rect 42705 5012 42717 5015
rect 41656 4984 42717 5012
rect 41656 4972 41662 4984
rect 42705 4981 42717 4984
rect 42751 4981 42763 5015
rect 42705 4975 42763 4981
rect 43714 4972 43720 5024
rect 43772 5012 43778 5024
rect 44821 5015 44879 5021
rect 44821 5012 44833 5015
rect 43772 4984 44833 5012
rect 43772 4972 43778 4984
rect 44821 4981 44833 4984
rect 44867 4981 44879 5015
rect 44821 4975 44879 4981
rect 45830 4972 45836 5024
rect 45888 5012 45894 5024
rect 46937 5015 46995 5021
rect 46937 5012 46949 5015
rect 45888 4984 46949 5012
rect 45888 4972 45894 4984
rect 46937 4981 46949 4984
rect 46983 4981 46995 5015
rect 46937 4975 46995 4981
rect 47946 4972 47952 5024
rect 48004 5012 48010 5024
rect 49053 5015 49111 5021
rect 49053 5012 49065 5015
rect 48004 4984 49065 5012
rect 48004 4972 48010 4984
rect 49053 4981 49065 4984
rect 49099 4981 49111 5015
rect 51166 5012 51172 5024
rect 51127 4984 51172 5012
rect 49053 4975 49111 4981
rect 51166 4972 51172 4984
rect 51224 4972 51230 5024
rect 52178 4972 52184 5024
rect 52236 5012 52242 5024
rect 53285 5015 53343 5021
rect 53285 5012 53297 5015
rect 52236 4984 53297 5012
rect 52236 4972 52242 4984
rect 53285 4981 53297 4984
rect 53331 4981 53343 5015
rect 53285 4975 53343 4981
rect 54294 4972 54300 5024
rect 54352 5012 54358 5024
rect 55401 5015 55459 5021
rect 55401 5012 55413 5015
rect 54352 4984 55413 5012
rect 54352 4972 54358 4984
rect 55401 4981 55413 4984
rect 55447 4981 55459 5015
rect 55401 4975 55459 4981
rect 56410 4972 56416 5024
rect 56468 5012 56474 5024
rect 57517 5015 57575 5021
rect 57517 5012 57529 5015
rect 56468 4984 57529 5012
rect 56468 4972 56474 4984
rect 57517 4981 57529 4984
rect 57563 4981 57575 5015
rect 57517 4975 57575 4981
rect 58526 4972 58532 5024
rect 58584 5012 58590 5024
rect 59633 5015 59691 5021
rect 59633 5012 59645 5015
rect 58584 4984 59645 5012
rect 58584 4972 58590 4984
rect 59633 4981 59645 4984
rect 59679 4981 59691 5015
rect 59633 4975 59691 4981
rect 60642 4972 60648 5024
rect 60700 5012 60706 5024
rect 61749 5015 61807 5021
rect 61749 5012 61761 5015
rect 60700 4984 61761 5012
rect 60700 4972 60706 4984
rect 61749 4981 61761 4984
rect 61795 4981 61807 5015
rect 61749 4975 61807 4981
rect 62758 4972 62764 5024
rect 62816 5012 62822 5024
rect 63865 5015 63923 5021
rect 63865 5012 63877 5015
rect 62816 4984 63877 5012
rect 62816 4972 62822 4984
rect 63865 4981 63877 4984
rect 63911 4981 63923 5015
rect 63865 4975 63923 4981
rect 64874 4972 64880 5024
rect 64932 5012 64938 5024
rect 65981 5015 66039 5021
rect 65981 5012 65993 5015
rect 64932 4984 65993 5012
rect 64932 4972 64938 4984
rect 65981 4981 65993 4984
rect 66027 4981 66039 5015
rect 65981 4975 66039 4981
rect 66990 4972 66996 5024
rect 67048 5012 67054 5024
rect 68097 5015 68155 5021
rect 68097 5012 68109 5015
rect 67048 4984 68109 5012
rect 67048 4972 67054 4984
rect 68097 4981 68109 4984
rect 68143 4981 68155 5015
rect 68097 4975 68155 4981
rect 69106 4972 69112 5024
rect 69164 5012 69170 5024
rect 70213 5015 70271 5021
rect 70213 5012 70225 5015
rect 69164 4984 70225 5012
rect 69164 4972 69170 4984
rect 70213 4981 70225 4984
rect 70259 4981 70271 5015
rect 70213 4975 70271 4981
rect 71222 4972 71228 5024
rect 71280 5012 71286 5024
rect 72329 5015 72387 5021
rect 72329 5012 72341 5015
rect 71280 4984 72341 5012
rect 71280 4972 71286 4984
rect 72329 4981 72341 4984
rect 72375 4981 72387 5015
rect 72329 4975 72387 4981
rect 73338 4972 73344 5024
rect 73396 5012 73402 5024
rect 74445 5015 74503 5021
rect 74445 5012 74457 5015
rect 73396 4984 74457 5012
rect 73396 4972 73402 4984
rect 74445 4981 74457 4984
rect 74491 4981 74503 5015
rect 74445 4975 74503 4981
rect 75454 4972 75460 5024
rect 75512 5012 75518 5024
rect 76561 5015 76619 5021
rect 76561 5012 76573 5015
rect 75512 4984 76573 5012
rect 75512 4972 75518 4984
rect 76561 4981 76573 4984
rect 76607 4981 76619 5015
rect 76561 4975 76619 4981
rect 77570 4972 77576 5024
rect 77628 5012 77634 5024
rect 78677 5015 78735 5021
rect 78677 5012 78689 5015
rect 77628 4984 78689 5012
rect 77628 4972 77634 4984
rect 78677 4981 78689 4984
rect 78723 4981 78735 5015
rect 78677 4975 78735 4981
rect 79686 4972 79692 5024
rect 79744 5012 79750 5024
rect 80793 5015 80851 5021
rect 80793 5012 80805 5015
rect 79744 4984 80805 5012
rect 79744 4972 79750 4984
rect 80793 4981 80805 4984
rect 80839 4981 80851 5015
rect 80793 4975 80851 4981
rect 81802 4972 81808 5024
rect 81860 5012 81866 5024
rect 82909 5015 82967 5021
rect 82909 5012 82921 5015
rect 81860 4984 82921 5012
rect 81860 4972 81866 4984
rect 82909 4981 82921 4984
rect 82955 4981 82967 5015
rect 82909 4975 82967 4981
rect 83918 4972 83924 5024
rect 83976 5012 83982 5024
rect 85025 5015 85083 5021
rect 85025 5012 85037 5015
rect 83976 4984 85037 5012
rect 83976 4972 83982 4984
rect 85025 4981 85037 4984
rect 85071 4981 85083 5015
rect 85025 4975 85083 4981
rect 86034 4972 86040 5024
rect 86092 5012 86098 5024
rect 87141 5015 87199 5021
rect 87141 5012 87153 5015
rect 86092 4984 87153 5012
rect 86092 4972 86098 4984
rect 87141 4981 87153 4984
rect 87187 4981 87199 5015
rect 87141 4975 87199 4981
rect 88150 4972 88156 5024
rect 88208 5012 88214 5024
rect 89257 5015 89315 5021
rect 89257 5012 89269 5015
rect 88208 4984 89269 5012
rect 88208 4972 88214 4984
rect 89257 4981 89269 4984
rect 89303 4981 89315 5015
rect 89257 4975 89315 4981
rect 90266 4972 90272 5024
rect 90324 5012 90330 5024
rect 91373 5015 91431 5021
rect 91373 5012 91385 5015
rect 90324 4984 91385 5012
rect 90324 4972 90330 4984
rect 91373 4981 91385 4984
rect 91419 4981 91431 5015
rect 91373 4975 91431 4981
rect 92382 4972 92388 5024
rect 92440 5012 92446 5024
rect 93489 5015 93547 5021
rect 93489 5012 93501 5015
rect 92440 4984 93501 5012
rect 92440 4972 92446 4984
rect 93489 4981 93501 4984
rect 93535 4981 93547 5015
rect 93489 4975 93547 4981
rect 94498 4972 94504 5024
rect 94556 5012 94562 5024
rect 95605 5015 95663 5021
rect 95605 5012 95617 5015
rect 94556 4984 95617 5012
rect 94556 4972 94562 4984
rect 95605 4981 95617 4984
rect 95651 4981 95663 5015
rect 95605 4975 95663 4981
rect 96614 4972 96620 5024
rect 96672 5012 96678 5024
rect 97721 5015 97779 5021
rect 97721 5012 97733 5015
rect 96672 4984 97733 5012
rect 96672 4972 96678 4984
rect 97721 4981 97733 4984
rect 97767 4981 97779 5015
rect 97721 4975 97779 4981
rect 98730 4972 98736 5024
rect 98788 5012 98794 5024
rect 99837 5015 99895 5021
rect 99837 5012 99849 5015
rect 98788 4984 99849 5012
rect 98788 4972 98794 4984
rect 99837 4981 99849 4984
rect 99883 4981 99895 5015
rect 99837 4975 99895 4981
rect 100846 4972 100852 5024
rect 100904 5012 100910 5024
rect 101953 5015 102011 5021
rect 101953 5012 101965 5015
rect 100904 4984 101965 5012
rect 100904 4972 100910 4984
rect 101953 4981 101965 4984
rect 101999 4981 102011 5015
rect 101953 4975 102011 4981
rect 102962 4972 102968 5024
rect 103020 5012 103026 5024
rect 104069 5015 104127 5021
rect 104069 5012 104081 5015
rect 103020 4984 104081 5012
rect 103020 4972 103026 4984
rect 104069 4981 104081 4984
rect 104115 4981 104127 5015
rect 104069 4975 104127 4981
rect 105078 4972 105084 5024
rect 105136 5012 105142 5024
rect 106185 5015 106243 5021
rect 106185 5012 106197 5015
rect 105136 4984 106197 5012
rect 105136 4972 105142 4984
rect 106185 4981 106197 4984
rect 106231 4981 106243 5015
rect 106185 4975 106243 4981
rect 1104 4922 106904 4944
rect 1104 4870 19402 4922
rect 19454 4870 19466 4922
rect 19518 4870 19530 4922
rect 19582 4870 19594 4922
rect 19646 4870 50122 4922
rect 50174 4870 50186 4922
rect 50238 4870 50250 4922
rect 50302 4870 50314 4922
rect 50366 4870 80842 4922
rect 80894 4870 80906 4922
rect 80958 4870 80970 4922
rect 81022 4870 81034 4922
rect 81086 4870 106904 4922
rect 1104 4848 106904 4870
rect 1397 4675 1455 4681
rect 1397 4672 1409 4675
rect 1044 4644 1409 4672
rect 1397 4641 1409 4644
rect 1443 4641 1455 4675
rect 3234 4672 3240 4684
rect 3195 4644 3240 4672
rect 1397 4635 1455 4641
rect 3234 4632 3240 4644
rect 3292 4632 3298 4684
rect 3510 4672 3516 4684
rect 3471 4644 3516 4672
rect 3510 4632 3516 4644
rect 3568 4632 3574 4684
rect 5258 4632 5264 4684
rect 5316 4672 5322 4684
rect 5353 4675 5411 4681
rect 5353 4672 5365 4675
rect 5316 4644 5365 4672
rect 5316 4632 5322 4644
rect 5353 4641 5365 4644
rect 5399 4641 5411 4675
rect 5626 4672 5632 4684
rect 5587 4644 5632 4672
rect 5353 4635 5411 4641
rect 5626 4632 5632 4644
rect 5684 4632 5690 4684
rect 7374 4632 7380 4684
rect 7432 4672 7438 4684
rect 7469 4675 7527 4681
rect 7469 4672 7481 4675
rect 7432 4644 7481 4672
rect 7432 4632 7438 4644
rect 7469 4641 7481 4644
rect 7515 4641 7527 4675
rect 7742 4672 7748 4684
rect 7703 4644 7748 4672
rect 7469 4635 7527 4641
rect 7742 4632 7748 4644
rect 7800 4632 7806 4684
rect 9582 4672 9588 4684
rect 9543 4644 9588 4672
rect 9582 4632 9588 4644
rect 9640 4632 9646 4684
rect 9858 4672 9864 4684
rect 9819 4644 9864 4672
rect 9858 4632 9864 4644
rect 9916 4632 9922 4684
rect 11698 4672 11704 4684
rect 11659 4644 11704 4672
rect 11698 4632 11704 4644
rect 11756 4632 11762 4684
rect 11974 4672 11980 4684
rect 11935 4644 11980 4672
rect 11974 4632 11980 4644
rect 12032 4632 12038 4684
rect 13814 4672 13820 4684
rect 13775 4644 13820 4672
rect 13814 4632 13820 4644
rect 13872 4632 13878 4684
rect 14090 4672 14096 4684
rect 14051 4644 14096 4672
rect 14090 4632 14096 4644
rect 14148 4632 14154 4684
rect 15930 4672 15936 4684
rect 15891 4644 15936 4672
rect 15930 4632 15936 4644
rect 15988 4632 15994 4684
rect 16206 4672 16212 4684
rect 16167 4644 16212 4672
rect 16206 4632 16212 4644
rect 16264 4632 16270 4684
rect 18046 4672 18052 4684
rect 18007 4644 18052 4672
rect 18046 4632 18052 4644
rect 18104 4632 18110 4684
rect 18322 4672 18328 4684
rect 18283 4644 18328 4672
rect 18322 4632 18328 4644
rect 18380 4632 18386 4684
rect 20070 4632 20076 4684
rect 20128 4672 20134 4684
rect 20165 4675 20223 4681
rect 20165 4672 20177 4675
rect 20128 4644 20177 4672
rect 20128 4632 20134 4644
rect 20165 4641 20177 4644
rect 20211 4641 20223 4675
rect 20438 4672 20444 4684
rect 20399 4644 20444 4672
rect 20165 4635 20223 4641
rect 20438 4632 20444 4644
rect 20496 4632 20502 4684
rect 22186 4632 22192 4684
rect 22244 4672 22250 4684
rect 22281 4675 22339 4681
rect 22281 4672 22293 4675
rect 22244 4644 22293 4672
rect 22244 4632 22250 4644
rect 22281 4641 22293 4644
rect 22327 4641 22339 4675
rect 22554 4672 22560 4684
rect 22515 4644 22560 4672
rect 22281 4635 22339 4641
rect 22554 4632 22560 4644
rect 22612 4632 22618 4684
rect 24394 4672 24400 4684
rect 24355 4644 24400 4672
rect 24394 4632 24400 4644
rect 24452 4632 24458 4684
rect 24670 4672 24676 4684
rect 24631 4644 24676 4672
rect 24670 4632 24676 4644
rect 24728 4632 24734 4684
rect 26510 4672 26516 4684
rect 26471 4644 26516 4672
rect 26510 4632 26516 4644
rect 26568 4632 26574 4684
rect 26786 4672 26792 4684
rect 26747 4644 26792 4672
rect 26786 4632 26792 4644
rect 26844 4632 26850 4684
rect 28626 4672 28632 4684
rect 28587 4644 28632 4672
rect 28626 4632 28632 4644
rect 28684 4632 28690 4684
rect 28902 4672 28908 4684
rect 28863 4644 28908 4672
rect 28902 4632 28908 4644
rect 28960 4632 28966 4684
rect 30742 4672 30748 4684
rect 30703 4644 30748 4672
rect 30742 4632 30748 4644
rect 30800 4632 30806 4684
rect 31018 4672 31024 4684
rect 30979 4644 31024 4672
rect 31018 4632 31024 4644
rect 31076 4632 31082 4684
rect 32858 4672 32864 4684
rect 32819 4644 32864 4672
rect 32858 4632 32864 4644
rect 32916 4632 32922 4684
rect 33134 4672 33140 4684
rect 33095 4644 33140 4672
rect 33134 4632 33140 4644
rect 33192 4632 33198 4684
rect 34977 4675 35035 4681
rect 34977 4641 34989 4675
rect 35023 4672 35035 4675
rect 35066 4672 35072 4684
rect 35023 4644 35072 4672
rect 35023 4641 35035 4644
rect 34977 4635 35035 4641
rect 35066 4632 35072 4644
rect 35124 4632 35130 4684
rect 35250 4672 35256 4684
rect 35211 4644 35256 4672
rect 35250 4632 35256 4644
rect 35308 4632 35314 4684
rect 37090 4672 37096 4684
rect 37051 4644 37096 4672
rect 37090 4632 37096 4644
rect 37148 4632 37154 4684
rect 37366 4672 37372 4684
rect 37327 4644 37372 4672
rect 37366 4632 37372 4644
rect 37424 4632 37430 4684
rect 39206 4672 39212 4684
rect 39167 4644 39212 4672
rect 39206 4632 39212 4644
rect 39264 4632 39270 4684
rect 39482 4672 39488 4684
rect 39443 4644 39488 4672
rect 39482 4632 39488 4644
rect 39540 4632 39546 4684
rect 41230 4632 41236 4684
rect 41288 4672 41294 4684
rect 41325 4675 41383 4681
rect 41325 4672 41337 4675
rect 41288 4644 41337 4672
rect 41288 4632 41294 4644
rect 41325 4641 41337 4644
rect 41371 4641 41383 4675
rect 41598 4672 41604 4684
rect 41559 4644 41604 4672
rect 41325 4635 41383 4641
rect 41598 4632 41604 4644
rect 41656 4632 41662 4684
rect 43438 4672 43444 4684
rect 43399 4644 43444 4672
rect 43438 4632 43444 4644
rect 43496 4632 43502 4684
rect 43714 4672 43720 4684
rect 43675 4644 43720 4672
rect 43714 4632 43720 4644
rect 43772 4632 43778 4684
rect 45554 4672 45560 4684
rect 45515 4644 45560 4672
rect 45554 4632 45560 4644
rect 45612 4632 45618 4684
rect 45830 4672 45836 4684
rect 45791 4644 45836 4672
rect 45830 4632 45836 4644
rect 45888 4632 45894 4684
rect 47670 4672 47676 4684
rect 47631 4644 47676 4672
rect 47670 4632 47676 4644
rect 47728 4632 47734 4684
rect 47946 4672 47952 4684
rect 47907 4644 47952 4672
rect 47946 4632 47952 4644
rect 48004 4632 48010 4684
rect 49786 4672 49792 4684
rect 49747 4644 49792 4672
rect 49786 4632 49792 4644
rect 49844 4632 49850 4684
rect 50065 4675 50123 4681
rect 50065 4641 50077 4675
rect 50111 4672 50123 4675
rect 51166 4672 51172 4684
rect 50111 4644 51172 4672
rect 50111 4641 50123 4644
rect 50065 4635 50123 4641
rect 51166 4632 51172 4644
rect 51224 4632 51230 4684
rect 51902 4672 51908 4684
rect 51863 4644 51908 4672
rect 51902 4632 51908 4644
rect 51960 4632 51966 4684
rect 52178 4672 52184 4684
rect 52139 4644 52184 4672
rect 52178 4632 52184 4644
rect 52236 4632 52242 4684
rect 54018 4672 54024 4684
rect 53979 4644 54024 4672
rect 54018 4632 54024 4644
rect 54076 4632 54082 4684
rect 54294 4672 54300 4684
rect 54255 4644 54300 4672
rect 54294 4632 54300 4644
rect 54352 4632 54358 4684
rect 56042 4632 56048 4684
rect 56100 4672 56106 4684
rect 56137 4675 56195 4681
rect 56137 4672 56149 4675
rect 56100 4644 56149 4672
rect 56100 4632 56106 4644
rect 56137 4641 56149 4644
rect 56183 4641 56195 4675
rect 56410 4672 56416 4684
rect 56371 4644 56416 4672
rect 56137 4635 56195 4641
rect 56410 4632 56416 4644
rect 56468 4632 56474 4684
rect 58158 4632 58164 4684
rect 58216 4672 58222 4684
rect 58253 4675 58311 4681
rect 58253 4672 58265 4675
rect 58216 4644 58265 4672
rect 58216 4632 58222 4644
rect 58253 4641 58265 4644
rect 58299 4641 58311 4675
rect 58526 4672 58532 4684
rect 58487 4644 58532 4672
rect 58253 4635 58311 4641
rect 58526 4632 58532 4644
rect 58584 4632 58590 4684
rect 60642 4672 60648 4684
rect 60603 4644 60648 4672
rect 60642 4632 60648 4644
rect 60700 4632 60706 4684
rect 62482 4672 62488 4684
rect 62443 4644 62488 4672
rect 62482 4632 62488 4644
rect 62540 4632 62546 4684
rect 62758 4672 62764 4684
rect 62719 4644 62764 4672
rect 62758 4632 62764 4644
rect 62816 4632 62822 4684
rect 64598 4672 64604 4684
rect 64559 4644 64604 4672
rect 64598 4632 64604 4644
rect 64656 4632 64662 4684
rect 64874 4672 64880 4684
rect 64835 4644 64880 4672
rect 64874 4632 64880 4644
rect 64932 4632 64938 4684
rect 66714 4672 66720 4684
rect 66675 4644 66720 4672
rect 66714 4632 66720 4644
rect 66772 4632 66778 4684
rect 66990 4672 66996 4684
rect 66951 4644 66996 4672
rect 66990 4632 66996 4644
rect 67048 4632 67054 4684
rect 68830 4672 68836 4684
rect 68791 4644 68836 4672
rect 68830 4632 68836 4644
rect 68888 4632 68894 4684
rect 69106 4672 69112 4684
rect 69067 4644 69112 4672
rect 69106 4632 69112 4644
rect 69164 4632 69170 4684
rect 70854 4632 70860 4684
rect 70912 4672 70918 4684
rect 70949 4675 71007 4681
rect 70949 4672 70961 4675
rect 70912 4644 70961 4672
rect 70912 4632 70918 4644
rect 70949 4641 70961 4644
rect 70995 4641 71007 4675
rect 71222 4672 71228 4684
rect 71183 4644 71228 4672
rect 70949 4635 71007 4641
rect 71222 4632 71228 4644
rect 71280 4632 71286 4684
rect 72970 4632 72976 4684
rect 73028 4672 73034 4684
rect 73065 4675 73123 4681
rect 73065 4672 73077 4675
rect 73028 4644 73077 4672
rect 73028 4632 73034 4644
rect 73065 4641 73077 4644
rect 73111 4641 73123 4675
rect 73338 4672 73344 4684
rect 73299 4644 73344 4672
rect 73065 4635 73123 4641
rect 73338 4632 73344 4644
rect 73396 4632 73402 4684
rect 75086 4632 75092 4684
rect 75144 4672 75150 4684
rect 75181 4675 75239 4681
rect 75181 4672 75193 4675
rect 75144 4644 75193 4672
rect 75144 4632 75150 4644
rect 75181 4641 75193 4644
rect 75227 4641 75239 4675
rect 75454 4672 75460 4684
rect 75415 4644 75460 4672
rect 75181 4635 75239 4641
rect 75454 4632 75460 4644
rect 75512 4632 75518 4684
rect 77570 4672 77576 4684
rect 77531 4644 77576 4672
rect 77570 4632 77576 4644
rect 77628 4632 77634 4684
rect 79318 4632 79324 4684
rect 79376 4672 79382 4684
rect 79413 4675 79471 4681
rect 79413 4672 79425 4675
rect 79376 4644 79425 4672
rect 79376 4632 79382 4644
rect 79413 4641 79425 4644
rect 79459 4641 79471 4675
rect 79686 4672 79692 4684
rect 79647 4644 79692 4672
rect 79413 4635 79471 4641
rect 79686 4632 79692 4644
rect 79744 4632 79750 4684
rect 81434 4632 81440 4684
rect 81492 4672 81498 4684
rect 81529 4675 81587 4681
rect 81529 4672 81541 4675
rect 81492 4644 81541 4672
rect 81492 4632 81498 4644
rect 81529 4641 81541 4644
rect 81575 4641 81587 4675
rect 81802 4672 81808 4684
rect 81763 4644 81808 4672
rect 81529 4635 81587 4641
rect 81802 4632 81808 4644
rect 81860 4632 81866 4684
rect 83550 4632 83556 4684
rect 83608 4672 83614 4684
rect 83645 4675 83703 4681
rect 83645 4672 83657 4675
rect 83608 4644 83657 4672
rect 83608 4632 83614 4644
rect 83645 4641 83657 4644
rect 83691 4641 83703 4675
rect 83918 4672 83924 4684
rect 83879 4644 83924 4672
rect 83645 4635 83703 4641
rect 83918 4632 83924 4644
rect 83976 4632 83982 4684
rect 85666 4632 85672 4684
rect 85724 4672 85730 4684
rect 85761 4675 85819 4681
rect 85761 4672 85773 4675
rect 85724 4644 85773 4672
rect 85724 4632 85730 4644
rect 85761 4641 85773 4644
rect 85807 4641 85819 4675
rect 86034 4672 86040 4684
rect 85995 4644 86040 4672
rect 85761 4635 85819 4641
rect 86034 4632 86040 4644
rect 86092 4632 86098 4684
rect 87782 4632 87788 4684
rect 87840 4672 87846 4684
rect 87877 4675 87935 4681
rect 87877 4672 87889 4675
rect 87840 4644 87889 4672
rect 87840 4632 87846 4644
rect 87877 4641 87889 4644
rect 87923 4641 87935 4675
rect 88150 4672 88156 4684
rect 88111 4644 88156 4672
rect 87877 4635 87935 4641
rect 88150 4632 88156 4644
rect 88208 4632 88214 4684
rect 89898 4632 89904 4684
rect 89956 4672 89962 4684
rect 89993 4675 90051 4681
rect 89993 4672 90005 4675
rect 89956 4644 90005 4672
rect 89956 4632 89962 4644
rect 89993 4641 90005 4644
rect 90039 4641 90051 4675
rect 90266 4672 90272 4684
rect 90227 4644 90272 4672
rect 89993 4635 90051 4641
rect 90266 4632 90272 4644
rect 90324 4632 90330 4684
rect 92014 4632 92020 4684
rect 92072 4672 92078 4684
rect 92109 4675 92167 4681
rect 92109 4672 92121 4675
rect 92072 4644 92121 4672
rect 92072 4632 92078 4644
rect 92109 4641 92121 4644
rect 92155 4641 92167 4675
rect 92382 4672 92388 4684
rect 92343 4644 92388 4672
rect 92109 4635 92167 4641
rect 92382 4632 92388 4644
rect 92440 4632 92446 4684
rect 94222 4672 94228 4684
rect 94183 4644 94228 4672
rect 94222 4632 94228 4644
rect 94280 4632 94286 4684
rect 94498 4672 94504 4684
rect 94459 4644 94504 4672
rect 94498 4632 94504 4644
rect 94556 4632 94562 4684
rect 96062 4632 96068 4684
rect 96120 4672 96126 4684
rect 96341 4675 96399 4681
rect 96341 4672 96353 4675
rect 96120 4644 96353 4672
rect 96120 4632 96126 4644
rect 96341 4641 96353 4644
rect 96387 4641 96399 4675
rect 96614 4672 96620 4684
rect 96575 4644 96620 4672
rect 96341 4635 96399 4641
rect 96614 4632 96620 4644
rect 96672 4632 96678 4684
rect 98362 4632 98368 4684
rect 98420 4672 98426 4684
rect 98457 4675 98515 4681
rect 98457 4672 98469 4675
rect 98420 4644 98469 4672
rect 98420 4632 98426 4644
rect 98457 4641 98469 4644
rect 98503 4641 98515 4675
rect 98730 4672 98736 4684
rect 98691 4644 98736 4672
rect 98457 4635 98515 4641
rect 98730 4632 98736 4644
rect 98788 4632 98794 4684
rect 100478 4632 100484 4684
rect 100536 4672 100542 4684
rect 100573 4675 100631 4681
rect 100573 4672 100585 4675
rect 100536 4644 100585 4672
rect 100536 4632 100542 4644
rect 100573 4641 100585 4644
rect 100619 4641 100631 4675
rect 100846 4672 100852 4684
rect 100807 4644 100852 4672
rect 100573 4635 100631 4641
rect 100846 4632 100852 4644
rect 100904 4632 100910 4684
rect 102686 4672 102692 4684
rect 102647 4644 102692 4672
rect 102686 4632 102692 4644
rect 102744 4632 102750 4684
rect 102962 4672 102968 4684
rect 102923 4644 102968 4672
rect 102962 4632 102968 4644
rect 103020 4632 103026 4684
rect 104802 4672 104808 4684
rect 104763 4644 104808 4672
rect 104802 4632 104808 4644
rect 104860 4632 104866 4684
rect 105078 4672 105084 4684
rect 105039 4644 105084 4672
rect 105078 4632 105084 4644
rect 105136 4632 105142 4684
rect 1118 4604 1124 4616
rect 1079 4576 1124 4604
rect 1118 4564 1124 4576
rect 1176 4564 1182 4616
rect 6270 4564 6276 4616
rect 6328 4604 6334 4616
rect 6733 4607 6791 4613
rect 6733 4604 6745 4607
rect 6328 4576 6745 4604
rect 6328 4564 6334 4576
rect 6733 4573 6745 4576
rect 6779 4573 6791 4607
rect 6733 4567 6791 4573
rect 27430 4564 27436 4616
rect 27488 4604 27494 4616
rect 27893 4607 27951 4613
rect 27893 4604 27905 4607
rect 27488 4576 27905 4604
rect 27488 4564 27494 4576
rect 27893 4573 27905 4576
rect 27939 4573 27951 4607
rect 27893 4567 27951 4573
rect 29546 4564 29552 4616
rect 29604 4604 29610 4616
rect 30009 4607 30067 4613
rect 30009 4604 30021 4607
rect 29604 4576 30021 4604
rect 29604 4564 29610 4576
rect 30009 4573 30021 4576
rect 30055 4573 30067 4607
rect 30009 4567 30067 4573
rect 38010 4564 38016 4616
rect 38068 4604 38074 4616
rect 38473 4607 38531 4613
rect 38473 4604 38485 4607
rect 38068 4576 38485 4604
rect 38068 4564 38074 4576
rect 38473 4573 38485 4576
rect 38519 4573 38531 4607
rect 38473 4567 38531 4573
rect 60366 4564 60372 4616
rect 60424 4604 60430 4616
rect 60424 4576 60469 4604
rect 60424 4564 60430 4576
rect 77294 4564 77300 4616
rect 77352 4604 77358 4616
rect 77352 4576 77397 4604
rect 77352 4564 77358 4576
rect 2222 4428 2228 4480
rect 2280 4468 2286 4480
rect 2501 4471 2559 4477
rect 2501 4468 2513 4471
rect 2280 4440 2513 4468
rect 2280 4428 2286 4440
rect 2501 4437 2513 4440
rect 2547 4437 2559 4471
rect 2501 4431 2559 4437
rect 4338 4428 4344 4480
rect 4396 4468 4402 4480
rect 4617 4471 4675 4477
rect 4617 4468 4629 4471
rect 4396 4440 4629 4468
rect 4396 4428 4402 4440
rect 4617 4437 4629 4440
rect 4663 4437 4675 4471
rect 4617 4431 4675 4437
rect 8202 4428 8208 4480
rect 8260 4468 8266 4480
rect 8849 4471 8907 4477
rect 8849 4468 8861 4471
rect 8260 4440 8861 4468
rect 8260 4428 8266 4440
rect 8849 4437 8861 4440
rect 8895 4437 8907 4471
rect 8849 4431 8907 4437
rect 10502 4428 10508 4480
rect 10560 4468 10566 4480
rect 10965 4471 11023 4477
rect 10965 4468 10977 4471
rect 10560 4440 10977 4468
rect 10560 4428 10566 4440
rect 10965 4437 10977 4440
rect 11011 4437 11023 4471
rect 10965 4431 11023 4437
rect 12618 4428 12624 4480
rect 12676 4468 12682 4480
rect 13081 4471 13139 4477
rect 13081 4468 13093 4471
rect 12676 4440 13093 4468
rect 12676 4428 12682 4440
rect 13081 4437 13093 4440
rect 13127 4437 13139 4471
rect 13081 4431 13139 4437
rect 14550 4428 14556 4480
rect 14608 4468 14614 4480
rect 15197 4471 15255 4477
rect 15197 4468 15209 4471
rect 14608 4440 15209 4468
rect 14608 4428 14614 4440
rect 15197 4437 15209 4440
rect 15243 4437 15255 4471
rect 15197 4431 15255 4437
rect 16850 4428 16856 4480
rect 16908 4468 16914 4480
rect 17313 4471 17371 4477
rect 17313 4468 17325 4471
rect 16908 4440 17325 4468
rect 16908 4428 16914 4440
rect 17313 4437 17325 4440
rect 17359 4437 17371 4471
rect 17313 4431 17371 4437
rect 18966 4428 18972 4480
rect 19024 4468 19030 4480
rect 19429 4471 19487 4477
rect 19429 4468 19441 4471
rect 19024 4440 19441 4468
rect 19024 4428 19030 4440
rect 19429 4437 19441 4440
rect 19475 4437 19487 4471
rect 19429 4431 19487 4437
rect 21082 4428 21088 4480
rect 21140 4468 21146 4480
rect 21545 4471 21603 4477
rect 21545 4468 21557 4471
rect 21140 4440 21557 4468
rect 21140 4428 21146 4440
rect 21545 4437 21557 4440
rect 21591 4437 21603 4471
rect 21545 4431 21603 4437
rect 23198 4428 23204 4480
rect 23256 4468 23262 4480
rect 23661 4471 23719 4477
rect 23661 4468 23673 4471
rect 23256 4440 23673 4468
rect 23256 4428 23262 4440
rect 23661 4437 23673 4440
rect 23707 4437 23719 4471
rect 23661 4431 23719 4437
rect 25314 4428 25320 4480
rect 25372 4468 25378 4480
rect 25777 4471 25835 4477
rect 25777 4468 25789 4471
rect 25372 4440 25789 4468
rect 25372 4428 25378 4440
rect 25777 4437 25789 4440
rect 25823 4437 25835 4471
rect 25777 4431 25835 4437
rect 31478 4428 31484 4480
rect 31536 4468 31542 4480
rect 32125 4471 32183 4477
rect 32125 4468 32137 4471
rect 31536 4440 32137 4468
rect 31536 4428 31542 4440
rect 32125 4437 32137 4440
rect 32171 4437 32183 4471
rect 32125 4431 32183 4437
rect 33778 4428 33784 4480
rect 33836 4468 33842 4480
rect 34241 4471 34299 4477
rect 34241 4468 34253 4471
rect 33836 4440 34253 4468
rect 33836 4428 33842 4440
rect 34241 4437 34253 4440
rect 34287 4437 34299 4471
rect 34241 4431 34299 4437
rect 35894 4428 35900 4480
rect 35952 4468 35958 4480
rect 36357 4471 36415 4477
rect 36357 4468 36369 4471
rect 35952 4440 36369 4468
rect 35952 4428 35958 4440
rect 36357 4437 36369 4440
rect 36403 4437 36415 4471
rect 36357 4431 36415 4437
rect 40126 4428 40132 4480
rect 40184 4468 40190 4480
rect 40589 4471 40647 4477
rect 40589 4468 40601 4471
rect 40184 4440 40601 4468
rect 40184 4428 40190 4440
rect 40589 4437 40601 4440
rect 40635 4437 40647 4471
rect 40589 4431 40647 4437
rect 42242 4428 42248 4480
rect 42300 4468 42306 4480
rect 42705 4471 42763 4477
rect 42705 4468 42717 4471
rect 42300 4440 42717 4468
rect 42300 4428 42306 4440
rect 42705 4437 42717 4440
rect 42751 4437 42763 4471
rect 42705 4431 42763 4437
rect 44358 4428 44364 4480
rect 44416 4468 44422 4480
rect 44821 4471 44879 4477
rect 44821 4468 44833 4471
rect 44416 4440 44833 4468
rect 44416 4428 44422 4440
rect 44821 4437 44833 4440
rect 44867 4437 44879 4471
rect 44821 4431 44879 4437
rect 46474 4428 46480 4480
rect 46532 4468 46538 4480
rect 46937 4471 46995 4477
rect 46937 4468 46949 4471
rect 46532 4440 46949 4468
rect 46532 4428 46538 4440
rect 46937 4437 46949 4440
rect 46983 4437 46995 4471
rect 46937 4431 46995 4437
rect 48406 4428 48412 4480
rect 48464 4468 48470 4480
rect 49053 4471 49111 4477
rect 49053 4468 49065 4471
rect 48464 4440 49065 4468
rect 48464 4428 48470 4440
rect 49053 4437 49065 4440
rect 49099 4437 49111 4471
rect 49053 4431 49111 4437
rect 50706 4428 50712 4480
rect 50764 4468 50770 4480
rect 51169 4471 51227 4477
rect 51169 4468 51181 4471
rect 50764 4440 51181 4468
rect 50764 4428 50770 4440
rect 51169 4437 51181 4440
rect 51215 4437 51227 4471
rect 51169 4431 51227 4437
rect 52822 4428 52828 4480
rect 52880 4468 52886 4480
rect 53285 4471 53343 4477
rect 53285 4468 53297 4471
rect 52880 4440 53297 4468
rect 52880 4428 52886 4440
rect 53285 4437 53297 4440
rect 53331 4437 53343 4471
rect 53285 4431 53343 4437
rect 54938 4428 54944 4480
rect 54996 4468 55002 4480
rect 55401 4471 55459 4477
rect 55401 4468 55413 4471
rect 54996 4440 55413 4468
rect 54996 4428 55002 4440
rect 55401 4437 55413 4440
rect 55447 4437 55459 4471
rect 55401 4431 55459 4437
rect 57054 4428 57060 4480
rect 57112 4468 57118 4480
rect 57517 4471 57575 4477
rect 57517 4468 57529 4471
rect 57112 4440 57529 4468
rect 57112 4428 57118 4440
rect 57517 4437 57529 4440
rect 57563 4437 57575 4471
rect 57517 4431 57575 4437
rect 59170 4428 59176 4480
rect 59228 4468 59234 4480
rect 59633 4471 59691 4477
rect 59633 4468 59645 4471
rect 59228 4440 59645 4468
rect 59228 4428 59234 4440
rect 59633 4437 59645 4440
rect 59679 4437 59691 4471
rect 59633 4431 59691 4437
rect 61286 4428 61292 4480
rect 61344 4468 61350 4480
rect 61749 4471 61807 4477
rect 61749 4468 61761 4471
rect 61344 4440 61761 4468
rect 61344 4428 61350 4440
rect 61749 4437 61761 4440
rect 61795 4437 61807 4471
rect 61749 4431 61807 4437
rect 63402 4428 63408 4480
rect 63460 4468 63466 4480
rect 63865 4471 63923 4477
rect 63865 4468 63877 4471
rect 63460 4440 63877 4468
rect 63460 4428 63466 4440
rect 63865 4437 63877 4440
rect 63911 4437 63923 4471
rect 63865 4431 63923 4437
rect 65334 4428 65340 4480
rect 65392 4468 65398 4480
rect 65981 4471 66039 4477
rect 65981 4468 65993 4471
rect 65392 4440 65993 4468
rect 65392 4428 65398 4440
rect 65981 4437 65993 4440
rect 66027 4437 66039 4471
rect 65981 4431 66039 4437
rect 67634 4428 67640 4480
rect 67692 4468 67698 4480
rect 68097 4471 68155 4477
rect 68097 4468 68109 4471
rect 67692 4440 68109 4468
rect 67692 4428 67698 4440
rect 68097 4437 68109 4440
rect 68143 4437 68155 4471
rect 68097 4431 68155 4437
rect 69750 4428 69756 4480
rect 69808 4468 69814 4480
rect 70213 4471 70271 4477
rect 70213 4468 70225 4471
rect 69808 4440 70225 4468
rect 69808 4428 69814 4440
rect 70213 4437 70225 4440
rect 70259 4437 70271 4471
rect 70213 4431 70271 4437
rect 71866 4428 71872 4480
rect 71924 4468 71930 4480
rect 72329 4471 72387 4477
rect 72329 4468 72341 4471
rect 71924 4440 72341 4468
rect 71924 4428 71930 4440
rect 72329 4437 72341 4440
rect 72375 4437 72387 4471
rect 72329 4431 72387 4437
rect 73982 4428 73988 4480
rect 74040 4468 74046 4480
rect 74445 4471 74503 4477
rect 74445 4468 74457 4471
rect 74040 4440 74457 4468
rect 74040 4428 74046 4440
rect 74445 4437 74457 4440
rect 74491 4437 74503 4471
rect 76558 4468 76564 4480
rect 76519 4440 76564 4468
rect 74445 4431 74503 4437
rect 76558 4428 76564 4440
rect 76616 4428 76622 4480
rect 78858 4468 78864 4480
rect 78819 4440 78864 4468
rect 78858 4428 78864 4440
rect 78916 4428 78922 4480
rect 80977 4471 81035 4477
rect 80977 4437 80989 4471
rect 81023 4468 81035 4471
rect 81158 4468 81164 4480
rect 81023 4440 81164 4468
rect 81023 4437 81035 4440
rect 80977 4431 81035 4437
rect 81158 4428 81164 4440
rect 81216 4428 81222 4480
rect 82630 4428 82636 4480
rect 82688 4468 82694 4480
rect 82909 4471 82967 4477
rect 82909 4468 82921 4471
rect 82688 4440 82921 4468
rect 82688 4428 82694 4440
rect 82909 4437 82921 4440
rect 82955 4437 82967 4471
rect 82909 4431 82967 4437
rect 84654 4428 84660 4480
rect 84712 4468 84718 4480
rect 85025 4471 85083 4477
rect 85025 4468 85037 4471
rect 84712 4440 85037 4468
rect 84712 4428 84718 4440
rect 85025 4437 85037 4440
rect 85071 4437 85083 4471
rect 85025 4431 85083 4437
rect 86862 4428 86868 4480
rect 86920 4468 86926 4480
rect 87141 4471 87199 4477
rect 87141 4468 87153 4471
rect 86920 4440 87153 4468
rect 86920 4428 86926 4440
rect 87141 4437 87153 4440
rect 87187 4437 87199 4471
rect 89254 4468 89260 4480
rect 89215 4440 89260 4468
rect 87141 4431 87199 4437
rect 89254 4428 89260 4440
rect 89312 4428 89318 4480
rect 91278 4428 91284 4480
rect 91336 4468 91342 4480
rect 91373 4471 91431 4477
rect 91373 4468 91385 4471
rect 91336 4440 91385 4468
rect 91336 4428 91342 4440
rect 91373 4437 91385 4440
rect 91419 4437 91431 4471
rect 93670 4468 93676 4480
rect 93631 4440 93676 4468
rect 91373 4431 91431 4437
rect 93670 4428 93676 4440
rect 93728 4428 93734 4480
rect 95786 4468 95792 4480
rect 95747 4440 95792 4468
rect 95786 4428 95792 4440
rect 95844 4428 95850 4480
rect 97905 4471 97963 4477
rect 97905 4437 97917 4471
rect 97951 4468 97963 4471
rect 97994 4468 98000 4480
rect 97951 4440 98000 4468
rect 97951 4437 97963 4440
rect 97905 4431 97963 4437
rect 97994 4428 98000 4440
rect 98052 4428 98058 4480
rect 99374 4428 99380 4480
rect 99432 4468 99438 4480
rect 99837 4471 99895 4477
rect 99837 4468 99849 4471
rect 99432 4440 99849 4468
rect 99432 4428 99438 4440
rect 99837 4437 99849 4440
rect 99883 4437 99895 4471
rect 99837 4431 99895 4437
rect 101582 4428 101588 4480
rect 101640 4468 101646 4480
rect 101953 4471 102011 4477
rect 101953 4468 101965 4471
rect 101640 4440 101965 4468
rect 101640 4428 101646 4440
rect 101953 4437 101965 4440
rect 101999 4437 102011 4471
rect 101953 4431 102011 4437
rect 103790 4428 103796 4480
rect 103848 4468 103854 4480
rect 104069 4471 104127 4477
rect 104069 4468 104081 4471
rect 103848 4440 104081 4468
rect 103848 4428 103854 4440
rect 104069 4437 104081 4440
rect 104115 4437 104127 4471
rect 104069 4431 104127 4437
rect 105998 4428 106004 4480
rect 106056 4468 106062 4480
rect 106185 4471 106243 4477
rect 106185 4468 106197 4471
rect 106056 4440 106197 4468
rect 106056 4428 106062 4440
rect 106185 4437 106197 4440
rect 106231 4437 106243 4471
rect 106185 4431 106243 4437
rect 1104 4378 106904 4400
rect 1104 4326 4042 4378
rect 4094 4326 4106 4378
rect 4158 4326 4170 4378
rect 4222 4326 4234 4378
rect 4286 4326 34762 4378
rect 34814 4326 34826 4378
rect 34878 4326 34890 4378
rect 34942 4326 34954 4378
rect 35006 4326 65482 4378
rect 65534 4326 65546 4378
rect 65598 4326 65610 4378
rect 65662 4326 65674 4378
rect 65726 4326 96202 4378
rect 96254 4326 96266 4378
rect 96318 4326 96330 4378
rect 96382 4326 96394 4378
rect 96446 4326 106904 4378
rect 1104 4304 106904 4326
rect 20070 4156 20076 4208
rect 20128 4196 20134 4208
rect 20128 4168 20208 4196
rect 20128 4156 20134 4168
rect 1118 4128 1124 4140
rect 1079 4100 1124 4128
rect 1118 4088 1124 4100
rect 1176 4088 1182 4140
rect 3234 4128 3240 4140
rect 3195 4100 3240 4128
rect 3234 4088 3240 4100
rect 3292 4088 3298 4140
rect 5258 4088 5264 4140
rect 5316 4128 5322 4140
rect 5353 4131 5411 4137
rect 5353 4128 5365 4131
rect 5316 4100 5365 4128
rect 5316 4088 5322 4100
rect 5353 4097 5365 4100
rect 5399 4097 5411 4131
rect 5353 4091 5411 4097
rect 7374 4088 7380 4140
rect 7432 4128 7438 4140
rect 7469 4131 7527 4137
rect 7469 4128 7481 4131
rect 7432 4100 7481 4128
rect 7432 4088 7438 4100
rect 7469 4097 7481 4100
rect 7515 4097 7527 4131
rect 9582 4128 9588 4140
rect 9543 4100 9588 4128
rect 7469 4091 7527 4097
rect 9582 4088 9588 4100
rect 9640 4088 9646 4140
rect 11698 4128 11704 4140
rect 11659 4100 11704 4128
rect 11698 4088 11704 4100
rect 11756 4088 11762 4140
rect 13814 4128 13820 4140
rect 13775 4100 13820 4128
rect 13814 4088 13820 4100
rect 13872 4088 13878 4140
rect 15930 4128 15936 4140
rect 15891 4100 15936 4128
rect 15930 4088 15936 4100
rect 15988 4088 15994 4140
rect 18046 4128 18052 4140
rect 18007 4100 18052 4128
rect 18046 4088 18052 4100
rect 18104 4088 18110 4140
rect 20180 4137 20208 4168
rect 58158 4156 58164 4208
rect 58216 4196 58222 4208
rect 58216 4168 58296 4196
rect 58216 4156 58222 4168
rect 20165 4131 20223 4137
rect 20165 4097 20177 4131
rect 20211 4097 20223 4131
rect 20165 4091 20223 4097
rect 22186 4088 22192 4140
rect 22244 4128 22250 4140
rect 22281 4131 22339 4137
rect 22281 4128 22293 4131
rect 22244 4100 22293 4128
rect 22244 4088 22250 4100
rect 22281 4097 22293 4100
rect 22327 4097 22339 4131
rect 24394 4128 24400 4140
rect 24355 4100 24400 4128
rect 22281 4091 22339 4097
rect 24394 4088 24400 4100
rect 24452 4088 24458 4140
rect 26510 4128 26516 4140
rect 26471 4100 26516 4128
rect 26510 4088 26516 4100
rect 26568 4088 26574 4140
rect 28626 4128 28632 4140
rect 28587 4100 28632 4128
rect 28626 4088 28632 4100
rect 28684 4088 28690 4140
rect 30742 4128 30748 4140
rect 30703 4100 30748 4128
rect 30742 4088 30748 4100
rect 30800 4088 30806 4140
rect 32858 4128 32864 4140
rect 32819 4100 32864 4128
rect 32858 4088 32864 4100
rect 32916 4088 32922 4140
rect 37090 4128 37096 4140
rect 37051 4100 37096 4128
rect 37090 4088 37096 4100
rect 37148 4088 37154 4140
rect 39206 4128 39212 4140
rect 39167 4100 39212 4128
rect 39206 4088 39212 4100
rect 39264 4088 39270 4140
rect 41230 4088 41236 4140
rect 41288 4128 41294 4140
rect 41325 4131 41383 4137
rect 41325 4128 41337 4131
rect 41288 4100 41337 4128
rect 41288 4088 41294 4100
rect 41325 4097 41337 4100
rect 41371 4097 41383 4131
rect 43438 4128 43444 4140
rect 43399 4100 43444 4128
rect 41325 4091 41383 4097
rect 43438 4088 43444 4100
rect 43496 4088 43502 4140
rect 45554 4128 45560 4140
rect 45515 4100 45560 4128
rect 45554 4088 45560 4100
rect 45612 4088 45618 4140
rect 47670 4128 47676 4140
rect 47631 4100 47676 4128
rect 47670 4088 47676 4100
rect 47728 4088 47734 4140
rect 49786 4128 49792 4140
rect 49747 4100 49792 4128
rect 49786 4088 49792 4100
rect 49844 4088 49850 4140
rect 51902 4128 51908 4140
rect 51863 4100 51908 4128
rect 51902 4088 51908 4100
rect 51960 4088 51966 4140
rect 54018 4128 54024 4140
rect 53979 4100 54024 4128
rect 54018 4088 54024 4100
rect 54076 4088 54082 4140
rect 58268 4137 58296 4168
rect 70854 4156 70860 4208
rect 70912 4196 70918 4208
rect 70912 4168 70992 4196
rect 70912 4156 70918 4168
rect 58253 4131 58311 4137
rect 58253 4097 58265 4131
rect 58299 4097 58311 4131
rect 62482 4128 62488 4140
rect 62443 4100 62488 4128
rect 58253 4091 58311 4097
rect 62482 4088 62488 4100
rect 62540 4088 62546 4140
rect 64598 4128 64604 4140
rect 64559 4100 64604 4128
rect 64598 4088 64604 4100
rect 64656 4088 64662 4140
rect 66714 4128 66720 4140
rect 66675 4100 66720 4128
rect 66714 4088 66720 4100
rect 66772 4088 66778 4140
rect 68830 4128 68836 4140
rect 68791 4100 68836 4128
rect 68830 4088 68836 4100
rect 68888 4088 68894 4140
rect 70964 4137 70992 4168
rect 75086 4156 75092 4208
rect 75144 4196 75150 4208
rect 75144 4168 75224 4196
rect 75144 4156 75150 4168
rect 70949 4131 71007 4137
rect 70949 4097 70961 4131
rect 70995 4097 71007 4131
rect 73062 4128 73068 4140
rect 73023 4100 73068 4128
rect 70949 4091 71007 4097
rect 73062 4088 73068 4100
rect 73120 4088 73126 4140
rect 75196 4137 75224 4168
rect 83550 4156 83556 4208
rect 83608 4196 83614 4208
rect 83608 4168 83688 4196
rect 83608 4156 83614 4168
rect 75181 4131 75239 4137
rect 75181 4097 75193 4131
rect 75227 4097 75239 4131
rect 75181 4091 75239 4097
rect 79318 4088 79324 4140
rect 79376 4128 79382 4140
rect 79413 4131 79471 4137
rect 79413 4128 79425 4131
rect 79376 4100 79425 4128
rect 79376 4088 79382 4100
rect 79413 4097 79425 4100
rect 79459 4097 79471 4131
rect 81526 4128 81532 4140
rect 81487 4100 81532 4128
rect 79413 4091 79471 4097
rect 81526 4088 81532 4100
rect 81584 4088 81590 4140
rect 83660 4137 83688 4168
rect 87782 4156 87788 4208
rect 87840 4196 87846 4208
rect 87840 4168 87920 4196
rect 87840 4156 87846 4168
rect 83645 4131 83703 4137
rect 83645 4097 83657 4131
rect 83691 4097 83703 4131
rect 85758 4128 85764 4140
rect 85719 4100 85764 4128
rect 83645 4091 83703 4097
rect 85758 4088 85764 4100
rect 85816 4088 85822 4140
rect 87892 4137 87920 4168
rect 87877 4131 87935 4137
rect 87877 4097 87889 4131
rect 87923 4097 87935 4131
rect 87877 4091 87935 4097
rect 92014 4088 92020 4140
rect 92072 4128 92078 4140
rect 92109 4131 92167 4137
rect 92109 4128 92121 4131
rect 92072 4100 92121 4128
rect 92072 4088 92078 4100
rect 92109 4097 92121 4100
rect 92155 4097 92167 4131
rect 94222 4128 94228 4140
rect 94183 4100 94228 4128
rect 92109 4091 92167 4097
rect 94222 4088 94228 4100
rect 94280 4088 94286 4140
rect 96062 4088 96068 4140
rect 96120 4128 96126 4140
rect 96341 4131 96399 4137
rect 96341 4128 96353 4131
rect 96120 4100 96353 4128
rect 96120 4088 96126 4100
rect 96341 4097 96353 4100
rect 96387 4097 96399 4131
rect 96341 4091 96399 4097
rect 98362 4088 98368 4140
rect 98420 4128 98426 4140
rect 98457 4131 98515 4137
rect 98457 4128 98469 4131
rect 98420 4100 98469 4128
rect 98420 4088 98426 4100
rect 98457 4097 98469 4100
rect 98503 4097 98515 4131
rect 98457 4091 98515 4097
rect 100478 4088 100484 4140
rect 100536 4128 100542 4140
rect 100573 4131 100631 4137
rect 100573 4128 100585 4131
rect 100536 4100 100585 4128
rect 100536 4088 100542 4100
rect 100573 4097 100585 4100
rect 100619 4097 100631 4131
rect 102686 4128 102692 4140
rect 102647 4100 102692 4128
rect 100573 4091 100631 4097
rect 102686 4088 102692 4100
rect 102744 4088 102750 4140
rect 104802 4128 104808 4140
rect 104763 4100 104808 4128
rect 104802 4088 104808 4100
rect 104860 4088 104866 4140
rect 1397 4063 1455 4069
rect 1397 4029 1409 4063
rect 1443 4060 1455 4063
rect 2498 4060 2504 4072
rect 1443 4032 2504 4060
rect 1443 4029 1455 4032
rect 1397 4023 1455 4029
rect 2498 4020 2504 4032
rect 2556 4020 2562 4072
rect 3513 4063 3571 4069
rect 3513 4029 3525 4063
rect 3559 4060 3571 4063
rect 3878 4060 3884 4072
rect 3559 4032 3884 4060
rect 3559 4029 3571 4032
rect 3513 4023 3571 4029
rect 3878 4020 3884 4032
rect 3936 4020 3942 4072
rect 5629 4063 5687 4069
rect 5629 4029 5641 4063
rect 5675 4060 5687 4063
rect 5994 4060 6000 4072
rect 5675 4032 6000 4060
rect 5675 4029 5687 4032
rect 5629 4023 5687 4029
rect 5994 4020 6000 4032
rect 6052 4020 6058 4072
rect 7745 4063 7803 4069
rect 7745 4029 7757 4063
rect 7791 4060 7803 4063
rect 8110 4060 8116 4072
rect 7791 4032 8116 4060
rect 7791 4029 7803 4032
rect 7745 4023 7803 4029
rect 8110 4020 8116 4032
rect 8168 4020 8174 4072
rect 9861 4063 9919 4069
rect 9861 4029 9873 4063
rect 9907 4060 9919 4063
rect 10962 4060 10968 4072
rect 9907 4032 10968 4060
rect 9907 4029 9919 4032
rect 9861 4023 9919 4029
rect 10962 4020 10968 4032
rect 11020 4020 11026 4072
rect 11977 4063 12035 4069
rect 11977 4029 11989 4063
rect 12023 4060 12035 4063
rect 13078 4060 13084 4072
rect 12023 4032 13084 4060
rect 12023 4029 12035 4032
rect 11977 4023 12035 4029
rect 13078 4020 13084 4032
rect 13136 4020 13142 4072
rect 14093 4063 14151 4069
rect 14093 4029 14105 4063
rect 14139 4060 14151 4063
rect 15194 4060 15200 4072
rect 14139 4032 15200 4060
rect 14139 4029 14151 4032
rect 14093 4023 14151 4029
rect 15194 4020 15200 4032
rect 15252 4020 15258 4072
rect 16209 4063 16267 4069
rect 16209 4029 16221 4063
rect 16255 4060 16267 4063
rect 17310 4060 17316 4072
rect 16255 4032 17316 4060
rect 16255 4029 16267 4032
rect 16209 4023 16267 4029
rect 17310 4020 17316 4032
rect 17368 4020 17374 4072
rect 18325 4063 18383 4069
rect 18325 4029 18337 4063
rect 18371 4060 18383 4063
rect 18414 4060 18420 4072
rect 18371 4032 18420 4060
rect 18371 4029 18383 4032
rect 18325 4023 18383 4029
rect 18414 4020 18420 4032
rect 18472 4020 18478 4072
rect 20441 4063 20499 4069
rect 20441 4029 20453 4063
rect 20487 4060 20499 4063
rect 21082 4060 21088 4072
rect 20487 4032 21088 4060
rect 20487 4029 20499 4032
rect 20441 4023 20499 4029
rect 21082 4020 21088 4032
rect 21140 4020 21146 4072
rect 22557 4063 22615 4069
rect 22557 4029 22569 4063
rect 22603 4060 22615 4063
rect 22922 4060 22928 4072
rect 22603 4032 22928 4060
rect 22603 4029 22615 4032
rect 22557 4023 22615 4029
rect 22922 4020 22928 4032
rect 22980 4020 22986 4072
rect 24673 4063 24731 4069
rect 24673 4029 24685 4063
rect 24719 4060 24731 4063
rect 25038 4060 25044 4072
rect 24719 4032 25044 4060
rect 24719 4029 24731 4032
rect 24673 4023 24731 4029
rect 25038 4020 25044 4032
rect 25096 4020 25102 4072
rect 26789 4063 26847 4069
rect 26789 4029 26801 4063
rect 26835 4060 26847 4063
rect 27890 4060 27896 4072
rect 26835 4032 27896 4060
rect 26835 4029 26847 4032
rect 26789 4023 26847 4029
rect 27890 4020 27896 4032
rect 27948 4020 27954 4072
rect 28905 4063 28963 4069
rect 28905 4029 28917 4063
rect 28951 4060 28963 4063
rect 30006 4060 30012 4072
rect 28951 4032 30012 4060
rect 28951 4029 28963 4032
rect 28905 4023 28963 4029
rect 30006 4020 30012 4032
rect 30064 4020 30070 4072
rect 31021 4063 31079 4069
rect 31021 4029 31033 4063
rect 31067 4060 31079 4063
rect 32122 4060 32128 4072
rect 31067 4032 32128 4060
rect 31067 4029 31079 4032
rect 31021 4023 31079 4029
rect 32122 4020 32128 4032
rect 32180 4020 32186 4072
rect 33137 4063 33195 4069
rect 33137 4029 33149 4063
rect 33183 4060 33195 4063
rect 34238 4060 34244 4072
rect 33183 4032 34244 4060
rect 33183 4029 33195 4032
rect 33137 4023 33195 4029
rect 34238 4020 34244 4032
rect 34296 4020 34302 4072
rect 34977 4063 35035 4069
rect 34977 4029 34989 4063
rect 35023 4060 35035 4063
rect 35066 4060 35072 4072
rect 35023 4032 35072 4060
rect 35023 4029 35035 4032
rect 34977 4023 35035 4029
rect 35066 4020 35072 4032
rect 35124 4020 35130 4072
rect 35253 4063 35311 4069
rect 35253 4029 35265 4063
rect 35299 4060 35311 4063
rect 35618 4060 35624 4072
rect 35299 4032 35624 4060
rect 35299 4029 35311 4032
rect 35253 4023 35311 4029
rect 35618 4020 35624 4032
rect 35676 4020 35682 4072
rect 37369 4063 37427 4069
rect 37369 4029 37381 4063
rect 37415 4060 37427 4063
rect 37734 4060 37740 4072
rect 37415 4032 37740 4060
rect 37415 4029 37427 4032
rect 37369 4023 37427 4029
rect 37734 4020 37740 4032
rect 37792 4020 37798 4072
rect 39485 4063 39543 4069
rect 39485 4029 39497 4063
rect 39531 4060 39543 4063
rect 39942 4060 39948 4072
rect 39531 4032 39948 4060
rect 39531 4029 39543 4032
rect 39485 4023 39543 4029
rect 39942 4020 39948 4032
rect 40000 4020 40006 4072
rect 41601 4063 41659 4069
rect 41601 4029 41613 4063
rect 41647 4060 41659 4063
rect 41966 4060 41972 4072
rect 41647 4032 41972 4060
rect 41647 4029 41659 4032
rect 41601 4023 41659 4029
rect 41966 4020 41972 4032
rect 42024 4020 42030 4072
rect 43717 4063 43775 4069
rect 43717 4029 43729 4063
rect 43763 4060 43775 4063
rect 44818 4060 44824 4072
rect 43763 4032 44824 4060
rect 43763 4029 43775 4032
rect 43717 4023 43775 4029
rect 44818 4020 44824 4032
rect 44876 4020 44882 4072
rect 45833 4063 45891 4069
rect 45833 4029 45845 4063
rect 45879 4060 45891 4063
rect 46934 4060 46940 4072
rect 45879 4032 46940 4060
rect 45879 4029 45891 4032
rect 45833 4023 45891 4029
rect 46934 4020 46940 4032
rect 46992 4020 46998 4072
rect 47949 4063 48007 4069
rect 47949 4029 47961 4063
rect 47995 4060 48007 4063
rect 49050 4060 49056 4072
rect 47995 4032 49056 4060
rect 47995 4029 48007 4032
rect 47949 4023 48007 4029
rect 49050 4020 49056 4032
rect 49108 4020 49114 4072
rect 50065 4063 50123 4069
rect 50065 4029 50077 4063
rect 50111 4060 50123 4063
rect 51166 4060 51172 4072
rect 50111 4032 51172 4060
rect 50111 4029 50123 4032
rect 50065 4023 50123 4029
rect 51166 4020 51172 4032
rect 51224 4020 51230 4072
rect 52181 4063 52239 4069
rect 52181 4029 52193 4063
rect 52227 4060 52239 4063
rect 52270 4060 52276 4072
rect 52227 4032 52276 4060
rect 52227 4029 52239 4032
rect 52181 4023 52239 4029
rect 52270 4020 52276 4032
rect 52328 4020 52334 4072
rect 54297 4063 54355 4069
rect 54297 4029 54309 4063
rect 54343 4060 54355 4063
rect 54662 4060 54668 4072
rect 54343 4032 54668 4060
rect 54343 4029 54355 4032
rect 54297 4023 54355 4029
rect 54662 4020 54668 4032
rect 54720 4020 54726 4072
rect 56134 4060 56140 4072
rect 56095 4032 56140 4060
rect 56134 4020 56140 4032
rect 56192 4020 56198 4072
rect 56413 4063 56471 4069
rect 56413 4029 56425 4063
rect 56459 4060 56471 4063
rect 57146 4060 57152 4072
rect 56459 4032 57152 4060
rect 56459 4029 56471 4032
rect 56413 4023 56471 4029
rect 57146 4020 57152 4032
rect 57204 4020 57210 4072
rect 58529 4063 58587 4069
rect 58529 4029 58541 4063
rect 58575 4060 58587 4063
rect 58986 4060 58992 4072
rect 58575 4032 58992 4060
rect 58575 4029 58587 4032
rect 58529 4023 58587 4029
rect 58986 4020 58992 4032
rect 59044 4020 59050 4072
rect 60366 4020 60372 4072
rect 60424 4060 60430 4072
rect 60645 4063 60703 4069
rect 60424 4032 60469 4060
rect 60424 4020 60430 4032
rect 60645 4029 60657 4063
rect 60691 4060 60703 4063
rect 61286 4060 61292 4072
rect 60691 4032 61292 4060
rect 60691 4029 60703 4032
rect 60645 4023 60703 4029
rect 61286 4020 61292 4032
rect 61344 4020 61350 4072
rect 62761 4063 62819 4069
rect 62761 4029 62773 4063
rect 62807 4060 62819 4063
rect 63862 4060 63868 4072
rect 62807 4032 63868 4060
rect 62807 4029 62819 4032
rect 62761 4023 62819 4029
rect 63862 4020 63868 4032
rect 63920 4020 63926 4072
rect 64877 4063 64935 4069
rect 64877 4029 64889 4063
rect 64923 4060 64935 4063
rect 65978 4060 65984 4072
rect 64923 4032 65984 4060
rect 64923 4029 64935 4032
rect 64877 4023 64935 4029
rect 65978 4020 65984 4032
rect 66036 4020 66042 4072
rect 66993 4063 67051 4069
rect 66993 4029 67005 4063
rect 67039 4060 67051 4063
rect 68094 4060 68100 4072
rect 67039 4032 68100 4060
rect 67039 4029 67051 4032
rect 66993 4023 67051 4029
rect 68094 4020 68100 4032
rect 68152 4020 68158 4072
rect 69109 4063 69167 4069
rect 69109 4029 69121 4063
rect 69155 4060 69167 4063
rect 69198 4060 69204 4072
rect 69155 4032 69204 4060
rect 69155 4029 69167 4032
rect 69109 4023 69167 4029
rect 69198 4020 69204 4032
rect 69256 4020 69262 4072
rect 71225 4063 71283 4069
rect 71225 4029 71237 4063
rect 71271 4060 71283 4063
rect 71682 4060 71688 4072
rect 71271 4032 71688 4060
rect 71271 4029 71283 4032
rect 71225 4023 71283 4029
rect 71682 4020 71688 4032
rect 71740 4020 71746 4072
rect 73341 4063 73399 4069
rect 73341 4029 73353 4063
rect 73387 4060 73399 4063
rect 73706 4060 73712 4072
rect 73387 4032 73712 4060
rect 73387 4029 73399 4032
rect 73341 4023 73399 4029
rect 73706 4020 73712 4032
rect 73764 4020 73770 4072
rect 75457 4063 75515 4069
rect 75457 4029 75469 4063
rect 75503 4060 75515 4063
rect 75822 4060 75828 4072
rect 75503 4032 75828 4060
rect 75503 4029 75515 4032
rect 75457 4023 75515 4029
rect 75822 4020 75828 4032
rect 75880 4020 75886 4072
rect 77294 4020 77300 4072
rect 77352 4060 77358 4072
rect 77573 4063 77631 4069
rect 77352 4032 77397 4060
rect 77352 4020 77358 4032
rect 77573 4029 77585 4063
rect 77619 4060 77631 4063
rect 78674 4060 78680 4072
rect 77619 4032 78680 4060
rect 77619 4029 77631 4032
rect 77573 4023 77631 4029
rect 78674 4020 78680 4032
rect 78732 4020 78738 4072
rect 79689 4063 79747 4069
rect 79689 4029 79701 4063
rect 79735 4060 79747 4063
rect 80698 4060 80704 4072
rect 79735 4032 80704 4060
rect 79735 4029 79747 4032
rect 79689 4023 79747 4029
rect 80698 4020 80704 4032
rect 80756 4020 80762 4072
rect 81805 4063 81863 4069
rect 81805 4029 81817 4063
rect 81851 4060 81863 4063
rect 82906 4060 82912 4072
rect 81851 4032 82912 4060
rect 81851 4029 81863 4032
rect 81805 4023 81863 4029
rect 82906 4020 82912 4032
rect 82964 4020 82970 4072
rect 83921 4063 83979 4069
rect 83921 4029 83933 4063
rect 83967 4060 83979 4063
rect 85022 4060 85028 4072
rect 83967 4032 85028 4060
rect 83967 4029 83979 4032
rect 83921 4023 83979 4029
rect 85022 4020 85028 4032
rect 85080 4020 85086 4072
rect 86037 4063 86095 4069
rect 86037 4029 86049 4063
rect 86083 4060 86095 4063
rect 86126 4060 86132 4072
rect 86083 4032 86132 4060
rect 86083 4029 86095 4032
rect 86037 4023 86095 4029
rect 86126 4020 86132 4032
rect 86184 4020 86190 4072
rect 88153 4063 88211 4069
rect 88153 4029 88165 4063
rect 88199 4060 88211 4063
rect 88518 4060 88524 4072
rect 88199 4032 88524 4060
rect 88199 4029 88211 4032
rect 88153 4023 88211 4029
rect 88518 4020 88524 4032
rect 88576 4020 88582 4072
rect 89990 4060 89996 4072
rect 89951 4032 89996 4060
rect 89990 4020 89996 4032
rect 90048 4020 90054 4072
rect 90269 4063 90327 4069
rect 90269 4029 90281 4063
rect 90315 4060 90327 4063
rect 90634 4060 90640 4072
rect 90315 4032 90640 4060
rect 90315 4029 90327 4032
rect 90269 4023 90327 4029
rect 90634 4020 90640 4032
rect 90692 4020 90698 4072
rect 92385 4063 92443 4069
rect 92385 4029 92397 4063
rect 92431 4060 92443 4063
rect 93118 4060 93124 4072
rect 92431 4032 93124 4060
rect 92431 4029 92443 4032
rect 92385 4023 92443 4029
rect 93118 4020 93124 4032
rect 93176 4020 93182 4072
rect 94501 4063 94559 4069
rect 94501 4029 94513 4063
rect 94547 4060 94559 4063
rect 95602 4060 95608 4072
rect 94547 4032 95608 4060
rect 94547 4029 94559 4032
rect 94501 4023 94559 4029
rect 95602 4020 95608 4032
rect 95660 4020 95666 4072
rect 96617 4063 96675 4069
rect 96617 4029 96629 4063
rect 96663 4060 96675 4063
rect 97258 4060 97264 4072
rect 96663 4032 97264 4060
rect 96663 4029 96675 4032
rect 96617 4023 96675 4029
rect 97258 4020 97264 4032
rect 97316 4020 97322 4072
rect 98733 4063 98791 4069
rect 98733 4029 98745 4063
rect 98779 4060 98791 4063
rect 99834 4060 99840 4072
rect 98779 4032 99840 4060
rect 98779 4029 98791 4032
rect 98733 4023 98791 4029
rect 99834 4020 99840 4032
rect 99892 4020 99898 4072
rect 100849 4063 100907 4069
rect 100849 4029 100861 4063
rect 100895 4060 100907 4063
rect 101950 4060 101956 4072
rect 100895 4032 101956 4060
rect 100895 4029 100907 4032
rect 100849 4023 100907 4029
rect 101950 4020 101956 4032
rect 102008 4020 102014 4072
rect 102965 4063 103023 4069
rect 102965 4029 102977 4063
rect 103011 4060 103023 4063
rect 103606 4060 103612 4072
rect 103011 4032 103612 4060
rect 103011 4029 103023 4032
rect 102965 4023 103023 4029
rect 103606 4020 103612 4032
rect 103664 4020 103670 4072
rect 105081 4063 105139 4069
rect 105081 4029 105093 4063
rect 105127 4060 105139 4063
rect 105446 4060 105452 4072
rect 105127 4032 105452 4060
rect 105127 4029 105139 4032
rect 105081 4023 105139 4029
rect 105446 4020 105452 4032
rect 105504 4020 105510 4072
rect 81069 3995 81127 4001
rect 81069 3961 81081 3995
rect 81115 3992 81127 3995
rect 81250 3992 81256 4004
rect 81115 3964 81256 3992
rect 81115 3961 81127 3964
rect 81069 3955 81127 3961
rect 81250 3952 81256 3964
rect 81308 3952 81314 4004
rect 1486 3884 1492 3936
rect 1544 3924 1550 3936
rect 2501 3927 2559 3933
rect 2501 3924 2513 3927
rect 1544 3896 2513 3924
rect 1544 3884 1550 3896
rect 2501 3893 2513 3896
rect 2547 3893 2559 3927
rect 4614 3924 4620 3936
rect 4575 3896 4620 3924
rect 2501 3887 2559 3893
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 6730 3924 6736 3936
rect 6691 3896 6736 3924
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 8846 3884 8852 3936
rect 8904 3924 8910 3936
rect 11146 3924 11152 3936
rect 8904 3896 8949 3924
rect 11107 3896 11152 3924
rect 8904 3884 8910 3896
rect 11146 3884 11152 3896
rect 11204 3884 11210 3936
rect 13262 3924 13268 3936
rect 13223 3896 13268 3924
rect 13262 3884 13268 3896
rect 13320 3884 13326 3936
rect 14182 3884 14188 3936
rect 14240 3924 14246 3936
rect 15197 3927 15255 3933
rect 15197 3924 15209 3927
rect 14240 3896 15209 3924
rect 14240 3884 14246 3896
rect 15197 3893 15209 3896
rect 15243 3893 15255 3927
rect 15197 3887 15255 3893
rect 16298 3884 16304 3936
rect 16356 3924 16362 3936
rect 17313 3927 17371 3933
rect 17313 3924 17325 3927
rect 16356 3896 17325 3924
rect 16356 3884 16362 3896
rect 17313 3893 17325 3896
rect 17359 3893 17371 3927
rect 17313 3887 17371 3893
rect 18690 3884 18696 3936
rect 18748 3924 18754 3936
rect 19429 3927 19487 3933
rect 19429 3924 19441 3927
rect 18748 3896 19441 3924
rect 18748 3884 18754 3896
rect 19429 3893 19441 3896
rect 19475 3893 19487 3927
rect 21542 3924 21548 3936
rect 21503 3896 21548 3924
rect 19429 3887 19487 3893
rect 21542 3884 21548 3896
rect 21600 3884 21606 3936
rect 23658 3924 23664 3936
rect 23619 3896 23664 3924
rect 23658 3884 23664 3896
rect 23716 3884 23722 3936
rect 25774 3924 25780 3936
rect 25735 3896 25780 3924
rect 25774 3884 25780 3896
rect 25832 3884 25838 3936
rect 28074 3924 28080 3936
rect 28035 3896 28080 3924
rect 28074 3884 28080 3896
rect 28132 3884 28138 3936
rect 30190 3924 30196 3936
rect 30151 3896 30196 3924
rect 30190 3884 30196 3896
rect 30248 3884 30254 3936
rect 31110 3884 31116 3936
rect 31168 3924 31174 3936
rect 32125 3927 32183 3933
rect 32125 3924 32137 3927
rect 31168 3896 32137 3924
rect 31168 3884 31174 3896
rect 32125 3893 32137 3896
rect 32171 3893 32183 3927
rect 32125 3887 32183 3893
rect 33226 3884 33232 3936
rect 33284 3924 33290 3936
rect 34241 3927 34299 3933
rect 34241 3924 34253 3927
rect 33284 3896 34253 3924
rect 33284 3884 33290 3896
rect 34241 3893 34253 3896
rect 34287 3893 34299 3927
rect 34241 3887 34299 3893
rect 35342 3884 35348 3936
rect 35400 3924 35406 3936
rect 36357 3927 36415 3933
rect 36357 3924 36369 3927
rect 35400 3896 36369 3924
rect 35400 3884 35406 3896
rect 36357 3893 36369 3896
rect 36403 3893 36415 3927
rect 38470 3924 38476 3936
rect 38431 3896 38476 3924
rect 36357 3887 36415 3893
rect 38470 3884 38476 3896
rect 38528 3884 38534 3936
rect 40586 3924 40592 3936
rect 40547 3896 40592 3924
rect 40586 3884 40592 3896
rect 40644 3884 40650 3936
rect 42702 3924 42708 3936
rect 42663 3896 42708 3924
rect 42702 3884 42708 3896
rect 42760 3884 42766 3936
rect 45002 3924 45008 3936
rect 44963 3896 45008 3924
rect 45002 3884 45008 3896
rect 45060 3884 45066 3936
rect 47118 3924 47124 3936
rect 47079 3896 47124 3924
rect 47118 3884 47124 3896
rect 47176 3884 47182 3936
rect 48038 3884 48044 3936
rect 48096 3924 48102 3936
rect 49053 3927 49111 3933
rect 49053 3924 49065 3927
rect 48096 3896 49065 3924
rect 48096 3884 48102 3896
rect 49053 3893 49065 3896
rect 49099 3893 49111 3927
rect 49053 3887 49111 3893
rect 50522 3884 50528 3936
rect 50580 3924 50586 3936
rect 51169 3927 51227 3933
rect 51169 3924 51181 3927
rect 50580 3896 51181 3924
rect 50580 3884 50586 3896
rect 51169 3893 51181 3896
rect 51215 3893 51227 3927
rect 51169 3887 51227 3893
rect 52546 3884 52552 3936
rect 52604 3924 52610 3936
rect 53285 3927 53343 3933
rect 53285 3924 53297 3927
rect 52604 3896 53297 3924
rect 52604 3884 52610 3896
rect 53285 3893 53297 3896
rect 53331 3893 53343 3927
rect 55398 3924 55404 3936
rect 55359 3896 55404 3924
rect 53285 3887 53343 3893
rect 55398 3884 55404 3896
rect 55456 3884 55462 3936
rect 57514 3924 57520 3936
rect 57475 3896 57520 3924
rect 57514 3884 57520 3896
rect 57572 3884 57578 3936
rect 59630 3924 59636 3936
rect 59591 3896 59636 3924
rect 59630 3884 59636 3896
rect 59688 3884 59694 3936
rect 61930 3924 61936 3936
rect 61891 3896 61936 3924
rect 61930 3884 61936 3896
rect 61988 3884 61994 3936
rect 64046 3924 64052 3936
rect 64007 3896 64052 3924
rect 64046 3884 64052 3896
rect 64104 3884 64110 3936
rect 64966 3884 64972 3936
rect 65024 3924 65030 3936
rect 65981 3927 66039 3933
rect 65981 3924 65993 3927
rect 65024 3896 65993 3924
rect 65024 3884 65030 3896
rect 65981 3893 65993 3896
rect 66027 3893 66039 3927
rect 65981 3887 66039 3893
rect 67082 3884 67088 3936
rect 67140 3924 67146 3936
rect 68097 3927 68155 3933
rect 68097 3924 68109 3927
rect 67140 3896 68109 3924
rect 67140 3884 67146 3896
rect 68097 3893 68109 3896
rect 68143 3893 68155 3927
rect 68097 3887 68155 3893
rect 69474 3884 69480 3936
rect 69532 3924 69538 3936
rect 70213 3927 70271 3933
rect 70213 3924 70225 3927
rect 69532 3896 70225 3924
rect 69532 3884 69538 3896
rect 70213 3893 70225 3896
rect 70259 3893 70271 3927
rect 72326 3924 72332 3936
rect 72287 3896 72332 3924
rect 70213 3887 70271 3893
rect 72326 3884 72332 3896
rect 72384 3884 72390 3936
rect 74442 3924 74448 3936
rect 74403 3896 74448 3924
rect 74442 3884 74448 3896
rect 74500 3884 74506 3936
rect 76742 3924 76748 3936
rect 76703 3896 76748 3924
rect 76742 3884 76748 3896
rect 76800 3884 76806 3936
rect 78766 3884 78772 3936
rect 78824 3924 78830 3936
rect 78861 3927 78919 3933
rect 78861 3924 78873 3927
rect 78824 3896 78873 3924
rect 78824 3884 78830 3896
rect 78861 3893 78873 3896
rect 78907 3893 78919 3927
rect 78861 3887 78919 3893
rect 81894 3884 81900 3936
rect 81952 3924 81958 3936
rect 82909 3927 82967 3933
rect 82909 3924 82921 3927
rect 81952 3896 82921 3924
rect 81952 3884 81958 3896
rect 82909 3893 82921 3896
rect 82955 3893 82967 3927
rect 82909 3887 82967 3893
rect 84010 3884 84016 3936
rect 84068 3924 84074 3936
rect 85025 3927 85083 3933
rect 85025 3924 85037 3927
rect 84068 3896 85037 3924
rect 84068 3884 84074 3896
rect 85025 3893 85037 3896
rect 85071 3893 85083 3927
rect 85025 3887 85083 3893
rect 86402 3884 86408 3936
rect 86460 3924 86466 3936
rect 87141 3927 87199 3933
rect 87141 3924 87153 3927
rect 86460 3896 87153 3924
rect 86460 3884 86466 3896
rect 87141 3893 87153 3896
rect 87187 3893 87199 3927
rect 89438 3924 89444 3936
rect 89399 3896 89444 3924
rect 87141 3887 87199 3893
rect 89438 3884 89444 3896
rect 89496 3884 89502 3936
rect 91370 3924 91376 3936
rect 91331 3896 91376 3924
rect 91370 3884 91376 3896
rect 91428 3884 91434 3936
rect 93486 3924 93492 3936
rect 93447 3896 93492 3924
rect 93486 3884 93492 3896
rect 93544 3884 93550 3936
rect 95694 3884 95700 3936
rect 95752 3924 95758 3936
rect 95789 3927 95847 3933
rect 95789 3924 95801 3927
rect 95752 3896 95801 3924
rect 95752 3884 95758 3896
rect 95789 3893 95801 3896
rect 95835 3893 95847 3927
rect 97902 3924 97908 3936
rect 97863 3896 97908 3924
rect 95789 3887 95847 3893
rect 97902 3884 97908 3896
rect 97960 3884 97966 3936
rect 98822 3884 98828 3936
rect 98880 3924 98886 3936
rect 99837 3927 99895 3933
rect 99837 3924 99849 3927
rect 98880 3896 99849 3924
rect 98880 3884 98886 3896
rect 99837 3893 99849 3896
rect 99883 3893 99895 3927
rect 99837 3887 99895 3893
rect 100938 3884 100944 3936
rect 100996 3924 101002 3936
rect 101953 3927 102011 3933
rect 101953 3924 101965 3927
rect 100996 3896 101965 3924
rect 100996 3884 101002 3896
rect 101953 3893 101965 3896
rect 101999 3893 102011 3927
rect 101953 3887 102011 3893
rect 103054 3884 103060 3936
rect 103112 3924 103118 3936
rect 104069 3927 104127 3933
rect 104069 3924 104081 3927
rect 103112 3896 104081 3924
rect 103112 3884 103118 3896
rect 104069 3893 104081 3896
rect 104115 3893 104127 3927
rect 104069 3887 104127 3893
rect 105170 3884 105176 3936
rect 105228 3924 105234 3936
rect 106185 3927 106243 3933
rect 106185 3924 106197 3927
rect 105228 3896 106197 3924
rect 105228 3884 105234 3896
rect 106185 3893 106197 3896
rect 106231 3893 106243 3927
rect 106185 3887 106243 3893
rect 1104 3834 106904 3856
rect 1104 3782 19402 3834
rect 19454 3782 19466 3834
rect 19518 3782 19530 3834
rect 19582 3782 19594 3834
rect 19646 3782 50122 3834
rect 50174 3782 50186 3834
rect 50238 3782 50250 3834
rect 50302 3782 50314 3834
rect 50366 3782 80842 3834
rect 80894 3782 80906 3834
rect 80958 3782 80970 3834
rect 81022 3782 81034 3834
rect 81086 3782 106904 3834
rect 1104 3760 106904 3782
rect 2498 3720 2504 3732
rect 2459 3692 2504 3720
rect 2498 3680 2504 3692
rect 2556 3680 2562 3732
rect 10962 3720 10968 3732
rect 10923 3692 10968 3720
rect 10962 3680 10968 3692
rect 11020 3680 11026 3732
rect 13078 3720 13084 3732
rect 13039 3692 13084 3720
rect 13078 3680 13084 3692
rect 13136 3680 13142 3732
rect 15194 3720 15200 3732
rect 15155 3692 15200 3720
rect 15194 3680 15200 3692
rect 15252 3680 15258 3732
rect 17310 3720 17316 3732
rect 17271 3692 17316 3720
rect 17310 3680 17316 3692
rect 17368 3680 17374 3732
rect 27890 3720 27896 3732
rect 27851 3692 27896 3720
rect 27890 3680 27896 3692
rect 27948 3680 27954 3732
rect 30006 3720 30012 3732
rect 29967 3692 30012 3720
rect 30006 3680 30012 3692
rect 30064 3680 30070 3732
rect 32122 3720 32128 3732
rect 32083 3692 32128 3720
rect 32122 3680 32128 3692
rect 32180 3680 32186 3732
rect 34238 3720 34244 3732
rect 34199 3692 34244 3720
rect 34238 3680 34244 3692
rect 34296 3680 34302 3732
rect 44818 3720 44824 3732
rect 44779 3692 44824 3720
rect 44818 3680 44824 3692
rect 44876 3680 44882 3732
rect 46934 3720 46940 3732
rect 46895 3692 46940 3720
rect 46934 3680 46940 3692
rect 46992 3680 46998 3732
rect 49050 3720 49056 3732
rect 49011 3692 49056 3720
rect 49050 3680 49056 3692
rect 49108 3680 49114 3732
rect 51166 3720 51172 3732
rect 51127 3692 51172 3720
rect 51166 3680 51172 3692
rect 51224 3680 51230 3732
rect 63862 3720 63868 3732
rect 63823 3692 63868 3720
rect 63862 3680 63868 3692
rect 63920 3680 63926 3732
rect 65978 3720 65984 3732
rect 65939 3692 65984 3720
rect 65978 3680 65984 3692
rect 66036 3680 66042 3732
rect 68094 3720 68100 3732
rect 68055 3692 68100 3720
rect 68094 3680 68100 3692
rect 68152 3680 68158 3732
rect 78674 3720 78680 3732
rect 78635 3692 78680 3720
rect 78674 3680 78680 3692
rect 78732 3680 78738 3732
rect 80698 3680 80704 3732
rect 80756 3720 80762 3732
rect 80793 3723 80851 3729
rect 80793 3720 80805 3723
rect 80756 3692 80805 3720
rect 80756 3680 80762 3692
rect 80793 3689 80805 3692
rect 80839 3689 80851 3723
rect 82906 3720 82912 3732
rect 82867 3692 82912 3720
rect 80793 3683 80851 3689
rect 82906 3680 82912 3692
rect 82964 3680 82970 3732
rect 85022 3720 85028 3732
rect 84983 3692 85028 3720
rect 85022 3680 85028 3692
rect 85080 3680 85086 3732
rect 95602 3720 95608 3732
rect 95563 3692 95608 3720
rect 95602 3680 95608 3692
rect 95660 3680 95666 3732
rect 99834 3720 99840 3732
rect 99795 3692 99840 3720
rect 99834 3680 99840 3692
rect 99892 3680 99898 3732
rect 101950 3720 101956 3732
rect 101911 3692 101956 3720
rect 101950 3680 101956 3692
rect 102008 3680 102014 3732
rect 1118 3584 1124 3596
rect 1079 3556 1124 3584
rect 1118 3544 1124 3556
rect 1176 3544 1182 3596
rect 3234 3584 3240 3596
rect 3195 3556 3240 3584
rect 3234 3544 3240 3556
rect 3292 3544 3298 3596
rect 5350 3584 5356 3596
rect 5311 3556 5356 3584
rect 5350 3544 5356 3556
rect 5408 3544 5414 3596
rect 7466 3584 7472 3596
rect 7427 3556 7472 3584
rect 7466 3544 7472 3556
rect 7524 3544 7530 3596
rect 9582 3584 9588 3596
rect 9543 3556 9588 3584
rect 9582 3544 9588 3556
rect 9640 3544 9646 3596
rect 11698 3584 11704 3596
rect 11659 3556 11704 3584
rect 11698 3544 11704 3556
rect 11756 3544 11762 3596
rect 13814 3584 13820 3596
rect 13775 3556 13820 3584
rect 13814 3544 13820 3556
rect 13872 3544 13878 3596
rect 15930 3584 15936 3596
rect 15891 3556 15936 3584
rect 15930 3544 15936 3556
rect 15988 3544 15994 3596
rect 18046 3584 18052 3596
rect 18007 3556 18052 3584
rect 18046 3544 18052 3556
rect 18104 3544 18110 3596
rect 20162 3584 20168 3596
rect 20123 3556 20168 3584
rect 20162 3544 20168 3556
rect 20220 3544 20226 3596
rect 22186 3544 22192 3596
rect 22244 3584 22250 3596
rect 22281 3587 22339 3593
rect 22281 3584 22293 3587
rect 22244 3556 22293 3584
rect 22244 3544 22250 3556
rect 22281 3553 22293 3556
rect 22327 3553 22339 3587
rect 24394 3584 24400 3596
rect 24355 3556 24400 3584
rect 22281 3547 22339 3553
rect 24394 3544 24400 3556
rect 24452 3544 24458 3596
rect 26510 3584 26516 3596
rect 26471 3556 26516 3584
rect 26510 3544 26516 3556
rect 26568 3544 26574 3596
rect 28626 3584 28632 3596
rect 28587 3556 28632 3584
rect 28626 3544 28632 3556
rect 28684 3544 28690 3596
rect 30742 3584 30748 3596
rect 30703 3556 30748 3584
rect 30742 3544 30748 3556
rect 30800 3544 30806 3596
rect 32858 3584 32864 3596
rect 32819 3556 32864 3584
rect 32858 3544 32864 3556
rect 32916 3544 32922 3596
rect 34977 3587 35035 3593
rect 34977 3553 34989 3587
rect 35023 3584 35035 3587
rect 35066 3584 35072 3596
rect 35023 3556 35072 3584
rect 35023 3553 35035 3556
rect 34977 3547 35035 3553
rect 35066 3544 35072 3556
rect 35124 3544 35130 3596
rect 37090 3584 37096 3596
rect 37051 3556 37096 3584
rect 37090 3544 37096 3556
rect 37148 3544 37154 3596
rect 39206 3584 39212 3596
rect 39167 3556 39212 3584
rect 39206 3544 39212 3556
rect 39264 3544 39270 3596
rect 39482 3584 39488 3596
rect 39443 3556 39488 3584
rect 39482 3544 39488 3556
rect 39540 3584 39546 3596
rect 40402 3584 40408 3596
rect 39540 3556 40408 3584
rect 39540 3544 39546 3556
rect 40402 3544 40408 3556
rect 40460 3544 40466 3596
rect 41322 3584 41328 3596
rect 41283 3556 41328 3584
rect 41322 3544 41328 3556
rect 41380 3544 41386 3596
rect 43438 3584 43444 3596
rect 43399 3556 43444 3584
rect 43438 3544 43444 3556
rect 43496 3544 43502 3596
rect 45554 3584 45560 3596
rect 45515 3556 45560 3584
rect 45554 3544 45560 3556
rect 45612 3544 45618 3596
rect 47670 3584 47676 3596
rect 47631 3556 47676 3584
rect 47670 3544 47676 3556
rect 47728 3544 47734 3596
rect 49786 3584 49792 3596
rect 49747 3556 49792 3584
rect 49786 3544 49792 3556
rect 49844 3544 49850 3596
rect 51902 3584 51908 3596
rect 51863 3556 51908 3584
rect 51902 3544 51908 3556
rect 51960 3544 51966 3596
rect 54018 3584 54024 3596
rect 53979 3556 54024 3584
rect 54018 3544 54024 3556
rect 54076 3544 54082 3596
rect 56134 3584 56140 3596
rect 56095 3556 56140 3584
rect 56134 3544 56140 3556
rect 56192 3544 56198 3596
rect 58250 3584 58256 3596
rect 58211 3556 58256 3584
rect 58250 3544 58256 3556
rect 58308 3544 58314 3596
rect 60366 3544 60372 3596
rect 60424 3584 60430 3596
rect 62482 3584 62488 3596
rect 60424 3556 60469 3584
rect 62443 3556 62488 3584
rect 60424 3544 60430 3556
rect 62482 3544 62488 3556
rect 62540 3544 62546 3596
rect 64598 3584 64604 3596
rect 64559 3556 64604 3584
rect 64598 3544 64604 3556
rect 64656 3544 64662 3596
rect 66714 3584 66720 3596
rect 66675 3556 66720 3584
rect 66714 3544 66720 3556
rect 66772 3544 66778 3596
rect 68830 3584 68836 3596
rect 68791 3556 68836 3584
rect 68830 3544 68836 3556
rect 68888 3544 68894 3596
rect 70946 3584 70952 3596
rect 70907 3556 70952 3584
rect 70946 3544 70952 3556
rect 71004 3544 71010 3596
rect 73062 3584 73068 3596
rect 73023 3556 73068 3584
rect 73062 3544 73068 3556
rect 73120 3544 73126 3596
rect 75178 3584 75184 3596
rect 75139 3556 75184 3584
rect 75178 3544 75184 3556
rect 75236 3544 75242 3596
rect 77386 3584 77392 3596
rect 75472 3556 77392 3584
rect 1394 3516 1400 3528
rect 1355 3488 1400 3516
rect 1394 3476 1400 3488
rect 1452 3476 1458 3528
rect 3510 3516 3516 3528
rect 3471 3488 3516 3516
rect 3510 3476 3516 3488
rect 3568 3476 3574 3528
rect 3878 3476 3884 3528
rect 3936 3516 3942 3528
rect 4617 3519 4675 3525
rect 4617 3516 4629 3519
rect 3936 3488 4629 3516
rect 3936 3476 3942 3488
rect 4617 3485 4629 3488
rect 4663 3485 4675 3519
rect 5626 3516 5632 3528
rect 5587 3488 5632 3516
rect 4617 3479 4675 3485
rect 5626 3476 5632 3488
rect 5684 3476 5690 3528
rect 5994 3476 6000 3528
rect 6052 3516 6058 3528
rect 6733 3519 6791 3525
rect 6733 3516 6745 3519
rect 6052 3488 6745 3516
rect 6052 3476 6058 3488
rect 6733 3485 6745 3488
rect 6779 3485 6791 3519
rect 7742 3516 7748 3528
rect 7703 3488 7748 3516
rect 6733 3479 6791 3485
rect 7742 3476 7748 3488
rect 7800 3476 7806 3528
rect 8110 3476 8116 3528
rect 8168 3516 8174 3528
rect 8849 3519 8907 3525
rect 8849 3516 8861 3519
rect 8168 3488 8861 3516
rect 8168 3476 8174 3488
rect 8849 3485 8861 3488
rect 8895 3485 8907 3519
rect 9858 3516 9864 3528
rect 9819 3488 9864 3516
rect 8849 3479 8907 3485
rect 9858 3476 9864 3488
rect 9916 3476 9922 3528
rect 11974 3516 11980 3528
rect 11935 3488 11980 3516
rect 11974 3476 11980 3488
rect 12032 3476 12038 3528
rect 14090 3516 14096 3528
rect 14051 3488 14096 3516
rect 14090 3476 14096 3488
rect 14148 3476 14154 3528
rect 16206 3516 16212 3528
rect 16167 3488 16212 3516
rect 16206 3476 16212 3488
rect 16264 3476 16270 3528
rect 18322 3516 18328 3528
rect 18283 3488 18328 3516
rect 18322 3476 18328 3488
rect 18380 3476 18386 3528
rect 18414 3476 18420 3528
rect 18472 3516 18478 3528
rect 19429 3519 19487 3525
rect 19429 3516 19441 3519
rect 18472 3488 19441 3516
rect 18472 3476 18478 3488
rect 19429 3485 19441 3488
rect 19475 3485 19487 3519
rect 20438 3516 20444 3528
rect 20399 3488 20444 3516
rect 19429 3479 19487 3485
rect 20438 3476 20444 3488
rect 20496 3476 20502 3528
rect 21082 3476 21088 3528
rect 21140 3516 21146 3528
rect 21545 3519 21603 3525
rect 21545 3516 21557 3519
rect 21140 3488 21557 3516
rect 21140 3476 21146 3488
rect 21545 3485 21557 3488
rect 21591 3485 21603 3519
rect 22554 3516 22560 3528
rect 22515 3488 22560 3516
rect 21545 3479 21603 3485
rect 22554 3476 22560 3488
rect 22612 3476 22618 3528
rect 22922 3476 22928 3528
rect 22980 3516 22986 3528
rect 23661 3519 23719 3525
rect 23661 3516 23673 3519
rect 22980 3488 23673 3516
rect 22980 3476 22986 3488
rect 23661 3485 23673 3488
rect 23707 3485 23719 3519
rect 24670 3516 24676 3528
rect 24631 3488 24676 3516
rect 23661 3479 23719 3485
rect 24670 3476 24676 3488
rect 24728 3476 24734 3528
rect 25038 3476 25044 3528
rect 25096 3516 25102 3528
rect 25777 3519 25835 3525
rect 25777 3516 25789 3519
rect 25096 3488 25789 3516
rect 25096 3476 25102 3488
rect 25777 3485 25789 3488
rect 25823 3485 25835 3519
rect 26786 3516 26792 3528
rect 26747 3488 26792 3516
rect 25777 3479 25835 3485
rect 26786 3476 26792 3488
rect 26844 3476 26850 3528
rect 28902 3516 28908 3528
rect 28863 3488 28908 3516
rect 28902 3476 28908 3488
rect 28960 3476 28966 3528
rect 31018 3516 31024 3528
rect 30979 3488 31024 3516
rect 31018 3476 31024 3488
rect 31076 3476 31082 3528
rect 33134 3516 33140 3528
rect 33095 3488 33140 3516
rect 33134 3476 33140 3488
rect 33192 3476 33198 3528
rect 35250 3516 35256 3528
rect 35211 3488 35256 3516
rect 35250 3476 35256 3488
rect 35308 3476 35314 3528
rect 35618 3476 35624 3528
rect 35676 3516 35682 3528
rect 36357 3519 36415 3525
rect 36357 3516 36369 3519
rect 35676 3488 36369 3516
rect 35676 3476 35682 3488
rect 36357 3485 36369 3488
rect 36403 3485 36415 3519
rect 37366 3516 37372 3528
rect 37327 3488 37372 3516
rect 36357 3479 36415 3485
rect 37366 3476 37372 3488
rect 37424 3476 37430 3528
rect 37734 3476 37740 3528
rect 37792 3516 37798 3528
rect 38473 3519 38531 3525
rect 38473 3516 38485 3519
rect 37792 3488 38485 3516
rect 37792 3476 37798 3488
rect 38473 3485 38485 3488
rect 38519 3485 38531 3519
rect 38473 3479 38531 3485
rect 39942 3476 39948 3528
rect 40000 3516 40006 3528
rect 40681 3519 40739 3525
rect 40681 3516 40693 3519
rect 40000 3488 40693 3516
rect 40000 3476 40006 3488
rect 40681 3485 40693 3488
rect 40727 3485 40739 3519
rect 41598 3516 41604 3528
rect 41559 3488 41604 3516
rect 40681 3479 40739 3485
rect 41598 3476 41604 3488
rect 41656 3476 41662 3528
rect 41966 3476 41972 3528
rect 42024 3516 42030 3528
rect 42705 3519 42763 3525
rect 42705 3516 42717 3519
rect 42024 3488 42717 3516
rect 42024 3476 42030 3488
rect 42705 3485 42717 3488
rect 42751 3485 42763 3519
rect 43714 3516 43720 3528
rect 43675 3488 43720 3516
rect 42705 3479 42763 3485
rect 43714 3476 43720 3488
rect 43772 3476 43778 3528
rect 45830 3516 45836 3528
rect 45791 3488 45836 3516
rect 45830 3476 45836 3488
rect 45888 3476 45894 3528
rect 47946 3516 47952 3528
rect 47907 3488 47952 3516
rect 47946 3476 47952 3488
rect 48004 3476 48010 3528
rect 50062 3476 50068 3528
rect 50120 3516 50126 3528
rect 52178 3516 52184 3528
rect 50120 3488 50165 3516
rect 52139 3488 52184 3516
rect 50120 3476 50126 3488
rect 52178 3476 52184 3488
rect 52236 3476 52242 3528
rect 52270 3476 52276 3528
rect 52328 3516 52334 3528
rect 53285 3519 53343 3525
rect 53285 3516 53297 3519
rect 52328 3488 53297 3516
rect 52328 3476 52334 3488
rect 53285 3485 53297 3488
rect 53331 3485 53343 3519
rect 54294 3516 54300 3528
rect 54255 3488 54300 3516
rect 53285 3479 53343 3485
rect 54294 3476 54300 3488
rect 54352 3476 54358 3528
rect 54662 3476 54668 3528
rect 54720 3516 54726 3528
rect 55401 3519 55459 3525
rect 55401 3516 55413 3519
rect 54720 3488 55413 3516
rect 54720 3476 54726 3488
rect 55401 3485 55413 3488
rect 55447 3485 55459 3519
rect 56410 3516 56416 3528
rect 56371 3488 56416 3516
rect 55401 3479 55459 3485
rect 56410 3476 56416 3488
rect 56468 3476 56474 3528
rect 57146 3476 57152 3528
rect 57204 3516 57210 3528
rect 57517 3519 57575 3525
rect 57517 3516 57529 3519
rect 57204 3488 57529 3516
rect 57204 3476 57210 3488
rect 57517 3485 57529 3488
rect 57563 3485 57575 3519
rect 58526 3516 58532 3528
rect 58487 3488 58532 3516
rect 57517 3479 57575 3485
rect 58526 3476 58532 3488
rect 58584 3476 58590 3528
rect 58986 3476 58992 3528
rect 59044 3516 59050 3528
rect 59633 3519 59691 3525
rect 59633 3516 59645 3519
rect 59044 3488 59645 3516
rect 59044 3476 59050 3488
rect 59633 3485 59645 3488
rect 59679 3485 59691 3519
rect 60642 3516 60648 3528
rect 60603 3488 60648 3516
rect 59633 3479 59691 3485
rect 60642 3476 60648 3488
rect 60700 3476 60706 3528
rect 61286 3476 61292 3528
rect 61344 3516 61350 3528
rect 61749 3519 61807 3525
rect 61749 3516 61761 3519
rect 61344 3488 61761 3516
rect 61344 3476 61350 3488
rect 61749 3485 61761 3488
rect 61795 3485 61807 3519
rect 62758 3516 62764 3528
rect 62719 3488 62764 3516
rect 61749 3479 61807 3485
rect 62758 3476 62764 3488
rect 62816 3476 62822 3528
rect 64874 3516 64880 3528
rect 64835 3488 64880 3516
rect 64874 3476 64880 3488
rect 64932 3476 64938 3528
rect 66990 3516 66996 3528
rect 66951 3488 66996 3516
rect 66990 3476 66996 3488
rect 67048 3476 67054 3528
rect 69106 3516 69112 3528
rect 69067 3488 69112 3516
rect 69106 3476 69112 3488
rect 69164 3476 69170 3528
rect 69198 3476 69204 3528
rect 69256 3516 69262 3528
rect 70213 3519 70271 3525
rect 70213 3516 70225 3519
rect 69256 3488 70225 3516
rect 69256 3476 69262 3488
rect 70213 3485 70225 3488
rect 70259 3485 70271 3519
rect 71222 3516 71228 3528
rect 71183 3488 71228 3516
rect 70213 3479 70271 3485
rect 71222 3476 71228 3488
rect 71280 3476 71286 3528
rect 71682 3476 71688 3528
rect 71740 3516 71746 3528
rect 72329 3519 72387 3525
rect 72329 3516 72341 3519
rect 71740 3488 72341 3516
rect 71740 3476 71746 3488
rect 72329 3485 72341 3488
rect 72375 3485 72387 3519
rect 73338 3516 73344 3528
rect 73299 3488 73344 3516
rect 72329 3479 72387 3485
rect 73338 3476 73344 3488
rect 73396 3476 73402 3528
rect 73706 3476 73712 3528
rect 73764 3516 73770 3528
rect 74445 3519 74503 3525
rect 74445 3516 74457 3519
rect 73764 3488 74457 3516
rect 73764 3476 73770 3488
rect 74445 3485 74457 3488
rect 74491 3485 74503 3519
rect 74445 3479 74503 3485
rect 75362 3476 75368 3528
rect 75420 3516 75426 3528
rect 75472 3525 75500 3556
rect 77386 3544 77392 3556
rect 77444 3544 77450 3596
rect 79410 3584 79416 3596
rect 79371 3556 79416 3584
rect 79410 3544 79416 3556
rect 79468 3544 79474 3596
rect 81526 3584 81532 3596
rect 81487 3556 81532 3584
rect 81526 3544 81532 3556
rect 81584 3544 81590 3596
rect 83642 3584 83648 3596
rect 83603 3556 83648 3584
rect 83642 3544 83648 3556
rect 83700 3544 83706 3596
rect 85758 3584 85764 3596
rect 85719 3556 85764 3584
rect 85758 3544 85764 3556
rect 85816 3544 85822 3596
rect 87046 3584 87052 3596
rect 86052 3556 87052 3584
rect 75457 3519 75515 3525
rect 75457 3516 75469 3519
rect 75420 3488 75469 3516
rect 75420 3476 75426 3488
rect 75457 3485 75469 3488
rect 75503 3485 75515 3519
rect 75457 3479 75515 3485
rect 75822 3476 75828 3528
rect 75880 3516 75886 3528
rect 76561 3519 76619 3525
rect 76561 3516 76573 3519
rect 75880 3488 76573 3516
rect 75880 3476 75886 3488
rect 76561 3485 76573 3488
rect 76607 3485 76619 3519
rect 76561 3479 76619 3485
rect 77294 3476 77300 3528
rect 77352 3516 77358 3528
rect 77570 3516 77576 3528
rect 77352 3488 77397 3516
rect 77531 3488 77576 3516
rect 77352 3476 77358 3488
rect 77570 3476 77576 3488
rect 77628 3476 77634 3528
rect 79686 3516 79692 3528
rect 79647 3488 79692 3516
rect 79686 3476 79692 3488
rect 79744 3476 79750 3528
rect 81802 3516 81808 3528
rect 81763 3488 81808 3516
rect 81802 3476 81808 3488
rect 81860 3476 81866 3528
rect 83918 3516 83924 3528
rect 83879 3488 83924 3516
rect 83918 3476 83924 3488
rect 83976 3476 83982 3528
rect 85942 3476 85948 3528
rect 86000 3516 86006 3528
rect 86052 3525 86080 3556
rect 87046 3544 87052 3556
rect 87104 3544 87110 3596
rect 87874 3584 87880 3596
rect 87835 3556 87880 3584
rect 87874 3544 87880 3556
rect 87932 3544 87938 3596
rect 89990 3584 89996 3596
rect 89951 3556 89996 3584
rect 89990 3544 89996 3556
rect 90048 3544 90054 3596
rect 92106 3584 92112 3596
rect 92067 3556 92112 3584
rect 92106 3544 92112 3556
rect 92164 3544 92170 3596
rect 94222 3584 94228 3596
rect 94183 3556 94228 3584
rect 94222 3544 94228 3556
rect 94280 3544 94286 3596
rect 96062 3544 96068 3596
rect 96120 3584 96126 3596
rect 96341 3587 96399 3593
rect 96341 3584 96353 3587
rect 96120 3556 96353 3584
rect 96120 3544 96126 3556
rect 96341 3553 96353 3556
rect 96387 3553 96399 3587
rect 98454 3584 98460 3596
rect 98415 3556 98460 3584
rect 96341 3547 96399 3553
rect 98454 3544 98460 3556
rect 98512 3544 98518 3596
rect 100570 3584 100576 3596
rect 100531 3556 100576 3584
rect 100570 3544 100576 3556
rect 100628 3544 100634 3596
rect 102686 3584 102692 3596
rect 102647 3556 102692 3584
rect 102686 3544 102692 3556
rect 102744 3544 102750 3596
rect 104802 3584 104808 3596
rect 104763 3556 104808 3584
rect 104802 3544 104808 3556
rect 104860 3544 104866 3596
rect 86037 3519 86095 3525
rect 86037 3516 86049 3519
rect 86000 3488 86049 3516
rect 86000 3476 86006 3488
rect 86037 3485 86049 3488
rect 86083 3485 86095 3519
rect 86037 3479 86095 3485
rect 86126 3476 86132 3528
rect 86184 3516 86190 3528
rect 87141 3519 87199 3525
rect 87141 3516 87153 3519
rect 86184 3488 87153 3516
rect 86184 3476 86190 3488
rect 87141 3485 87153 3488
rect 87187 3485 87199 3519
rect 88150 3516 88156 3528
rect 88111 3488 88156 3516
rect 87141 3479 87199 3485
rect 88150 3476 88156 3488
rect 88208 3476 88214 3528
rect 88518 3476 88524 3528
rect 88576 3516 88582 3528
rect 89257 3519 89315 3525
rect 89257 3516 89269 3519
rect 88576 3488 89269 3516
rect 88576 3476 88582 3488
rect 89257 3485 89269 3488
rect 89303 3485 89315 3519
rect 90266 3516 90272 3528
rect 90227 3488 90272 3516
rect 89257 3479 89315 3485
rect 90266 3476 90272 3488
rect 90324 3476 90330 3528
rect 90634 3476 90640 3528
rect 90692 3516 90698 3528
rect 91373 3519 91431 3525
rect 91373 3516 91385 3519
rect 90692 3488 91385 3516
rect 90692 3476 90698 3488
rect 91373 3485 91385 3488
rect 91419 3485 91431 3519
rect 92382 3516 92388 3528
rect 92343 3488 92388 3516
rect 91373 3479 91431 3485
rect 92382 3476 92388 3488
rect 92440 3476 92446 3528
rect 93118 3476 93124 3528
rect 93176 3516 93182 3528
rect 93489 3519 93547 3525
rect 93489 3516 93501 3519
rect 93176 3488 93501 3516
rect 93176 3476 93182 3488
rect 93489 3485 93501 3488
rect 93535 3485 93547 3519
rect 94498 3516 94504 3528
rect 94459 3488 94504 3516
rect 93489 3479 93547 3485
rect 94498 3476 94504 3488
rect 94556 3476 94562 3528
rect 96614 3516 96620 3528
rect 96575 3488 96620 3516
rect 96614 3476 96620 3488
rect 96672 3476 96678 3528
rect 97258 3476 97264 3528
rect 97316 3516 97322 3528
rect 97721 3519 97779 3525
rect 97721 3516 97733 3519
rect 97316 3488 97733 3516
rect 97316 3476 97322 3488
rect 97721 3485 97733 3488
rect 97767 3485 97779 3519
rect 98730 3516 98736 3528
rect 98691 3488 98736 3516
rect 97721 3479 97779 3485
rect 98730 3476 98736 3488
rect 98788 3476 98794 3528
rect 100846 3516 100852 3528
rect 100807 3488 100852 3516
rect 100846 3476 100852 3488
rect 100904 3476 100910 3528
rect 102962 3516 102968 3528
rect 102923 3488 102968 3516
rect 102962 3476 102968 3488
rect 103020 3476 103026 3528
rect 103606 3476 103612 3528
rect 103664 3516 103670 3528
rect 104069 3519 104127 3525
rect 104069 3516 104081 3519
rect 103664 3488 104081 3516
rect 103664 3476 103670 3488
rect 104069 3485 104081 3488
rect 104115 3485 104127 3519
rect 105078 3516 105084 3528
rect 105039 3488 105084 3516
rect 104069 3479 104127 3485
rect 105078 3476 105084 3488
rect 105136 3476 105142 3528
rect 105446 3476 105452 3528
rect 105504 3516 105510 3528
rect 106185 3519 106243 3525
rect 106185 3516 106197 3519
rect 105504 3488 106197 3516
rect 105504 3476 105510 3488
rect 106185 3485 106197 3488
rect 106231 3485 106243 3519
rect 106185 3479 106243 3485
rect 1104 3290 106904 3312
rect 1104 3238 4042 3290
rect 4094 3238 4106 3290
rect 4158 3238 4170 3290
rect 4222 3238 4234 3290
rect 4286 3238 34762 3290
rect 34814 3238 34826 3290
rect 34878 3238 34890 3290
rect 34942 3238 34954 3290
rect 35006 3238 65482 3290
rect 65534 3238 65546 3290
rect 65598 3238 65610 3290
rect 65662 3238 65674 3290
rect 65726 3238 96202 3290
rect 96254 3238 96266 3290
rect 96318 3238 96330 3290
rect 96382 3238 96394 3290
rect 96446 3238 106904 3290
rect 1104 3216 106904 3238
rect 1213 3179 1271 3185
rect 1213 3145 1225 3179
rect 1259 3176 1271 3179
rect 1302 3176 1308 3188
rect 1259 3148 1308 3176
rect 1259 3145 1271 3148
rect 1213 3139 1271 3145
rect 1302 3136 1308 3148
rect 1360 3136 1366 3188
rect 40402 3136 40408 3188
rect 40460 3176 40466 3188
rect 41417 3179 41475 3185
rect 41417 3176 41429 3179
rect 40460 3148 41429 3176
rect 40460 3136 40466 3148
rect 41417 3145 41429 3148
rect 41463 3145 41475 3179
rect 77386 3176 77392 3188
rect 77347 3148 77392 3176
rect 41417 3139 41475 3145
rect 77386 3136 77392 3148
rect 77444 3136 77450 3188
rect 87046 3136 87052 3188
rect 87104 3176 87110 3188
rect 87969 3179 88027 3185
rect 87969 3176 87981 3179
rect 87104 3148 87981 3176
rect 87104 3136 87110 3148
rect 87969 3145 87981 3148
rect 88015 3145 88027 3179
rect 87969 3139 88027 3145
rect 50709 3043 50767 3049
rect 50709 3009 50721 3043
rect 50755 3040 50767 3043
rect 51905 3043 51963 3049
rect 51905 3040 51917 3043
rect 50755 3012 51917 3040
rect 50755 3009 50767 3012
rect 50709 3003 50767 3009
rect 51905 3009 51917 3012
rect 51951 3009 51963 3043
rect 51905 3003 51963 3009
rect 1305 2975 1363 2981
rect 1305 2941 1317 2975
rect 1351 2972 1363 2975
rect 1394 2972 1400 2984
rect 1351 2944 1400 2972
rect 1351 2941 1363 2944
rect 1305 2935 1363 2941
rect 1394 2932 1400 2944
rect 1452 2972 1458 2984
rect 3237 2975 3295 2981
rect 3237 2972 3249 2975
rect 1452 2944 3249 2972
rect 1452 2932 1458 2944
rect 3237 2941 3249 2944
rect 3283 2941 3295 2975
rect 3237 2935 3295 2941
rect 3421 2975 3479 2981
rect 3421 2941 3433 2975
rect 3467 2972 3479 2975
rect 3510 2972 3516 2984
rect 3467 2944 3516 2972
rect 3467 2941 3479 2944
rect 3421 2935 3479 2941
rect 3510 2932 3516 2944
rect 3568 2972 3574 2984
rect 5353 2975 5411 2981
rect 5353 2972 5365 2975
rect 3568 2944 5365 2972
rect 3568 2932 3574 2944
rect 5353 2941 5365 2944
rect 5399 2941 5411 2975
rect 5353 2935 5411 2941
rect 5537 2975 5595 2981
rect 5537 2941 5549 2975
rect 5583 2972 5595 2975
rect 5626 2972 5632 2984
rect 5583 2944 5632 2972
rect 5583 2941 5595 2944
rect 5537 2935 5595 2941
rect 5626 2932 5632 2944
rect 5684 2972 5690 2984
rect 7469 2975 7527 2981
rect 7469 2972 7481 2975
rect 5684 2944 7481 2972
rect 5684 2932 5690 2944
rect 7469 2941 7481 2944
rect 7515 2941 7527 2975
rect 7469 2935 7527 2941
rect 7653 2975 7711 2981
rect 7653 2941 7665 2975
rect 7699 2972 7711 2975
rect 7742 2972 7748 2984
rect 7699 2944 7748 2972
rect 7699 2941 7711 2944
rect 7653 2935 7711 2941
rect 7742 2932 7748 2944
rect 7800 2972 7806 2984
rect 9585 2975 9643 2981
rect 9585 2972 9597 2975
rect 7800 2944 9597 2972
rect 7800 2932 7806 2944
rect 9585 2941 9597 2944
rect 9631 2941 9643 2975
rect 9585 2935 9643 2941
rect 9769 2975 9827 2981
rect 9769 2941 9781 2975
rect 9815 2972 9827 2975
rect 9858 2972 9864 2984
rect 9815 2944 9864 2972
rect 9815 2941 9827 2944
rect 9769 2935 9827 2941
rect 9858 2932 9864 2944
rect 9916 2972 9922 2984
rect 11701 2975 11759 2981
rect 11701 2972 11713 2975
rect 9916 2944 11713 2972
rect 9916 2932 9922 2944
rect 11701 2941 11713 2944
rect 11747 2941 11759 2975
rect 11701 2935 11759 2941
rect 11885 2975 11943 2981
rect 11885 2941 11897 2975
rect 11931 2972 11943 2975
rect 11974 2972 11980 2984
rect 11931 2944 11980 2972
rect 11931 2941 11943 2944
rect 11885 2935 11943 2941
rect 11974 2932 11980 2944
rect 12032 2972 12038 2984
rect 13817 2975 13875 2981
rect 13817 2972 13829 2975
rect 12032 2944 13829 2972
rect 12032 2932 12038 2944
rect 13817 2941 13829 2944
rect 13863 2941 13875 2975
rect 13817 2935 13875 2941
rect 14001 2975 14059 2981
rect 14001 2941 14013 2975
rect 14047 2972 14059 2975
rect 14090 2972 14096 2984
rect 14047 2944 14096 2972
rect 14047 2941 14059 2944
rect 14001 2935 14059 2941
rect 14090 2932 14096 2944
rect 14148 2972 14154 2984
rect 15933 2975 15991 2981
rect 15933 2972 15945 2975
rect 14148 2944 15945 2972
rect 14148 2932 14154 2944
rect 15933 2941 15945 2944
rect 15979 2941 15991 2975
rect 18049 2975 18107 2981
rect 18049 2972 18061 2975
rect 15933 2935 15991 2941
rect 16868 2944 18061 2972
rect 16117 2907 16175 2913
rect 16117 2873 16129 2907
rect 16163 2904 16175 2907
rect 16206 2904 16212 2916
rect 16163 2876 16212 2904
rect 16163 2873 16175 2876
rect 16117 2867 16175 2873
rect 16206 2864 16212 2876
rect 16264 2904 16270 2916
rect 16868 2904 16896 2944
rect 18049 2941 18061 2944
rect 18095 2941 18107 2975
rect 18049 2935 18107 2941
rect 18233 2975 18291 2981
rect 18233 2941 18245 2975
rect 18279 2972 18291 2975
rect 18322 2972 18328 2984
rect 18279 2944 18328 2972
rect 18279 2941 18291 2944
rect 18233 2935 18291 2941
rect 18322 2932 18328 2944
rect 18380 2972 18386 2984
rect 20165 2975 20223 2981
rect 20165 2972 20177 2975
rect 18380 2944 20177 2972
rect 18380 2932 18386 2944
rect 20165 2941 20177 2944
rect 20211 2941 20223 2975
rect 20165 2935 20223 2941
rect 20349 2975 20407 2981
rect 20349 2941 20361 2975
rect 20395 2972 20407 2975
rect 20438 2972 20444 2984
rect 20395 2944 20444 2972
rect 20395 2941 20407 2944
rect 20349 2935 20407 2941
rect 20438 2932 20444 2944
rect 20496 2972 20502 2984
rect 22281 2975 22339 2981
rect 22281 2972 22293 2975
rect 20496 2944 22293 2972
rect 20496 2932 20502 2944
rect 22281 2941 22293 2944
rect 22327 2941 22339 2975
rect 22281 2935 22339 2941
rect 22465 2975 22523 2981
rect 22465 2941 22477 2975
rect 22511 2972 22523 2975
rect 22554 2972 22560 2984
rect 22511 2944 22560 2972
rect 22511 2941 22523 2944
rect 22465 2935 22523 2941
rect 22554 2932 22560 2944
rect 22612 2972 22618 2984
rect 24397 2975 24455 2981
rect 24397 2972 24409 2975
rect 22612 2944 24409 2972
rect 22612 2932 22618 2944
rect 24397 2941 24409 2944
rect 24443 2941 24455 2975
rect 24397 2935 24455 2941
rect 24581 2975 24639 2981
rect 24581 2941 24593 2975
rect 24627 2972 24639 2975
rect 24670 2972 24676 2984
rect 24627 2944 24676 2972
rect 24627 2941 24639 2944
rect 24581 2935 24639 2941
rect 24670 2932 24676 2944
rect 24728 2972 24734 2984
rect 26513 2975 26571 2981
rect 26513 2972 26525 2975
rect 24728 2944 26525 2972
rect 24728 2932 24734 2944
rect 26513 2941 26525 2944
rect 26559 2941 26571 2975
rect 26513 2935 26571 2941
rect 26697 2975 26755 2981
rect 26697 2941 26709 2975
rect 26743 2972 26755 2975
rect 26786 2972 26792 2984
rect 26743 2944 26792 2972
rect 26743 2941 26755 2944
rect 26697 2935 26755 2941
rect 26786 2932 26792 2944
rect 26844 2972 26850 2984
rect 28629 2975 28687 2981
rect 28629 2972 28641 2975
rect 26844 2944 28641 2972
rect 26844 2932 26850 2944
rect 28629 2941 28641 2944
rect 28675 2941 28687 2975
rect 28629 2935 28687 2941
rect 28813 2975 28871 2981
rect 28813 2941 28825 2975
rect 28859 2972 28871 2975
rect 28902 2972 28908 2984
rect 28859 2944 28908 2972
rect 28859 2941 28871 2944
rect 28813 2935 28871 2941
rect 28902 2932 28908 2944
rect 28960 2972 28966 2984
rect 30745 2975 30803 2981
rect 30745 2972 30757 2975
rect 28960 2944 30757 2972
rect 28960 2932 28966 2944
rect 30745 2941 30757 2944
rect 30791 2941 30803 2975
rect 30745 2935 30803 2941
rect 30929 2975 30987 2981
rect 30929 2941 30941 2975
rect 30975 2972 30987 2975
rect 31018 2972 31024 2984
rect 30975 2944 31024 2972
rect 30975 2941 30987 2944
rect 30929 2935 30987 2941
rect 31018 2932 31024 2944
rect 31076 2972 31082 2984
rect 32861 2975 32919 2981
rect 32861 2972 32873 2975
rect 31076 2944 32873 2972
rect 31076 2932 31082 2944
rect 32861 2941 32873 2944
rect 32907 2941 32919 2975
rect 34977 2975 35035 2981
rect 34977 2972 34989 2975
rect 32861 2935 32919 2941
rect 33612 2944 34989 2972
rect 16264 2876 16896 2904
rect 33045 2907 33103 2913
rect 16264 2864 16270 2876
rect 33045 2873 33057 2907
rect 33091 2904 33103 2907
rect 33134 2904 33140 2916
rect 33091 2876 33140 2904
rect 33091 2873 33103 2876
rect 33045 2867 33103 2873
rect 33134 2864 33140 2876
rect 33192 2904 33198 2916
rect 33612 2904 33640 2944
rect 34977 2941 34989 2944
rect 35023 2941 35035 2975
rect 34977 2935 35035 2941
rect 35161 2975 35219 2981
rect 35161 2941 35173 2975
rect 35207 2972 35219 2975
rect 35250 2972 35256 2984
rect 35207 2944 35256 2972
rect 35207 2941 35219 2944
rect 35161 2935 35219 2941
rect 35250 2932 35256 2944
rect 35308 2972 35314 2984
rect 37093 2975 37151 2981
rect 37093 2972 37105 2975
rect 35308 2944 37105 2972
rect 35308 2932 35314 2944
rect 37093 2941 37105 2944
rect 37139 2941 37151 2975
rect 37093 2935 37151 2941
rect 37277 2975 37335 2981
rect 37277 2941 37289 2975
rect 37323 2972 37335 2975
rect 37366 2972 37372 2984
rect 37323 2944 37372 2972
rect 37323 2941 37335 2944
rect 37277 2935 37335 2941
rect 37366 2932 37372 2944
rect 37424 2972 37430 2984
rect 39209 2975 39267 2981
rect 39209 2972 39221 2975
rect 37424 2944 39221 2972
rect 37424 2932 37430 2944
rect 39209 2941 39221 2944
rect 39255 2941 39267 2975
rect 39209 2935 39267 2941
rect 39393 2975 39451 2981
rect 39393 2941 39405 2975
rect 39439 2972 39451 2975
rect 39482 2972 39488 2984
rect 39439 2944 39488 2972
rect 39439 2941 39451 2944
rect 39393 2935 39451 2941
rect 39482 2932 39488 2944
rect 39540 2932 39546 2984
rect 41509 2975 41567 2981
rect 41509 2941 41521 2975
rect 41555 2972 41567 2975
rect 41598 2972 41604 2984
rect 41555 2944 41604 2972
rect 41555 2941 41567 2944
rect 41509 2935 41567 2941
rect 41598 2932 41604 2944
rect 41656 2972 41662 2984
rect 43441 2975 43499 2981
rect 43441 2972 43453 2975
rect 41656 2944 43453 2972
rect 41656 2932 41662 2944
rect 43441 2941 43453 2944
rect 43487 2941 43499 2975
rect 43441 2935 43499 2941
rect 43625 2975 43683 2981
rect 43625 2941 43637 2975
rect 43671 2972 43683 2975
rect 43714 2972 43720 2984
rect 43671 2944 43720 2972
rect 43671 2941 43683 2944
rect 43625 2935 43683 2941
rect 43714 2932 43720 2944
rect 43772 2972 43778 2984
rect 45557 2975 45615 2981
rect 45557 2972 45569 2975
rect 43772 2944 45569 2972
rect 43772 2932 43778 2944
rect 45557 2941 45569 2944
rect 45603 2941 45615 2975
rect 45557 2935 45615 2941
rect 45741 2975 45799 2981
rect 45741 2941 45753 2975
rect 45787 2972 45799 2975
rect 45830 2972 45836 2984
rect 45787 2944 45836 2972
rect 45787 2941 45799 2944
rect 45741 2935 45799 2941
rect 45830 2932 45836 2944
rect 45888 2972 45894 2984
rect 47673 2975 47731 2981
rect 47673 2972 47685 2975
rect 45888 2944 47685 2972
rect 45888 2932 45894 2944
rect 47673 2941 47685 2944
rect 47719 2941 47731 2975
rect 47673 2935 47731 2941
rect 47857 2975 47915 2981
rect 47857 2941 47869 2975
rect 47903 2972 47915 2975
rect 47946 2972 47952 2984
rect 47903 2944 47952 2972
rect 47903 2941 47915 2944
rect 47857 2935 47915 2941
rect 47946 2932 47952 2944
rect 48004 2972 48010 2984
rect 49789 2975 49847 2981
rect 49789 2972 49801 2975
rect 48004 2944 49801 2972
rect 48004 2932 48010 2944
rect 49789 2941 49801 2944
rect 49835 2941 49847 2975
rect 49789 2935 49847 2941
rect 52089 2975 52147 2981
rect 52089 2941 52101 2975
rect 52135 2972 52147 2975
rect 52178 2972 52184 2984
rect 52135 2944 52184 2972
rect 52135 2941 52147 2944
rect 52089 2935 52147 2941
rect 52178 2932 52184 2944
rect 52236 2972 52242 2984
rect 54021 2975 54079 2981
rect 54021 2972 54033 2975
rect 52236 2944 54033 2972
rect 52236 2932 52242 2944
rect 54021 2941 54033 2944
rect 54067 2941 54079 2975
rect 54021 2935 54079 2941
rect 54205 2975 54263 2981
rect 54205 2941 54217 2975
rect 54251 2972 54263 2975
rect 54294 2972 54300 2984
rect 54251 2944 54300 2972
rect 54251 2941 54263 2944
rect 54205 2935 54263 2941
rect 54294 2932 54300 2944
rect 54352 2972 54358 2984
rect 56137 2975 56195 2981
rect 56137 2972 56149 2975
rect 54352 2944 56149 2972
rect 54352 2932 54358 2944
rect 56137 2941 56149 2944
rect 56183 2941 56195 2975
rect 56137 2935 56195 2941
rect 56321 2975 56379 2981
rect 56321 2941 56333 2975
rect 56367 2972 56379 2975
rect 56410 2972 56416 2984
rect 56367 2944 56416 2972
rect 56367 2941 56379 2944
rect 56321 2935 56379 2941
rect 56410 2932 56416 2944
rect 56468 2972 56474 2984
rect 58253 2975 58311 2981
rect 58253 2972 58265 2975
rect 56468 2944 58265 2972
rect 56468 2932 56474 2944
rect 58253 2941 58265 2944
rect 58299 2941 58311 2975
rect 58253 2935 58311 2941
rect 58437 2975 58495 2981
rect 58437 2941 58449 2975
rect 58483 2972 58495 2975
rect 58526 2972 58532 2984
rect 58483 2944 58532 2972
rect 58483 2941 58495 2944
rect 58437 2935 58495 2941
rect 58526 2932 58532 2944
rect 58584 2972 58590 2984
rect 60369 2975 60427 2981
rect 60369 2972 60381 2975
rect 58584 2944 60381 2972
rect 58584 2932 58590 2944
rect 60369 2941 60381 2944
rect 60415 2941 60427 2975
rect 60369 2935 60427 2941
rect 60553 2975 60611 2981
rect 60553 2941 60565 2975
rect 60599 2972 60611 2975
rect 60642 2972 60648 2984
rect 60599 2944 60648 2972
rect 60599 2941 60611 2944
rect 60553 2935 60611 2941
rect 60642 2932 60648 2944
rect 60700 2972 60706 2984
rect 62485 2975 62543 2981
rect 62485 2972 62497 2975
rect 60700 2944 62497 2972
rect 60700 2932 60706 2944
rect 62485 2941 62497 2944
rect 62531 2941 62543 2975
rect 62485 2935 62543 2941
rect 62669 2975 62727 2981
rect 62669 2941 62681 2975
rect 62715 2972 62727 2975
rect 62758 2972 62764 2984
rect 62715 2944 62764 2972
rect 62715 2941 62727 2944
rect 62669 2935 62727 2941
rect 62758 2932 62764 2944
rect 62816 2972 62822 2984
rect 64601 2975 64659 2981
rect 64601 2972 64613 2975
rect 62816 2944 64613 2972
rect 62816 2932 62822 2944
rect 64601 2941 64613 2944
rect 64647 2941 64659 2975
rect 64601 2935 64659 2941
rect 64785 2975 64843 2981
rect 64785 2941 64797 2975
rect 64831 2972 64843 2975
rect 64874 2972 64880 2984
rect 64831 2944 64880 2972
rect 64831 2941 64843 2944
rect 64785 2935 64843 2941
rect 64874 2932 64880 2944
rect 64932 2972 64938 2984
rect 66717 2975 66775 2981
rect 66717 2972 66729 2975
rect 64932 2944 66729 2972
rect 64932 2932 64938 2944
rect 66717 2941 66729 2944
rect 66763 2941 66775 2975
rect 68833 2975 68891 2981
rect 68833 2972 68845 2975
rect 66717 2935 66775 2941
rect 67652 2944 68845 2972
rect 33192 2876 33640 2904
rect 49973 2907 50031 2913
rect 33192 2864 33198 2876
rect 49973 2873 49985 2907
rect 50019 2904 50031 2907
rect 50062 2904 50068 2916
rect 50019 2876 50068 2904
rect 50019 2873 50031 2876
rect 49973 2867 50031 2873
rect 50062 2864 50068 2876
rect 50120 2904 50126 2916
rect 50709 2907 50767 2913
rect 50709 2904 50721 2907
rect 50120 2876 50721 2904
rect 50120 2864 50126 2876
rect 50709 2873 50721 2876
rect 50755 2873 50767 2907
rect 50709 2867 50767 2873
rect 66901 2907 66959 2913
rect 66901 2873 66913 2907
rect 66947 2904 66959 2907
rect 66990 2904 66996 2916
rect 66947 2876 66996 2904
rect 66947 2873 66959 2876
rect 66901 2867 66959 2873
rect 66990 2864 66996 2876
rect 67048 2904 67054 2916
rect 67652 2904 67680 2944
rect 68833 2941 68845 2944
rect 68879 2941 68891 2975
rect 68833 2935 68891 2941
rect 69017 2975 69075 2981
rect 69017 2941 69029 2975
rect 69063 2972 69075 2975
rect 69106 2972 69112 2984
rect 69063 2944 69112 2972
rect 69063 2941 69075 2944
rect 69017 2935 69075 2941
rect 69106 2932 69112 2944
rect 69164 2972 69170 2984
rect 70949 2975 71007 2981
rect 70949 2972 70961 2975
rect 69164 2944 70961 2972
rect 69164 2932 69170 2944
rect 70949 2941 70961 2944
rect 70995 2941 71007 2975
rect 70949 2935 71007 2941
rect 71133 2975 71191 2981
rect 71133 2941 71145 2975
rect 71179 2972 71191 2975
rect 71222 2972 71228 2984
rect 71179 2944 71228 2972
rect 71179 2941 71191 2944
rect 71133 2935 71191 2941
rect 71222 2932 71228 2944
rect 71280 2972 71286 2984
rect 73065 2975 73123 2981
rect 73065 2972 73077 2975
rect 71280 2944 73077 2972
rect 71280 2932 71286 2944
rect 73065 2941 73077 2944
rect 73111 2941 73123 2975
rect 73065 2935 73123 2941
rect 73249 2975 73307 2981
rect 73249 2941 73261 2975
rect 73295 2972 73307 2975
rect 73338 2972 73344 2984
rect 73295 2944 73344 2972
rect 73295 2941 73307 2944
rect 73249 2935 73307 2941
rect 73338 2932 73344 2944
rect 73396 2972 73402 2984
rect 75181 2975 75239 2981
rect 75181 2972 75193 2975
rect 73396 2944 75193 2972
rect 73396 2932 73402 2944
rect 75181 2941 75193 2944
rect 75227 2941 75239 2975
rect 75362 2972 75368 2984
rect 75323 2944 75368 2972
rect 75181 2935 75239 2941
rect 75362 2932 75368 2944
rect 75420 2932 75426 2984
rect 77481 2975 77539 2981
rect 77481 2941 77493 2975
rect 77527 2972 77539 2975
rect 77570 2972 77576 2984
rect 77527 2944 77576 2972
rect 77527 2941 77539 2944
rect 77481 2935 77539 2941
rect 77570 2932 77576 2944
rect 77628 2972 77634 2984
rect 79413 2975 79471 2981
rect 79413 2972 79425 2975
rect 77628 2944 79425 2972
rect 77628 2932 77634 2944
rect 79413 2941 79425 2944
rect 79459 2941 79471 2975
rect 79413 2935 79471 2941
rect 79597 2975 79655 2981
rect 79597 2941 79609 2975
rect 79643 2972 79655 2975
rect 79686 2972 79692 2984
rect 79643 2944 79692 2972
rect 79643 2941 79655 2944
rect 79597 2935 79655 2941
rect 79686 2932 79692 2944
rect 79744 2972 79750 2984
rect 81529 2975 81587 2981
rect 81529 2972 81541 2975
rect 79744 2944 81541 2972
rect 79744 2932 79750 2944
rect 81529 2941 81541 2944
rect 81575 2941 81587 2975
rect 81529 2935 81587 2941
rect 81713 2975 81771 2981
rect 81713 2941 81725 2975
rect 81759 2972 81771 2975
rect 81802 2972 81808 2984
rect 81759 2944 81808 2972
rect 81759 2941 81771 2944
rect 81713 2935 81771 2941
rect 81802 2932 81808 2944
rect 81860 2972 81866 2984
rect 83645 2975 83703 2981
rect 83645 2972 83657 2975
rect 81860 2944 83657 2972
rect 81860 2932 81866 2944
rect 83645 2941 83657 2944
rect 83691 2941 83703 2975
rect 85761 2975 85819 2981
rect 85761 2972 85773 2975
rect 83645 2935 83703 2941
rect 84580 2944 85773 2972
rect 67048 2876 67680 2904
rect 83829 2907 83887 2913
rect 67048 2864 67054 2876
rect 83829 2873 83841 2907
rect 83875 2904 83887 2907
rect 83918 2904 83924 2916
rect 83875 2876 83924 2904
rect 83875 2873 83887 2876
rect 83829 2867 83887 2873
rect 83918 2864 83924 2876
rect 83976 2904 83982 2916
rect 84580 2904 84608 2944
rect 85761 2941 85773 2944
rect 85807 2941 85819 2975
rect 85942 2972 85948 2984
rect 85903 2944 85948 2972
rect 85761 2935 85819 2941
rect 85942 2932 85948 2944
rect 86000 2932 86006 2984
rect 88061 2975 88119 2981
rect 88061 2941 88073 2975
rect 88107 2972 88119 2975
rect 88150 2972 88156 2984
rect 88107 2944 88156 2972
rect 88107 2941 88119 2944
rect 88061 2935 88119 2941
rect 88150 2932 88156 2944
rect 88208 2972 88214 2984
rect 89993 2975 90051 2981
rect 89993 2972 90005 2975
rect 88208 2944 90005 2972
rect 88208 2932 88214 2944
rect 89993 2941 90005 2944
rect 90039 2941 90051 2975
rect 89993 2935 90051 2941
rect 90177 2975 90235 2981
rect 90177 2941 90189 2975
rect 90223 2972 90235 2975
rect 90266 2972 90272 2984
rect 90223 2944 90272 2972
rect 90223 2941 90235 2944
rect 90177 2935 90235 2941
rect 90266 2932 90272 2944
rect 90324 2972 90330 2984
rect 92109 2975 92167 2981
rect 92109 2972 92121 2975
rect 90324 2944 92121 2972
rect 90324 2932 90330 2944
rect 92109 2941 92121 2944
rect 92155 2941 92167 2975
rect 92109 2935 92167 2941
rect 92293 2975 92351 2981
rect 92293 2941 92305 2975
rect 92339 2972 92351 2975
rect 92382 2972 92388 2984
rect 92339 2944 92388 2972
rect 92339 2941 92351 2944
rect 92293 2935 92351 2941
rect 92382 2932 92388 2944
rect 92440 2972 92446 2984
rect 94225 2975 94283 2981
rect 94225 2972 94237 2975
rect 92440 2944 94237 2972
rect 92440 2932 92446 2944
rect 94225 2941 94237 2944
rect 94271 2941 94283 2975
rect 94225 2935 94283 2941
rect 94409 2975 94467 2981
rect 94409 2941 94421 2975
rect 94455 2972 94467 2975
rect 94498 2972 94504 2984
rect 94455 2944 94504 2972
rect 94455 2941 94467 2944
rect 94409 2935 94467 2941
rect 94498 2932 94504 2944
rect 94556 2972 94562 2984
rect 96341 2975 96399 2981
rect 96341 2972 96353 2975
rect 94556 2944 96353 2972
rect 94556 2932 94562 2944
rect 96341 2941 96353 2944
rect 96387 2941 96399 2975
rect 96341 2935 96399 2941
rect 96525 2975 96583 2981
rect 96525 2941 96537 2975
rect 96571 2972 96583 2975
rect 96614 2972 96620 2984
rect 96571 2944 96620 2972
rect 96571 2941 96583 2944
rect 96525 2935 96583 2941
rect 96614 2932 96620 2944
rect 96672 2972 96678 2984
rect 98457 2975 98515 2981
rect 98457 2972 98469 2975
rect 96672 2944 98469 2972
rect 96672 2932 96678 2944
rect 98457 2941 98469 2944
rect 98503 2941 98515 2975
rect 98457 2935 98515 2941
rect 98641 2975 98699 2981
rect 98641 2941 98653 2975
rect 98687 2972 98699 2975
rect 98730 2972 98736 2984
rect 98687 2944 98736 2972
rect 98687 2941 98699 2944
rect 98641 2935 98699 2941
rect 98730 2932 98736 2944
rect 98788 2972 98794 2984
rect 100573 2975 100631 2981
rect 100573 2972 100585 2975
rect 98788 2944 100585 2972
rect 98788 2932 98794 2944
rect 100573 2941 100585 2944
rect 100619 2941 100631 2975
rect 100573 2935 100631 2941
rect 100757 2975 100815 2981
rect 100757 2941 100769 2975
rect 100803 2972 100815 2975
rect 100846 2972 100852 2984
rect 100803 2944 100852 2972
rect 100803 2941 100815 2944
rect 100757 2935 100815 2941
rect 100846 2932 100852 2944
rect 100904 2972 100910 2984
rect 102689 2975 102747 2981
rect 102689 2972 102701 2975
rect 100904 2944 102701 2972
rect 100904 2932 100910 2944
rect 102689 2941 102701 2944
rect 102735 2941 102747 2975
rect 102689 2935 102747 2941
rect 102873 2975 102931 2981
rect 102873 2941 102885 2975
rect 102919 2972 102931 2975
rect 102962 2972 102968 2984
rect 102919 2944 102968 2972
rect 102919 2941 102931 2944
rect 102873 2935 102931 2941
rect 102962 2932 102968 2944
rect 103020 2972 103026 2984
rect 104805 2975 104863 2981
rect 104805 2972 104817 2975
rect 103020 2944 104817 2972
rect 103020 2932 103026 2944
rect 104805 2941 104817 2944
rect 104851 2941 104863 2975
rect 104805 2935 104863 2941
rect 104989 2975 105047 2981
rect 104989 2941 105001 2975
rect 105035 2972 105047 2975
rect 105078 2972 105084 2984
rect 105035 2944 105084 2972
rect 105035 2941 105047 2944
rect 104989 2935 105047 2941
rect 105078 2932 105084 2944
rect 105136 2932 105142 2984
rect 83976 2876 84608 2904
rect 83976 2864 83982 2876
rect 1104 2746 106904 2768
rect 1104 2694 19402 2746
rect 19454 2694 19466 2746
rect 19518 2694 19530 2746
rect 19582 2694 19594 2746
rect 19646 2694 50122 2746
rect 50174 2694 50186 2746
rect 50238 2694 50250 2746
rect 50302 2694 50314 2746
rect 50366 2694 80842 2746
rect 80894 2694 80906 2746
rect 80958 2694 80970 2746
rect 81022 2694 81034 2746
rect 81086 2694 106904 2746
rect 1104 2672 106904 2694
rect 5537 2635 5595 2641
rect 5537 2601 5549 2635
rect 5583 2601 5595 2635
rect 5537 2595 5595 2601
rect 20349 2635 20407 2641
rect 20349 2601 20361 2635
rect 20395 2632 20407 2635
rect 22465 2635 22523 2641
rect 20395 2604 22416 2632
rect 20395 2601 20407 2604
rect 20349 2595 20407 2601
rect 5552 2564 5580 2595
rect 22388 2576 22416 2604
rect 22465 2601 22477 2635
rect 22511 2601 22523 2635
rect 22465 2595 22523 2601
rect 7561 2567 7619 2573
rect 7561 2564 7573 2567
rect 5552 2536 7573 2564
rect 7561 2533 7573 2536
rect 7607 2564 7619 2567
rect 7742 2564 7748 2576
rect 7607 2536 7748 2564
rect 7607 2533 7619 2536
rect 7561 2527 7619 2533
rect 7742 2524 7748 2536
rect 7800 2524 7806 2576
rect 9861 2567 9919 2573
rect 9861 2533 9873 2567
rect 9907 2564 9919 2567
rect 11793 2567 11851 2573
rect 11793 2564 11805 2567
rect 9907 2536 11805 2564
rect 9907 2533 9919 2536
rect 9861 2527 9919 2533
rect 11793 2533 11805 2536
rect 11839 2564 11851 2567
rect 11882 2564 11888 2576
rect 11839 2536 11888 2564
rect 11839 2533 11851 2536
rect 11793 2527 11851 2533
rect 11882 2524 11888 2536
rect 11940 2524 11946 2576
rect 11977 2567 12035 2573
rect 11977 2533 11989 2567
rect 12023 2564 12035 2567
rect 13909 2567 13967 2573
rect 13909 2564 13921 2567
rect 12023 2536 13921 2564
rect 12023 2533 12035 2536
rect 11977 2527 12035 2533
rect 13909 2533 13921 2536
rect 13955 2564 13967 2567
rect 14090 2564 14096 2576
rect 13955 2536 14096 2564
rect 13955 2533 13967 2536
rect 13909 2527 13967 2533
rect 14090 2524 14096 2536
rect 14148 2524 14154 2576
rect 22370 2564 22376 2576
rect 22331 2536 22376 2564
rect 22370 2524 22376 2536
rect 22428 2524 22434 2576
rect 22480 2564 22508 2595
rect 23382 2592 23388 2644
rect 23440 2632 23446 2644
rect 23750 2632 23756 2644
rect 23440 2604 23756 2632
rect 23440 2592 23446 2604
rect 23750 2592 23756 2604
rect 23808 2592 23814 2644
rect 30929 2635 30987 2641
rect 30929 2601 30941 2635
rect 30975 2601 30987 2635
rect 33134 2632 33140 2644
rect 30929 2595 30987 2601
rect 32968 2604 33140 2632
rect 24489 2567 24547 2573
rect 24489 2564 24501 2567
rect 22480 2536 24501 2564
rect 24489 2533 24501 2536
rect 24535 2564 24547 2567
rect 24670 2564 24676 2576
rect 24535 2536 24676 2564
rect 24535 2533 24547 2536
rect 24489 2527 24547 2533
rect 24670 2524 24676 2536
rect 24728 2524 24734 2576
rect 30944 2564 30972 2595
rect 32968 2573 32996 2604
rect 33134 2592 33140 2604
rect 33192 2592 33198 2644
rect 35161 2635 35219 2641
rect 35161 2601 35173 2635
rect 35207 2632 35219 2635
rect 41509 2635 41567 2641
rect 35207 2604 37228 2632
rect 35207 2601 35219 2604
rect 35161 2595 35219 2601
rect 37200 2573 37228 2604
rect 41509 2601 41521 2635
rect 41555 2601 41567 2635
rect 41509 2595 41567 2601
rect 60553 2635 60611 2641
rect 60553 2601 60565 2635
rect 60599 2601 60611 2635
rect 60553 2595 60611 2601
rect 71133 2635 71191 2641
rect 71133 2601 71145 2635
rect 71179 2632 71191 2635
rect 77481 2635 77539 2641
rect 71179 2604 73200 2632
rect 71179 2601 71191 2604
rect 71133 2595 71191 2601
rect 32953 2567 33011 2573
rect 32953 2564 32965 2567
rect 30944 2536 32965 2564
rect 32953 2533 32965 2536
rect 32999 2533 33011 2567
rect 32953 2527 33011 2533
rect 37185 2567 37243 2573
rect 37185 2533 37197 2567
rect 37231 2564 37243 2567
rect 37366 2564 37372 2576
rect 37231 2536 37372 2564
rect 37231 2533 37243 2536
rect 37185 2527 37243 2533
rect 37366 2524 37372 2536
rect 37424 2524 37430 2576
rect 41524 2564 41552 2595
rect 43533 2567 43591 2573
rect 43533 2564 43545 2567
rect 41524 2536 43545 2564
rect 43533 2533 43545 2536
rect 43579 2564 43591 2567
rect 43714 2564 43720 2576
rect 43579 2536 43720 2564
rect 43579 2533 43591 2536
rect 43533 2527 43591 2533
rect 43714 2524 43720 2536
rect 43772 2524 43778 2576
rect 45833 2567 45891 2573
rect 45833 2533 45845 2567
rect 45879 2564 45891 2567
rect 47765 2567 47823 2573
rect 47765 2564 47777 2567
rect 45879 2536 47777 2564
rect 45879 2533 45891 2536
rect 45833 2527 45891 2533
rect 47765 2533 47777 2536
rect 47811 2564 47823 2567
rect 47854 2564 47860 2576
rect 47811 2536 47860 2564
rect 47811 2533 47823 2536
rect 47765 2527 47823 2533
rect 47854 2524 47860 2536
rect 47912 2524 47918 2576
rect 56413 2567 56471 2573
rect 56413 2533 56425 2567
rect 56459 2564 56471 2567
rect 58345 2567 58403 2573
rect 58345 2564 58357 2567
rect 56459 2536 58357 2564
rect 56459 2533 56471 2536
rect 56413 2527 56471 2533
rect 58345 2533 58357 2536
rect 58391 2564 58403 2567
rect 58434 2564 58440 2576
rect 58391 2536 58440 2564
rect 58391 2533 58403 2536
rect 58345 2527 58403 2533
rect 58434 2524 58440 2536
rect 58492 2524 58498 2576
rect 58529 2567 58587 2573
rect 58529 2533 58541 2567
rect 58575 2564 58587 2567
rect 60458 2564 60464 2576
rect 58575 2536 60464 2564
rect 58575 2533 58587 2536
rect 58529 2527 58587 2533
rect 60458 2524 60464 2536
rect 60516 2524 60522 2576
rect 60568 2564 60596 2595
rect 62577 2567 62635 2573
rect 62577 2564 62589 2567
rect 60568 2536 62589 2564
rect 62577 2533 62589 2536
rect 62623 2564 62635 2567
rect 62758 2564 62764 2576
rect 62623 2536 62764 2564
rect 62623 2533 62635 2536
rect 62577 2527 62635 2533
rect 62758 2524 62764 2536
rect 62816 2524 62822 2576
rect 73172 2573 73200 2604
rect 77481 2601 77493 2635
rect 77527 2601 77539 2635
rect 77481 2595 77539 2601
rect 96525 2635 96583 2641
rect 96525 2601 96537 2635
rect 96571 2632 96583 2635
rect 102873 2635 102931 2641
rect 96571 2604 98592 2632
rect 96571 2601 96583 2604
rect 96525 2595 96583 2601
rect 73157 2567 73215 2573
rect 73157 2533 73169 2567
rect 73203 2564 73215 2567
rect 73338 2564 73344 2576
rect 73203 2536 73344 2564
rect 73203 2533 73215 2536
rect 73157 2527 73215 2533
rect 73338 2524 73344 2536
rect 73396 2524 73402 2576
rect 77496 2564 77524 2595
rect 79505 2567 79563 2573
rect 79505 2564 79517 2567
rect 77496 2536 79517 2564
rect 79505 2533 79517 2536
rect 79551 2564 79563 2567
rect 79594 2564 79600 2576
rect 79551 2536 79600 2564
rect 79551 2533 79563 2536
rect 79505 2527 79563 2533
rect 79594 2524 79600 2536
rect 79652 2524 79658 2576
rect 88153 2567 88211 2573
rect 88153 2533 88165 2567
rect 88199 2564 88211 2567
rect 90085 2567 90143 2573
rect 90085 2564 90097 2567
rect 88199 2536 90097 2564
rect 88199 2533 88211 2536
rect 88153 2527 88211 2533
rect 90085 2533 90097 2536
rect 90131 2564 90143 2567
rect 90266 2564 90272 2576
rect 90131 2536 90272 2564
rect 90131 2533 90143 2536
rect 90085 2527 90143 2533
rect 90266 2524 90272 2536
rect 90324 2524 90330 2576
rect 92385 2567 92443 2573
rect 92385 2533 92397 2567
rect 92431 2564 92443 2567
rect 94317 2567 94375 2573
rect 94317 2564 94329 2567
rect 92431 2536 94329 2564
rect 92431 2533 92443 2536
rect 92385 2527 92443 2533
rect 94317 2533 94329 2536
rect 94363 2564 94375 2567
rect 94406 2564 94412 2576
rect 94363 2536 94412 2564
rect 94363 2533 94375 2536
rect 94317 2527 94375 2533
rect 94406 2524 94412 2536
rect 94464 2524 94470 2576
rect 94501 2567 94559 2573
rect 94501 2533 94513 2567
rect 94547 2564 94559 2567
rect 96433 2567 96491 2573
rect 96433 2564 96445 2567
rect 94547 2536 96445 2564
rect 94547 2533 94559 2536
rect 94501 2527 94559 2533
rect 96433 2533 96445 2536
rect 96479 2564 96491 2567
rect 96614 2564 96620 2576
rect 96479 2536 96620 2564
rect 96479 2533 96491 2536
rect 96433 2527 96491 2533
rect 96614 2524 96620 2536
rect 96672 2524 96678 2576
rect 98564 2573 98592 2604
rect 102873 2601 102885 2635
rect 102919 2632 102931 2635
rect 102919 2604 104940 2632
rect 102919 2601 102931 2604
rect 102873 2595 102931 2601
rect 104912 2576 104940 2604
rect 98549 2567 98607 2573
rect 98549 2533 98561 2567
rect 98595 2564 98607 2567
rect 98730 2564 98736 2576
rect 98595 2536 98736 2564
rect 98595 2533 98607 2536
rect 98549 2527 98607 2533
rect 98730 2524 98736 2536
rect 98788 2524 98794 2576
rect 102597 2567 102655 2573
rect 102597 2533 102609 2567
rect 102643 2564 102655 2567
rect 102781 2567 102839 2573
rect 102781 2564 102793 2567
rect 102643 2536 102793 2564
rect 102643 2533 102655 2536
rect 102597 2527 102655 2533
rect 102781 2533 102793 2536
rect 102827 2533 102839 2567
rect 104894 2564 104900 2576
rect 104807 2536 104900 2564
rect 102781 2527 102839 2533
rect 104894 2524 104900 2536
rect 104952 2524 104958 2576
rect 105078 2564 105084 2576
rect 105039 2536 105084 2564
rect 105078 2524 105084 2536
rect 105136 2524 105142 2576
rect 1210 2496 1216 2508
rect 1171 2468 1216 2496
rect 1210 2456 1216 2468
rect 1268 2456 1274 2508
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2496 1455 2499
rect 3329 2499 3387 2505
rect 3329 2496 3341 2499
rect 1443 2468 3341 2496
rect 1443 2465 1455 2468
rect 1397 2459 1455 2465
rect 3329 2465 3341 2468
rect 3375 2496 3387 2499
rect 3510 2496 3516 2508
rect 3375 2468 3516 2496
rect 3375 2465 3387 2468
rect 3329 2459 3387 2465
rect 3510 2456 3516 2468
rect 3568 2456 3574 2508
rect 5445 2499 5503 2505
rect 5445 2496 5457 2499
rect 4908 2468 5457 2496
rect 3421 2295 3479 2301
rect 3421 2261 3433 2295
rect 3467 2292 3479 2295
rect 4908 2292 4936 2468
rect 5445 2465 5457 2468
rect 5491 2496 5503 2499
rect 5626 2496 5632 2508
rect 5491 2468 5632 2496
rect 5491 2465 5503 2468
rect 5445 2459 5503 2465
rect 5626 2456 5632 2468
rect 5684 2456 5690 2508
rect 9677 2499 9735 2505
rect 9677 2465 9689 2499
rect 9723 2465 9735 2499
rect 16025 2499 16083 2505
rect 16025 2496 16037 2499
rect 9677 2459 9735 2465
rect 14108 2468 16037 2496
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2428 7803 2431
rect 9692 2428 9720 2459
rect 9858 2428 9864 2440
rect 7791 2400 9864 2428
rect 7791 2397 7803 2400
rect 7745 2391 7803 2397
rect 9858 2388 9864 2400
rect 9916 2388 9922 2440
rect 14108 2437 14136 2468
rect 16025 2465 16037 2468
rect 16071 2496 16083 2499
rect 16206 2496 16212 2508
rect 16071 2468 16212 2496
rect 16071 2465 16083 2468
rect 16025 2459 16083 2465
rect 16206 2456 16212 2468
rect 16264 2456 16270 2508
rect 18141 2499 18199 2505
rect 18141 2465 18153 2499
rect 18187 2465 18199 2499
rect 18141 2459 18199 2465
rect 18325 2499 18383 2505
rect 18325 2465 18337 2499
rect 18371 2496 18383 2499
rect 20257 2499 20315 2505
rect 20257 2496 20269 2499
rect 18371 2468 20269 2496
rect 18371 2465 18383 2468
rect 18325 2459 18383 2465
rect 20257 2465 20269 2468
rect 20303 2496 20315 2499
rect 20438 2496 20444 2508
rect 20303 2468 20444 2496
rect 20303 2465 20315 2468
rect 20257 2459 20315 2465
rect 14093 2431 14151 2437
rect 14093 2397 14105 2431
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 16209 2363 16267 2369
rect 16209 2329 16221 2363
rect 16255 2360 16267 2363
rect 18156 2360 18184 2459
rect 20438 2456 20444 2468
rect 20496 2456 20502 2508
rect 26605 2499 26663 2505
rect 26605 2465 26617 2499
rect 26651 2465 26663 2499
rect 26605 2459 26663 2465
rect 28721 2499 28779 2505
rect 28721 2465 28733 2499
rect 28767 2465 28779 2499
rect 28721 2459 28779 2465
rect 28905 2499 28963 2505
rect 28905 2465 28917 2499
rect 28951 2496 28963 2499
rect 30837 2499 30895 2505
rect 30837 2496 30849 2499
rect 28951 2468 30849 2496
rect 28951 2465 28963 2468
rect 28905 2459 28963 2465
rect 30837 2465 30849 2468
rect 30883 2496 30895 2499
rect 31018 2496 31024 2508
rect 30883 2468 31024 2496
rect 30883 2465 30895 2468
rect 30837 2459 30895 2465
rect 24673 2431 24731 2437
rect 24673 2397 24685 2431
rect 24719 2428 24731 2431
rect 26620 2428 26648 2459
rect 26694 2428 26700 2440
rect 24719 2400 26700 2428
rect 24719 2397 24731 2400
rect 24673 2391 24731 2397
rect 26694 2388 26700 2400
rect 26752 2388 26758 2440
rect 26789 2431 26847 2437
rect 26789 2397 26801 2431
rect 26835 2428 26847 2431
rect 28736 2428 28764 2459
rect 31018 2456 31024 2468
rect 31076 2456 31082 2508
rect 33137 2499 33195 2505
rect 33137 2465 33149 2499
rect 33183 2496 33195 2499
rect 35069 2499 35127 2505
rect 35069 2496 35081 2499
rect 33183 2468 35081 2496
rect 33183 2465 33195 2468
rect 33137 2459 33195 2465
rect 35069 2465 35081 2468
rect 35115 2496 35127 2499
rect 35250 2496 35256 2508
rect 35115 2468 35256 2496
rect 35115 2465 35127 2468
rect 35069 2459 35127 2465
rect 35250 2456 35256 2468
rect 35308 2456 35314 2508
rect 39301 2499 39359 2505
rect 39301 2465 39313 2499
rect 39347 2465 39359 2499
rect 41417 2499 41475 2505
rect 41417 2496 41429 2499
rect 39301 2459 39359 2465
rect 40880 2468 41429 2496
rect 28810 2428 28816 2440
rect 26835 2400 28816 2428
rect 26835 2397 26847 2400
rect 26789 2391 26847 2397
rect 28810 2388 28816 2400
rect 28868 2388 28874 2440
rect 37369 2431 37427 2437
rect 37369 2397 37381 2431
rect 37415 2428 37427 2431
rect 39316 2428 39344 2459
rect 39390 2428 39396 2440
rect 37415 2400 39396 2428
rect 37415 2397 37427 2400
rect 37369 2391 37427 2397
rect 39390 2388 39396 2400
rect 39448 2388 39454 2440
rect 18322 2360 18328 2372
rect 16255 2332 18328 2360
rect 16255 2329 16267 2332
rect 16209 2323 16267 2329
rect 18322 2320 18328 2332
rect 18380 2320 18386 2372
rect 39485 2363 39543 2369
rect 39485 2329 39497 2363
rect 39531 2360 39543 2363
rect 40880 2360 40908 2468
rect 41417 2465 41429 2468
rect 41463 2496 41475 2499
rect 41598 2496 41604 2508
rect 41463 2468 41604 2496
rect 41463 2465 41475 2468
rect 41417 2459 41475 2465
rect 41598 2456 41604 2468
rect 41656 2456 41662 2508
rect 45649 2499 45707 2505
rect 45649 2465 45661 2499
rect 45695 2465 45707 2499
rect 45649 2459 45707 2465
rect 47949 2499 48007 2505
rect 47949 2465 47961 2499
rect 47995 2496 48007 2499
rect 49881 2499 49939 2505
rect 49881 2496 49893 2499
rect 47995 2468 49893 2496
rect 47995 2465 48007 2468
rect 47949 2459 48007 2465
rect 49881 2465 49893 2468
rect 49927 2496 49939 2499
rect 50062 2496 50068 2508
rect 49927 2468 50068 2496
rect 49927 2465 49939 2468
rect 49881 2459 49939 2465
rect 43717 2431 43775 2437
rect 43717 2397 43729 2431
rect 43763 2428 43775 2431
rect 45664 2428 45692 2459
rect 50062 2456 50068 2468
rect 50120 2456 50126 2508
rect 51997 2499 52055 2505
rect 51997 2465 52009 2499
rect 52043 2465 52055 2499
rect 51997 2459 52055 2465
rect 52181 2499 52239 2505
rect 52181 2465 52193 2499
rect 52227 2496 52239 2499
rect 54113 2499 54171 2505
rect 54113 2496 54125 2499
rect 52227 2468 54125 2496
rect 52227 2465 52239 2468
rect 52181 2459 52239 2465
rect 54113 2465 54125 2468
rect 54159 2496 54171 2499
rect 54202 2496 54208 2508
rect 54159 2468 54208 2496
rect 54159 2465 54171 2468
rect 54113 2459 54171 2465
rect 45830 2428 45836 2440
rect 43763 2400 45836 2428
rect 43763 2397 43775 2400
rect 43717 2391 43775 2397
rect 45830 2388 45836 2400
rect 45888 2388 45894 2440
rect 39531 2332 40908 2360
rect 50065 2363 50123 2369
rect 39531 2329 39543 2332
rect 39485 2323 39543 2329
rect 50065 2329 50077 2363
rect 50111 2360 50123 2363
rect 52012 2360 52040 2459
rect 54202 2456 54208 2468
rect 54260 2456 54266 2508
rect 56229 2499 56287 2505
rect 56229 2465 56241 2499
rect 56275 2465 56287 2499
rect 64693 2499 64751 2505
rect 64693 2496 64705 2499
rect 56229 2459 56287 2465
rect 62776 2468 64705 2496
rect 54297 2431 54355 2437
rect 54297 2397 54309 2431
rect 54343 2428 54355 2431
rect 56244 2428 56272 2459
rect 56410 2428 56416 2440
rect 54343 2400 56416 2428
rect 54343 2397 54355 2400
rect 54297 2391 54355 2397
rect 56410 2388 56416 2400
rect 56468 2388 56474 2440
rect 62776 2437 62804 2468
rect 64693 2465 64705 2468
rect 64739 2496 64751 2499
rect 64782 2496 64788 2508
rect 64739 2468 64788 2496
rect 64739 2465 64751 2468
rect 64693 2459 64751 2465
rect 64782 2456 64788 2468
rect 64840 2456 64846 2508
rect 64877 2499 64935 2505
rect 64877 2465 64889 2499
rect 64923 2496 64935 2499
rect 66809 2499 66867 2505
rect 66809 2496 66821 2499
rect 64923 2468 66821 2496
rect 64923 2465 64935 2468
rect 64877 2459 64935 2465
rect 66809 2465 66821 2468
rect 66855 2496 66867 2499
rect 66990 2496 66996 2508
rect 66855 2468 66996 2496
rect 66855 2465 66867 2468
rect 66809 2459 66867 2465
rect 66990 2456 66996 2468
rect 67048 2456 67054 2508
rect 68925 2499 68983 2505
rect 68925 2465 68937 2499
rect 68971 2465 68983 2499
rect 68925 2459 68983 2465
rect 69109 2499 69167 2505
rect 69109 2465 69121 2499
rect 69155 2496 69167 2499
rect 71041 2499 71099 2505
rect 71041 2496 71053 2499
rect 69155 2468 71053 2496
rect 69155 2465 69167 2468
rect 69109 2459 69167 2465
rect 71041 2465 71053 2468
rect 71087 2496 71099 2499
rect 71222 2496 71228 2508
rect 71087 2468 71228 2496
rect 71087 2465 71099 2468
rect 71041 2459 71099 2465
rect 62761 2431 62819 2437
rect 62761 2397 62773 2431
rect 62807 2397 62819 2431
rect 62761 2391 62819 2397
rect 52178 2360 52184 2372
rect 50111 2332 52184 2360
rect 50111 2329 50123 2332
rect 50065 2323 50123 2329
rect 52178 2320 52184 2332
rect 52236 2320 52242 2372
rect 66993 2363 67051 2369
rect 66993 2329 67005 2363
rect 67039 2360 67051 2363
rect 68940 2360 68968 2459
rect 71222 2456 71228 2468
rect 71280 2456 71286 2508
rect 75273 2499 75331 2505
rect 75273 2465 75285 2499
rect 75319 2465 75331 2499
rect 75273 2459 75331 2465
rect 77389 2499 77447 2505
rect 77389 2465 77401 2499
rect 77435 2465 77447 2499
rect 77389 2459 77447 2465
rect 79689 2499 79747 2505
rect 79689 2465 79701 2499
rect 79735 2496 79747 2499
rect 81621 2499 81679 2505
rect 81621 2496 81633 2499
rect 79735 2468 81633 2496
rect 79735 2465 79747 2468
rect 79689 2459 79747 2465
rect 81621 2465 81633 2468
rect 81667 2496 81679 2499
rect 81710 2496 81716 2508
rect 81667 2468 81716 2496
rect 81667 2465 81679 2468
rect 81621 2459 81679 2465
rect 73341 2431 73399 2437
rect 73341 2397 73353 2431
rect 73387 2428 73399 2431
rect 75288 2428 75316 2459
rect 75454 2428 75460 2440
rect 73387 2400 75460 2428
rect 73387 2397 73399 2400
rect 73341 2391 73399 2397
rect 75454 2388 75460 2400
rect 75512 2388 75518 2440
rect 69106 2360 69112 2372
rect 67039 2332 69112 2360
rect 67039 2329 67051 2332
rect 66993 2323 67051 2329
rect 69106 2320 69112 2332
rect 69164 2320 69170 2372
rect 3467 2264 4936 2292
rect 75365 2295 75423 2301
rect 3467 2261 3479 2264
rect 3421 2255 3479 2261
rect 75365 2261 75377 2295
rect 75411 2292 75423 2295
rect 77404 2292 77432 2459
rect 81710 2456 81716 2468
rect 81768 2456 81774 2508
rect 81805 2499 81863 2505
rect 81805 2465 81817 2499
rect 81851 2496 81863 2499
rect 83737 2499 83795 2505
rect 83737 2496 83749 2499
rect 81851 2468 83749 2496
rect 81851 2465 81863 2468
rect 81805 2459 81863 2465
rect 83737 2465 83749 2468
rect 83783 2496 83795 2499
rect 83918 2496 83924 2508
rect 83783 2468 83924 2496
rect 83783 2465 83795 2468
rect 83737 2459 83795 2465
rect 83918 2456 83924 2468
rect 83976 2456 83982 2508
rect 85853 2499 85911 2505
rect 85853 2465 85865 2499
rect 85899 2465 85911 2499
rect 85853 2459 85911 2465
rect 87969 2499 88027 2505
rect 87969 2465 87981 2499
rect 88015 2465 88027 2499
rect 87969 2459 88027 2465
rect 92201 2499 92259 2505
rect 92201 2465 92213 2499
rect 92247 2465 92259 2499
rect 100665 2499 100723 2505
rect 100665 2496 100677 2499
rect 92201 2459 92259 2465
rect 98748 2468 100677 2496
rect 83921 2363 83979 2369
rect 83921 2329 83933 2363
rect 83967 2360 83979 2363
rect 85868 2360 85896 2459
rect 86037 2431 86095 2437
rect 86037 2397 86049 2431
rect 86083 2428 86095 2431
rect 87984 2428 88012 2459
rect 88150 2428 88156 2440
rect 86083 2400 88156 2428
rect 86083 2397 86095 2400
rect 86037 2391 86095 2397
rect 88150 2388 88156 2400
rect 88208 2388 88214 2440
rect 90269 2431 90327 2437
rect 90269 2397 90281 2431
rect 90315 2428 90327 2431
rect 92216 2428 92244 2459
rect 92382 2428 92388 2440
rect 90315 2400 92388 2428
rect 90315 2397 90327 2400
rect 90269 2391 90327 2397
rect 92382 2388 92388 2400
rect 92440 2388 92446 2440
rect 98748 2437 98776 2468
rect 100665 2465 100677 2468
rect 100711 2496 100723 2499
rect 100846 2496 100852 2508
rect 100711 2468 100852 2496
rect 100711 2465 100723 2468
rect 100665 2459 100723 2465
rect 100846 2456 100852 2468
rect 100904 2456 100910 2508
rect 98733 2431 98791 2437
rect 98733 2397 98745 2431
rect 98779 2397 98791 2431
rect 98733 2391 98791 2397
rect 85942 2360 85948 2372
rect 83967 2332 85948 2360
rect 83967 2329 83979 2332
rect 83921 2323 83979 2329
rect 85942 2320 85948 2332
rect 86000 2320 86006 2372
rect 100849 2363 100907 2369
rect 100849 2329 100861 2363
rect 100895 2360 100907 2363
rect 102597 2363 102655 2369
rect 102597 2360 102609 2363
rect 100895 2332 102609 2360
rect 100895 2329 100907 2332
rect 100849 2323 100907 2329
rect 102597 2329 102609 2332
rect 102643 2360 102655 2363
rect 102962 2360 102968 2372
rect 102643 2332 102968 2360
rect 102643 2329 102655 2332
rect 102597 2323 102655 2329
rect 102962 2320 102968 2332
rect 103020 2320 103026 2372
rect 77570 2292 77576 2304
rect 75411 2264 77576 2292
rect 75411 2261 75423 2264
rect 75365 2255 75423 2261
rect 77570 2252 77576 2264
rect 77628 2252 77634 2304
rect 1104 2202 106904 2224
rect 1104 2150 4042 2202
rect 4094 2150 4106 2202
rect 4158 2150 4170 2202
rect 4222 2150 4234 2202
rect 4286 2150 34762 2202
rect 34814 2150 34826 2202
rect 34878 2150 34890 2202
rect 34942 2150 34954 2202
rect 35006 2150 65482 2202
rect 65534 2150 65546 2202
rect 65598 2150 65610 2202
rect 65662 2150 65674 2202
rect 65726 2150 96202 2202
rect 96254 2150 96266 2202
rect 96318 2150 96330 2202
rect 96382 2150 96394 2202
rect 96446 2150 106904 2202
rect 1104 2128 106904 2150
rect 22646 2048 22652 2100
rect 22704 2088 22710 2100
rect 23658 2088 23664 2100
rect 22704 2060 23664 2088
rect 22704 2048 22710 2060
rect 23658 2048 23664 2060
rect 23716 2048 23722 2100
rect 24762 2048 24768 2100
rect 24820 2088 24826 2100
rect 25774 2088 25780 2100
rect 24820 2060 25780 2088
rect 24820 2048 24826 2060
rect 25774 2048 25780 2060
rect 25832 2048 25838 2100
rect 58618 2048 58624 2100
rect 58676 2088 58682 2100
rect 59630 2088 59636 2100
rect 58676 2060 59636 2088
rect 58676 2048 58682 2060
rect 59630 2048 59636 2060
rect 59688 2048 59694 2100
rect 77662 2048 77668 2100
rect 77720 2088 77726 2100
rect 78766 2088 78772 2100
rect 77720 2060 78772 2088
rect 77720 2048 77726 2060
rect 78766 2048 78772 2060
rect 78824 2048 78830 2100
rect 80330 2048 80336 2100
rect 80388 2088 80394 2100
rect 81158 2088 81164 2100
rect 80388 2060 81164 2088
rect 80388 2048 80394 2060
rect 81158 2048 81164 2060
rect 81216 2048 81222 2100
rect 96706 2048 96712 2100
rect 96764 2088 96770 2100
rect 97902 2088 97908 2100
rect 96764 2060 97908 2088
rect 96764 2048 96770 2060
rect 97902 2048 97908 2060
rect 97960 2048 97966 2100
rect 80606 1980 80612 2032
rect 80664 2020 80670 2032
rect 81342 2020 81348 2032
rect 80664 1992 81348 2020
rect 80664 1980 80670 1992
rect 81342 1980 81348 1992
rect 81400 1980 81406 2032
rect 1118 1952 1124 1964
rect 1079 1924 1124 1952
rect 1118 1912 1124 1924
rect 1176 1912 1182 1964
rect 3234 1952 3240 1964
rect 3195 1924 3240 1952
rect 3234 1912 3240 1924
rect 3292 1912 3298 1964
rect 3510 1952 3516 1964
rect 3471 1924 3516 1952
rect 3510 1912 3516 1924
rect 3568 1912 3574 1964
rect 3602 1912 3608 1964
rect 3660 1952 3666 1964
rect 4614 1952 4620 1964
rect 3660 1924 4620 1952
rect 3660 1912 3666 1924
rect 4614 1912 4620 1924
rect 4672 1912 4678 1964
rect 5350 1952 5356 1964
rect 5311 1924 5356 1952
rect 5350 1912 5356 1924
rect 5408 1912 5414 1964
rect 5626 1952 5632 1964
rect 5587 1924 5632 1952
rect 5626 1912 5632 1924
rect 5684 1912 5690 1964
rect 7466 1952 7472 1964
rect 7427 1924 7472 1952
rect 7466 1912 7472 1924
rect 7524 1912 7530 1964
rect 7742 1952 7748 1964
rect 7703 1924 7748 1952
rect 7742 1912 7748 1924
rect 7800 1912 7806 1964
rect 7834 1912 7840 1964
rect 7892 1952 7898 1964
rect 8846 1952 8852 1964
rect 7892 1924 8852 1952
rect 7892 1912 7898 1924
rect 8846 1912 8852 1924
rect 8904 1912 8910 1964
rect 9582 1952 9588 1964
rect 9543 1924 9588 1952
rect 9582 1912 9588 1924
rect 9640 1912 9646 1964
rect 9858 1952 9864 1964
rect 9819 1924 9864 1952
rect 9858 1912 9864 1924
rect 9916 1912 9922 1964
rect 9950 1912 9956 1964
rect 10008 1952 10014 1964
rect 11146 1952 11152 1964
rect 10008 1924 11152 1952
rect 10008 1912 10014 1924
rect 11146 1912 11152 1924
rect 11204 1912 11210 1964
rect 11698 1952 11704 1964
rect 11659 1924 11704 1952
rect 11698 1912 11704 1924
rect 11756 1912 11762 1964
rect 11882 1912 11888 1964
rect 11940 1952 11946 1964
rect 11977 1955 12035 1961
rect 11977 1952 11989 1955
rect 11940 1924 11989 1952
rect 11940 1912 11946 1924
rect 11977 1921 11989 1924
rect 12023 1921 12035 1955
rect 11977 1915 12035 1921
rect 12066 1912 12072 1964
rect 12124 1952 12130 1964
rect 13262 1952 13268 1964
rect 12124 1924 13268 1952
rect 12124 1912 12130 1924
rect 13262 1912 13268 1924
rect 13320 1912 13326 1964
rect 13814 1952 13820 1964
rect 13775 1924 13820 1952
rect 13814 1912 13820 1924
rect 13872 1912 13878 1964
rect 14090 1952 14096 1964
rect 14051 1924 14096 1952
rect 14090 1912 14096 1924
rect 14148 1912 14154 1964
rect 15930 1952 15936 1964
rect 15891 1924 15936 1952
rect 15930 1912 15936 1924
rect 15988 1912 15994 1964
rect 16206 1952 16212 1964
rect 16167 1924 16212 1952
rect 16206 1912 16212 1924
rect 16264 1912 16270 1964
rect 18046 1952 18052 1964
rect 18007 1924 18052 1952
rect 18046 1912 18052 1924
rect 18104 1912 18110 1964
rect 18322 1952 18328 1964
rect 18283 1924 18328 1952
rect 18322 1912 18328 1924
rect 18380 1912 18386 1964
rect 20162 1952 20168 1964
rect 20123 1924 20168 1952
rect 20162 1912 20168 1924
rect 20220 1912 20226 1964
rect 20438 1952 20444 1964
rect 20399 1924 20444 1952
rect 20438 1912 20444 1924
rect 20496 1912 20502 1964
rect 22186 1912 22192 1964
rect 22244 1952 22250 1964
rect 22281 1955 22339 1961
rect 22281 1952 22293 1955
rect 22244 1924 22293 1952
rect 22244 1912 22250 1924
rect 22281 1921 22293 1924
rect 22327 1921 22339 1955
rect 24394 1952 24400 1964
rect 24355 1924 24400 1952
rect 22281 1915 22339 1921
rect 24394 1912 24400 1924
rect 24452 1912 24458 1964
rect 24670 1952 24676 1964
rect 24631 1924 24676 1952
rect 24670 1912 24676 1924
rect 24728 1912 24734 1964
rect 26510 1952 26516 1964
rect 26471 1924 26516 1952
rect 26510 1912 26516 1924
rect 26568 1912 26574 1964
rect 26694 1912 26700 1964
rect 26752 1952 26758 1964
rect 26789 1955 26847 1961
rect 26789 1952 26801 1955
rect 26752 1924 26801 1952
rect 26752 1912 26758 1924
rect 26789 1921 26801 1924
rect 26835 1921 26847 1955
rect 28626 1952 28632 1964
rect 28587 1924 28632 1952
rect 26789 1915 26847 1921
rect 28626 1912 28632 1924
rect 28684 1912 28690 1964
rect 28810 1912 28816 1964
rect 28868 1952 28874 1964
rect 28905 1955 28963 1961
rect 28905 1952 28917 1955
rect 28868 1924 28917 1952
rect 28868 1912 28874 1924
rect 28905 1921 28917 1924
rect 28951 1921 28963 1955
rect 28905 1915 28963 1921
rect 28994 1912 29000 1964
rect 29052 1952 29058 1964
rect 30190 1952 30196 1964
rect 29052 1924 30196 1952
rect 29052 1912 29058 1924
rect 30190 1912 30196 1924
rect 30248 1912 30254 1964
rect 30742 1952 30748 1964
rect 30703 1924 30748 1952
rect 30742 1912 30748 1924
rect 30800 1912 30806 1964
rect 31018 1952 31024 1964
rect 30979 1924 31024 1952
rect 31018 1912 31024 1924
rect 31076 1912 31082 1964
rect 32858 1952 32864 1964
rect 32819 1924 32864 1952
rect 32858 1912 32864 1924
rect 32916 1912 32922 1964
rect 33134 1952 33140 1964
rect 33095 1924 33140 1952
rect 33134 1912 33140 1924
rect 33192 1912 33198 1964
rect 35250 1952 35256 1964
rect 35211 1924 35256 1952
rect 35250 1912 35256 1924
rect 35308 1912 35314 1964
rect 37090 1952 37096 1964
rect 37051 1924 37096 1952
rect 37090 1912 37096 1924
rect 37148 1912 37154 1964
rect 37366 1952 37372 1964
rect 37327 1924 37372 1952
rect 37366 1912 37372 1924
rect 37424 1912 37430 1964
rect 39206 1952 39212 1964
rect 39167 1924 39212 1952
rect 39206 1912 39212 1924
rect 39264 1912 39270 1964
rect 39390 1912 39396 1964
rect 39448 1952 39454 1964
rect 39485 1955 39543 1961
rect 39485 1952 39497 1955
rect 39448 1924 39497 1952
rect 39448 1912 39454 1924
rect 39485 1921 39497 1924
rect 39531 1921 39543 1955
rect 39485 1915 39543 1921
rect 39574 1912 39580 1964
rect 39632 1952 39638 1964
rect 40678 1952 40684 1964
rect 39632 1924 40684 1952
rect 39632 1912 39638 1924
rect 40678 1912 40684 1924
rect 40736 1912 40742 1964
rect 41322 1952 41328 1964
rect 41283 1924 41328 1952
rect 41322 1912 41328 1924
rect 41380 1912 41386 1964
rect 41598 1952 41604 1964
rect 41559 1924 41604 1952
rect 41598 1912 41604 1924
rect 41656 1912 41662 1964
rect 41690 1912 41696 1964
rect 41748 1952 41754 1964
rect 42702 1952 42708 1964
rect 41748 1924 42708 1952
rect 41748 1912 41754 1924
rect 42702 1912 42708 1924
rect 42760 1912 42766 1964
rect 43438 1952 43444 1964
rect 43399 1924 43444 1952
rect 43438 1912 43444 1924
rect 43496 1912 43502 1964
rect 43714 1952 43720 1964
rect 43675 1924 43720 1952
rect 43714 1912 43720 1924
rect 43772 1912 43778 1964
rect 43806 1912 43812 1964
rect 43864 1952 43870 1964
rect 45002 1952 45008 1964
rect 43864 1924 45008 1952
rect 43864 1912 43870 1924
rect 45002 1912 45008 1924
rect 45060 1912 45066 1964
rect 45554 1952 45560 1964
rect 45515 1924 45560 1952
rect 45554 1912 45560 1924
rect 45612 1912 45618 1964
rect 45830 1952 45836 1964
rect 45791 1924 45836 1952
rect 45830 1912 45836 1924
rect 45888 1912 45894 1964
rect 45922 1912 45928 1964
rect 45980 1952 45986 1964
rect 47118 1952 47124 1964
rect 45980 1924 47124 1952
rect 45980 1912 45986 1924
rect 47118 1912 47124 1924
rect 47176 1912 47182 1964
rect 47670 1952 47676 1964
rect 47631 1924 47676 1952
rect 47670 1912 47676 1924
rect 47728 1912 47734 1964
rect 47854 1912 47860 1964
rect 47912 1952 47918 1964
rect 47949 1955 48007 1961
rect 47949 1952 47961 1955
rect 47912 1924 47961 1952
rect 47912 1912 47918 1924
rect 47949 1921 47961 1924
rect 47995 1921 48007 1955
rect 49786 1952 49792 1964
rect 49747 1924 49792 1952
rect 47949 1915 48007 1921
rect 49786 1912 49792 1924
rect 49844 1912 49850 1964
rect 50062 1912 50068 1964
rect 50120 1952 50126 1964
rect 51902 1952 51908 1964
rect 50120 1924 50165 1952
rect 51863 1924 51908 1952
rect 50120 1912 50126 1924
rect 51902 1912 51908 1924
rect 51960 1912 51966 1964
rect 52178 1952 52184 1964
rect 52139 1924 52184 1952
rect 52178 1912 52184 1924
rect 52236 1912 52242 1964
rect 54018 1952 54024 1964
rect 53979 1924 54024 1952
rect 54018 1912 54024 1924
rect 54076 1912 54082 1964
rect 54202 1912 54208 1964
rect 54260 1952 54266 1964
rect 54297 1955 54355 1961
rect 54297 1952 54309 1955
rect 54260 1924 54309 1952
rect 54260 1912 54266 1924
rect 54297 1921 54309 1924
rect 54343 1921 54355 1955
rect 54297 1915 54355 1921
rect 54386 1912 54392 1964
rect 54444 1952 54450 1964
rect 55398 1952 55404 1964
rect 54444 1924 55404 1952
rect 54444 1912 54450 1924
rect 55398 1912 55404 1924
rect 55456 1912 55462 1964
rect 56134 1952 56140 1964
rect 56095 1924 56140 1952
rect 56134 1912 56140 1924
rect 56192 1912 56198 1964
rect 56410 1952 56416 1964
rect 56371 1924 56416 1952
rect 56410 1912 56416 1924
rect 56468 1912 56474 1964
rect 58250 1952 58256 1964
rect 58211 1924 58256 1952
rect 58250 1912 58256 1924
rect 58308 1912 58314 1964
rect 58434 1912 58440 1964
rect 58492 1952 58498 1964
rect 58529 1955 58587 1961
rect 58529 1952 58541 1955
rect 58492 1924 58541 1952
rect 58492 1912 58498 1924
rect 58529 1921 58541 1924
rect 58575 1921 58587 1955
rect 58529 1915 58587 1921
rect 60366 1912 60372 1964
rect 60424 1952 60430 1964
rect 62482 1952 62488 1964
rect 60424 1924 60469 1952
rect 62443 1924 62488 1952
rect 60424 1912 60430 1924
rect 62482 1912 62488 1924
rect 62540 1912 62546 1964
rect 62758 1952 62764 1964
rect 62719 1924 62764 1952
rect 62758 1912 62764 1924
rect 62816 1912 62822 1964
rect 62850 1912 62856 1964
rect 62908 1952 62914 1964
rect 64046 1952 64052 1964
rect 62908 1924 64052 1952
rect 62908 1912 62914 1924
rect 64046 1912 64052 1924
rect 64104 1912 64110 1964
rect 64598 1952 64604 1964
rect 64559 1924 64604 1952
rect 64598 1912 64604 1924
rect 64656 1912 64662 1964
rect 64782 1912 64788 1964
rect 64840 1952 64846 1964
rect 64877 1955 64935 1961
rect 64877 1952 64889 1955
rect 64840 1924 64889 1952
rect 64840 1912 64846 1924
rect 64877 1921 64889 1924
rect 64923 1921 64935 1955
rect 66714 1952 66720 1964
rect 66675 1924 66720 1952
rect 64877 1915 64935 1921
rect 66714 1912 66720 1924
rect 66772 1912 66778 1964
rect 66990 1952 66996 1964
rect 66951 1924 66996 1952
rect 66990 1912 66996 1924
rect 67048 1912 67054 1964
rect 68830 1952 68836 1964
rect 68791 1924 68836 1952
rect 68830 1912 68836 1924
rect 68888 1912 68894 1964
rect 69106 1952 69112 1964
rect 69067 1924 69112 1952
rect 69106 1912 69112 1924
rect 69164 1912 69170 1964
rect 70946 1952 70952 1964
rect 70907 1924 70952 1952
rect 70946 1912 70952 1924
rect 71004 1912 71010 1964
rect 71222 1952 71228 1964
rect 71183 1924 71228 1952
rect 71222 1912 71228 1924
rect 71280 1912 71286 1964
rect 73062 1952 73068 1964
rect 73023 1924 73068 1952
rect 73062 1912 73068 1924
rect 73120 1912 73126 1964
rect 73338 1952 73344 1964
rect 73299 1924 73344 1952
rect 73338 1912 73344 1924
rect 73396 1912 73402 1964
rect 75178 1952 75184 1964
rect 75139 1924 75184 1952
rect 75178 1912 75184 1924
rect 75236 1912 75242 1964
rect 75454 1952 75460 1964
rect 75415 1924 75460 1952
rect 75454 1912 75460 1924
rect 75512 1912 75518 1964
rect 75546 1912 75552 1964
rect 75604 1952 75610 1964
rect 76742 1952 76748 1964
rect 75604 1924 76748 1952
rect 75604 1912 75610 1924
rect 76742 1912 76748 1924
rect 76800 1912 76806 1964
rect 77570 1952 77576 1964
rect 77531 1924 77576 1952
rect 77570 1912 77576 1924
rect 77628 1912 77634 1964
rect 78214 1912 78220 1964
rect 78272 1952 78278 1964
rect 78858 1952 78864 1964
rect 78272 1924 78864 1952
rect 78272 1912 78278 1924
rect 78858 1912 78864 1924
rect 78916 1912 78922 1964
rect 79410 1952 79416 1964
rect 79371 1924 79416 1952
rect 79410 1912 79416 1924
rect 79468 1912 79474 1964
rect 79594 1912 79600 1964
rect 79652 1952 79658 1964
rect 79689 1955 79747 1961
rect 79689 1952 79701 1955
rect 79652 1924 79701 1952
rect 79652 1912 79658 1924
rect 79689 1921 79701 1924
rect 79735 1921 79747 1955
rect 79689 1915 79747 1921
rect 79778 1912 79784 1964
rect 79836 1952 79842 1964
rect 81250 1952 81256 1964
rect 79836 1924 81256 1952
rect 79836 1912 79842 1924
rect 81250 1912 81256 1924
rect 81308 1912 81314 1964
rect 81526 1952 81532 1964
rect 81487 1924 81532 1952
rect 81526 1912 81532 1924
rect 81584 1912 81590 1964
rect 81710 1912 81716 1964
rect 81768 1952 81774 1964
rect 81805 1955 81863 1961
rect 81805 1952 81817 1955
rect 81768 1924 81817 1952
rect 81768 1912 81774 1924
rect 81805 1921 81817 1924
rect 81851 1921 81863 1955
rect 83642 1952 83648 1964
rect 83603 1924 83648 1952
rect 81805 1915 81863 1921
rect 83642 1912 83648 1924
rect 83700 1912 83706 1964
rect 83918 1952 83924 1964
rect 83879 1924 83924 1952
rect 83918 1912 83924 1924
rect 83976 1912 83982 1964
rect 85758 1952 85764 1964
rect 85719 1924 85764 1952
rect 85758 1912 85764 1924
rect 85816 1912 85822 1964
rect 85942 1912 85948 1964
rect 86000 1952 86006 1964
rect 86037 1955 86095 1961
rect 86037 1952 86049 1955
rect 86000 1924 86049 1952
rect 86000 1912 86006 1924
rect 86037 1921 86049 1924
rect 86083 1921 86095 1955
rect 87874 1952 87880 1964
rect 87835 1924 87880 1952
rect 86037 1915 86095 1921
rect 87874 1912 87880 1924
rect 87932 1912 87938 1964
rect 88150 1952 88156 1964
rect 88111 1924 88156 1952
rect 88150 1912 88156 1924
rect 88208 1912 88214 1964
rect 88794 1912 88800 1964
rect 88852 1952 88858 1964
rect 89254 1952 89260 1964
rect 88852 1924 89260 1952
rect 88852 1912 88858 1924
rect 89254 1912 89260 1924
rect 89312 1912 89318 1964
rect 89990 1952 89996 1964
rect 89951 1924 89996 1952
rect 89990 1912 89996 1924
rect 90048 1912 90054 1964
rect 90266 1952 90272 1964
rect 90227 1924 90272 1952
rect 90266 1912 90272 1924
rect 90324 1912 90330 1964
rect 90358 1912 90364 1964
rect 90416 1952 90422 1964
rect 91370 1952 91376 1964
rect 90416 1924 91376 1952
rect 90416 1912 90422 1924
rect 91370 1912 91376 1924
rect 91428 1912 91434 1964
rect 92106 1952 92112 1964
rect 92067 1924 92112 1952
rect 92106 1912 92112 1924
rect 92164 1912 92170 1964
rect 92382 1952 92388 1964
rect 92343 1924 92388 1952
rect 92382 1912 92388 1924
rect 92440 1912 92446 1964
rect 92474 1912 92480 1964
rect 92532 1952 92538 1964
rect 93486 1952 93492 1964
rect 92532 1924 93492 1952
rect 92532 1912 92538 1924
rect 93486 1912 93492 1924
rect 93544 1912 93550 1964
rect 94222 1952 94228 1964
rect 94183 1924 94228 1952
rect 94222 1912 94228 1924
rect 94280 1912 94286 1964
rect 94406 1912 94412 1964
rect 94464 1952 94470 1964
rect 94501 1955 94559 1961
rect 94501 1952 94513 1955
rect 94464 1924 94513 1952
rect 94464 1912 94470 1924
rect 94501 1921 94513 1924
rect 94547 1921 94559 1955
rect 94501 1915 94559 1921
rect 95142 1912 95148 1964
rect 95200 1952 95206 1964
rect 95786 1952 95792 1964
rect 95200 1924 95792 1952
rect 95200 1912 95206 1924
rect 95786 1912 95792 1924
rect 95844 1912 95850 1964
rect 96062 1912 96068 1964
rect 96120 1952 96126 1964
rect 96341 1955 96399 1961
rect 96341 1952 96353 1955
rect 96120 1924 96353 1952
rect 96120 1912 96126 1924
rect 96341 1921 96353 1924
rect 96387 1921 96399 1955
rect 96614 1952 96620 1964
rect 96575 1924 96620 1952
rect 96341 1915 96399 1921
rect 96614 1912 96620 1924
rect 96672 1912 96678 1964
rect 97258 1912 97264 1964
rect 97316 1952 97322 1964
rect 97994 1952 98000 1964
rect 97316 1924 98000 1952
rect 97316 1912 97322 1924
rect 97994 1912 98000 1924
rect 98052 1912 98058 1964
rect 98454 1952 98460 1964
rect 98415 1924 98460 1952
rect 98454 1912 98460 1924
rect 98512 1912 98518 1964
rect 98730 1952 98736 1964
rect 98691 1924 98736 1952
rect 98730 1912 98736 1924
rect 98788 1912 98794 1964
rect 100570 1952 100576 1964
rect 100531 1924 100576 1952
rect 100570 1912 100576 1924
rect 100628 1912 100634 1964
rect 100846 1952 100852 1964
rect 100807 1924 100852 1952
rect 100846 1912 100852 1924
rect 100904 1912 100910 1964
rect 102686 1952 102692 1964
rect 102647 1924 102692 1952
rect 102686 1912 102692 1924
rect 102744 1912 102750 1964
rect 102962 1952 102968 1964
rect 102923 1924 102968 1952
rect 102962 1912 102968 1924
rect 103020 1912 103026 1964
rect 104802 1952 104808 1964
rect 104763 1924 104808 1952
rect 104802 1912 104808 1924
rect 104860 1912 104866 1964
rect 1210 1844 1216 1896
rect 1268 1884 1274 1896
rect 1397 1887 1455 1893
rect 1397 1884 1409 1887
rect 1268 1856 1409 1884
rect 1268 1844 1274 1856
rect 1397 1853 1409 1856
rect 1443 1853 1455 1887
rect 1397 1847 1455 1853
rect 5718 1844 5724 1896
rect 5776 1884 5782 1896
rect 6730 1884 6736 1896
rect 5776 1856 6736 1884
rect 5776 1844 5782 1856
rect 6730 1844 6736 1856
rect 6788 1844 6794 1896
rect 10778 1844 10784 1896
rect 10836 1884 10842 1896
rect 11238 1884 11244 1896
rect 10836 1856 11244 1884
rect 10836 1844 10842 1856
rect 11238 1844 11244 1856
rect 11296 1844 11302 1896
rect 18414 1844 18420 1896
rect 18472 1884 18478 1896
rect 18690 1884 18696 1896
rect 18472 1856 18696 1884
rect 18472 1844 18478 1856
rect 18690 1844 18696 1856
rect 18748 1844 18754 1896
rect 20530 1844 20536 1896
rect 20588 1884 20594 1896
rect 21542 1884 21548 1896
rect 20588 1856 21548 1884
rect 20588 1844 20594 1856
rect 21542 1844 21548 1856
rect 21600 1844 21606 1896
rect 22370 1844 22376 1896
rect 22428 1884 22434 1896
rect 22557 1887 22615 1893
rect 22557 1884 22569 1887
rect 22428 1856 22569 1884
rect 22428 1844 22434 1856
rect 22557 1853 22569 1856
rect 22603 1853 22615 1887
rect 22557 1847 22615 1853
rect 26878 1844 26884 1896
rect 26936 1884 26942 1896
rect 28074 1884 28080 1896
rect 26936 1856 28080 1884
rect 26936 1844 26942 1856
rect 28074 1844 28080 1856
rect 28132 1844 28138 1896
rect 34977 1887 35035 1893
rect 34977 1853 34989 1887
rect 35023 1884 35035 1887
rect 35066 1884 35072 1896
rect 35023 1856 35072 1884
rect 35023 1853 35035 1856
rect 34977 1847 35035 1853
rect 35066 1844 35072 1856
rect 35124 1844 35130 1896
rect 37458 1844 37464 1896
rect 37516 1884 37522 1896
rect 38470 1884 38476 1896
rect 37516 1856 38476 1884
rect 37516 1844 37522 1856
rect 38470 1844 38476 1856
rect 38528 1844 38534 1896
rect 56502 1844 56508 1896
rect 56560 1884 56566 1896
rect 57514 1884 57520 1896
rect 56560 1856 57520 1884
rect 56560 1844 56566 1856
rect 57514 1844 57520 1856
rect 57572 1844 57578 1896
rect 60458 1844 60464 1896
rect 60516 1884 60522 1896
rect 60645 1887 60703 1893
rect 60645 1884 60657 1887
rect 60516 1856 60657 1884
rect 60516 1844 60522 1856
rect 60645 1853 60657 1856
rect 60691 1853 60703 1887
rect 60645 1847 60703 1853
rect 60734 1844 60740 1896
rect 60792 1884 60798 1896
rect 61930 1884 61936 1896
rect 60792 1856 61936 1884
rect 60792 1844 60798 1856
rect 61930 1844 61936 1856
rect 61988 1844 61994 1896
rect 71314 1844 71320 1896
rect 71372 1884 71378 1896
rect 72326 1884 72332 1896
rect 71372 1856 72332 1884
rect 71372 1844 71378 1856
rect 72326 1844 72332 1856
rect 72384 1844 72390 1896
rect 73430 1844 73436 1896
rect 73488 1884 73494 1896
rect 74442 1884 74448 1896
rect 73488 1856 74448 1884
rect 73488 1844 73494 1856
rect 74442 1844 74448 1856
rect 74500 1844 74506 1896
rect 77294 1844 77300 1896
rect 77352 1884 77358 1896
rect 77352 1856 77397 1884
rect 77352 1844 77358 1856
rect 78490 1844 78496 1896
rect 78548 1884 78554 1896
rect 78950 1884 78956 1896
rect 78548 1856 78956 1884
rect 78548 1844 78554 1856
rect 78950 1844 78956 1856
rect 79008 1844 79014 1896
rect 88242 1844 88248 1896
rect 88300 1884 88306 1896
rect 89438 1884 89444 1896
rect 88300 1856 89444 1884
rect 88300 1844 88306 1856
rect 89438 1844 89444 1856
rect 89496 1844 89502 1896
rect 93026 1844 93032 1896
rect 93084 1884 93090 1896
rect 93670 1884 93676 1896
rect 93084 1856 93676 1884
rect 93084 1844 93090 1856
rect 93670 1844 93676 1856
rect 93728 1844 93734 1896
rect 94590 1844 94596 1896
rect 94648 1884 94654 1896
rect 95694 1884 95700 1896
rect 94648 1856 95700 1884
rect 94648 1844 94654 1856
rect 95694 1844 95700 1856
rect 95752 1844 95758 1896
rect 97534 1844 97540 1896
rect 97592 1884 97598 1896
rect 98086 1884 98092 1896
rect 97592 1856 98092 1884
rect 97592 1844 97598 1856
rect 98086 1844 98092 1856
rect 98144 1844 98150 1896
rect 104894 1844 104900 1896
rect 104952 1884 104958 1896
rect 105081 1887 105139 1893
rect 105081 1884 105093 1887
rect 104952 1856 105093 1884
rect 104952 1844 104958 1856
rect 105081 1853 105093 1856
rect 105127 1853 105139 1887
rect 105081 1847 105139 1853
rect 81069 1819 81127 1825
rect 81069 1785 81081 1819
rect 81115 1816 81127 1819
rect 81158 1816 81164 1828
rect 81115 1788 81164 1816
rect 81115 1785 81127 1788
rect 81069 1779 81127 1785
rect 81158 1776 81164 1788
rect 81216 1776 81222 1828
rect 95418 1776 95424 1828
rect 95476 1816 95482 1828
rect 95878 1816 95884 1828
rect 95476 1788 95884 1816
rect 95476 1776 95482 1788
rect 95878 1776 95884 1788
rect 95936 1776 95942 1828
rect 2498 1748 2504 1760
rect 2459 1720 2504 1748
rect 2498 1708 2504 1720
rect 2556 1708 2562 1760
rect 4154 1708 4160 1760
rect 4212 1748 4218 1760
rect 4617 1751 4675 1757
rect 4617 1748 4629 1751
rect 4212 1720 4629 1748
rect 4212 1708 4218 1720
rect 4617 1717 4629 1720
rect 4663 1717 4675 1751
rect 4617 1711 4675 1717
rect 5902 1708 5908 1760
rect 5960 1748 5966 1760
rect 6733 1751 6791 1757
rect 6733 1748 6745 1751
rect 5960 1720 6745 1748
rect 5960 1708 5966 1720
rect 6733 1717 6745 1720
rect 6779 1717 6791 1751
rect 6733 1711 6791 1717
rect 8202 1708 8208 1760
rect 8260 1748 8266 1760
rect 8849 1751 8907 1757
rect 8849 1748 8861 1751
rect 8260 1720 8861 1748
rect 8260 1708 8266 1720
rect 8849 1717 8861 1720
rect 8895 1717 8907 1751
rect 11146 1748 11152 1760
rect 11107 1720 11152 1748
rect 8849 1711 8907 1717
rect 11146 1708 11152 1720
rect 11204 1708 11210 1760
rect 13262 1748 13268 1760
rect 13223 1720 13268 1748
rect 13262 1708 13268 1720
rect 13320 1708 13326 1760
rect 15194 1748 15200 1760
rect 15155 1720 15200 1748
rect 15194 1708 15200 1720
rect 15252 1708 15258 1760
rect 17310 1748 17316 1760
rect 17271 1720 17316 1748
rect 17310 1708 17316 1720
rect 17368 1708 17374 1760
rect 18690 1708 18696 1760
rect 18748 1748 18754 1760
rect 19429 1751 19487 1757
rect 19429 1748 19441 1751
rect 18748 1720 19441 1748
rect 18748 1708 18754 1720
rect 19429 1717 19441 1720
rect 19475 1717 19487 1751
rect 19429 1711 19487 1717
rect 20714 1708 20720 1760
rect 20772 1748 20778 1760
rect 21545 1751 21603 1757
rect 21545 1748 21557 1751
rect 20772 1720 21557 1748
rect 20772 1708 20778 1720
rect 21545 1717 21557 1720
rect 21591 1717 21603 1751
rect 21545 1711 21603 1717
rect 22830 1708 22836 1760
rect 22888 1748 22894 1760
rect 23661 1751 23719 1757
rect 23661 1748 23673 1751
rect 22888 1720 23673 1748
rect 22888 1708 22894 1720
rect 23661 1717 23673 1720
rect 23707 1717 23719 1751
rect 23661 1711 23719 1717
rect 25038 1708 25044 1760
rect 25096 1748 25102 1760
rect 25777 1751 25835 1757
rect 25777 1748 25789 1751
rect 25096 1720 25789 1748
rect 25096 1708 25102 1720
rect 25777 1717 25789 1720
rect 25823 1717 25835 1751
rect 28074 1748 28080 1760
rect 28035 1720 28080 1748
rect 25777 1711 25835 1717
rect 28074 1708 28080 1720
rect 28132 1708 28138 1760
rect 30190 1748 30196 1760
rect 30151 1720 30196 1748
rect 30190 1708 30196 1720
rect 30248 1708 30254 1760
rect 32122 1748 32128 1760
rect 32083 1720 32128 1748
rect 32122 1708 32128 1720
rect 32180 1708 32186 1760
rect 34238 1748 34244 1760
rect 34199 1720 34244 1748
rect 34238 1708 34244 1720
rect 34296 1708 34302 1760
rect 35526 1708 35532 1760
rect 35584 1748 35590 1760
rect 36357 1751 36415 1757
rect 36357 1748 36369 1751
rect 35584 1720 36369 1748
rect 35584 1708 35590 1720
rect 36357 1717 36369 1720
rect 36403 1717 36415 1751
rect 36357 1711 36415 1717
rect 37642 1708 37648 1760
rect 37700 1748 37706 1760
rect 38473 1751 38531 1757
rect 38473 1748 38485 1751
rect 37700 1720 38485 1748
rect 37700 1708 37706 1720
rect 38473 1717 38485 1720
rect 38519 1717 38531 1751
rect 38473 1711 38531 1717
rect 40126 1708 40132 1760
rect 40184 1748 40190 1760
rect 40589 1751 40647 1757
rect 40589 1748 40601 1751
rect 40184 1720 40601 1748
rect 40184 1708 40190 1720
rect 40589 1717 40601 1720
rect 40635 1717 40647 1751
rect 40589 1711 40647 1717
rect 41966 1708 41972 1760
rect 42024 1748 42030 1760
rect 42705 1751 42763 1757
rect 42705 1748 42717 1751
rect 42024 1720 42717 1748
rect 42024 1708 42030 1720
rect 42705 1717 42717 1720
rect 42751 1717 42763 1751
rect 45002 1748 45008 1760
rect 44963 1720 45008 1748
rect 42705 1711 42763 1717
rect 45002 1708 45008 1720
rect 45060 1708 45066 1760
rect 47118 1748 47124 1760
rect 47079 1720 47124 1748
rect 47118 1708 47124 1720
rect 47176 1708 47182 1760
rect 49050 1748 49056 1760
rect 49011 1720 49056 1748
rect 49050 1708 49056 1720
rect 49108 1708 49114 1760
rect 51166 1748 51172 1760
rect 51127 1720 51172 1748
rect 51166 1708 51172 1720
rect 51224 1708 51230 1760
rect 52270 1708 52276 1760
rect 52328 1748 52334 1760
rect 53285 1751 53343 1757
rect 53285 1748 53297 1751
rect 52328 1720 53297 1748
rect 52328 1708 52334 1720
rect 53285 1717 53297 1720
rect 53331 1717 53343 1751
rect 53285 1711 53343 1717
rect 54754 1708 54760 1760
rect 54812 1748 54818 1760
rect 55401 1751 55459 1757
rect 55401 1748 55413 1751
rect 54812 1720 55413 1748
rect 54812 1708 54818 1720
rect 55401 1717 55413 1720
rect 55447 1717 55459 1751
rect 55401 1711 55459 1717
rect 56686 1708 56692 1760
rect 56744 1748 56750 1760
rect 57517 1751 57575 1757
rect 57517 1748 57529 1751
rect 56744 1720 57529 1748
rect 56744 1708 56750 1720
rect 57517 1717 57529 1720
rect 57563 1717 57575 1751
rect 57517 1711 57575 1717
rect 58894 1708 58900 1760
rect 58952 1748 58958 1760
rect 59633 1751 59691 1757
rect 59633 1748 59645 1751
rect 58952 1720 59645 1748
rect 58952 1708 58958 1720
rect 59633 1717 59645 1720
rect 59679 1717 59691 1751
rect 61930 1748 61936 1760
rect 61891 1720 61936 1748
rect 59633 1711 59691 1717
rect 61930 1708 61936 1720
rect 61988 1708 61994 1760
rect 64046 1748 64052 1760
rect 64007 1720 64052 1748
rect 64046 1708 64052 1720
rect 64104 1708 64110 1760
rect 65978 1748 65984 1760
rect 65939 1720 65984 1748
rect 65978 1708 65984 1720
rect 66036 1708 66042 1760
rect 68094 1748 68100 1760
rect 68055 1720 68100 1748
rect 68094 1708 68100 1720
rect 68152 1708 68158 1760
rect 69198 1708 69204 1760
rect 69256 1748 69262 1760
rect 70213 1751 70271 1757
rect 70213 1748 70225 1751
rect 69256 1720 70225 1748
rect 69256 1708 69262 1720
rect 70213 1717 70225 1720
rect 70259 1717 70271 1751
rect 70213 1711 70271 1717
rect 71498 1708 71504 1760
rect 71556 1748 71562 1760
rect 72329 1751 72387 1757
rect 72329 1748 72341 1751
rect 71556 1720 72341 1748
rect 71556 1708 71562 1720
rect 72329 1717 72341 1720
rect 72375 1717 72387 1751
rect 72329 1711 72387 1717
rect 73614 1708 73620 1760
rect 73672 1748 73678 1760
rect 74445 1751 74503 1757
rect 74445 1748 74457 1751
rect 73672 1720 74457 1748
rect 73672 1708 73678 1720
rect 74445 1717 74457 1720
rect 74491 1717 74503 1751
rect 74445 1711 74503 1717
rect 76190 1708 76196 1760
rect 76248 1748 76254 1760
rect 76561 1751 76619 1757
rect 76561 1748 76573 1751
rect 76248 1720 76573 1748
rect 76248 1708 76254 1720
rect 76561 1717 76573 1720
rect 76607 1717 76619 1751
rect 78858 1748 78864 1760
rect 78819 1720 78864 1748
rect 76561 1711 76619 1717
rect 78858 1708 78864 1720
rect 78916 1708 78922 1760
rect 82906 1748 82912 1760
rect 82867 1720 82912 1748
rect 82906 1708 82912 1720
rect 82964 1708 82970 1760
rect 85022 1748 85028 1760
rect 84983 1720 85028 1748
rect 85022 1708 85028 1720
rect 85080 1708 85086 1760
rect 86494 1708 86500 1760
rect 86552 1748 86558 1760
rect 87141 1751 87199 1757
rect 87141 1748 87153 1751
rect 86552 1720 87153 1748
rect 86552 1708 86558 1720
rect 87141 1717 87153 1720
rect 87187 1717 87199 1751
rect 87141 1711 87199 1717
rect 88426 1708 88432 1760
rect 88484 1748 88490 1760
rect 89257 1751 89315 1757
rect 89257 1748 89269 1751
rect 88484 1720 89269 1748
rect 88484 1708 88490 1720
rect 89257 1717 89269 1720
rect 89303 1717 89315 1751
rect 89257 1711 89315 1717
rect 90726 1708 90732 1760
rect 90784 1748 90790 1760
rect 91373 1751 91431 1757
rect 91373 1748 91385 1751
rect 90784 1720 91385 1748
rect 90784 1708 90790 1720
rect 91373 1717 91385 1720
rect 91419 1717 91431 1751
rect 91373 1711 91431 1717
rect 92750 1708 92756 1760
rect 92808 1748 92814 1760
rect 93489 1751 93547 1757
rect 93489 1748 93501 1751
rect 92808 1720 93501 1748
rect 92808 1708 92814 1720
rect 93489 1717 93501 1720
rect 93535 1717 93547 1751
rect 95786 1748 95792 1760
rect 95747 1720 95792 1748
rect 93489 1711 93547 1717
rect 95786 1708 95792 1720
rect 95844 1708 95850 1760
rect 97902 1748 97908 1760
rect 97863 1720 97908 1748
rect 97902 1708 97908 1720
rect 97960 1708 97966 1760
rect 99834 1748 99840 1760
rect 99795 1720 99840 1748
rect 99834 1708 99840 1720
rect 99892 1708 99898 1760
rect 101950 1748 101956 1760
rect 101911 1720 101956 1748
rect 101950 1708 101956 1720
rect 102008 1708 102014 1760
rect 103238 1708 103244 1760
rect 103296 1748 103302 1760
rect 104069 1751 104127 1757
rect 104069 1748 104081 1751
rect 103296 1720 104081 1748
rect 103296 1708 103302 1720
rect 104069 1717 104081 1720
rect 104115 1717 104127 1751
rect 104069 1711 104127 1717
rect 105354 1708 105360 1760
rect 105412 1748 105418 1760
rect 106185 1751 106243 1757
rect 106185 1748 106197 1751
rect 105412 1720 106197 1748
rect 105412 1708 105418 1720
rect 106185 1717 106197 1720
rect 106231 1717 106243 1751
rect 106185 1711 106243 1717
rect 1104 1658 106904 1680
rect 1104 1606 19402 1658
rect 19454 1606 19466 1658
rect 19518 1606 19530 1658
rect 19582 1606 19594 1658
rect 19646 1606 50122 1658
rect 50174 1606 50186 1658
rect 50238 1606 50250 1658
rect 50302 1606 50314 1658
rect 50366 1606 80842 1658
rect 80894 1606 80906 1658
rect 80958 1606 80970 1658
rect 81022 1606 81034 1658
rect 81086 1606 106904 1658
rect 1104 1584 106904 1606
rect 1026 1504 1032 1556
rect 1084 1544 1090 1556
rect 2501 1547 2559 1553
rect 2501 1544 2513 1547
rect 1084 1516 2513 1544
rect 1084 1504 1090 1516
rect 2501 1513 2513 1516
rect 2547 1513 2559 1547
rect 2501 1507 2559 1513
rect 7374 1504 7380 1556
rect 7432 1544 7438 1556
rect 8849 1547 8907 1553
rect 8849 1544 8861 1547
rect 7432 1516 8861 1544
rect 7432 1504 7438 1516
rect 8849 1513 8861 1516
rect 8895 1513 8907 1547
rect 8849 1507 8907 1513
rect 9490 1504 9496 1556
rect 9548 1544 9554 1556
rect 10965 1547 11023 1553
rect 10965 1544 10977 1547
rect 9548 1516 10977 1544
rect 9548 1504 9554 1516
rect 10965 1513 10977 1516
rect 11011 1513 11023 1547
rect 10965 1507 11023 1513
rect 13722 1504 13728 1556
rect 13780 1544 13786 1556
rect 15197 1547 15255 1553
rect 15197 1544 15209 1547
rect 13780 1516 15209 1544
rect 13780 1504 13786 1516
rect 15197 1513 15209 1516
rect 15243 1513 15255 1547
rect 15197 1507 15255 1513
rect 24302 1504 24308 1556
rect 24360 1544 24366 1556
rect 25777 1547 25835 1553
rect 25777 1544 25789 1547
rect 24360 1516 25789 1544
rect 24360 1504 24366 1516
rect 25777 1513 25789 1516
rect 25823 1513 25835 1547
rect 25777 1507 25835 1513
rect 26418 1504 26424 1556
rect 26476 1544 26482 1556
rect 27893 1547 27951 1553
rect 27893 1544 27905 1547
rect 26476 1516 27905 1544
rect 26476 1504 26482 1516
rect 27893 1513 27905 1516
rect 27939 1513 27951 1547
rect 27893 1507 27951 1513
rect 30650 1504 30656 1556
rect 30708 1544 30714 1556
rect 32125 1547 32183 1553
rect 32125 1544 32137 1547
rect 30708 1516 32137 1544
rect 30708 1504 30714 1516
rect 32125 1513 32137 1516
rect 32171 1513 32183 1547
rect 32125 1507 32183 1513
rect 41230 1504 41236 1556
rect 41288 1544 41294 1556
rect 42705 1547 42763 1553
rect 42705 1544 42717 1547
rect 41288 1516 42717 1544
rect 41288 1504 41294 1516
rect 42705 1513 42717 1516
rect 42751 1513 42763 1547
rect 42705 1507 42763 1513
rect 43346 1504 43352 1556
rect 43404 1544 43410 1556
rect 44821 1547 44879 1553
rect 44821 1544 44833 1547
rect 43404 1516 44833 1544
rect 43404 1504 43410 1516
rect 44821 1513 44833 1516
rect 44867 1513 44879 1547
rect 44821 1507 44879 1513
rect 47578 1504 47584 1556
rect 47636 1544 47642 1556
rect 49053 1547 49111 1553
rect 49053 1544 49065 1547
rect 47636 1516 49065 1544
rect 47636 1504 47642 1516
rect 49053 1513 49065 1516
rect 49099 1513 49111 1547
rect 49053 1507 49111 1513
rect 58158 1504 58164 1556
rect 58216 1544 58222 1556
rect 59633 1547 59691 1553
rect 59633 1544 59645 1547
rect 58216 1516 59645 1544
rect 58216 1504 58222 1516
rect 59633 1513 59645 1516
rect 59679 1513 59691 1547
rect 59633 1507 59691 1513
rect 64506 1504 64512 1556
rect 64564 1544 64570 1556
rect 65981 1547 66039 1553
rect 65981 1544 65993 1547
rect 64564 1516 65993 1544
rect 64564 1504 64570 1516
rect 65981 1513 65993 1516
rect 66027 1513 66039 1547
rect 65981 1507 66039 1513
rect 75086 1504 75092 1556
rect 75144 1544 75150 1556
rect 76561 1547 76619 1553
rect 76561 1544 76573 1547
rect 75144 1516 76573 1544
rect 75144 1504 75150 1516
rect 76561 1513 76573 1516
rect 76607 1513 76619 1547
rect 76561 1507 76619 1513
rect 77202 1504 77208 1556
rect 77260 1544 77266 1556
rect 78677 1547 78735 1553
rect 78677 1544 78689 1547
rect 77260 1516 78689 1544
rect 77260 1504 77266 1516
rect 78677 1513 78689 1516
rect 78723 1513 78735 1547
rect 78677 1507 78735 1513
rect 81434 1504 81440 1556
rect 81492 1544 81498 1556
rect 82909 1547 82967 1553
rect 82909 1544 82921 1547
rect 81492 1516 82921 1544
rect 81492 1504 81498 1516
rect 82909 1513 82921 1516
rect 82955 1513 82967 1547
rect 82909 1507 82967 1513
rect 92014 1504 92020 1556
rect 92072 1544 92078 1556
rect 93489 1547 93547 1553
rect 93489 1544 93501 1547
rect 92072 1516 93501 1544
rect 92072 1504 92078 1516
rect 93489 1513 93501 1516
rect 93535 1513 93547 1547
rect 93489 1507 93547 1513
rect 94130 1504 94136 1556
rect 94188 1544 94194 1556
rect 95605 1547 95663 1553
rect 95605 1544 95617 1547
rect 94188 1516 95617 1544
rect 94188 1504 94194 1516
rect 95605 1513 95617 1516
rect 95651 1513 95663 1547
rect 95605 1507 95663 1513
rect 98362 1504 98368 1556
rect 98420 1544 98426 1556
rect 99837 1547 99895 1553
rect 99837 1544 99849 1547
rect 98420 1516 99849 1544
rect 98420 1504 98426 1516
rect 99837 1513 99849 1516
rect 99883 1513 99895 1547
rect 99837 1507 99895 1513
rect 1118 1408 1124 1420
rect 1079 1380 1124 1408
rect 1118 1368 1124 1380
rect 1176 1368 1182 1420
rect 1397 1411 1455 1417
rect 1397 1377 1409 1411
rect 1443 1408 1455 1411
rect 2498 1408 2504 1420
rect 1443 1380 2504 1408
rect 1443 1377 1455 1380
rect 1397 1371 1455 1377
rect 2498 1368 2504 1380
rect 2556 1368 2562 1420
rect 3234 1408 3240 1420
rect 3195 1380 3240 1408
rect 3234 1368 3240 1380
rect 3292 1368 3298 1420
rect 3513 1411 3571 1417
rect 3513 1377 3525 1411
rect 3559 1408 3571 1411
rect 4154 1408 4160 1420
rect 3559 1380 4160 1408
rect 3559 1377 3571 1380
rect 3513 1371 3571 1377
rect 4154 1368 4160 1380
rect 4212 1368 4218 1420
rect 5350 1408 5356 1420
rect 5311 1380 5356 1408
rect 5350 1368 5356 1380
rect 5408 1368 5414 1420
rect 5629 1411 5687 1417
rect 5629 1377 5641 1411
rect 5675 1408 5687 1411
rect 5902 1408 5908 1420
rect 5675 1380 5908 1408
rect 5675 1377 5687 1380
rect 5629 1371 5687 1377
rect 5902 1368 5908 1380
rect 5960 1368 5966 1420
rect 7466 1408 7472 1420
rect 7427 1380 7472 1408
rect 7466 1368 7472 1380
rect 7524 1368 7530 1420
rect 7745 1411 7803 1417
rect 7745 1377 7757 1411
rect 7791 1408 7803 1411
rect 8202 1408 8208 1420
rect 7791 1380 8208 1408
rect 7791 1377 7803 1380
rect 7745 1371 7803 1377
rect 8202 1368 8208 1380
rect 8260 1368 8266 1420
rect 9582 1408 9588 1420
rect 9543 1380 9588 1408
rect 9582 1368 9588 1380
rect 9640 1368 9646 1420
rect 9861 1411 9919 1417
rect 9861 1377 9873 1411
rect 9907 1408 9919 1411
rect 11146 1408 11152 1420
rect 9907 1380 11152 1408
rect 9907 1377 9919 1380
rect 9861 1371 9919 1377
rect 11146 1368 11152 1380
rect 11204 1368 11210 1420
rect 11698 1408 11704 1420
rect 11659 1380 11704 1408
rect 11698 1368 11704 1380
rect 11756 1368 11762 1420
rect 11977 1411 12035 1417
rect 11977 1377 11989 1411
rect 12023 1408 12035 1411
rect 13262 1408 13268 1420
rect 12023 1380 13268 1408
rect 12023 1377 12035 1380
rect 11977 1371 12035 1377
rect 13262 1368 13268 1380
rect 13320 1368 13326 1420
rect 13814 1408 13820 1420
rect 13775 1380 13820 1408
rect 13814 1368 13820 1380
rect 13872 1368 13878 1420
rect 14093 1411 14151 1417
rect 14093 1377 14105 1411
rect 14139 1408 14151 1411
rect 15194 1408 15200 1420
rect 14139 1380 15200 1408
rect 14139 1377 14151 1380
rect 14093 1371 14151 1377
rect 15194 1368 15200 1380
rect 15252 1368 15258 1420
rect 15930 1408 15936 1420
rect 15891 1380 15936 1408
rect 15930 1368 15936 1380
rect 15988 1368 15994 1420
rect 16209 1411 16267 1417
rect 16209 1377 16221 1411
rect 16255 1408 16267 1411
rect 17310 1408 17316 1420
rect 16255 1380 17316 1408
rect 16255 1377 16267 1380
rect 16209 1371 16267 1377
rect 17310 1368 17316 1380
rect 17368 1368 17374 1420
rect 18046 1408 18052 1420
rect 18007 1380 18052 1408
rect 18046 1368 18052 1380
rect 18104 1368 18110 1420
rect 18325 1411 18383 1417
rect 18325 1377 18337 1411
rect 18371 1408 18383 1411
rect 18690 1408 18696 1420
rect 18371 1380 18696 1408
rect 18371 1377 18383 1380
rect 18325 1371 18383 1377
rect 18690 1368 18696 1380
rect 18748 1368 18754 1420
rect 20162 1408 20168 1420
rect 20123 1380 20168 1408
rect 20162 1368 20168 1380
rect 20220 1368 20226 1420
rect 20441 1411 20499 1417
rect 20441 1377 20453 1411
rect 20487 1408 20499 1411
rect 20714 1408 20720 1420
rect 20487 1380 20720 1408
rect 20487 1377 20499 1380
rect 20441 1371 20499 1377
rect 20714 1368 20720 1380
rect 20772 1368 20778 1420
rect 22278 1408 22284 1420
rect 22239 1380 22284 1408
rect 22278 1368 22284 1380
rect 22336 1368 22342 1420
rect 22557 1411 22615 1417
rect 22557 1377 22569 1411
rect 22603 1408 22615 1411
rect 22830 1408 22836 1420
rect 22603 1380 22836 1408
rect 22603 1377 22615 1380
rect 22557 1371 22615 1377
rect 22830 1368 22836 1380
rect 22888 1368 22894 1420
rect 24394 1408 24400 1420
rect 24355 1380 24400 1408
rect 24394 1368 24400 1380
rect 24452 1368 24458 1420
rect 24673 1411 24731 1417
rect 24673 1377 24685 1411
rect 24719 1408 24731 1411
rect 25038 1408 25044 1420
rect 24719 1380 25044 1408
rect 24719 1377 24731 1380
rect 24673 1371 24731 1377
rect 25038 1368 25044 1380
rect 25096 1368 25102 1420
rect 26510 1408 26516 1420
rect 26471 1380 26516 1408
rect 26510 1368 26516 1380
rect 26568 1368 26574 1420
rect 26789 1411 26847 1417
rect 26789 1377 26801 1411
rect 26835 1408 26847 1411
rect 28074 1408 28080 1420
rect 26835 1380 28080 1408
rect 26835 1377 26847 1380
rect 26789 1371 26847 1377
rect 28074 1368 28080 1380
rect 28132 1368 28138 1420
rect 28626 1408 28632 1420
rect 28587 1380 28632 1408
rect 28626 1368 28632 1380
rect 28684 1368 28690 1420
rect 28905 1411 28963 1417
rect 28905 1377 28917 1411
rect 28951 1408 28963 1411
rect 30190 1408 30196 1420
rect 28951 1380 30196 1408
rect 28951 1377 28963 1380
rect 28905 1371 28963 1377
rect 30190 1368 30196 1380
rect 30248 1368 30254 1420
rect 30742 1408 30748 1420
rect 30703 1380 30748 1408
rect 30742 1368 30748 1380
rect 30800 1368 30806 1420
rect 31021 1411 31079 1417
rect 31021 1377 31033 1411
rect 31067 1408 31079 1411
rect 32122 1408 32128 1420
rect 31067 1380 32128 1408
rect 31067 1377 31079 1380
rect 31021 1371 31079 1377
rect 32122 1368 32128 1380
rect 32180 1368 32186 1420
rect 32858 1408 32864 1420
rect 32819 1380 32864 1408
rect 32858 1368 32864 1380
rect 32916 1368 32922 1420
rect 33137 1411 33195 1417
rect 33137 1377 33149 1411
rect 33183 1408 33195 1411
rect 34238 1408 34244 1420
rect 33183 1380 34244 1408
rect 33183 1377 33195 1380
rect 33137 1371 33195 1377
rect 34238 1368 34244 1380
rect 34296 1368 34302 1420
rect 34977 1411 35035 1417
rect 34977 1377 34989 1411
rect 35023 1408 35035 1411
rect 35066 1408 35072 1420
rect 35023 1380 35072 1408
rect 35023 1377 35035 1380
rect 34977 1371 35035 1377
rect 35066 1368 35072 1380
rect 35124 1368 35130 1420
rect 35253 1411 35311 1417
rect 35253 1377 35265 1411
rect 35299 1408 35311 1411
rect 35526 1408 35532 1420
rect 35299 1380 35532 1408
rect 35299 1377 35311 1380
rect 35253 1371 35311 1377
rect 35526 1368 35532 1380
rect 35584 1368 35590 1420
rect 37090 1408 37096 1420
rect 37051 1380 37096 1408
rect 37090 1368 37096 1380
rect 37148 1368 37154 1420
rect 37369 1411 37427 1417
rect 37369 1377 37381 1411
rect 37415 1408 37427 1411
rect 37642 1408 37648 1420
rect 37415 1380 37648 1408
rect 37415 1377 37427 1380
rect 37369 1371 37427 1377
rect 37642 1368 37648 1380
rect 37700 1368 37706 1420
rect 39206 1408 39212 1420
rect 39167 1380 39212 1408
rect 39206 1368 39212 1380
rect 39264 1368 39270 1420
rect 39485 1411 39543 1417
rect 39485 1377 39497 1411
rect 39531 1408 39543 1411
rect 40126 1408 40132 1420
rect 39531 1380 40132 1408
rect 39531 1377 39543 1380
rect 39485 1371 39543 1377
rect 40126 1368 40132 1380
rect 40184 1368 40190 1420
rect 41322 1408 41328 1420
rect 41283 1380 41328 1408
rect 41322 1368 41328 1380
rect 41380 1368 41386 1420
rect 41601 1411 41659 1417
rect 41601 1377 41613 1411
rect 41647 1408 41659 1411
rect 41966 1408 41972 1420
rect 41647 1380 41972 1408
rect 41647 1377 41659 1380
rect 41601 1371 41659 1377
rect 41966 1368 41972 1380
rect 42024 1368 42030 1420
rect 43438 1408 43444 1420
rect 43399 1380 43444 1408
rect 43438 1368 43444 1380
rect 43496 1368 43502 1420
rect 43717 1411 43775 1417
rect 43717 1377 43729 1411
rect 43763 1408 43775 1411
rect 45002 1408 45008 1420
rect 43763 1380 45008 1408
rect 43763 1377 43775 1380
rect 43717 1371 43775 1377
rect 45002 1368 45008 1380
rect 45060 1368 45066 1420
rect 45554 1408 45560 1420
rect 45515 1380 45560 1408
rect 45554 1368 45560 1380
rect 45612 1368 45618 1420
rect 45833 1411 45891 1417
rect 45833 1377 45845 1411
rect 45879 1408 45891 1411
rect 47118 1408 47124 1420
rect 45879 1380 47124 1408
rect 45879 1377 45891 1380
rect 45833 1371 45891 1377
rect 47118 1368 47124 1380
rect 47176 1368 47182 1420
rect 47670 1408 47676 1420
rect 47631 1380 47676 1408
rect 47670 1368 47676 1380
rect 47728 1368 47734 1420
rect 47949 1411 48007 1417
rect 47949 1377 47961 1411
rect 47995 1408 48007 1411
rect 49050 1408 49056 1420
rect 47995 1380 49056 1408
rect 47995 1377 48007 1380
rect 47949 1371 48007 1377
rect 49050 1368 49056 1380
rect 49108 1368 49114 1420
rect 49786 1408 49792 1420
rect 49747 1380 49792 1408
rect 49786 1368 49792 1380
rect 49844 1368 49850 1420
rect 50065 1411 50123 1417
rect 50065 1377 50077 1411
rect 50111 1408 50123 1411
rect 51166 1408 51172 1420
rect 50111 1380 51172 1408
rect 50111 1377 50123 1380
rect 50065 1371 50123 1377
rect 51166 1368 51172 1380
rect 51224 1368 51230 1420
rect 51902 1408 51908 1420
rect 51863 1380 51908 1408
rect 51902 1368 51908 1380
rect 51960 1368 51966 1420
rect 52181 1411 52239 1417
rect 52181 1377 52193 1411
rect 52227 1408 52239 1411
rect 52270 1408 52276 1420
rect 52227 1380 52276 1408
rect 52227 1377 52239 1380
rect 52181 1371 52239 1377
rect 52270 1368 52276 1380
rect 52328 1368 52334 1420
rect 54018 1408 54024 1420
rect 53979 1380 54024 1408
rect 54018 1368 54024 1380
rect 54076 1368 54082 1420
rect 54297 1411 54355 1417
rect 54297 1377 54309 1411
rect 54343 1408 54355 1411
rect 54754 1408 54760 1420
rect 54343 1380 54760 1408
rect 54343 1377 54355 1380
rect 54297 1371 54355 1377
rect 54754 1368 54760 1380
rect 54812 1368 54818 1420
rect 56134 1408 56140 1420
rect 56095 1380 56140 1408
rect 56134 1368 56140 1380
rect 56192 1368 56198 1420
rect 56413 1411 56471 1417
rect 56413 1377 56425 1411
rect 56459 1408 56471 1411
rect 56686 1408 56692 1420
rect 56459 1380 56692 1408
rect 56459 1377 56471 1380
rect 56413 1371 56471 1377
rect 56686 1368 56692 1380
rect 56744 1368 56750 1420
rect 58250 1408 58256 1420
rect 58211 1380 58256 1408
rect 58250 1368 58256 1380
rect 58308 1368 58314 1420
rect 58529 1411 58587 1417
rect 58529 1377 58541 1411
rect 58575 1408 58587 1411
rect 58894 1408 58900 1420
rect 58575 1380 58900 1408
rect 58575 1377 58587 1380
rect 58529 1371 58587 1377
rect 58894 1368 58900 1380
rect 58952 1368 58958 1420
rect 60366 1368 60372 1420
rect 60424 1408 60430 1420
rect 60645 1411 60703 1417
rect 60424 1380 60469 1408
rect 60424 1368 60430 1380
rect 60645 1377 60657 1411
rect 60691 1408 60703 1411
rect 61930 1408 61936 1420
rect 60691 1380 61936 1408
rect 60691 1377 60703 1380
rect 60645 1371 60703 1377
rect 61930 1368 61936 1380
rect 61988 1368 61994 1420
rect 62482 1408 62488 1420
rect 62443 1380 62488 1408
rect 62482 1368 62488 1380
rect 62540 1368 62546 1420
rect 62761 1411 62819 1417
rect 62761 1377 62773 1411
rect 62807 1408 62819 1411
rect 64046 1408 64052 1420
rect 62807 1380 64052 1408
rect 62807 1377 62819 1380
rect 62761 1371 62819 1377
rect 64046 1368 64052 1380
rect 64104 1368 64110 1420
rect 64598 1408 64604 1420
rect 64559 1380 64604 1408
rect 64598 1368 64604 1380
rect 64656 1368 64662 1420
rect 64877 1411 64935 1417
rect 64877 1377 64889 1411
rect 64923 1408 64935 1411
rect 65978 1408 65984 1420
rect 64923 1380 65984 1408
rect 64923 1377 64935 1380
rect 64877 1371 64935 1377
rect 65978 1368 65984 1380
rect 66036 1368 66042 1420
rect 66714 1408 66720 1420
rect 66675 1380 66720 1408
rect 66714 1368 66720 1380
rect 66772 1368 66778 1420
rect 66993 1411 67051 1417
rect 66993 1377 67005 1411
rect 67039 1408 67051 1411
rect 68094 1408 68100 1420
rect 67039 1380 68100 1408
rect 67039 1377 67051 1380
rect 66993 1371 67051 1377
rect 68094 1368 68100 1380
rect 68152 1368 68158 1420
rect 68830 1408 68836 1420
rect 68791 1380 68836 1408
rect 68830 1368 68836 1380
rect 68888 1368 68894 1420
rect 69109 1411 69167 1417
rect 69109 1377 69121 1411
rect 69155 1408 69167 1411
rect 69198 1408 69204 1420
rect 69155 1380 69204 1408
rect 69155 1377 69167 1380
rect 69109 1371 69167 1377
rect 69198 1368 69204 1380
rect 69256 1368 69262 1420
rect 70946 1408 70952 1420
rect 70907 1380 70952 1408
rect 70946 1368 70952 1380
rect 71004 1368 71010 1420
rect 71225 1411 71283 1417
rect 71225 1377 71237 1411
rect 71271 1408 71283 1411
rect 71498 1408 71504 1420
rect 71271 1380 71504 1408
rect 71271 1377 71283 1380
rect 71225 1371 71283 1377
rect 71498 1368 71504 1380
rect 71556 1368 71562 1420
rect 73062 1408 73068 1420
rect 73023 1380 73068 1408
rect 73062 1368 73068 1380
rect 73120 1368 73126 1420
rect 73341 1411 73399 1417
rect 73341 1377 73353 1411
rect 73387 1408 73399 1411
rect 73614 1408 73620 1420
rect 73387 1380 73620 1408
rect 73387 1377 73399 1380
rect 73341 1371 73399 1377
rect 73614 1368 73620 1380
rect 73672 1368 73678 1420
rect 75178 1408 75184 1420
rect 75139 1380 75184 1408
rect 75178 1368 75184 1380
rect 75236 1368 75242 1420
rect 75457 1411 75515 1417
rect 75457 1377 75469 1411
rect 75503 1408 75515 1411
rect 76190 1408 76196 1420
rect 75503 1380 76196 1408
rect 75503 1377 75515 1380
rect 75457 1371 75515 1377
rect 76190 1368 76196 1380
rect 76248 1368 76254 1420
rect 77294 1368 77300 1420
rect 77352 1408 77358 1420
rect 77573 1411 77631 1417
rect 77352 1380 77397 1408
rect 77352 1368 77358 1380
rect 77573 1377 77585 1411
rect 77619 1408 77631 1411
rect 78858 1408 78864 1420
rect 77619 1380 78864 1408
rect 77619 1377 77631 1380
rect 77573 1371 77631 1377
rect 78858 1368 78864 1380
rect 78916 1368 78922 1420
rect 79410 1408 79416 1420
rect 79371 1380 79416 1408
rect 79410 1368 79416 1380
rect 79468 1368 79474 1420
rect 79689 1411 79747 1417
rect 79689 1377 79701 1411
rect 79735 1408 79747 1411
rect 81158 1408 81164 1420
rect 79735 1380 81164 1408
rect 79735 1377 79747 1380
rect 79689 1371 79747 1377
rect 81158 1368 81164 1380
rect 81216 1368 81222 1420
rect 81526 1408 81532 1420
rect 81487 1380 81532 1408
rect 81526 1368 81532 1380
rect 81584 1368 81590 1420
rect 81805 1411 81863 1417
rect 81805 1377 81817 1411
rect 81851 1408 81863 1411
rect 82906 1408 82912 1420
rect 81851 1380 82912 1408
rect 81851 1377 81863 1380
rect 81805 1371 81863 1377
rect 82906 1368 82912 1380
rect 82964 1368 82970 1420
rect 83642 1408 83648 1420
rect 83603 1380 83648 1408
rect 83642 1368 83648 1380
rect 83700 1368 83706 1420
rect 83921 1411 83979 1417
rect 83921 1377 83933 1411
rect 83967 1408 83979 1411
rect 85022 1408 85028 1420
rect 83967 1380 85028 1408
rect 83967 1377 83979 1380
rect 83921 1371 83979 1377
rect 85022 1368 85028 1380
rect 85080 1368 85086 1420
rect 85758 1408 85764 1420
rect 85719 1380 85764 1408
rect 85758 1368 85764 1380
rect 85816 1368 85822 1420
rect 86037 1411 86095 1417
rect 86037 1377 86049 1411
rect 86083 1408 86095 1411
rect 86494 1408 86500 1420
rect 86083 1380 86500 1408
rect 86083 1377 86095 1380
rect 86037 1371 86095 1377
rect 86494 1368 86500 1380
rect 86552 1368 86558 1420
rect 87874 1408 87880 1420
rect 87835 1380 87880 1408
rect 87874 1368 87880 1380
rect 87932 1368 87938 1420
rect 88153 1411 88211 1417
rect 88153 1377 88165 1411
rect 88199 1408 88211 1411
rect 88426 1408 88432 1420
rect 88199 1380 88432 1408
rect 88199 1377 88211 1380
rect 88153 1371 88211 1377
rect 88426 1368 88432 1380
rect 88484 1368 88490 1420
rect 89990 1408 89996 1420
rect 89951 1380 89996 1408
rect 89990 1368 89996 1380
rect 90048 1368 90054 1420
rect 90269 1411 90327 1417
rect 90269 1377 90281 1411
rect 90315 1408 90327 1411
rect 90726 1408 90732 1420
rect 90315 1380 90732 1408
rect 90315 1377 90327 1380
rect 90269 1371 90327 1377
rect 90726 1368 90732 1380
rect 90784 1368 90790 1420
rect 92106 1408 92112 1420
rect 92067 1380 92112 1408
rect 92106 1368 92112 1380
rect 92164 1368 92170 1420
rect 92385 1411 92443 1417
rect 92385 1377 92397 1411
rect 92431 1408 92443 1411
rect 92750 1408 92756 1420
rect 92431 1380 92756 1408
rect 92431 1377 92443 1380
rect 92385 1371 92443 1377
rect 92750 1368 92756 1380
rect 92808 1368 92814 1420
rect 94222 1408 94228 1420
rect 94183 1380 94228 1408
rect 94222 1368 94228 1380
rect 94280 1368 94286 1420
rect 94501 1411 94559 1417
rect 94501 1377 94513 1411
rect 94547 1408 94559 1411
rect 95786 1408 95792 1420
rect 94547 1380 95792 1408
rect 94547 1377 94559 1380
rect 94501 1371 94559 1377
rect 95786 1368 95792 1380
rect 95844 1368 95850 1420
rect 96062 1368 96068 1420
rect 96120 1408 96126 1420
rect 96341 1411 96399 1417
rect 96341 1408 96353 1411
rect 96120 1380 96353 1408
rect 96120 1368 96126 1380
rect 96341 1377 96353 1380
rect 96387 1377 96399 1411
rect 96341 1371 96399 1377
rect 96617 1411 96675 1417
rect 96617 1377 96629 1411
rect 96663 1408 96675 1411
rect 97902 1408 97908 1420
rect 96663 1380 97908 1408
rect 96663 1377 96675 1380
rect 96617 1371 96675 1377
rect 97902 1368 97908 1380
rect 97960 1368 97966 1420
rect 98454 1408 98460 1420
rect 98415 1380 98460 1408
rect 98454 1368 98460 1380
rect 98512 1368 98518 1420
rect 98733 1411 98791 1417
rect 98733 1377 98745 1411
rect 98779 1408 98791 1411
rect 99834 1408 99840 1420
rect 98779 1380 99840 1408
rect 98779 1377 98791 1380
rect 98733 1371 98791 1377
rect 99834 1368 99840 1380
rect 99892 1368 99898 1420
rect 100570 1408 100576 1420
rect 100531 1380 100576 1408
rect 100570 1368 100576 1380
rect 100628 1368 100634 1420
rect 100849 1411 100907 1417
rect 100849 1377 100861 1411
rect 100895 1408 100907 1411
rect 101950 1408 101956 1420
rect 100895 1380 101956 1408
rect 100895 1377 100907 1380
rect 100849 1371 100907 1377
rect 101950 1368 101956 1380
rect 102008 1368 102014 1420
rect 102686 1408 102692 1420
rect 102647 1380 102692 1408
rect 102686 1368 102692 1380
rect 102744 1368 102750 1420
rect 102965 1411 103023 1417
rect 102965 1377 102977 1411
rect 103011 1408 103023 1411
rect 103238 1408 103244 1420
rect 103011 1380 103244 1408
rect 103011 1377 103023 1380
rect 102965 1371 103023 1377
rect 103238 1368 103244 1380
rect 103296 1368 103302 1420
rect 104802 1408 104808 1420
rect 104763 1380 104808 1408
rect 104802 1368 104808 1380
rect 104860 1368 104866 1420
rect 105081 1411 105139 1417
rect 105081 1377 105093 1411
rect 105127 1408 105139 1411
rect 105354 1408 105360 1420
rect 105127 1380 105360 1408
rect 105127 1377 105139 1380
rect 105081 1371 105139 1377
rect 105354 1368 105360 1380
rect 105412 1368 105418 1420
rect 3418 1164 3424 1216
rect 3476 1204 3482 1216
rect 4617 1207 4675 1213
rect 4617 1204 4629 1207
rect 3476 1176 4629 1204
rect 3476 1164 3482 1176
rect 4617 1173 4629 1176
rect 4663 1173 4675 1207
rect 4617 1167 4675 1173
rect 5626 1164 5632 1216
rect 5684 1204 5690 1216
rect 6733 1207 6791 1213
rect 6733 1204 6745 1207
rect 5684 1176 6745 1204
rect 5684 1164 5690 1176
rect 6733 1173 6745 1176
rect 6779 1173 6791 1207
rect 6733 1167 6791 1173
rect 11606 1164 11612 1216
rect 11664 1204 11670 1216
rect 13081 1207 13139 1213
rect 13081 1204 13093 1207
rect 11664 1176 13093 1204
rect 11664 1164 11670 1176
rect 13081 1173 13093 1176
rect 13127 1173 13139 1207
rect 13081 1167 13139 1173
rect 16114 1164 16120 1216
rect 16172 1204 16178 1216
rect 17313 1207 17371 1213
rect 17313 1204 17325 1207
rect 16172 1176 17325 1204
rect 16172 1164 16178 1176
rect 17313 1173 17325 1176
rect 17359 1173 17371 1207
rect 17313 1167 17371 1173
rect 18322 1164 18328 1216
rect 18380 1204 18386 1216
rect 19429 1207 19487 1213
rect 19429 1204 19441 1207
rect 18380 1176 19441 1204
rect 18380 1164 18386 1176
rect 19429 1173 19441 1176
rect 19475 1173 19487 1207
rect 19429 1167 19487 1173
rect 20346 1164 20352 1216
rect 20404 1204 20410 1216
rect 21545 1207 21603 1213
rect 21545 1204 21557 1207
rect 20404 1176 21557 1204
rect 20404 1164 20410 1176
rect 21545 1173 21557 1176
rect 21591 1173 21603 1207
rect 21545 1167 21603 1173
rect 22554 1164 22560 1216
rect 22612 1204 22618 1216
rect 23661 1207 23719 1213
rect 23661 1204 23673 1207
rect 22612 1176 23673 1204
rect 22612 1164 22618 1176
rect 23661 1173 23673 1176
rect 23707 1173 23719 1207
rect 23661 1167 23719 1173
rect 28534 1164 28540 1216
rect 28592 1204 28598 1216
rect 30009 1207 30067 1213
rect 30009 1204 30021 1207
rect 28592 1176 30021 1204
rect 28592 1164 28598 1176
rect 30009 1173 30021 1176
rect 30055 1173 30067 1207
rect 30009 1167 30067 1173
rect 33042 1164 33048 1216
rect 33100 1204 33106 1216
rect 34241 1207 34299 1213
rect 34241 1204 34253 1207
rect 33100 1176 34253 1204
rect 33100 1164 33106 1176
rect 34241 1173 34253 1176
rect 34287 1173 34299 1207
rect 34241 1167 34299 1173
rect 35250 1164 35256 1216
rect 35308 1204 35314 1216
rect 36357 1207 36415 1213
rect 36357 1204 36369 1207
rect 35308 1176 36369 1204
rect 35308 1164 35314 1176
rect 36357 1173 36369 1176
rect 36403 1173 36415 1207
rect 36357 1167 36415 1173
rect 37274 1164 37280 1216
rect 37332 1204 37338 1216
rect 38473 1207 38531 1213
rect 38473 1204 38485 1207
rect 37332 1176 38485 1204
rect 37332 1164 37338 1176
rect 38473 1173 38485 1176
rect 38519 1173 38531 1207
rect 38473 1167 38531 1173
rect 39482 1164 39488 1216
rect 39540 1204 39546 1216
rect 40589 1207 40647 1213
rect 40589 1204 40601 1207
rect 39540 1176 40601 1204
rect 39540 1164 39546 1176
rect 40589 1173 40601 1176
rect 40635 1173 40647 1207
rect 40589 1167 40647 1173
rect 45462 1164 45468 1216
rect 45520 1204 45526 1216
rect 46937 1207 46995 1213
rect 46937 1204 46949 1207
rect 45520 1176 46949 1204
rect 45520 1164 45526 1176
rect 46937 1173 46949 1176
rect 46983 1173 46995 1207
rect 46937 1167 46995 1173
rect 49970 1164 49976 1216
rect 50028 1204 50034 1216
rect 51169 1207 51227 1213
rect 51169 1204 51181 1207
rect 50028 1176 51181 1204
rect 50028 1164 50034 1176
rect 51169 1173 51181 1176
rect 51215 1173 51227 1207
rect 51169 1167 51227 1173
rect 52178 1164 52184 1216
rect 52236 1204 52242 1216
rect 53285 1207 53343 1213
rect 53285 1204 53297 1207
rect 52236 1176 53297 1204
rect 52236 1164 52242 1176
rect 53285 1173 53297 1176
rect 53331 1173 53343 1207
rect 53285 1167 53343 1173
rect 54202 1164 54208 1216
rect 54260 1204 54266 1216
rect 55401 1207 55459 1213
rect 55401 1204 55413 1207
rect 54260 1176 55413 1204
rect 54260 1164 54266 1176
rect 55401 1173 55413 1176
rect 55447 1173 55459 1207
rect 55401 1167 55459 1173
rect 56410 1164 56416 1216
rect 56468 1204 56474 1216
rect 57517 1207 57575 1213
rect 57517 1204 57529 1207
rect 56468 1176 57529 1204
rect 56468 1164 56474 1176
rect 57517 1173 57529 1176
rect 57563 1173 57575 1207
rect 57517 1167 57575 1173
rect 60274 1164 60280 1216
rect 60332 1204 60338 1216
rect 61749 1207 61807 1213
rect 61749 1204 61761 1207
rect 60332 1176 61761 1204
rect 60332 1164 60338 1176
rect 61749 1173 61761 1176
rect 61795 1173 61807 1207
rect 61749 1167 61807 1173
rect 62390 1164 62396 1216
rect 62448 1204 62454 1216
rect 63865 1207 63923 1213
rect 63865 1204 63877 1207
rect 62448 1176 63877 1204
rect 62448 1164 62454 1176
rect 63865 1173 63877 1176
rect 63911 1173 63923 1207
rect 63865 1167 63923 1173
rect 66898 1164 66904 1216
rect 66956 1204 66962 1216
rect 68097 1207 68155 1213
rect 68097 1204 68109 1207
rect 66956 1176 68109 1204
rect 66956 1164 66962 1176
rect 68097 1173 68109 1176
rect 68143 1173 68155 1207
rect 68097 1167 68155 1173
rect 69106 1164 69112 1216
rect 69164 1204 69170 1216
rect 70213 1207 70271 1213
rect 70213 1204 70225 1207
rect 69164 1176 70225 1204
rect 69164 1164 69170 1176
rect 70213 1173 70225 1176
rect 70259 1173 70271 1207
rect 70213 1167 70271 1173
rect 71130 1164 71136 1216
rect 71188 1204 71194 1216
rect 72329 1207 72387 1213
rect 72329 1204 72341 1207
rect 71188 1176 72341 1204
rect 71188 1164 71194 1176
rect 72329 1173 72341 1176
rect 72375 1173 72387 1207
rect 72329 1167 72387 1173
rect 73338 1164 73344 1216
rect 73396 1204 73402 1216
rect 74445 1207 74503 1213
rect 74445 1204 74457 1207
rect 73396 1176 74457 1204
rect 73396 1164 73402 1176
rect 74445 1173 74457 1176
rect 74491 1173 74503 1207
rect 74445 1167 74503 1173
rect 79318 1164 79324 1216
rect 79376 1204 79382 1216
rect 80793 1207 80851 1213
rect 80793 1204 80805 1207
rect 79376 1176 80805 1204
rect 79376 1164 79382 1176
rect 80793 1173 80805 1176
rect 80839 1173 80851 1207
rect 80793 1167 80851 1173
rect 83826 1164 83832 1216
rect 83884 1204 83890 1216
rect 85025 1207 85083 1213
rect 85025 1204 85037 1207
rect 83884 1176 85037 1204
rect 83884 1164 83890 1176
rect 85025 1173 85037 1176
rect 85071 1173 85083 1207
rect 85025 1167 85083 1173
rect 86034 1164 86040 1216
rect 86092 1204 86098 1216
rect 87141 1207 87199 1213
rect 87141 1204 87153 1207
rect 86092 1176 87153 1204
rect 86092 1164 86098 1176
rect 87141 1173 87153 1176
rect 87187 1173 87199 1207
rect 87141 1167 87199 1173
rect 88058 1164 88064 1216
rect 88116 1204 88122 1216
rect 89257 1207 89315 1213
rect 89257 1204 89269 1207
rect 88116 1176 89269 1204
rect 88116 1164 88122 1176
rect 89257 1173 89269 1176
rect 89303 1173 89315 1207
rect 89257 1167 89315 1173
rect 90266 1164 90272 1216
rect 90324 1204 90330 1216
rect 91373 1207 91431 1213
rect 91373 1204 91385 1207
rect 90324 1176 91385 1204
rect 90324 1164 90330 1176
rect 91373 1173 91385 1176
rect 91419 1173 91431 1207
rect 91373 1167 91431 1173
rect 96522 1164 96528 1216
rect 96580 1204 96586 1216
rect 97721 1207 97779 1213
rect 97721 1204 97733 1207
rect 96580 1176 97733 1204
rect 96580 1164 96586 1176
rect 97721 1173 97733 1176
rect 97767 1173 97779 1207
rect 97721 1167 97779 1173
rect 100754 1164 100760 1216
rect 100812 1204 100818 1216
rect 101953 1207 102011 1213
rect 101953 1204 101965 1207
rect 100812 1176 101965 1204
rect 100812 1164 100818 1176
rect 101953 1173 101965 1176
rect 101999 1173 102011 1207
rect 101953 1167 102011 1173
rect 102962 1164 102968 1216
rect 103020 1204 103026 1216
rect 104069 1207 104127 1213
rect 104069 1204 104081 1207
rect 103020 1176 104081 1204
rect 103020 1164 103026 1176
rect 104069 1173 104081 1176
rect 104115 1173 104127 1207
rect 104069 1167 104127 1173
rect 104986 1164 104992 1216
rect 105044 1204 105050 1216
rect 106185 1207 106243 1213
rect 106185 1204 106197 1207
rect 105044 1176 106197 1204
rect 105044 1164 105050 1176
rect 106185 1173 106197 1176
rect 106231 1173 106243 1207
rect 106185 1167 106243 1173
rect 1104 1114 106904 1136
rect 1104 1062 4042 1114
rect 4094 1062 4106 1114
rect 4158 1062 4170 1114
rect 4222 1062 4234 1114
rect 4286 1062 34762 1114
rect 34814 1062 34826 1114
rect 34878 1062 34890 1114
rect 34942 1062 34954 1114
rect 35006 1062 65482 1114
rect 65534 1062 65546 1114
rect 65598 1062 65610 1114
rect 65662 1062 65674 1114
rect 65726 1062 96202 1114
rect 96254 1062 96266 1114
rect 96318 1062 96330 1114
rect 96382 1062 96394 1114
rect 96446 1062 106904 1114
rect 1104 1040 106904 1062
<< via1 >>
rect 4042 7590 4094 7642
rect 4106 7590 4158 7642
rect 4170 7590 4222 7642
rect 4234 7590 4286 7642
rect 34762 7590 34814 7642
rect 34826 7590 34878 7642
rect 34890 7590 34942 7642
rect 34954 7590 35006 7642
rect 65482 7590 65534 7642
rect 65546 7590 65598 7642
rect 65610 7590 65662 7642
rect 65674 7590 65726 7642
rect 96202 7590 96254 7642
rect 96266 7590 96318 7642
rect 96330 7590 96382 7642
rect 96394 7590 96446 7642
rect 1124 7327 1176 7336
rect 1124 7293 1133 7327
rect 1133 7293 1167 7327
rect 1167 7293 1176 7327
rect 1124 7284 1176 7293
rect 3240 7327 3292 7336
rect 3240 7293 3249 7327
rect 3249 7293 3283 7327
rect 3283 7293 3292 7327
rect 3240 7284 3292 7293
rect 3516 7327 3568 7336
rect 3516 7293 3525 7327
rect 3525 7293 3559 7327
rect 3559 7293 3568 7327
rect 3516 7284 3568 7293
rect 5264 7284 5316 7336
rect 5632 7327 5684 7336
rect 5632 7293 5641 7327
rect 5641 7293 5675 7327
rect 5675 7293 5684 7327
rect 5632 7284 5684 7293
rect 7380 7284 7432 7336
rect 7748 7327 7800 7336
rect 7748 7293 7757 7327
rect 7757 7293 7791 7327
rect 7791 7293 7800 7327
rect 7748 7284 7800 7293
rect 9588 7327 9640 7336
rect 9588 7293 9597 7327
rect 9597 7293 9631 7327
rect 9631 7293 9640 7327
rect 9588 7284 9640 7293
rect 9864 7327 9916 7336
rect 9864 7293 9873 7327
rect 9873 7293 9907 7327
rect 9907 7293 9916 7327
rect 9864 7284 9916 7293
rect 11704 7327 11756 7336
rect 11704 7293 11713 7327
rect 11713 7293 11747 7327
rect 11747 7293 11756 7327
rect 11704 7284 11756 7293
rect 11980 7327 12032 7336
rect 11980 7293 11989 7327
rect 11989 7293 12023 7327
rect 12023 7293 12032 7327
rect 11980 7284 12032 7293
rect 13820 7327 13872 7336
rect 13820 7293 13829 7327
rect 13829 7293 13863 7327
rect 13863 7293 13872 7327
rect 13820 7284 13872 7293
rect 14096 7327 14148 7336
rect 14096 7293 14105 7327
rect 14105 7293 14139 7327
rect 14139 7293 14148 7327
rect 14096 7284 14148 7293
rect 15936 7327 15988 7336
rect 15936 7293 15945 7327
rect 15945 7293 15979 7327
rect 15979 7293 15988 7327
rect 15936 7284 15988 7293
rect 16212 7327 16264 7336
rect 16212 7293 16221 7327
rect 16221 7293 16255 7327
rect 16255 7293 16264 7327
rect 16212 7284 16264 7293
rect 18052 7327 18104 7336
rect 18052 7293 18061 7327
rect 18061 7293 18095 7327
rect 18095 7293 18104 7327
rect 18052 7284 18104 7293
rect 18328 7327 18380 7336
rect 18328 7293 18337 7327
rect 18337 7293 18371 7327
rect 18371 7293 18380 7327
rect 18328 7284 18380 7293
rect 20076 7284 20128 7336
rect 20444 7327 20496 7336
rect 20444 7293 20453 7327
rect 20453 7293 20487 7327
rect 20487 7293 20496 7327
rect 20444 7284 20496 7293
rect 22192 7284 22244 7336
rect 22560 7327 22612 7336
rect 22560 7293 22569 7327
rect 22569 7293 22603 7327
rect 22603 7293 22612 7327
rect 22560 7284 22612 7293
rect 24400 7327 24452 7336
rect 24400 7293 24409 7327
rect 24409 7293 24443 7327
rect 24443 7293 24452 7327
rect 24400 7284 24452 7293
rect 24676 7327 24728 7336
rect 24676 7293 24685 7327
rect 24685 7293 24719 7327
rect 24719 7293 24728 7327
rect 24676 7284 24728 7293
rect 26516 7327 26568 7336
rect 26516 7293 26525 7327
rect 26525 7293 26559 7327
rect 26559 7293 26568 7327
rect 26516 7284 26568 7293
rect 26792 7327 26844 7336
rect 26792 7293 26801 7327
rect 26801 7293 26835 7327
rect 26835 7293 26844 7327
rect 26792 7284 26844 7293
rect 28632 7327 28684 7336
rect 28632 7293 28641 7327
rect 28641 7293 28675 7327
rect 28675 7293 28684 7327
rect 28632 7284 28684 7293
rect 28908 7327 28960 7336
rect 28908 7293 28917 7327
rect 28917 7293 28951 7327
rect 28951 7293 28960 7327
rect 28908 7284 28960 7293
rect 30748 7327 30800 7336
rect 30748 7293 30757 7327
rect 30757 7293 30791 7327
rect 30791 7293 30800 7327
rect 30748 7284 30800 7293
rect 31024 7327 31076 7336
rect 31024 7293 31033 7327
rect 31033 7293 31067 7327
rect 31067 7293 31076 7327
rect 31024 7284 31076 7293
rect 32864 7327 32916 7336
rect 32864 7293 32873 7327
rect 32873 7293 32907 7327
rect 32907 7293 32916 7327
rect 32864 7284 32916 7293
rect 33140 7327 33192 7336
rect 33140 7293 33149 7327
rect 33149 7293 33183 7327
rect 33183 7293 33192 7327
rect 33140 7284 33192 7293
rect 35072 7284 35124 7336
rect 35256 7327 35308 7336
rect 35256 7293 35265 7327
rect 35265 7293 35299 7327
rect 35299 7293 35308 7327
rect 35256 7284 35308 7293
rect 37096 7327 37148 7336
rect 37096 7293 37105 7327
rect 37105 7293 37139 7327
rect 37139 7293 37148 7327
rect 37096 7284 37148 7293
rect 37372 7327 37424 7336
rect 37372 7293 37381 7327
rect 37381 7293 37415 7327
rect 37415 7293 37424 7327
rect 37372 7284 37424 7293
rect 39212 7327 39264 7336
rect 39212 7293 39221 7327
rect 39221 7293 39255 7327
rect 39255 7293 39264 7327
rect 39212 7284 39264 7293
rect 39488 7327 39540 7336
rect 39488 7293 39497 7327
rect 39497 7293 39531 7327
rect 39531 7293 39540 7327
rect 39488 7284 39540 7293
rect 41236 7284 41288 7336
rect 41604 7327 41656 7336
rect 41604 7293 41613 7327
rect 41613 7293 41647 7327
rect 41647 7293 41656 7327
rect 41604 7284 41656 7293
rect 43444 7327 43496 7336
rect 43444 7293 43453 7327
rect 43453 7293 43487 7327
rect 43487 7293 43496 7327
rect 43444 7284 43496 7293
rect 43720 7327 43772 7336
rect 43720 7293 43729 7327
rect 43729 7293 43763 7327
rect 43763 7293 43772 7327
rect 43720 7284 43772 7293
rect 45560 7327 45612 7336
rect 45560 7293 45569 7327
rect 45569 7293 45603 7327
rect 45603 7293 45612 7327
rect 45560 7284 45612 7293
rect 45836 7327 45888 7336
rect 45836 7293 45845 7327
rect 45845 7293 45879 7327
rect 45879 7293 45888 7327
rect 45836 7284 45888 7293
rect 47676 7327 47728 7336
rect 47676 7293 47685 7327
rect 47685 7293 47719 7327
rect 47719 7293 47728 7327
rect 47676 7284 47728 7293
rect 47952 7327 48004 7336
rect 47952 7293 47961 7327
rect 47961 7293 47995 7327
rect 47995 7293 48004 7327
rect 47952 7284 48004 7293
rect 49792 7327 49844 7336
rect 49792 7293 49801 7327
rect 49801 7293 49835 7327
rect 49835 7293 49844 7327
rect 49792 7284 49844 7293
rect 51172 7284 51224 7336
rect 51908 7327 51960 7336
rect 51908 7293 51917 7327
rect 51917 7293 51951 7327
rect 51951 7293 51960 7327
rect 51908 7284 51960 7293
rect 52184 7327 52236 7336
rect 52184 7293 52193 7327
rect 52193 7293 52227 7327
rect 52227 7293 52236 7327
rect 52184 7284 52236 7293
rect 54024 7327 54076 7336
rect 54024 7293 54033 7327
rect 54033 7293 54067 7327
rect 54067 7293 54076 7327
rect 54024 7284 54076 7293
rect 54300 7327 54352 7336
rect 54300 7293 54309 7327
rect 54309 7293 54343 7327
rect 54343 7293 54352 7327
rect 54300 7284 54352 7293
rect 56048 7284 56100 7336
rect 56416 7327 56468 7336
rect 56416 7293 56425 7327
rect 56425 7293 56459 7327
rect 56459 7293 56468 7327
rect 56416 7284 56468 7293
rect 58164 7284 58216 7336
rect 58532 7327 58584 7336
rect 58532 7293 58541 7327
rect 58541 7293 58575 7327
rect 58575 7293 58584 7327
rect 58532 7284 58584 7293
rect 60372 7327 60424 7336
rect 60372 7293 60381 7327
rect 60381 7293 60415 7327
rect 60415 7293 60424 7327
rect 60648 7327 60700 7336
rect 60372 7284 60424 7293
rect 60648 7293 60657 7327
rect 60657 7293 60691 7327
rect 60691 7293 60700 7327
rect 60648 7284 60700 7293
rect 62488 7327 62540 7336
rect 62488 7293 62497 7327
rect 62497 7293 62531 7327
rect 62531 7293 62540 7327
rect 62488 7284 62540 7293
rect 62764 7327 62816 7336
rect 62764 7293 62773 7327
rect 62773 7293 62807 7327
rect 62807 7293 62816 7327
rect 62764 7284 62816 7293
rect 64604 7327 64656 7336
rect 64604 7293 64613 7327
rect 64613 7293 64647 7327
rect 64647 7293 64656 7327
rect 64604 7284 64656 7293
rect 64880 7327 64932 7336
rect 64880 7293 64889 7327
rect 64889 7293 64923 7327
rect 64923 7293 64932 7327
rect 64880 7284 64932 7293
rect 66720 7327 66772 7336
rect 66720 7293 66729 7327
rect 66729 7293 66763 7327
rect 66763 7293 66772 7327
rect 66720 7284 66772 7293
rect 66996 7327 67048 7336
rect 66996 7293 67005 7327
rect 67005 7293 67039 7327
rect 67039 7293 67048 7327
rect 66996 7284 67048 7293
rect 68836 7327 68888 7336
rect 68836 7293 68845 7327
rect 68845 7293 68879 7327
rect 68879 7293 68888 7327
rect 68836 7284 68888 7293
rect 69112 7327 69164 7336
rect 69112 7293 69121 7327
rect 69121 7293 69155 7327
rect 69155 7293 69164 7327
rect 69112 7284 69164 7293
rect 70860 7284 70912 7336
rect 71228 7327 71280 7336
rect 71228 7293 71237 7327
rect 71237 7293 71271 7327
rect 71271 7293 71280 7327
rect 71228 7284 71280 7293
rect 72976 7284 73028 7336
rect 73344 7327 73396 7336
rect 73344 7293 73353 7327
rect 73353 7293 73387 7327
rect 73387 7293 73396 7327
rect 73344 7284 73396 7293
rect 75092 7284 75144 7336
rect 75460 7327 75512 7336
rect 75460 7293 75469 7327
rect 75469 7293 75503 7327
rect 75503 7293 75512 7327
rect 75460 7284 75512 7293
rect 77208 7284 77260 7336
rect 77576 7327 77628 7336
rect 77576 7293 77585 7327
rect 77585 7293 77619 7327
rect 77619 7293 77628 7327
rect 77576 7284 77628 7293
rect 79324 7284 79376 7336
rect 79692 7327 79744 7336
rect 79692 7293 79701 7327
rect 79701 7293 79735 7327
rect 79735 7293 79744 7327
rect 79692 7284 79744 7293
rect 81440 7284 81492 7336
rect 81808 7327 81860 7336
rect 81808 7293 81817 7327
rect 81817 7293 81851 7327
rect 81851 7293 81860 7327
rect 81808 7284 81860 7293
rect 83556 7284 83608 7336
rect 83924 7327 83976 7336
rect 83924 7293 83933 7327
rect 83933 7293 83967 7327
rect 83967 7293 83976 7327
rect 83924 7284 83976 7293
rect 85672 7284 85724 7336
rect 86040 7327 86092 7336
rect 86040 7293 86049 7327
rect 86049 7293 86083 7327
rect 86083 7293 86092 7327
rect 86040 7284 86092 7293
rect 87788 7284 87840 7336
rect 88156 7327 88208 7336
rect 88156 7293 88165 7327
rect 88165 7293 88199 7327
rect 88199 7293 88208 7327
rect 88156 7284 88208 7293
rect 89904 7284 89956 7336
rect 90272 7327 90324 7336
rect 90272 7293 90281 7327
rect 90281 7293 90315 7327
rect 90315 7293 90324 7327
rect 90272 7284 90324 7293
rect 92020 7284 92072 7336
rect 92388 7327 92440 7336
rect 92388 7293 92397 7327
rect 92397 7293 92431 7327
rect 92431 7293 92440 7327
rect 92388 7284 92440 7293
rect 94228 7327 94280 7336
rect 94228 7293 94237 7327
rect 94237 7293 94271 7327
rect 94271 7293 94280 7327
rect 94228 7284 94280 7293
rect 94504 7327 94556 7336
rect 94504 7293 94513 7327
rect 94513 7293 94547 7327
rect 94547 7293 94556 7327
rect 94504 7284 94556 7293
rect 96068 7284 96120 7336
rect 96620 7327 96672 7336
rect 96620 7293 96629 7327
rect 96629 7293 96663 7327
rect 96663 7293 96672 7327
rect 96620 7284 96672 7293
rect 98368 7284 98420 7336
rect 98736 7327 98788 7336
rect 98736 7293 98745 7327
rect 98745 7293 98779 7327
rect 98779 7293 98788 7327
rect 98736 7284 98788 7293
rect 100484 7284 100536 7336
rect 100852 7327 100904 7336
rect 100852 7293 100861 7327
rect 100861 7293 100895 7327
rect 100895 7293 100904 7327
rect 100852 7284 100904 7293
rect 102692 7327 102744 7336
rect 102692 7293 102701 7327
rect 102701 7293 102735 7327
rect 102735 7293 102744 7327
rect 102692 7284 102744 7293
rect 102968 7327 103020 7336
rect 102968 7293 102977 7327
rect 102977 7293 103011 7327
rect 103011 7293 103020 7327
rect 102968 7284 103020 7293
rect 104808 7327 104860 7336
rect 104808 7293 104817 7327
rect 104817 7293 104851 7327
rect 104851 7293 104860 7327
rect 104808 7284 104860 7293
rect 105084 7327 105136 7336
rect 105084 7293 105093 7327
rect 105093 7293 105127 7327
rect 105127 7293 105136 7327
rect 105084 7284 105136 7293
rect 11244 7259 11296 7268
rect 11244 7225 11253 7259
rect 11253 7225 11287 7259
rect 11287 7225 11296 7259
rect 11244 7216 11296 7225
rect 13360 7259 13412 7268
rect 13360 7225 13369 7259
rect 13369 7225 13403 7259
rect 13403 7225 13412 7259
rect 13360 7216 13412 7225
rect 23940 7259 23992 7268
rect 23940 7225 23949 7259
rect 23949 7225 23983 7259
rect 23983 7225 23992 7259
rect 23940 7216 23992 7225
rect 30288 7259 30340 7268
rect 30288 7225 30297 7259
rect 30297 7225 30331 7259
rect 30331 7225 30340 7259
rect 30288 7216 30340 7225
rect 47216 7259 47268 7268
rect 47216 7225 47225 7259
rect 47225 7225 47259 7259
rect 47259 7225 47268 7259
rect 47216 7216 47268 7225
rect 64144 7259 64196 7268
rect 64144 7225 64153 7259
rect 64153 7225 64187 7259
rect 64187 7225 64196 7259
rect 64144 7216 64196 7225
rect 78956 7259 79008 7268
rect 78956 7225 78965 7259
rect 78965 7225 78999 7259
rect 78999 7225 79008 7259
rect 78956 7216 79008 7225
rect 81348 7216 81400 7268
rect 95884 7259 95936 7268
rect 95884 7225 95893 7259
rect 95893 7225 95927 7259
rect 95927 7225 95936 7259
rect 95884 7216 95936 7225
rect 98092 7216 98144 7268
rect 2596 7148 2648 7200
rect 4528 7148 4580 7200
rect 6644 7148 6696 7200
rect 8944 7148 8996 7200
rect 15108 7148 15160 7200
rect 17224 7148 17276 7200
rect 19248 7148 19300 7200
rect 21456 7148 21508 7200
rect 25872 7148 25924 7200
rect 27988 7148 28040 7200
rect 32036 7148 32088 7200
rect 34152 7148 34204 7200
rect 36176 7148 36228 7200
rect 38384 7148 38436 7200
rect 40500 7148 40552 7200
rect 42892 7191 42944 7200
rect 42892 7157 42901 7191
rect 42901 7157 42935 7191
rect 42935 7157 42944 7191
rect 42892 7148 42944 7157
rect 44916 7148 44968 7200
rect 48964 7148 49016 7200
rect 51080 7148 51132 7200
rect 53288 7191 53340 7200
rect 53288 7157 53297 7191
rect 53297 7157 53331 7191
rect 53331 7157 53340 7191
rect 53288 7148 53340 7157
rect 55312 7148 55364 7200
rect 57428 7148 57480 7200
rect 59728 7148 59780 7200
rect 61844 7148 61896 7200
rect 65892 7148 65944 7200
rect 68008 7148 68060 7200
rect 70216 7191 70268 7200
rect 70216 7157 70225 7191
rect 70225 7157 70259 7191
rect 70259 7157 70268 7191
rect 70216 7148 70268 7157
rect 72240 7148 72292 7200
rect 74356 7148 74408 7200
rect 76656 7148 76708 7200
rect 82820 7148 82872 7200
rect 85120 7148 85172 7200
rect 87144 7191 87196 7200
rect 87144 7157 87153 7191
rect 87153 7157 87187 7191
rect 87187 7157 87196 7191
rect 87144 7148 87196 7157
rect 89168 7148 89220 7200
rect 91468 7148 91520 7200
rect 93584 7148 93636 7200
rect 99748 7148 99800 7200
rect 101864 7148 101916 7200
rect 103888 7148 103940 7200
rect 106188 7191 106240 7200
rect 106188 7157 106197 7191
rect 106197 7157 106231 7191
rect 106231 7157 106240 7191
rect 106188 7148 106240 7157
rect 19402 7046 19454 7098
rect 19466 7046 19518 7098
rect 19530 7046 19582 7098
rect 19594 7046 19646 7098
rect 50122 7046 50174 7098
rect 50186 7046 50238 7098
rect 50250 7046 50302 7098
rect 50314 7046 50366 7098
rect 80842 7046 80894 7098
rect 80906 7046 80958 7098
rect 80970 7046 81022 7098
rect 81034 7046 81086 7098
rect 3516 6944 3568 6996
rect 5632 6944 5684 6996
rect 7748 6944 7800 6996
rect 9864 6944 9916 6996
rect 11980 6944 12032 6996
rect 14096 6944 14148 6996
rect 16212 6944 16264 6996
rect 18328 6944 18380 6996
rect 20444 6944 20496 6996
rect 22560 6944 22612 6996
rect 24676 6944 24728 6996
rect 26792 6944 26844 6996
rect 28908 6944 28960 6996
rect 31024 6944 31076 6996
rect 33140 6944 33192 6996
rect 35256 6944 35308 6996
rect 37372 6944 37424 6996
rect 39488 6944 39540 6996
rect 41604 6944 41656 6996
rect 43720 6944 43772 6996
rect 45836 6944 45888 6996
rect 47952 6944 48004 6996
rect 51172 6987 51224 6996
rect 51172 6953 51181 6987
rect 51181 6953 51215 6987
rect 51215 6953 51224 6987
rect 51172 6944 51224 6953
rect 52184 6944 52236 6996
rect 54300 6944 54352 6996
rect 56416 6944 56468 6996
rect 58532 6944 58584 6996
rect 60648 6944 60700 6996
rect 62764 6944 62816 6996
rect 64880 6944 64932 6996
rect 66996 6944 67048 6996
rect 69112 6944 69164 6996
rect 71228 6944 71280 6996
rect 73344 6944 73396 6996
rect 75460 6944 75512 6996
rect 77576 6944 77628 6996
rect 79692 6944 79744 6996
rect 81808 6944 81860 6996
rect 83924 6944 83976 6996
rect 86040 6944 86092 6996
rect 88156 6944 88208 6996
rect 90272 6944 90324 6996
rect 92388 6944 92440 6996
rect 94504 6944 94556 6996
rect 96620 6944 96672 6996
rect 98736 6944 98788 6996
rect 100852 6944 100904 6996
rect 102968 6944 103020 6996
rect 105084 6944 105136 6996
rect 1124 6851 1176 6860
rect 1124 6817 1133 6851
rect 1133 6817 1167 6851
rect 1167 6817 1176 6851
rect 1124 6808 1176 6817
rect 3240 6851 3292 6860
rect 3240 6817 3249 6851
rect 3249 6817 3283 6851
rect 3283 6817 3292 6851
rect 3240 6808 3292 6817
rect 5264 6808 5316 6860
rect 7380 6808 7432 6860
rect 9588 6851 9640 6860
rect 9588 6817 9597 6851
rect 9597 6817 9631 6851
rect 9631 6817 9640 6851
rect 9588 6808 9640 6817
rect 11704 6851 11756 6860
rect 11704 6817 11713 6851
rect 11713 6817 11747 6851
rect 11747 6817 11756 6851
rect 11704 6808 11756 6817
rect 13820 6851 13872 6860
rect 13820 6817 13829 6851
rect 13829 6817 13863 6851
rect 13863 6817 13872 6851
rect 13820 6808 13872 6817
rect 15936 6851 15988 6860
rect 15936 6817 15945 6851
rect 15945 6817 15979 6851
rect 15979 6817 15988 6851
rect 15936 6808 15988 6817
rect 18052 6851 18104 6860
rect 18052 6817 18061 6851
rect 18061 6817 18095 6851
rect 18095 6817 18104 6851
rect 18052 6808 18104 6817
rect 20076 6808 20128 6860
rect 22192 6808 22244 6860
rect 24400 6851 24452 6860
rect 24400 6817 24409 6851
rect 24409 6817 24443 6851
rect 24443 6817 24452 6851
rect 24400 6808 24452 6817
rect 26516 6851 26568 6860
rect 26516 6817 26525 6851
rect 26525 6817 26559 6851
rect 26559 6817 26568 6851
rect 26516 6808 26568 6817
rect 28632 6851 28684 6860
rect 28632 6817 28641 6851
rect 28641 6817 28675 6851
rect 28675 6817 28684 6851
rect 28632 6808 28684 6817
rect 30748 6851 30800 6860
rect 30748 6817 30757 6851
rect 30757 6817 30791 6851
rect 30791 6817 30800 6851
rect 30748 6808 30800 6817
rect 32864 6851 32916 6860
rect 32864 6817 32873 6851
rect 32873 6817 32907 6851
rect 32907 6817 32916 6851
rect 32864 6808 32916 6817
rect 35072 6808 35124 6860
rect 37096 6851 37148 6860
rect 37096 6817 37105 6851
rect 37105 6817 37139 6851
rect 37139 6817 37148 6851
rect 37096 6808 37148 6817
rect 39212 6851 39264 6860
rect 39212 6817 39221 6851
rect 39221 6817 39255 6851
rect 39255 6817 39264 6851
rect 39212 6808 39264 6817
rect 41236 6808 41288 6860
rect 43444 6851 43496 6860
rect 43444 6817 43453 6851
rect 43453 6817 43487 6851
rect 43487 6817 43496 6851
rect 43444 6808 43496 6817
rect 45560 6851 45612 6860
rect 45560 6817 45569 6851
rect 45569 6817 45603 6851
rect 45603 6817 45612 6851
rect 45560 6808 45612 6817
rect 47676 6851 47728 6860
rect 47676 6817 47685 6851
rect 47685 6817 47719 6851
rect 47719 6817 47728 6851
rect 47676 6808 47728 6817
rect 49792 6851 49844 6860
rect 49792 6817 49801 6851
rect 49801 6817 49835 6851
rect 49835 6817 49844 6851
rect 49792 6808 49844 6817
rect 51908 6851 51960 6860
rect 51908 6817 51917 6851
rect 51917 6817 51951 6851
rect 51951 6817 51960 6851
rect 51908 6808 51960 6817
rect 54024 6851 54076 6860
rect 54024 6817 54033 6851
rect 54033 6817 54067 6851
rect 54067 6817 54076 6851
rect 54024 6808 54076 6817
rect 56048 6808 56100 6860
rect 58164 6808 58216 6860
rect 62488 6851 62540 6860
rect 62488 6817 62497 6851
rect 62497 6817 62531 6851
rect 62531 6817 62540 6851
rect 62488 6808 62540 6817
rect 64604 6851 64656 6860
rect 64604 6817 64613 6851
rect 64613 6817 64647 6851
rect 64647 6817 64656 6851
rect 64604 6808 64656 6817
rect 66720 6851 66772 6860
rect 66720 6817 66729 6851
rect 66729 6817 66763 6851
rect 66763 6817 66772 6851
rect 66720 6808 66772 6817
rect 68836 6851 68888 6860
rect 68836 6817 68845 6851
rect 68845 6817 68879 6851
rect 68879 6817 68888 6851
rect 68836 6808 68888 6817
rect 70860 6808 70912 6860
rect 72976 6808 73028 6860
rect 75092 6808 75144 6860
rect 79324 6808 79376 6860
rect 81440 6808 81492 6860
rect 83556 6808 83608 6860
rect 85672 6808 85724 6860
rect 87788 6808 87840 6860
rect 89904 6808 89956 6860
rect 92020 6808 92072 6860
rect 94228 6851 94280 6860
rect 94228 6817 94237 6851
rect 94237 6817 94271 6851
rect 94271 6817 94280 6851
rect 94228 6808 94280 6817
rect 96068 6808 96120 6860
rect 98368 6808 98420 6860
rect 100484 6808 100536 6860
rect 102692 6851 102744 6860
rect 102692 6817 102701 6851
rect 102701 6817 102735 6851
rect 102735 6817 102744 6851
rect 102692 6808 102744 6817
rect 104808 6851 104860 6860
rect 104808 6817 104817 6851
rect 104817 6817 104851 6851
rect 104851 6817 104860 6851
rect 104808 6808 104860 6817
rect 2136 6740 2188 6792
rect 3516 6783 3568 6792
rect 3516 6749 3525 6783
rect 3525 6749 3559 6783
rect 3559 6749 3568 6783
rect 3516 6740 3568 6749
rect 5632 6783 5684 6792
rect 5632 6749 5641 6783
rect 5641 6749 5675 6783
rect 5675 6749 5684 6783
rect 5632 6740 5684 6749
rect 7748 6783 7800 6792
rect 7748 6749 7757 6783
rect 7757 6749 7791 6783
rect 7791 6749 7800 6783
rect 7748 6740 7800 6749
rect 9864 6783 9916 6792
rect 9864 6749 9873 6783
rect 9873 6749 9907 6783
rect 9907 6749 9916 6783
rect 9864 6740 9916 6749
rect 11980 6783 12032 6792
rect 11980 6749 11989 6783
rect 11989 6749 12023 6783
rect 12023 6749 12032 6783
rect 11980 6740 12032 6749
rect 14096 6783 14148 6792
rect 14096 6749 14105 6783
rect 14105 6749 14139 6783
rect 14139 6749 14148 6783
rect 14096 6740 14148 6749
rect 16212 6783 16264 6792
rect 16212 6749 16221 6783
rect 16221 6749 16255 6783
rect 16255 6749 16264 6783
rect 16212 6740 16264 6749
rect 18328 6783 18380 6792
rect 18328 6749 18337 6783
rect 18337 6749 18371 6783
rect 18371 6749 18380 6783
rect 18328 6740 18380 6749
rect 20444 6783 20496 6792
rect 20444 6749 20453 6783
rect 20453 6749 20487 6783
rect 20487 6749 20496 6783
rect 20444 6740 20496 6749
rect 22560 6783 22612 6792
rect 22560 6749 22569 6783
rect 22569 6749 22603 6783
rect 22603 6749 22612 6783
rect 22560 6740 22612 6749
rect 24676 6783 24728 6792
rect 24676 6749 24685 6783
rect 24685 6749 24719 6783
rect 24719 6749 24728 6783
rect 24676 6740 24728 6749
rect 26792 6783 26844 6792
rect 26792 6749 26801 6783
rect 26801 6749 26835 6783
rect 26835 6749 26844 6783
rect 26792 6740 26844 6749
rect 28908 6783 28960 6792
rect 28908 6749 28917 6783
rect 28917 6749 28951 6783
rect 28951 6749 28960 6783
rect 28908 6740 28960 6749
rect 31024 6783 31076 6792
rect 31024 6749 31033 6783
rect 31033 6749 31067 6783
rect 31067 6749 31076 6783
rect 31024 6740 31076 6749
rect 33140 6783 33192 6792
rect 33140 6749 33149 6783
rect 33149 6749 33183 6783
rect 33183 6749 33192 6783
rect 33140 6740 33192 6749
rect 35256 6783 35308 6792
rect 35256 6749 35265 6783
rect 35265 6749 35299 6783
rect 35299 6749 35308 6783
rect 35256 6740 35308 6749
rect 37372 6783 37424 6792
rect 37372 6749 37381 6783
rect 37381 6749 37415 6783
rect 37415 6749 37424 6783
rect 37372 6740 37424 6749
rect 39396 6740 39448 6792
rect 41604 6783 41656 6792
rect 41604 6749 41613 6783
rect 41613 6749 41647 6783
rect 41647 6749 41656 6783
rect 41604 6740 41656 6749
rect 43720 6783 43772 6792
rect 43720 6749 43729 6783
rect 43729 6749 43763 6783
rect 43763 6749 43772 6783
rect 43720 6740 43772 6749
rect 45836 6783 45888 6792
rect 45836 6749 45845 6783
rect 45845 6749 45879 6783
rect 45879 6749 45888 6783
rect 45836 6740 45888 6749
rect 47952 6783 48004 6792
rect 47952 6749 47961 6783
rect 47961 6749 47995 6783
rect 47995 6749 48004 6783
rect 47952 6740 48004 6749
rect 50068 6783 50120 6792
rect 50068 6749 50077 6783
rect 50077 6749 50111 6783
rect 50111 6749 50120 6783
rect 52184 6783 52236 6792
rect 50068 6740 50120 6749
rect 52184 6749 52193 6783
rect 52193 6749 52227 6783
rect 52227 6749 52236 6783
rect 52184 6740 52236 6749
rect 54300 6783 54352 6792
rect 54300 6749 54309 6783
rect 54309 6749 54343 6783
rect 54343 6749 54352 6783
rect 54300 6740 54352 6749
rect 56416 6783 56468 6792
rect 56416 6749 56425 6783
rect 56425 6749 56459 6783
rect 56459 6749 56468 6783
rect 56416 6740 56468 6749
rect 58532 6783 58584 6792
rect 58532 6749 58541 6783
rect 58541 6749 58575 6783
rect 58575 6749 58584 6783
rect 58532 6740 58584 6749
rect 60372 6783 60424 6792
rect 60372 6749 60381 6783
rect 60381 6749 60415 6783
rect 60415 6749 60424 6783
rect 60648 6783 60700 6792
rect 60372 6740 60424 6749
rect 60648 6749 60657 6783
rect 60657 6749 60691 6783
rect 60691 6749 60700 6783
rect 60648 6740 60700 6749
rect 62764 6783 62816 6792
rect 62764 6749 62773 6783
rect 62773 6749 62807 6783
rect 62807 6749 62816 6783
rect 62764 6740 62816 6749
rect 64880 6783 64932 6792
rect 64880 6749 64889 6783
rect 64889 6749 64923 6783
rect 64923 6749 64932 6783
rect 64880 6740 64932 6749
rect 66996 6783 67048 6792
rect 66996 6749 67005 6783
rect 67005 6749 67039 6783
rect 67039 6749 67048 6783
rect 66996 6740 67048 6749
rect 69112 6783 69164 6792
rect 69112 6749 69121 6783
rect 69121 6749 69155 6783
rect 69155 6749 69164 6783
rect 69112 6740 69164 6749
rect 71228 6783 71280 6792
rect 71228 6749 71237 6783
rect 71237 6749 71271 6783
rect 71271 6749 71280 6783
rect 71228 6740 71280 6749
rect 73344 6783 73396 6792
rect 73344 6749 73353 6783
rect 73353 6749 73387 6783
rect 73387 6749 73396 6783
rect 73344 6740 73396 6749
rect 75368 6740 75420 6792
rect 77300 6783 77352 6792
rect 77300 6749 77309 6783
rect 77309 6749 77343 6783
rect 77343 6749 77352 6783
rect 77300 6740 77352 6749
rect 77576 6783 77628 6792
rect 77576 6749 77585 6783
rect 77585 6749 77619 6783
rect 77619 6749 77628 6783
rect 77576 6740 77628 6749
rect 79692 6783 79744 6792
rect 79692 6749 79701 6783
rect 79701 6749 79735 6783
rect 79735 6749 79744 6783
rect 79692 6740 79744 6749
rect 81808 6783 81860 6792
rect 81808 6749 81817 6783
rect 81817 6749 81851 6783
rect 81851 6749 81860 6783
rect 81808 6740 81860 6749
rect 83924 6783 83976 6792
rect 83924 6749 83933 6783
rect 83933 6749 83967 6783
rect 83967 6749 83976 6783
rect 83924 6740 83976 6749
rect 85948 6740 86000 6792
rect 88156 6783 88208 6792
rect 88156 6749 88165 6783
rect 88165 6749 88199 6783
rect 88199 6749 88208 6783
rect 88156 6740 88208 6749
rect 90272 6783 90324 6792
rect 90272 6749 90281 6783
rect 90281 6749 90315 6783
rect 90315 6749 90324 6783
rect 90272 6740 90324 6749
rect 92388 6783 92440 6792
rect 92388 6749 92397 6783
rect 92397 6749 92431 6783
rect 92431 6749 92440 6783
rect 92388 6740 92440 6749
rect 94504 6783 94556 6792
rect 94504 6749 94513 6783
rect 94513 6749 94547 6783
rect 94547 6749 94556 6783
rect 94504 6740 94556 6749
rect 96620 6783 96672 6792
rect 96620 6749 96629 6783
rect 96629 6749 96663 6783
rect 96663 6749 96672 6783
rect 96620 6740 96672 6749
rect 98736 6783 98788 6792
rect 98736 6749 98745 6783
rect 98745 6749 98779 6783
rect 98779 6749 98788 6783
rect 98736 6740 98788 6749
rect 100852 6783 100904 6792
rect 100852 6749 100861 6783
rect 100861 6749 100895 6783
rect 100895 6749 100904 6783
rect 100852 6740 100904 6749
rect 102968 6783 103020 6792
rect 102968 6749 102977 6783
rect 102977 6749 103011 6783
rect 103011 6749 103020 6783
rect 102968 6740 103020 6749
rect 105084 6783 105136 6792
rect 105084 6749 105093 6783
rect 105093 6749 105127 6783
rect 105127 6749 105136 6783
rect 105084 6740 105136 6749
rect 4042 6502 4094 6554
rect 4106 6502 4158 6554
rect 4170 6502 4222 6554
rect 4234 6502 4286 6554
rect 34762 6502 34814 6554
rect 34826 6502 34878 6554
rect 34890 6502 34942 6554
rect 34954 6502 35006 6554
rect 65482 6502 65534 6554
rect 65546 6502 65598 6554
rect 65610 6502 65662 6554
rect 65674 6502 65726 6554
rect 96202 6502 96254 6554
rect 96266 6502 96318 6554
rect 96330 6502 96382 6554
rect 96394 6502 96446 6554
rect 2136 6332 2188 6384
rect 3516 6196 3568 6248
rect 5632 6196 5684 6248
rect 7748 6196 7800 6248
rect 9864 6196 9916 6248
rect 11980 6196 12032 6248
rect 14096 6196 14148 6248
rect 16212 6196 16264 6248
rect 18328 6196 18380 6248
rect 20444 6196 20496 6248
rect 22560 6196 22612 6248
rect 24676 6196 24728 6248
rect 26792 6196 26844 6248
rect 28908 6196 28960 6248
rect 31024 6196 31076 6248
rect 33140 6196 33192 6248
rect 35256 6196 35308 6248
rect 37372 6196 37424 6248
rect 41604 6196 41656 6248
rect 43720 6196 43772 6248
rect 45836 6196 45888 6248
rect 47952 6196 48004 6248
rect 39396 6171 39448 6180
rect 39396 6137 39405 6171
rect 39405 6137 39439 6171
rect 39439 6137 39448 6171
rect 39396 6128 39448 6137
rect 52184 6196 52236 6248
rect 54300 6196 54352 6248
rect 56416 6196 56468 6248
rect 58532 6196 58584 6248
rect 60648 6196 60700 6248
rect 62764 6196 62816 6248
rect 64880 6196 64932 6248
rect 66996 6196 67048 6248
rect 69112 6196 69164 6248
rect 71228 6196 71280 6248
rect 73344 6196 73396 6248
rect 77576 6196 77628 6248
rect 79692 6196 79744 6248
rect 81808 6196 81860 6248
rect 83924 6196 83976 6248
rect 88156 6196 88208 6248
rect 90272 6196 90324 6248
rect 92388 6196 92440 6248
rect 94504 6196 94556 6248
rect 96620 6196 96672 6248
rect 98736 6196 98788 6248
rect 100852 6196 100904 6248
rect 102968 6196 103020 6248
rect 105084 6196 105136 6248
rect 50068 6128 50120 6180
rect 75368 6171 75420 6180
rect 75368 6137 75377 6171
rect 75377 6137 75411 6171
rect 75411 6137 75420 6171
rect 75368 6128 75420 6137
rect 85948 6171 86000 6180
rect 85948 6137 85957 6171
rect 85957 6137 85991 6171
rect 85991 6137 86000 6171
rect 85948 6128 86000 6137
rect 19402 5958 19454 6010
rect 19466 5958 19518 6010
rect 19530 5958 19582 6010
rect 19594 5958 19646 6010
rect 50122 5958 50174 6010
rect 50186 5958 50238 6010
rect 50250 5958 50302 6010
rect 50314 5958 50366 6010
rect 80842 5958 80894 6010
rect 80906 5958 80958 6010
rect 80970 5958 81022 6010
rect 81034 5958 81086 6010
rect 11888 5788 11940 5840
rect 14096 5788 14148 5840
rect 22376 5831 22428 5840
rect 22376 5797 22385 5831
rect 22385 5797 22419 5831
rect 22419 5797 22428 5831
rect 22376 5788 22428 5797
rect 24676 5788 24728 5840
rect 33048 5788 33100 5840
rect 37372 5788 37424 5840
rect 43720 5788 43772 5840
rect 47860 5788 47912 5840
rect 58440 5788 58492 5840
rect 60464 5831 60516 5840
rect 60464 5797 60473 5831
rect 60473 5797 60507 5831
rect 60507 5797 60516 5831
rect 60464 5788 60516 5797
rect 62764 5788 62816 5840
rect 73344 5788 73396 5840
rect 1308 5720 1360 5772
rect 3516 5720 3568 5772
rect 7656 5720 7708 5772
rect 9864 5652 9916 5704
rect 16212 5720 16264 5772
rect 5632 5584 5684 5636
rect 20444 5720 20496 5772
rect 26700 5652 26752 5704
rect 31024 5720 31076 5772
rect 35256 5720 35308 5772
rect 28816 5652 28868 5704
rect 39488 5652 39540 5704
rect 50068 5720 50120 5772
rect 45836 5652 45888 5704
rect 18328 5584 18380 5636
rect 54208 5720 54260 5772
rect 56416 5652 56468 5704
rect 64788 5720 64840 5772
rect 66996 5720 67048 5772
rect 52184 5584 52236 5636
rect 71228 5720 71280 5772
rect 75460 5652 75512 5704
rect 69112 5584 69164 5636
rect 41604 5516 41656 5568
rect 79600 5788 79652 5840
rect 83924 5788 83976 5840
rect 90272 5788 90324 5840
rect 94412 5788 94464 5840
rect 96436 5831 96488 5840
rect 96436 5797 96445 5831
rect 96445 5797 96479 5831
rect 96479 5797 96488 5831
rect 96436 5788 96488 5797
rect 105084 5831 105136 5840
rect 81808 5720 81860 5772
rect 86040 5720 86092 5772
rect 98644 5720 98696 5772
rect 92388 5652 92440 5704
rect 100760 5720 100812 5772
rect 102968 5720 103020 5772
rect 105084 5797 105093 5831
rect 105093 5797 105127 5831
rect 105127 5797 105136 5831
rect 105084 5788 105136 5797
rect 104992 5720 105044 5772
rect 77576 5516 77628 5568
rect 88156 5516 88208 5568
rect 4042 5414 4094 5466
rect 4106 5414 4158 5466
rect 4170 5414 4222 5466
rect 4234 5414 4286 5466
rect 34762 5414 34814 5466
rect 34826 5414 34878 5466
rect 34890 5414 34942 5466
rect 34954 5414 35006 5466
rect 65482 5414 65534 5466
rect 65546 5414 65598 5466
rect 65610 5414 65662 5466
rect 65674 5414 65726 5466
rect 96202 5414 96254 5466
rect 96266 5414 96318 5466
rect 96330 5414 96382 5466
rect 96394 5414 96446 5466
rect 1124 5219 1176 5228
rect 1124 5185 1133 5219
rect 1133 5185 1167 5219
rect 1167 5185 1176 5219
rect 1124 5176 1176 5185
rect 1308 5176 1360 5228
rect 3240 5219 3292 5228
rect 3240 5185 3249 5219
rect 3249 5185 3283 5219
rect 3283 5185 3292 5219
rect 3240 5176 3292 5185
rect 3516 5219 3568 5228
rect 3516 5185 3525 5219
rect 3525 5185 3559 5219
rect 3559 5185 3568 5219
rect 3516 5176 3568 5185
rect 5264 5176 5316 5228
rect 5632 5219 5684 5228
rect 5632 5185 5641 5219
rect 5641 5185 5675 5219
rect 5675 5185 5684 5219
rect 5632 5176 5684 5185
rect 7380 5176 7432 5228
rect 7656 5176 7708 5228
rect 9588 5219 9640 5228
rect 9588 5185 9597 5219
rect 9597 5185 9631 5219
rect 9631 5185 9640 5219
rect 9588 5176 9640 5185
rect 9864 5219 9916 5228
rect 9864 5185 9873 5219
rect 9873 5185 9907 5219
rect 9907 5185 9916 5219
rect 9864 5176 9916 5185
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 11888 5176 11940 5228
rect 13820 5219 13872 5228
rect 13820 5185 13829 5219
rect 13829 5185 13863 5219
rect 13863 5185 13872 5219
rect 13820 5176 13872 5185
rect 14096 5219 14148 5228
rect 14096 5185 14105 5219
rect 14105 5185 14139 5219
rect 14139 5185 14148 5219
rect 14096 5176 14148 5185
rect 15936 5219 15988 5228
rect 15936 5185 15945 5219
rect 15945 5185 15979 5219
rect 15979 5185 15988 5219
rect 15936 5176 15988 5185
rect 16212 5219 16264 5228
rect 16212 5185 16221 5219
rect 16221 5185 16255 5219
rect 16255 5185 16264 5219
rect 16212 5176 16264 5185
rect 18052 5219 18104 5228
rect 18052 5185 18061 5219
rect 18061 5185 18095 5219
rect 18095 5185 18104 5219
rect 18052 5176 18104 5185
rect 18328 5219 18380 5228
rect 18328 5185 18337 5219
rect 18337 5185 18371 5219
rect 18371 5185 18380 5219
rect 18328 5176 18380 5185
rect 20076 5176 20128 5228
rect 20444 5219 20496 5228
rect 20444 5185 20453 5219
rect 20453 5185 20487 5219
rect 20487 5185 20496 5219
rect 20444 5176 20496 5185
rect 22192 5176 22244 5228
rect 22468 5176 22520 5228
rect 23756 5176 23808 5228
rect 23940 5176 23992 5228
rect 24400 5219 24452 5228
rect 24400 5185 24409 5219
rect 24409 5185 24443 5219
rect 24443 5185 24452 5219
rect 24400 5176 24452 5185
rect 24676 5219 24728 5228
rect 24676 5185 24685 5219
rect 24685 5185 24719 5219
rect 24719 5185 24728 5219
rect 24676 5176 24728 5185
rect 26516 5219 26568 5228
rect 26516 5185 26525 5219
rect 26525 5185 26559 5219
rect 26559 5185 26568 5219
rect 26516 5176 26568 5185
rect 26700 5176 26752 5228
rect 28632 5219 28684 5228
rect 28632 5185 28641 5219
rect 28641 5185 28675 5219
rect 28675 5185 28684 5219
rect 28632 5176 28684 5185
rect 28816 5176 28868 5228
rect 30748 5219 30800 5228
rect 30748 5185 30757 5219
rect 30757 5185 30791 5219
rect 30791 5185 30800 5219
rect 30748 5176 30800 5185
rect 31024 5219 31076 5228
rect 31024 5185 31033 5219
rect 31033 5185 31067 5219
rect 31067 5185 31076 5219
rect 31024 5176 31076 5185
rect 32864 5219 32916 5228
rect 32864 5185 32873 5219
rect 32873 5185 32907 5219
rect 32907 5185 32916 5219
rect 32864 5176 32916 5185
rect 33048 5176 33100 5228
rect 35256 5219 35308 5228
rect 35256 5185 35265 5219
rect 35265 5185 35299 5219
rect 35299 5185 35308 5219
rect 35256 5176 35308 5185
rect 37096 5219 37148 5228
rect 37096 5185 37105 5219
rect 37105 5185 37139 5219
rect 37139 5185 37148 5219
rect 37096 5176 37148 5185
rect 37372 5219 37424 5228
rect 37372 5185 37381 5219
rect 37381 5185 37415 5219
rect 37415 5185 37424 5219
rect 37372 5176 37424 5185
rect 39212 5219 39264 5228
rect 39212 5185 39221 5219
rect 39221 5185 39255 5219
rect 39255 5185 39264 5219
rect 39212 5176 39264 5185
rect 39488 5219 39540 5228
rect 39488 5185 39497 5219
rect 39497 5185 39531 5219
rect 39531 5185 39540 5219
rect 39488 5176 39540 5185
rect 41236 5176 41288 5228
rect 41604 5219 41656 5228
rect 41604 5185 41613 5219
rect 41613 5185 41647 5219
rect 41647 5185 41656 5219
rect 41604 5176 41656 5185
rect 43444 5219 43496 5228
rect 43444 5185 43453 5219
rect 43453 5185 43487 5219
rect 43487 5185 43496 5219
rect 43444 5176 43496 5185
rect 43720 5219 43772 5228
rect 43720 5185 43729 5219
rect 43729 5185 43763 5219
rect 43763 5185 43772 5219
rect 43720 5176 43772 5185
rect 45560 5219 45612 5228
rect 45560 5185 45569 5219
rect 45569 5185 45603 5219
rect 45603 5185 45612 5219
rect 45560 5176 45612 5185
rect 45836 5219 45888 5228
rect 45836 5185 45845 5219
rect 45845 5185 45879 5219
rect 45879 5185 45888 5219
rect 45836 5176 45888 5185
rect 47676 5219 47728 5228
rect 47676 5185 47685 5219
rect 47685 5185 47719 5219
rect 47719 5185 47728 5219
rect 47676 5176 47728 5185
rect 47860 5176 47912 5228
rect 49792 5219 49844 5228
rect 49792 5185 49801 5219
rect 49801 5185 49835 5219
rect 49835 5185 49844 5219
rect 49792 5176 49844 5185
rect 50068 5219 50120 5228
rect 50068 5185 50077 5219
rect 50077 5185 50111 5219
rect 50111 5185 50120 5219
rect 51908 5219 51960 5228
rect 50068 5176 50120 5185
rect 51908 5185 51917 5219
rect 51917 5185 51951 5219
rect 51951 5185 51960 5219
rect 51908 5176 51960 5185
rect 52184 5219 52236 5228
rect 52184 5185 52193 5219
rect 52193 5185 52227 5219
rect 52227 5185 52236 5219
rect 52184 5176 52236 5185
rect 54024 5219 54076 5228
rect 54024 5185 54033 5219
rect 54033 5185 54067 5219
rect 54067 5185 54076 5219
rect 54024 5176 54076 5185
rect 54208 5176 54260 5228
rect 56048 5176 56100 5228
rect 56416 5219 56468 5228
rect 56416 5185 56425 5219
rect 56425 5185 56459 5219
rect 56459 5185 56468 5219
rect 56416 5176 56468 5185
rect 58164 5176 58216 5228
rect 58440 5176 58492 5228
rect 60556 5176 60608 5228
rect 62488 5219 62540 5228
rect 62488 5185 62497 5219
rect 62497 5185 62531 5219
rect 62531 5185 62540 5219
rect 62488 5176 62540 5185
rect 62764 5219 62816 5228
rect 62764 5185 62773 5219
rect 62773 5185 62807 5219
rect 62807 5185 62816 5219
rect 62764 5176 62816 5185
rect 64604 5219 64656 5228
rect 64604 5185 64613 5219
rect 64613 5185 64647 5219
rect 64647 5185 64656 5219
rect 64604 5176 64656 5185
rect 64788 5176 64840 5228
rect 66720 5219 66772 5228
rect 66720 5185 66729 5219
rect 66729 5185 66763 5219
rect 66763 5185 66772 5219
rect 66720 5176 66772 5185
rect 66996 5219 67048 5228
rect 66996 5185 67005 5219
rect 67005 5185 67039 5219
rect 67039 5185 67048 5219
rect 66996 5176 67048 5185
rect 68836 5219 68888 5228
rect 68836 5185 68845 5219
rect 68845 5185 68879 5219
rect 68879 5185 68888 5219
rect 68836 5176 68888 5185
rect 69112 5219 69164 5228
rect 69112 5185 69121 5219
rect 69121 5185 69155 5219
rect 69155 5185 69164 5219
rect 69112 5176 69164 5185
rect 70860 5176 70912 5228
rect 71228 5219 71280 5228
rect 71228 5185 71237 5219
rect 71237 5185 71271 5219
rect 71271 5185 71280 5219
rect 71228 5176 71280 5185
rect 72976 5176 73028 5228
rect 73344 5219 73396 5228
rect 73344 5185 73353 5219
rect 73353 5185 73387 5219
rect 73387 5185 73396 5219
rect 73344 5176 73396 5185
rect 75092 5176 75144 5228
rect 75460 5219 75512 5228
rect 75460 5185 75469 5219
rect 75469 5185 75503 5219
rect 75503 5185 75512 5219
rect 75460 5176 75512 5185
rect 77576 5219 77628 5228
rect 77576 5185 77585 5219
rect 77585 5185 77619 5219
rect 77619 5185 77628 5219
rect 77576 5176 77628 5185
rect 79324 5176 79376 5228
rect 79600 5176 79652 5228
rect 81440 5176 81492 5228
rect 81808 5219 81860 5228
rect 81808 5185 81817 5219
rect 81817 5185 81851 5219
rect 81851 5185 81860 5219
rect 81808 5176 81860 5185
rect 83556 5176 83608 5228
rect 83924 5219 83976 5228
rect 83924 5185 83933 5219
rect 83933 5185 83967 5219
rect 83967 5185 83976 5219
rect 83924 5176 83976 5185
rect 85672 5176 85724 5228
rect 86040 5219 86092 5228
rect 86040 5185 86049 5219
rect 86049 5185 86083 5219
rect 86083 5185 86092 5219
rect 86040 5176 86092 5185
rect 87788 5176 87840 5228
rect 88156 5219 88208 5228
rect 88156 5185 88165 5219
rect 88165 5185 88199 5219
rect 88199 5185 88208 5219
rect 88156 5176 88208 5185
rect 89904 5176 89956 5228
rect 90272 5219 90324 5228
rect 90272 5185 90281 5219
rect 90281 5185 90315 5219
rect 90315 5185 90324 5219
rect 90272 5176 90324 5185
rect 92020 5176 92072 5228
rect 92388 5219 92440 5228
rect 92388 5185 92397 5219
rect 92397 5185 92431 5219
rect 92431 5185 92440 5219
rect 92388 5176 92440 5185
rect 94228 5219 94280 5228
rect 94228 5185 94237 5219
rect 94237 5185 94271 5219
rect 94271 5185 94280 5219
rect 94228 5176 94280 5185
rect 94412 5176 94464 5228
rect 96068 5176 96120 5228
rect 96528 5176 96580 5228
rect 98368 5176 98420 5228
rect 98644 5176 98696 5228
rect 100484 5176 100536 5228
rect 100760 5176 100812 5228
rect 102692 5219 102744 5228
rect 102692 5185 102701 5219
rect 102701 5185 102735 5219
rect 102735 5185 102744 5219
rect 102692 5176 102744 5185
rect 102968 5219 103020 5228
rect 102968 5185 102977 5219
rect 102977 5185 103011 5219
rect 103011 5185 103020 5219
rect 102968 5176 103020 5185
rect 104808 5219 104860 5228
rect 104808 5185 104817 5219
rect 104817 5185 104851 5219
rect 104851 5185 104860 5219
rect 104808 5176 104860 5185
rect 104992 5176 105044 5228
rect 35072 5108 35124 5160
rect 60372 5151 60424 5160
rect 60372 5117 60381 5151
rect 60381 5117 60415 5151
rect 60415 5117 60424 5151
rect 60372 5108 60424 5117
rect 77300 5151 77352 5160
rect 77300 5117 77309 5151
rect 77309 5117 77343 5151
rect 77343 5117 77352 5151
rect 77300 5108 77352 5117
rect 3516 4972 3568 5024
rect 5632 4972 5684 5024
rect 7748 4972 7800 5024
rect 9864 4972 9916 5024
rect 11980 4972 12032 5024
rect 14096 4972 14148 5024
rect 16212 4972 16264 5024
rect 18328 4972 18380 5024
rect 20444 4972 20496 5024
rect 22560 4972 22612 5024
rect 24676 4972 24728 5024
rect 26792 4972 26844 5024
rect 28908 4972 28960 5024
rect 31024 4972 31076 5024
rect 33140 4972 33192 5024
rect 35256 4972 35308 5024
rect 37372 4972 37424 5024
rect 39488 4972 39540 5024
rect 41604 4972 41656 5024
rect 43720 4972 43772 5024
rect 45836 4972 45888 5024
rect 47952 4972 48004 5024
rect 51172 5015 51224 5024
rect 51172 4981 51181 5015
rect 51181 4981 51215 5015
rect 51215 4981 51224 5015
rect 51172 4972 51224 4981
rect 52184 4972 52236 5024
rect 54300 4972 54352 5024
rect 56416 4972 56468 5024
rect 58532 4972 58584 5024
rect 60648 4972 60700 5024
rect 62764 4972 62816 5024
rect 64880 4972 64932 5024
rect 66996 4972 67048 5024
rect 69112 4972 69164 5024
rect 71228 4972 71280 5024
rect 73344 4972 73396 5024
rect 75460 4972 75512 5024
rect 77576 4972 77628 5024
rect 79692 4972 79744 5024
rect 81808 4972 81860 5024
rect 83924 4972 83976 5024
rect 86040 4972 86092 5024
rect 88156 4972 88208 5024
rect 90272 4972 90324 5024
rect 92388 4972 92440 5024
rect 94504 4972 94556 5024
rect 96620 4972 96672 5024
rect 98736 4972 98788 5024
rect 100852 4972 100904 5024
rect 102968 4972 103020 5024
rect 105084 4972 105136 5024
rect 19402 4870 19454 4922
rect 19466 4870 19518 4922
rect 19530 4870 19582 4922
rect 19594 4870 19646 4922
rect 50122 4870 50174 4922
rect 50186 4870 50238 4922
rect 50250 4870 50302 4922
rect 50314 4870 50366 4922
rect 80842 4870 80894 4922
rect 80906 4870 80958 4922
rect 80970 4870 81022 4922
rect 81034 4870 81086 4922
rect 3240 4675 3292 4684
rect 3240 4641 3249 4675
rect 3249 4641 3283 4675
rect 3283 4641 3292 4675
rect 3240 4632 3292 4641
rect 3516 4675 3568 4684
rect 3516 4641 3525 4675
rect 3525 4641 3559 4675
rect 3559 4641 3568 4675
rect 3516 4632 3568 4641
rect 5264 4632 5316 4684
rect 5632 4675 5684 4684
rect 5632 4641 5641 4675
rect 5641 4641 5675 4675
rect 5675 4641 5684 4675
rect 5632 4632 5684 4641
rect 7380 4632 7432 4684
rect 7748 4675 7800 4684
rect 7748 4641 7757 4675
rect 7757 4641 7791 4675
rect 7791 4641 7800 4675
rect 7748 4632 7800 4641
rect 9588 4675 9640 4684
rect 9588 4641 9597 4675
rect 9597 4641 9631 4675
rect 9631 4641 9640 4675
rect 9588 4632 9640 4641
rect 9864 4675 9916 4684
rect 9864 4641 9873 4675
rect 9873 4641 9907 4675
rect 9907 4641 9916 4675
rect 9864 4632 9916 4641
rect 11704 4675 11756 4684
rect 11704 4641 11713 4675
rect 11713 4641 11747 4675
rect 11747 4641 11756 4675
rect 11704 4632 11756 4641
rect 11980 4675 12032 4684
rect 11980 4641 11989 4675
rect 11989 4641 12023 4675
rect 12023 4641 12032 4675
rect 11980 4632 12032 4641
rect 13820 4675 13872 4684
rect 13820 4641 13829 4675
rect 13829 4641 13863 4675
rect 13863 4641 13872 4675
rect 13820 4632 13872 4641
rect 14096 4675 14148 4684
rect 14096 4641 14105 4675
rect 14105 4641 14139 4675
rect 14139 4641 14148 4675
rect 14096 4632 14148 4641
rect 15936 4675 15988 4684
rect 15936 4641 15945 4675
rect 15945 4641 15979 4675
rect 15979 4641 15988 4675
rect 15936 4632 15988 4641
rect 16212 4675 16264 4684
rect 16212 4641 16221 4675
rect 16221 4641 16255 4675
rect 16255 4641 16264 4675
rect 16212 4632 16264 4641
rect 18052 4675 18104 4684
rect 18052 4641 18061 4675
rect 18061 4641 18095 4675
rect 18095 4641 18104 4675
rect 18052 4632 18104 4641
rect 18328 4675 18380 4684
rect 18328 4641 18337 4675
rect 18337 4641 18371 4675
rect 18371 4641 18380 4675
rect 18328 4632 18380 4641
rect 20076 4632 20128 4684
rect 20444 4675 20496 4684
rect 20444 4641 20453 4675
rect 20453 4641 20487 4675
rect 20487 4641 20496 4675
rect 20444 4632 20496 4641
rect 22192 4632 22244 4684
rect 22560 4675 22612 4684
rect 22560 4641 22569 4675
rect 22569 4641 22603 4675
rect 22603 4641 22612 4675
rect 22560 4632 22612 4641
rect 24400 4675 24452 4684
rect 24400 4641 24409 4675
rect 24409 4641 24443 4675
rect 24443 4641 24452 4675
rect 24400 4632 24452 4641
rect 24676 4675 24728 4684
rect 24676 4641 24685 4675
rect 24685 4641 24719 4675
rect 24719 4641 24728 4675
rect 24676 4632 24728 4641
rect 26516 4675 26568 4684
rect 26516 4641 26525 4675
rect 26525 4641 26559 4675
rect 26559 4641 26568 4675
rect 26516 4632 26568 4641
rect 26792 4675 26844 4684
rect 26792 4641 26801 4675
rect 26801 4641 26835 4675
rect 26835 4641 26844 4675
rect 26792 4632 26844 4641
rect 28632 4675 28684 4684
rect 28632 4641 28641 4675
rect 28641 4641 28675 4675
rect 28675 4641 28684 4675
rect 28632 4632 28684 4641
rect 28908 4675 28960 4684
rect 28908 4641 28917 4675
rect 28917 4641 28951 4675
rect 28951 4641 28960 4675
rect 28908 4632 28960 4641
rect 30748 4675 30800 4684
rect 30748 4641 30757 4675
rect 30757 4641 30791 4675
rect 30791 4641 30800 4675
rect 30748 4632 30800 4641
rect 31024 4675 31076 4684
rect 31024 4641 31033 4675
rect 31033 4641 31067 4675
rect 31067 4641 31076 4675
rect 31024 4632 31076 4641
rect 32864 4675 32916 4684
rect 32864 4641 32873 4675
rect 32873 4641 32907 4675
rect 32907 4641 32916 4675
rect 32864 4632 32916 4641
rect 33140 4675 33192 4684
rect 33140 4641 33149 4675
rect 33149 4641 33183 4675
rect 33183 4641 33192 4675
rect 33140 4632 33192 4641
rect 35072 4632 35124 4684
rect 35256 4675 35308 4684
rect 35256 4641 35265 4675
rect 35265 4641 35299 4675
rect 35299 4641 35308 4675
rect 35256 4632 35308 4641
rect 37096 4675 37148 4684
rect 37096 4641 37105 4675
rect 37105 4641 37139 4675
rect 37139 4641 37148 4675
rect 37096 4632 37148 4641
rect 37372 4675 37424 4684
rect 37372 4641 37381 4675
rect 37381 4641 37415 4675
rect 37415 4641 37424 4675
rect 37372 4632 37424 4641
rect 39212 4675 39264 4684
rect 39212 4641 39221 4675
rect 39221 4641 39255 4675
rect 39255 4641 39264 4675
rect 39212 4632 39264 4641
rect 39488 4675 39540 4684
rect 39488 4641 39497 4675
rect 39497 4641 39531 4675
rect 39531 4641 39540 4675
rect 39488 4632 39540 4641
rect 41236 4632 41288 4684
rect 41604 4675 41656 4684
rect 41604 4641 41613 4675
rect 41613 4641 41647 4675
rect 41647 4641 41656 4675
rect 41604 4632 41656 4641
rect 43444 4675 43496 4684
rect 43444 4641 43453 4675
rect 43453 4641 43487 4675
rect 43487 4641 43496 4675
rect 43444 4632 43496 4641
rect 43720 4675 43772 4684
rect 43720 4641 43729 4675
rect 43729 4641 43763 4675
rect 43763 4641 43772 4675
rect 43720 4632 43772 4641
rect 45560 4675 45612 4684
rect 45560 4641 45569 4675
rect 45569 4641 45603 4675
rect 45603 4641 45612 4675
rect 45560 4632 45612 4641
rect 45836 4675 45888 4684
rect 45836 4641 45845 4675
rect 45845 4641 45879 4675
rect 45879 4641 45888 4675
rect 45836 4632 45888 4641
rect 47676 4675 47728 4684
rect 47676 4641 47685 4675
rect 47685 4641 47719 4675
rect 47719 4641 47728 4675
rect 47676 4632 47728 4641
rect 47952 4675 48004 4684
rect 47952 4641 47961 4675
rect 47961 4641 47995 4675
rect 47995 4641 48004 4675
rect 47952 4632 48004 4641
rect 49792 4675 49844 4684
rect 49792 4641 49801 4675
rect 49801 4641 49835 4675
rect 49835 4641 49844 4675
rect 49792 4632 49844 4641
rect 51172 4632 51224 4684
rect 51908 4675 51960 4684
rect 51908 4641 51917 4675
rect 51917 4641 51951 4675
rect 51951 4641 51960 4675
rect 51908 4632 51960 4641
rect 52184 4675 52236 4684
rect 52184 4641 52193 4675
rect 52193 4641 52227 4675
rect 52227 4641 52236 4675
rect 52184 4632 52236 4641
rect 54024 4675 54076 4684
rect 54024 4641 54033 4675
rect 54033 4641 54067 4675
rect 54067 4641 54076 4675
rect 54024 4632 54076 4641
rect 54300 4675 54352 4684
rect 54300 4641 54309 4675
rect 54309 4641 54343 4675
rect 54343 4641 54352 4675
rect 54300 4632 54352 4641
rect 56048 4632 56100 4684
rect 56416 4675 56468 4684
rect 56416 4641 56425 4675
rect 56425 4641 56459 4675
rect 56459 4641 56468 4675
rect 56416 4632 56468 4641
rect 58164 4632 58216 4684
rect 58532 4675 58584 4684
rect 58532 4641 58541 4675
rect 58541 4641 58575 4675
rect 58575 4641 58584 4675
rect 58532 4632 58584 4641
rect 60648 4675 60700 4684
rect 60648 4641 60657 4675
rect 60657 4641 60691 4675
rect 60691 4641 60700 4675
rect 60648 4632 60700 4641
rect 62488 4675 62540 4684
rect 62488 4641 62497 4675
rect 62497 4641 62531 4675
rect 62531 4641 62540 4675
rect 62488 4632 62540 4641
rect 62764 4675 62816 4684
rect 62764 4641 62773 4675
rect 62773 4641 62807 4675
rect 62807 4641 62816 4675
rect 62764 4632 62816 4641
rect 64604 4675 64656 4684
rect 64604 4641 64613 4675
rect 64613 4641 64647 4675
rect 64647 4641 64656 4675
rect 64604 4632 64656 4641
rect 64880 4675 64932 4684
rect 64880 4641 64889 4675
rect 64889 4641 64923 4675
rect 64923 4641 64932 4675
rect 64880 4632 64932 4641
rect 66720 4675 66772 4684
rect 66720 4641 66729 4675
rect 66729 4641 66763 4675
rect 66763 4641 66772 4675
rect 66720 4632 66772 4641
rect 66996 4675 67048 4684
rect 66996 4641 67005 4675
rect 67005 4641 67039 4675
rect 67039 4641 67048 4675
rect 66996 4632 67048 4641
rect 68836 4675 68888 4684
rect 68836 4641 68845 4675
rect 68845 4641 68879 4675
rect 68879 4641 68888 4675
rect 68836 4632 68888 4641
rect 69112 4675 69164 4684
rect 69112 4641 69121 4675
rect 69121 4641 69155 4675
rect 69155 4641 69164 4675
rect 69112 4632 69164 4641
rect 70860 4632 70912 4684
rect 71228 4675 71280 4684
rect 71228 4641 71237 4675
rect 71237 4641 71271 4675
rect 71271 4641 71280 4675
rect 71228 4632 71280 4641
rect 72976 4632 73028 4684
rect 73344 4675 73396 4684
rect 73344 4641 73353 4675
rect 73353 4641 73387 4675
rect 73387 4641 73396 4675
rect 73344 4632 73396 4641
rect 75092 4632 75144 4684
rect 75460 4675 75512 4684
rect 75460 4641 75469 4675
rect 75469 4641 75503 4675
rect 75503 4641 75512 4675
rect 75460 4632 75512 4641
rect 77576 4675 77628 4684
rect 77576 4641 77585 4675
rect 77585 4641 77619 4675
rect 77619 4641 77628 4675
rect 77576 4632 77628 4641
rect 79324 4632 79376 4684
rect 79692 4675 79744 4684
rect 79692 4641 79701 4675
rect 79701 4641 79735 4675
rect 79735 4641 79744 4675
rect 79692 4632 79744 4641
rect 81440 4632 81492 4684
rect 81808 4675 81860 4684
rect 81808 4641 81817 4675
rect 81817 4641 81851 4675
rect 81851 4641 81860 4675
rect 81808 4632 81860 4641
rect 83556 4632 83608 4684
rect 83924 4675 83976 4684
rect 83924 4641 83933 4675
rect 83933 4641 83967 4675
rect 83967 4641 83976 4675
rect 83924 4632 83976 4641
rect 85672 4632 85724 4684
rect 86040 4675 86092 4684
rect 86040 4641 86049 4675
rect 86049 4641 86083 4675
rect 86083 4641 86092 4675
rect 86040 4632 86092 4641
rect 87788 4632 87840 4684
rect 88156 4675 88208 4684
rect 88156 4641 88165 4675
rect 88165 4641 88199 4675
rect 88199 4641 88208 4675
rect 88156 4632 88208 4641
rect 89904 4632 89956 4684
rect 90272 4675 90324 4684
rect 90272 4641 90281 4675
rect 90281 4641 90315 4675
rect 90315 4641 90324 4675
rect 90272 4632 90324 4641
rect 92020 4632 92072 4684
rect 92388 4675 92440 4684
rect 92388 4641 92397 4675
rect 92397 4641 92431 4675
rect 92431 4641 92440 4675
rect 92388 4632 92440 4641
rect 94228 4675 94280 4684
rect 94228 4641 94237 4675
rect 94237 4641 94271 4675
rect 94271 4641 94280 4675
rect 94228 4632 94280 4641
rect 94504 4675 94556 4684
rect 94504 4641 94513 4675
rect 94513 4641 94547 4675
rect 94547 4641 94556 4675
rect 94504 4632 94556 4641
rect 96068 4632 96120 4684
rect 96620 4675 96672 4684
rect 96620 4641 96629 4675
rect 96629 4641 96663 4675
rect 96663 4641 96672 4675
rect 96620 4632 96672 4641
rect 98368 4632 98420 4684
rect 98736 4675 98788 4684
rect 98736 4641 98745 4675
rect 98745 4641 98779 4675
rect 98779 4641 98788 4675
rect 98736 4632 98788 4641
rect 100484 4632 100536 4684
rect 100852 4675 100904 4684
rect 100852 4641 100861 4675
rect 100861 4641 100895 4675
rect 100895 4641 100904 4675
rect 100852 4632 100904 4641
rect 102692 4675 102744 4684
rect 102692 4641 102701 4675
rect 102701 4641 102735 4675
rect 102735 4641 102744 4675
rect 102692 4632 102744 4641
rect 102968 4675 103020 4684
rect 102968 4641 102977 4675
rect 102977 4641 103011 4675
rect 103011 4641 103020 4675
rect 102968 4632 103020 4641
rect 104808 4675 104860 4684
rect 104808 4641 104817 4675
rect 104817 4641 104851 4675
rect 104851 4641 104860 4675
rect 104808 4632 104860 4641
rect 105084 4675 105136 4684
rect 105084 4641 105093 4675
rect 105093 4641 105127 4675
rect 105127 4641 105136 4675
rect 105084 4632 105136 4641
rect 1124 4607 1176 4616
rect 1124 4573 1133 4607
rect 1133 4573 1167 4607
rect 1167 4573 1176 4607
rect 1124 4564 1176 4573
rect 6276 4564 6328 4616
rect 27436 4564 27488 4616
rect 29552 4564 29604 4616
rect 38016 4564 38068 4616
rect 60372 4607 60424 4616
rect 60372 4573 60381 4607
rect 60381 4573 60415 4607
rect 60415 4573 60424 4607
rect 60372 4564 60424 4573
rect 77300 4607 77352 4616
rect 77300 4573 77309 4607
rect 77309 4573 77343 4607
rect 77343 4573 77352 4607
rect 77300 4564 77352 4573
rect 2228 4428 2280 4480
rect 4344 4428 4396 4480
rect 8208 4428 8260 4480
rect 10508 4428 10560 4480
rect 12624 4428 12676 4480
rect 14556 4428 14608 4480
rect 16856 4428 16908 4480
rect 18972 4428 19024 4480
rect 21088 4428 21140 4480
rect 23204 4428 23256 4480
rect 25320 4428 25372 4480
rect 31484 4428 31536 4480
rect 33784 4428 33836 4480
rect 35900 4428 35952 4480
rect 40132 4428 40184 4480
rect 42248 4428 42300 4480
rect 44364 4428 44416 4480
rect 46480 4428 46532 4480
rect 48412 4428 48464 4480
rect 50712 4428 50764 4480
rect 52828 4428 52880 4480
rect 54944 4428 54996 4480
rect 57060 4428 57112 4480
rect 59176 4428 59228 4480
rect 61292 4428 61344 4480
rect 63408 4428 63460 4480
rect 65340 4428 65392 4480
rect 67640 4428 67692 4480
rect 69756 4428 69808 4480
rect 71872 4428 71924 4480
rect 73988 4428 74040 4480
rect 76564 4471 76616 4480
rect 76564 4437 76573 4471
rect 76573 4437 76607 4471
rect 76607 4437 76616 4471
rect 76564 4428 76616 4437
rect 78864 4471 78916 4480
rect 78864 4437 78873 4471
rect 78873 4437 78907 4471
rect 78907 4437 78916 4471
rect 78864 4428 78916 4437
rect 81164 4428 81216 4480
rect 82636 4428 82688 4480
rect 84660 4428 84712 4480
rect 86868 4428 86920 4480
rect 89260 4471 89312 4480
rect 89260 4437 89269 4471
rect 89269 4437 89303 4471
rect 89303 4437 89312 4471
rect 89260 4428 89312 4437
rect 91284 4428 91336 4480
rect 93676 4471 93728 4480
rect 93676 4437 93685 4471
rect 93685 4437 93719 4471
rect 93719 4437 93728 4471
rect 93676 4428 93728 4437
rect 95792 4471 95844 4480
rect 95792 4437 95801 4471
rect 95801 4437 95835 4471
rect 95835 4437 95844 4471
rect 95792 4428 95844 4437
rect 98000 4428 98052 4480
rect 99380 4428 99432 4480
rect 101588 4428 101640 4480
rect 103796 4428 103848 4480
rect 106004 4428 106056 4480
rect 4042 4326 4094 4378
rect 4106 4326 4158 4378
rect 4170 4326 4222 4378
rect 4234 4326 4286 4378
rect 34762 4326 34814 4378
rect 34826 4326 34878 4378
rect 34890 4326 34942 4378
rect 34954 4326 35006 4378
rect 65482 4326 65534 4378
rect 65546 4326 65598 4378
rect 65610 4326 65662 4378
rect 65674 4326 65726 4378
rect 96202 4326 96254 4378
rect 96266 4326 96318 4378
rect 96330 4326 96382 4378
rect 96394 4326 96446 4378
rect 20076 4156 20128 4208
rect 1124 4131 1176 4140
rect 1124 4097 1133 4131
rect 1133 4097 1167 4131
rect 1167 4097 1176 4131
rect 1124 4088 1176 4097
rect 3240 4131 3292 4140
rect 3240 4097 3249 4131
rect 3249 4097 3283 4131
rect 3283 4097 3292 4131
rect 3240 4088 3292 4097
rect 5264 4088 5316 4140
rect 7380 4088 7432 4140
rect 9588 4131 9640 4140
rect 9588 4097 9597 4131
rect 9597 4097 9631 4131
rect 9631 4097 9640 4131
rect 9588 4088 9640 4097
rect 11704 4131 11756 4140
rect 11704 4097 11713 4131
rect 11713 4097 11747 4131
rect 11747 4097 11756 4131
rect 11704 4088 11756 4097
rect 13820 4131 13872 4140
rect 13820 4097 13829 4131
rect 13829 4097 13863 4131
rect 13863 4097 13872 4131
rect 13820 4088 13872 4097
rect 15936 4131 15988 4140
rect 15936 4097 15945 4131
rect 15945 4097 15979 4131
rect 15979 4097 15988 4131
rect 15936 4088 15988 4097
rect 18052 4131 18104 4140
rect 18052 4097 18061 4131
rect 18061 4097 18095 4131
rect 18095 4097 18104 4131
rect 18052 4088 18104 4097
rect 58164 4156 58216 4208
rect 22192 4088 22244 4140
rect 24400 4131 24452 4140
rect 24400 4097 24409 4131
rect 24409 4097 24443 4131
rect 24443 4097 24452 4131
rect 24400 4088 24452 4097
rect 26516 4131 26568 4140
rect 26516 4097 26525 4131
rect 26525 4097 26559 4131
rect 26559 4097 26568 4131
rect 26516 4088 26568 4097
rect 28632 4131 28684 4140
rect 28632 4097 28641 4131
rect 28641 4097 28675 4131
rect 28675 4097 28684 4131
rect 28632 4088 28684 4097
rect 30748 4131 30800 4140
rect 30748 4097 30757 4131
rect 30757 4097 30791 4131
rect 30791 4097 30800 4131
rect 30748 4088 30800 4097
rect 32864 4131 32916 4140
rect 32864 4097 32873 4131
rect 32873 4097 32907 4131
rect 32907 4097 32916 4131
rect 32864 4088 32916 4097
rect 37096 4131 37148 4140
rect 37096 4097 37105 4131
rect 37105 4097 37139 4131
rect 37139 4097 37148 4131
rect 37096 4088 37148 4097
rect 39212 4131 39264 4140
rect 39212 4097 39221 4131
rect 39221 4097 39255 4131
rect 39255 4097 39264 4131
rect 39212 4088 39264 4097
rect 41236 4088 41288 4140
rect 43444 4131 43496 4140
rect 43444 4097 43453 4131
rect 43453 4097 43487 4131
rect 43487 4097 43496 4131
rect 43444 4088 43496 4097
rect 45560 4131 45612 4140
rect 45560 4097 45569 4131
rect 45569 4097 45603 4131
rect 45603 4097 45612 4131
rect 45560 4088 45612 4097
rect 47676 4131 47728 4140
rect 47676 4097 47685 4131
rect 47685 4097 47719 4131
rect 47719 4097 47728 4131
rect 47676 4088 47728 4097
rect 49792 4131 49844 4140
rect 49792 4097 49801 4131
rect 49801 4097 49835 4131
rect 49835 4097 49844 4131
rect 49792 4088 49844 4097
rect 51908 4131 51960 4140
rect 51908 4097 51917 4131
rect 51917 4097 51951 4131
rect 51951 4097 51960 4131
rect 51908 4088 51960 4097
rect 54024 4131 54076 4140
rect 54024 4097 54033 4131
rect 54033 4097 54067 4131
rect 54067 4097 54076 4131
rect 54024 4088 54076 4097
rect 70860 4156 70912 4208
rect 62488 4131 62540 4140
rect 62488 4097 62497 4131
rect 62497 4097 62531 4131
rect 62531 4097 62540 4131
rect 62488 4088 62540 4097
rect 64604 4131 64656 4140
rect 64604 4097 64613 4131
rect 64613 4097 64647 4131
rect 64647 4097 64656 4131
rect 64604 4088 64656 4097
rect 66720 4131 66772 4140
rect 66720 4097 66729 4131
rect 66729 4097 66763 4131
rect 66763 4097 66772 4131
rect 66720 4088 66772 4097
rect 68836 4131 68888 4140
rect 68836 4097 68845 4131
rect 68845 4097 68879 4131
rect 68879 4097 68888 4131
rect 68836 4088 68888 4097
rect 75092 4156 75144 4208
rect 73068 4131 73120 4140
rect 73068 4097 73077 4131
rect 73077 4097 73111 4131
rect 73111 4097 73120 4131
rect 73068 4088 73120 4097
rect 83556 4156 83608 4208
rect 79324 4088 79376 4140
rect 81532 4131 81584 4140
rect 81532 4097 81541 4131
rect 81541 4097 81575 4131
rect 81575 4097 81584 4131
rect 81532 4088 81584 4097
rect 87788 4156 87840 4208
rect 85764 4131 85816 4140
rect 85764 4097 85773 4131
rect 85773 4097 85807 4131
rect 85807 4097 85816 4131
rect 85764 4088 85816 4097
rect 92020 4088 92072 4140
rect 94228 4131 94280 4140
rect 94228 4097 94237 4131
rect 94237 4097 94271 4131
rect 94271 4097 94280 4131
rect 94228 4088 94280 4097
rect 96068 4088 96120 4140
rect 98368 4088 98420 4140
rect 100484 4088 100536 4140
rect 102692 4131 102744 4140
rect 102692 4097 102701 4131
rect 102701 4097 102735 4131
rect 102735 4097 102744 4131
rect 102692 4088 102744 4097
rect 104808 4131 104860 4140
rect 104808 4097 104817 4131
rect 104817 4097 104851 4131
rect 104851 4097 104860 4131
rect 104808 4088 104860 4097
rect 2504 4020 2556 4072
rect 3884 4020 3936 4072
rect 6000 4020 6052 4072
rect 8116 4020 8168 4072
rect 10968 4020 11020 4072
rect 13084 4020 13136 4072
rect 15200 4020 15252 4072
rect 17316 4020 17368 4072
rect 18420 4020 18472 4072
rect 21088 4020 21140 4072
rect 22928 4020 22980 4072
rect 25044 4020 25096 4072
rect 27896 4020 27948 4072
rect 30012 4020 30064 4072
rect 32128 4020 32180 4072
rect 34244 4020 34296 4072
rect 35072 4020 35124 4072
rect 35624 4020 35676 4072
rect 37740 4020 37792 4072
rect 39948 4020 40000 4072
rect 41972 4020 42024 4072
rect 44824 4020 44876 4072
rect 46940 4020 46992 4072
rect 49056 4020 49108 4072
rect 51172 4020 51224 4072
rect 52276 4020 52328 4072
rect 54668 4020 54720 4072
rect 56140 4063 56192 4072
rect 56140 4029 56149 4063
rect 56149 4029 56183 4063
rect 56183 4029 56192 4063
rect 56140 4020 56192 4029
rect 57152 4020 57204 4072
rect 58992 4020 59044 4072
rect 60372 4063 60424 4072
rect 60372 4029 60381 4063
rect 60381 4029 60415 4063
rect 60415 4029 60424 4063
rect 60372 4020 60424 4029
rect 61292 4020 61344 4072
rect 63868 4020 63920 4072
rect 65984 4020 66036 4072
rect 68100 4020 68152 4072
rect 69204 4020 69256 4072
rect 71688 4020 71740 4072
rect 73712 4020 73764 4072
rect 75828 4020 75880 4072
rect 77300 4063 77352 4072
rect 77300 4029 77309 4063
rect 77309 4029 77343 4063
rect 77343 4029 77352 4063
rect 77300 4020 77352 4029
rect 78680 4020 78732 4072
rect 80704 4020 80756 4072
rect 82912 4020 82964 4072
rect 85028 4020 85080 4072
rect 86132 4020 86184 4072
rect 88524 4020 88576 4072
rect 89996 4063 90048 4072
rect 89996 4029 90005 4063
rect 90005 4029 90039 4063
rect 90039 4029 90048 4063
rect 89996 4020 90048 4029
rect 90640 4020 90692 4072
rect 93124 4020 93176 4072
rect 95608 4020 95660 4072
rect 97264 4020 97316 4072
rect 99840 4020 99892 4072
rect 101956 4020 102008 4072
rect 103612 4020 103664 4072
rect 105452 4020 105504 4072
rect 81256 3952 81308 4004
rect 1492 3884 1544 3936
rect 4620 3927 4672 3936
rect 4620 3893 4629 3927
rect 4629 3893 4663 3927
rect 4663 3893 4672 3927
rect 4620 3884 4672 3893
rect 6736 3927 6788 3936
rect 6736 3893 6745 3927
rect 6745 3893 6779 3927
rect 6779 3893 6788 3927
rect 6736 3884 6788 3893
rect 8852 3927 8904 3936
rect 8852 3893 8861 3927
rect 8861 3893 8895 3927
rect 8895 3893 8904 3927
rect 11152 3927 11204 3936
rect 8852 3884 8904 3893
rect 11152 3893 11161 3927
rect 11161 3893 11195 3927
rect 11195 3893 11204 3927
rect 11152 3884 11204 3893
rect 13268 3927 13320 3936
rect 13268 3893 13277 3927
rect 13277 3893 13311 3927
rect 13311 3893 13320 3927
rect 13268 3884 13320 3893
rect 14188 3884 14240 3936
rect 16304 3884 16356 3936
rect 18696 3884 18748 3936
rect 21548 3927 21600 3936
rect 21548 3893 21557 3927
rect 21557 3893 21591 3927
rect 21591 3893 21600 3927
rect 21548 3884 21600 3893
rect 23664 3927 23716 3936
rect 23664 3893 23673 3927
rect 23673 3893 23707 3927
rect 23707 3893 23716 3927
rect 23664 3884 23716 3893
rect 25780 3927 25832 3936
rect 25780 3893 25789 3927
rect 25789 3893 25823 3927
rect 25823 3893 25832 3927
rect 25780 3884 25832 3893
rect 28080 3927 28132 3936
rect 28080 3893 28089 3927
rect 28089 3893 28123 3927
rect 28123 3893 28132 3927
rect 28080 3884 28132 3893
rect 30196 3927 30248 3936
rect 30196 3893 30205 3927
rect 30205 3893 30239 3927
rect 30239 3893 30248 3927
rect 30196 3884 30248 3893
rect 31116 3884 31168 3936
rect 33232 3884 33284 3936
rect 35348 3884 35400 3936
rect 38476 3927 38528 3936
rect 38476 3893 38485 3927
rect 38485 3893 38519 3927
rect 38519 3893 38528 3927
rect 38476 3884 38528 3893
rect 40592 3927 40644 3936
rect 40592 3893 40601 3927
rect 40601 3893 40635 3927
rect 40635 3893 40644 3927
rect 40592 3884 40644 3893
rect 42708 3927 42760 3936
rect 42708 3893 42717 3927
rect 42717 3893 42751 3927
rect 42751 3893 42760 3927
rect 42708 3884 42760 3893
rect 45008 3927 45060 3936
rect 45008 3893 45017 3927
rect 45017 3893 45051 3927
rect 45051 3893 45060 3927
rect 45008 3884 45060 3893
rect 47124 3927 47176 3936
rect 47124 3893 47133 3927
rect 47133 3893 47167 3927
rect 47167 3893 47176 3927
rect 47124 3884 47176 3893
rect 48044 3884 48096 3936
rect 50528 3884 50580 3936
rect 52552 3884 52604 3936
rect 55404 3927 55456 3936
rect 55404 3893 55413 3927
rect 55413 3893 55447 3927
rect 55447 3893 55456 3927
rect 55404 3884 55456 3893
rect 57520 3927 57572 3936
rect 57520 3893 57529 3927
rect 57529 3893 57563 3927
rect 57563 3893 57572 3927
rect 57520 3884 57572 3893
rect 59636 3927 59688 3936
rect 59636 3893 59645 3927
rect 59645 3893 59679 3927
rect 59679 3893 59688 3927
rect 59636 3884 59688 3893
rect 61936 3927 61988 3936
rect 61936 3893 61945 3927
rect 61945 3893 61979 3927
rect 61979 3893 61988 3927
rect 61936 3884 61988 3893
rect 64052 3927 64104 3936
rect 64052 3893 64061 3927
rect 64061 3893 64095 3927
rect 64095 3893 64104 3927
rect 64052 3884 64104 3893
rect 64972 3884 65024 3936
rect 67088 3884 67140 3936
rect 69480 3884 69532 3936
rect 72332 3927 72384 3936
rect 72332 3893 72341 3927
rect 72341 3893 72375 3927
rect 72375 3893 72384 3927
rect 72332 3884 72384 3893
rect 74448 3927 74500 3936
rect 74448 3893 74457 3927
rect 74457 3893 74491 3927
rect 74491 3893 74500 3927
rect 74448 3884 74500 3893
rect 76748 3927 76800 3936
rect 76748 3893 76757 3927
rect 76757 3893 76791 3927
rect 76791 3893 76800 3927
rect 76748 3884 76800 3893
rect 78772 3884 78824 3936
rect 81900 3884 81952 3936
rect 84016 3884 84068 3936
rect 86408 3884 86460 3936
rect 89444 3927 89496 3936
rect 89444 3893 89453 3927
rect 89453 3893 89487 3927
rect 89487 3893 89496 3927
rect 89444 3884 89496 3893
rect 91376 3927 91428 3936
rect 91376 3893 91385 3927
rect 91385 3893 91419 3927
rect 91419 3893 91428 3927
rect 91376 3884 91428 3893
rect 93492 3927 93544 3936
rect 93492 3893 93501 3927
rect 93501 3893 93535 3927
rect 93535 3893 93544 3927
rect 93492 3884 93544 3893
rect 95700 3884 95752 3936
rect 97908 3927 97960 3936
rect 97908 3893 97917 3927
rect 97917 3893 97951 3927
rect 97951 3893 97960 3927
rect 97908 3884 97960 3893
rect 98828 3884 98880 3936
rect 100944 3884 100996 3936
rect 103060 3884 103112 3936
rect 105176 3884 105228 3936
rect 19402 3782 19454 3834
rect 19466 3782 19518 3834
rect 19530 3782 19582 3834
rect 19594 3782 19646 3834
rect 50122 3782 50174 3834
rect 50186 3782 50238 3834
rect 50250 3782 50302 3834
rect 50314 3782 50366 3834
rect 80842 3782 80894 3834
rect 80906 3782 80958 3834
rect 80970 3782 81022 3834
rect 81034 3782 81086 3834
rect 2504 3723 2556 3732
rect 2504 3689 2513 3723
rect 2513 3689 2547 3723
rect 2547 3689 2556 3723
rect 2504 3680 2556 3689
rect 10968 3723 11020 3732
rect 10968 3689 10977 3723
rect 10977 3689 11011 3723
rect 11011 3689 11020 3723
rect 10968 3680 11020 3689
rect 13084 3723 13136 3732
rect 13084 3689 13093 3723
rect 13093 3689 13127 3723
rect 13127 3689 13136 3723
rect 13084 3680 13136 3689
rect 15200 3723 15252 3732
rect 15200 3689 15209 3723
rect 15209 3689 15243 3723
rect 15243 3689 15252 3723
rect 15200 3680 15252 3689
rect 17316 3723 17368 3732
rect 17316 3689 17325 3723
rect 17325 3689 17359 3723
rect 17359 3689 17368 3723
rect 17316 3680 17368 3689
rect 27896 3723 27948 3732
rect 27896 3689 27905 3723
rect 27905 3689 27939 3723
rect 27939 3689 27948 3723
rect 27896 3680 27948 3689
rect 30012 3723 30064 3732
rect 30012 3689 30021 3723
rect 30021 3689 30055 3723
rect 30055 3689 30064 3723
rect 30012 3680 30064 3689
rect 32128 3723 32180 3732
rect 32128 3689 32137 3723
rect 32137 3689 32171 3723
rect 32171 3689 32180 3723
rect 32128 3680 32180 3689
rect 34244 3723 34296 3732
rect 34244 3689 34253 3723
rect 34253 3689 34287 3723
rect 34287 3689 34296 3723
rect 34244 3680 34296 3689
rect 44824 3723 44876 3732
rect 44824 3689 44833 3723
rect 44833 3689 44867 3723
rect 44867 3689 44876 3723
rect 44824 3680 44876 3689
rect 46940 3723 46992 3732
rect 46940 3689 46949 3723
rect 46949 3689 46983 3723
rect 46983 3689 46992 3723
rect 46940 3680 46992 3689
rect 49056 3723 49108 3732
rect 49056 3689 49065 3723
rect 49065 3689 49099 3723
rect 49099 3689 49108 3723
rect 49056 3680 49108 3689
rect 51172 3723 51224 3732
rect 51172 3689 51181 3723
rect 51181 3689 51215 3723
rect 51215 3689 51224 3723
rect 51172 3680 51224 3689
rect 63868 3723 63920 3732
rect 63868 3689 63877 3723
rect 63877 3689 63911 3723
rect 63911 3689 63920 3723
rect 63868 3680 63920 3689
rect 65984 3723 66036 3732
rect 65984 3689 65993 3723
rect 65993 3689 66027 3723
rect 66027 3689 66036 3723
rect 65984 3680 66036 3689
rect 68100 3723 68152 3732
rect 68100 3689 68109 3723
rect 68109 3689 68143 3723
rect 68143 3689 68152 3723
rect 68100 3680 68152 3689
rect 78680 3723 78732 3732
rect 78680 3689 78689 3723
rect 78689 3689 78723 3723
rect 78723 3689 78732 3723
rect 78680 3680 78732 3689
rect 80704 3680 80756 3732
rect 82912 3723 82964 3732
rect 82912 3689 82921 3723
rect 82921 3689 82955 3723
rect 82955 3689 82964 3723
rect 82912 3680 82964 3689
rect 85028 3723 85080 3732
rect 85028 3689 85037 3723
rect 85037 3689 85071 3723
rect 85071 3689 85080 3723
rect 85028 3680 85080 3689
rect 95608 3723 95660 3732
rect 95608 3689 95617 3723
rect 95617 3689 95651 3723
rect 95651 3689 95660 3723
rect 95608 3680 95660 3689
rect 99840 3723 99892 3732
rect 99840 3689 99849 3723
rect 99849 3689 99883 3723
rect 99883 3689 99892 3723
rect 99840 3680 99892 3689
rect 101956 3723 102008 3732
rect 101956 3689 101965 3723
rect 101965 3689 101999 3723
rect 101999 3689 102008 3723
rect 101956 3680 102008 3689
rect 1124 3587 1176 3596
rect 1124 3553 1133 3587
rect 1133 3553 1167 3587
rect 1167 3553 1176 3587
rect 1124 3544 1176 3553
rect 3240 3587 3292 3596
rect 3240 3553 3249 3587
rect 3249 3553 3283 3587
rect 3283 3553 3292 3587
rect 3240 3544 3292 3553
rect 5356 3587 5408 3596
rect 5356 3553 5365 3587
rect 5365 3553 5399 3587
rect 5399 3553 5408 3587
rect 5356 3544 5408 3553
rect 7472 3587 7524 3596
rect 7472 3553 7481 3587
rect 7481 3553 7515 3587
rect 7515 3553 7524 3587
rect 7472 3544 7524 3553
rect 9588 3587 9640 3596
rect 9588 3553 9597 3587
rect 9597 3553 9631 3587
rect 9631 3553 9640 3587
rect 9588 3544 9640 3553
rect 11704 3587 11756 3596
rect 11704 3553 11713 3587
rect 11713 3553 11747 3587
rect 11747 3553 11756 3587
rect 11704 3544 11756 3553
rect 13820 3587 13872 3596
rect 13820 3553 13829 3587
rect 13829 3553 13863 3587
rect 13863 3553 13872 3587
rect 13820 3544 13872 3553
rect 15936 3587 15988 3596
rect 15936 3553 15945 3587
rect 15945 3553 15979 3587
rect 15979 3553 15988 3587
rect 15936 3544 15988 3553
rect 18052 3587 18104 3596
rect 18052 3553 18061 3587
rect 18061 3553 18095 3587
rect 18095 3553 18104 3587
rect 18052 3544 18104 3553
rect 20168 3587 20220 3596
rect 20168 3553 20177 3587
rect 20177 3553 20211 3587
rect 20211 3553 20220 3587
rect 20168 3544 20220 3553
rect 22192 3544 22244 3596
rect 24400 3587 24452 3596
rect 24400 3553 24409 3587
rect 24409 3553 24443 3587
rect 24443 3553 24452 3587
rect 24400 3544 24452 3553
rect 26516 3587 26568 3596
rect 26516 3553 26525 3587
rect 26525 3553 26559 3587
rect 26559 3553 26568 3587
rect 26516 3544 26568 3553
rect 28632 3587 28684 3596
rect 28632 3553 28641 3587
rect 28641 3553 28675 3587
rect 28675 3553 28684 3587
rect 28632 3544 28684 3553
rect 30748 3587 30800 3596
rect 30748 3553 30757 3587
rect 30757 3553 30791 3587
rect 30791 3553 30800 3587
rect 30748 3544 30800 3553
rect 32864 3587 32916 3596
rect 32864 3553 32873 3587
rect 32873 3553 32907 3587
rect 32907 3553 32916 3587
rect 32864 3544 32916 3553
rect 35072 3544 35124 3596
rect 37096 3587 37148 3596
rect 37096 3553 37105 3587
rect 37105 3553 37139 3587
rect 37139 3553 37148 3587
rect 37096 3544 37148 3553
rect 39212 3587 39264 3596
rect 39212 3553 39221 3587
rect 39221 3553 39255 3587
rect 39255 3553 39264 3587
rect 39212 3544 39264 3553
rect 39488 3587 39540 3596
rect 39488 3553 39497 3587
rect 39497 3553 39531 3587
rect 39531 3553 39540 3587
rect 39488 3544 39540 3553
rect 40408 3544 40460 3596
rect 41328 3587 41380 3596
rect 41328 3553 41337 3587
rect 41337 3553 41371 3587
rect 41371 3553 41380 3587
rect 41328 3544 41380 3553
rect 43444 3587 43496 3596
rect 43444 3553 43453 3587
rect 43453 3553 43487 3587
rect 43487 3553 43496 3587
rect 43444 3544 43496 3553
rect 45560 3587 45612 3596
rect 45560 3553 45569 3587
rect 45569 3553 45603 3587
rect 45603 3553 45612 3587
rect 45560 3544 45612 3553
rect 47676 3587 47728 3596
rect 47676 3553 47685 3587
rect 47685 3553 47719 3587
rect 47719 3553 47728 3587
rect 47676 3544 47728 3553
rect 49792 3587 49844 3596
rect 49792 3553 49801 3587
rect 49801 3553 49835 3587
rect 49835 3553 49844 3587
rect 49792 3544 49844 3553
rect 51908 3587 51960 3596
rect 51908 3553 51917 3587
rect 51917 3553 51951 3587
rect 51951 3553 51960 3587
rect 51908 3544 51960 3553
rect 54024 3587 54076 3596
rect 54024 3553 54033 3587
rect 54033 3553 54067 3587
rect 54067 3553 54076 3587
rect 54024 3544 54076 3553
rect 56140 3587 56192 3596
rect 56140 3553 56149 3587
rect 56149 3553 56183 3587
rect 56183 3553 56192 3587
rect 56140 3544 56192 3553
rect 58256 3587 58308 3596
rect 58256 3553 58265 3587
rect 58265 3553 58299 3587
rect 58299 3553 58308 3587
rect 58256 3544 58308 3553
rect 60372 3587 60424 3596
rect 60372 3553 60381 3587
rect 60381 3553 60415 3587
rect 60415 3553 60424 3587
rect 62488 3587 62540 3596
rect 60372 3544 60424 3553
rect 62488 3553 62497 3587
rect 62497 3553 62531 3587
rect 62531 3553 62540 3587
rect 62488 3544 62540 3553
rect 64604 3587 64656 3596
rect 64604 3553 64613 3587
rect 64613 3553 64647 3587
rect 64647 3553 64656 3587
rect 64604 3544 64656 3553
rect 66720 3587 66772 3596
rect 66720 3553 66729 3587
rect 66729 3553 66763 3587
rect 66763 3553 66772 3587
rect 66720 3544 66772 3553
rect 68836 3587 68888 3596
rect 68836 3553 68845 3587
rect 68845 3553 68879 3587
rect 68879 3553 68888 3587
rect 68836 3544 68888 3553
rect 70952 3587 71004 3596
rect 70952 3553 70961 3587
rect 70961 3553 70995 3587
rect 70995 3553 71004 3587
rect 70952 3544 71004 3553
rect 73068 3587 73120 3596
rect 73068 3553 73077 3587
rect 73077 3553 73111 3587
rect 73111 3553 73120 3587
rect 73068 3544 73120 3553
rect 75184 3587 75236 3596
rect 75184 3553 75193 3587
rect 75193 3553 75227 3587
rect 75227 3553 75236 3587
rect 75184 3544 75236 3553
rect 1400 3519 1452 3528
rect 1400 3485 1409 3519
rect 1409 3485 1443 3519
rect 1443 3485 1452 3519
rect 1400 3476 1452 3485
rect 3516 3519 3568 3528
rect 3516 3485 3525 3519
rect 3525 3485 3559 3519
rect 3559 3485 3568 3519
rect 3516 3476 3568 3485
rect 3884 3476 3936 3528
rect 5632 3519 5684 3528
rect 5632 3485 5641 3519
rect 5641 3485 5675 3519
rect 5675 3485 5684 3519
rect 5632 3476 5684 3485
rect 6000 3476 6052 3528
rect 7748 3519 7800 3528
rect 7748 3485 7757 3519
rect 7757 3485 7791 3519
rect 7791 3485 7800 3519
rect 7748 3476 7800 3485
rect 8116 3476 8168 3528
rect 9864 3519 9916 3528
rect 9864 3485 9873 3519
rect 9873 3485 9907 3519
rect 9907 3485 9916 3519
rect 9864 3476 9916 3485
rect 11980 3519 12032 3528
rect 11980 3485 11989 3519
rect 11989 3485 12023 3519
rect 12023 3485 12032 3519
rect 11980 3476 12032 3485
rect 14096 3519 14148 3528
rect 14096 3485 14105 3519
rect 14105 3485 14139 3519
rect 14139 3485 14148 3519
rect 14096 3476 14148 3485
rect 16212 3519 16264 3528
rect 16212 3485 16221 3519
rect 16221 3485 16255 3519
rect 16255 3485 16264 3519
rect 16212 3476 16264 3485
rect 18328 3519 18380 3528
rect 18328 3485 18337 3519
rect 18337 3485 18371 3519
rect 18371 3485 18380 3519
rect 18328 3476 18380 3485
rect 18420 3476 18472 3528
rect 20444 3519 20496 3528
rect 20444 3485 20453 3519
rect 20453 3485 20487 3519
rect 20487 3485 20496 3519
rect 20444 3476 20496 3485
rect 21088 3476 21140 3528
rect 22560 3519 22612 3528
rect 22560 3485 22569 3519
rect 22569 3485 22603 3519
rect 22603 3485 22612 3519
rect 22560 3476 22612 3485
rect 22928 3476 22980 3528
rect 24676 3519 24728 3528
rect 24676 3485 24685 3519
rect 24685 3485 24719 3519
rect 24719 3485 24728 3519
rect 24676 3476 24728 3485
rect 25044 3476 25096 3528
rect 26792 3519 26844 3528
rect 26792 3485 26801 3519
rect 26801 3485 26835 3519
rect 26835 3485 26844 3519
rect 26792 3476 26844 3485
rect 28908 3519 28960 3528
rect 28908 3485 28917 3519
rect 28917 3485 28951 3519
rect 28951 3485 28960 3519
rect 28908 3476 28960 3485
rect 31024 3519 31076 3528
rect 31024 3485 31033 3519
rect 31033 3485 31067 3519
rect 31067 3485 31076 3519
rect 31024 3476 31076 3485
rect 33140 3519 33192 3528
rect 33140 3485 33149 3519
rect 33149 3485 33183 3519
rect 33183 3485 33192 3519
rect 33140 3476 33192 3485
rect 35256 3519 35308 3528
rect 35256 3485 35265 3519
rect 35265 3485 35299 3519
rect 35299 3485 35308 3519
rect 35256 3476 35308 3485
rect 35624 3476 35676 3528
rect 37372 3519 37424 3528
rect 37372 3485 37381 3519
rect 37381 3485 37415 3519
rect 37415 3485 37424 3519
rect 37372 3476 37424 3485
rect 37740 3476 37792 3528
rect 39948 3476 40000 3528
rect 41604 3519 41656 3528
rect 41604 3485 41613 3519
rect 41613 3485 41647 3519
rect 41647 3485 41656 3519
rect 41604 3476 41656 3485
rect 41972 3476 42024 3528
rect 43720 3519 43772 3528
rect 43720 3485 43729 3519
rect 43729 3485 43763 3519
rect 43763 3485 43772 3519
rect 43720 3476 43772 3485
rect 45836 3519 45888 3528
rect 45836 3485 45845 3519
rect 45845 3485 45879 3519
rect 45879 3485 45888 3519
rect 45836 3476 45888 3485
rect 47952 3519 48004 3528
rect 47952 3485 47961 3519
rect 47961 3485 47995 3519
rect 47995 3485 48004 3519
rect 47952 3476 48004 3485
rect 50068 3519 50120 3528
rect 50068 3485 50077 3519
rect 50077 3485 50111 3519
rect 50111 3485 50120 3519
rect 52184 3519 52236 3528
rect 50068 3476 50120 3485
rect 52184 3485 52193 3519
rect 52193 3485 52227 3519
rect 52227 3485 52236 3519
rect 52184 3476 52236 3485
rect 52276 3476 52328 3528
rect 54300 3519 54352 3528
rect 54300 3485 54309 3519
rect 54309 3485 54343 3519
rect 54343 3485 54352 3519
rect 54300 3476 54352 3485
rect 54668 3476 54720 3528
rect 56416 3519 56468 3528
rect 56416 3485 56425 3519
rect 56425 3485 56459 3519
rect 56459 3485 56468 3519
rect 56416 3476 56468 3485
rect 57152 3476 57204 3528
rect 58532 3519 58584 3528
rect 58532 3485 58541 3519
rect 58541 3485 58575 3519
rect 58575 3485 58584 3519
rect 58532 3476 58584 3485
rect 58992 3476 59044 3528
rect 60648 3519 60700 3528
rect 60648 3485 60657 3519
rect 60657 3485 60691 3519
rect 60691 3485 60700 3519
rect 60648 3476 60700 3485
rect 61292 3476 61344 3528
rect 62764 3519 62816 3528
rect 62764 3485 62773 3519
rect 62773 3485 62807 3519
rect 62807 3485 62816 3519
rect 62764 3476 62816 3485
rect 64880 3519 64932 3528
rect 64880 3485 64889 3519
rect 64889 3485 64923 3519
rect 64923 3485 64932 3519
rect 64880 3476 64932 3485
rect 66996 3519 67048 3528
rect 66996 3485 67005 3519
rect 67005 3485 67039 3519
rect 67039 3485 67048 3519
rect 66996 3476 67048 3485
rect 69112 3519 69164 3528
rect 69112 3485 69121 3519
rect 69121 3485 69155 3519
rect 69155 3485 69164 3519
rect 69112 3476 69164 3485
rect 69204 3476 69256 3528
rect 71228 3519 71280 3528
rect 71228 3485 71237 3519
rect 71237 3485 71271 3519
rect 71271 3485 71280 3519
rect 71228 3476 71280 3485
rect 71688 3476 71740 3528
rect 73344 3519 73396 3528
rect 73344 3485 73353 3519
rect 73353 3485 73387 3519
rect 73387 3485 73396 3519
rect 73344 3476 73396 3485
rect 73712 3476 73764 3528
rect 75368 3476 75420 3528
rect 77392 3544 77444 3596
rect 79416 3587 79468 3596
rect 79416 3553 79425 3587
rect 79425 3553 79459 3587
rect 79459 3553 79468 3587
rect 79416 3544 79468 3553
rect 81532 3587 81584 3596
rect 81532 3553 81541 3587
rect 81541 3553 81575 3587
rect 81575 3553 81584 3587
rect 81532 3544 81584 3553
rect 83648 3587 83700 3596
rect 83648 3553 83657 3587
rect 83657 3553 83691 3587
rect 83691 3553 83700 3587
rect 83648 3544 83700 3553
rect 85764 3587 85816 3596
rect 85764 3553 85773 3587
rect 85773 3553 85807 3587
rect 85807 3553 85816 3587
rect 85764 3544 85816 3553
rect 75828 3476 75880 3528
rect 77300 3519 77352 3528
rect 77300 3485 77309 3519
rect 77309 3485 77343 3519
rect 77343 3485 77352 3519
rect 77576 3519 77628 3528
rect 77300 3476 77352 3485
rect 77576 3485 77585 3519
rect 77585 3485 77619 3519
rect 77619 3485 77628 3519
rect 77576 3476 77628 3485
rect 79692 3519 79744 3528
rect 79692 3485 79701 3519
rect 79701 3485 79735 3519
rect 79735 3485 79744 3519
rect 79692 3476 79744 3485
rect 81808 3519 81860 3528
rect 81808 3485 81817 3519
rect 81817 3485 81851 3519
rect 81851 3485 81860 3519
rect 81808 3476 81860 3485
rect 83924 3519 83976 3528
rect 83924 3485 83933 3519
rect 83933 3485 83967 3519
rect 83967 3485 83976 3519
rect 83924 3476 83976 3485
rect 85948 3476 86000 3528
rect 87052 3544 87104 3596
rect 87880 3587 87932 3596
rect 87880 3553 87889 3587
rect 87889 3553 87923 3587
rect 87923 3553 87932 3587
rect 87880 3544 87932 3553
rect 89996 3587 90048 3596
rect 89996 3553 90005 3587
rect 90005 3553 90039 3587
rect 90039 3553 90048 3587
rect 89996 3544 90048 3553
rect 92112 3587 92164 3596
rect 92112 3553 92121 3587
rect 92121 3553 92155 3587
rect 92155 3553 92164 3587
rect 92112 3544 92164 3553
rect 94228 3587 94280 3596
rect 94228 3553 94237 3587
rect 94237 3553 94271 3587
rect 94271 3553 94280 3587
rect 94228 3544 94280 3553
rect 96068 3544 96120 3596
rect 98460 3587 98512 3596
rect 98460 3553 98469 3587
rect 98469 3553 98503 3587
rect 98503 3553 98512 3587
rect 98460 3544 98512 3553
rect 100576 3587 100628 3596
rect 100576 3553 100585 3587
rect 100585 3553 100619 3587
rect 100619 3553 100628 3587
rect 100576 3544 100628 3553
rect 102692 3587 102744 3596
rect 102692 3553 102701 3587
rect 102701 3553 102735 3587
rect 102735 3553 102744 3587
rect 102692 3544 102744 3553
rect 104808 3587 104860 3596
rect 104808 3553 104817 3587
rect 104817 3553 104851 3587
rect 104851 3553 104860 3587
rect 104808 3544 104860 3553
rect 86132 3476 86184 3528
rect 88156 3519 88208 3528
rect 88156 3485 88165 3519
rect 88165 3485 88199 3519
rect 88199 3485 88208 3519
rect 88156 3476 88208 3485
rect 88524 3476 88576 3528
rect 90272 3519 90324 3528
rect 90272 3485 90281 3519
rect 90281 3485 90315 3519
rect 90315 3485 90324 3519
rect 90272 3476 90324 3485
rect 90640 3476 90692 3528
rect 92388 3519 92440 3528
rect 92388 3485 92397 3519
rect 92397 3485 92431 3519
rect 92431 3485 92440 3519
rect 92388 3476 92440 3485
rect 93124 3476 93176 3528
rect 94504 3519 94556 3528
rect 94504 3485 94513 3519
rect 94513 3485 94547 3519
rect 94547 3485 94556 3519
rect 94504 3476 94556 3485
rect 96620 3519 96672 3528
rect 96620 3485 96629 3519
rect 96629 3485 96663 3519
rect 96663 3485 96672 3519
rect 96620 3476 96672 3485
rect 97264 3476 97316 3528
rect 98736 3519 98788 3528
rect 98736 3485 98745 3519
rect 98745 3485 98779 3519
rect 98779 3485 98788 3519
rect 98736 3476 98788 3485
rect 100852 3519 100904 3528
rect 100852 3485 100861 3519
rect 100861 3485 100895 3519
rect 100895 3485 100904 3519
rect 100852 3476 100904 3485
rect 102968 3519 103020 3528
rect 102968 3485 102977 3519
rect 102977 3485 103011 3519
rect 103011 3485 103020 3519
rect 102968 3476 103020 3485
rect 103612 3476 103664 3528
rect 105084 3519 105136 3528
rect 105084 3485 105093 3519
rect 105093 3485 105127 3519
rect 105127 3485 105136 3519
rect 105084 3476 105136 3485
rect 105452 3476 105504 3528
rect 4042 3238 4094 3290
rect 4106 3238 4158 3290
rect 4170 3238 4222 3290
rect 4234 3238 4286 3290
rect 34762 3238 34814 3290
rect 34826 3238 34878 3290
rect 34890 3238 34942 3290
rect 34954 3238 35006 3290
rect 65482 3238 65534 3290
rect 65546 3238 65598 3290
rect 65610 3238 65662 3290
rect 65674 3238 65726 3290
rect 96202 3238 96254 3290
rect 96266 3238 96318 3290
rect 96330 3238 96382 3290
rect 96394 3238 96446 3290
rect 1308 3136 1360 3188
rect 40408 3136 40460 3188
rect 77392 3179 77444 3188
rect 77392 3145 77401 3179
rect 77401 3145 77435 3179
rect 77435 3145 77444 3179
rect 77392 3136 77444 3145
rect 87052 3136 87104 3188
rect 1400 2932 1452 2984
rect 3516 2932 3568 2984
rect 5632 2932 5684 2984
rect 7748 2932 7800 2984
rect 9864 2932 9916 2984
rect 11980 2932 12032 2984
rect 14096 2932 14148 2984
rect 16212 2864 16264 2916
rect 18328 2932 18380 2984
rect 20444 2932 20496 2984
rect 22560 2932 22612 2984
rect 24676 2932 24728 2984
rect 26792 2932 26844 2984
rect 28908 2932 28960 2984
rect 31024 2932 31076 2984
rect 33140 2864 33192 2916
rect 35256 2932 35308 2984
rect 37372 2932 37424 2984
rect 39488 2932 39540 2984
rect 41604 2932 41656 2984
rect 43720 2932 43772 2984
rect 45836 2932 45888 2984
rect 47952 2932 48004 2984
rect 52184 2932 52236 2984
rect 54300 2932 54352 2984
rect 56416 2932 56468 2984
rect 58532 2932 58584 2984
rect 60648 2932 60700 2984
rect 62764 2932 62816 2984
rect 64880 2932 64932 2984
rect 50068 2864 50120 2916
rect 66996 2864 67048 2916
rect 69112 2932 69164 2984
rect 71228 2932 71280 2984
rect 73344 2932 73396 2984
rect 75368 2975 75420 2984
rect 75368 2941 75377 2975
rect 75377 2941 75411 2975
rect 75411 2941 75420 2975
rect 75368 2932 75420 2941
rect 77576 2932 77628 2984
rect 79692 2932 79744 2984
rect 81808 2932 81860 2984
rect 83924 2864 83976 2916
rect 85948 2975 86000 2984
rect 85948 2941 85957 2975
rect 85957 2941 85991 2975
rect 85991 2941 86000 2975
rect 85948 2932 86000 2941
rect 88156 2932 88208 2984
rect 90272 2932 90324 2984
rect 92388 2932 92440 2984
rect 94504 2932 94556 2984
rect 96620 2932 96672 2984
rect 98736 2932 98788 2984
rect 100852 2932 100904 2984
rect 102968 2932 103020 2984
rect 105084 2932 105136 2984
rect 19402 2694 19454 2746
rect 19466 2694 19518 2746
rect 19530 2694 19582 2746
rect 19594 2694 19646 2746
rect 50122 2694 50174 2746
rect 50186 2694 50238 2746
rect 50250 2694 50302 2746
rect 50314 2694 50366 2746
rect 80842 2694 80894 2746
rect 80906 2694 80958 2746
rect 80970 2694 81022 2746
rect 81034 2694 81086 2746
rect 7748 2524 7800 2576
rect 11888 2524 11940 2576
rect 14096 2524 14148 2576
rect 22376 2567 22428 2576
rect 22376 2533 22385 2567
rect 22385 2533 22419 2567
rect 22419 2533 22428 2567
rect 22376 2524 22428 2533
rect 23388 2592 23440 2644
rect 23756 2592 23808 2644
rect 24676 2524 24728 2576
rect 33140 2592 33192 2644
rect 37372 2524 37424 2576
rect 43720 2524 43772 2576
rect 47860 2524 47912 2576
rect 58440 2524 58492 2576
rect 60464 2567 60516 2576
rect 60464 2533 60473 2567
rect 60473 2533 60507 2567
rect 60507 2533 60516 2567
rect 60464 2524 60516 2533
rect 62764 2524 62816 2576
rect 73344 2524 73396 2576
rect 79600 2524 79652 2576
rect 90272 2524 90324 2576
rect 94412 2524 94464 2576
rect 96620 2524 96672 2576
rect 98736 2524 98788 2576
rect 104900 2567 104952 2576
rect 104900 2533 104909 2567
rect 104909 2533 104943 2567
rect 104943 2533 104952 2567
rect 104900 2524 104952 2533
rect 105084 2567 105136 2576
rect 105084 2533 105093 2567
rect 105093 2533 105127 2567
rect 105127 2533 105136 2567
rect 105084 2524 105136 2533
rect 1216 2499 1268 2508
rect 1216 2465 1225 2499
rect 1225 2465 1259 2499
rect 1259 2465 1268 2499
rect 1216 2456 1268 2465
rect 3516 2456 3568 2508
rect 5632 2456 5684 2508
rect 9864 2388 9916 2440
rect 16212 2456 16264 2508
rect 20444 2456 20496 2508
rect 26700 2388 26752 2440
rect 31024 2456 31076 2508
rect 35256 2456 35308 2508
rect 28816 2388 28868 2440
rect 39396 2388 39448 2440
rect 18328 2320 18380 2372
rect 41604 2456 41656 2508
rect 50068 2456 50120 2508
rect 45836 2388 45888 2440
rect 54208 2456 54260 2508
rect 56416 2388 56468 2440
rect 64788 2456 64840 2508
rect 66996 2456 67048 2508
rect 52184 2320 52236 2372
rect 71228 2456 71280 2508
rect 75460 2388 75512 2440
rect 69112 2320 69164 2372
rect 81716 2456 81768 2508
rect 83924 2456 83976 2508
rect 88156 2388 88208 2440
rect 92388 2388 92440 2440
rect 100852 2456 100904 2508
rect 85948 2320 86000 2372
rect 102968 2320 103020 2372
rect 77576 2252 77628 2304
rect 4042 2150 4094 2202
rect 4106 2150 4158 2202
rect 4170 2150 4222 2202
rect 4234 2150 4286 2202
rect 34762 2150 34814 2202
rect 34826 2150 34878 2202
rect 34890 2150 34942 2202
rect 34954 2150 35006 2202
rect 65482 2150 65534 2202
rect 65546 2150 65598 2202
rect 65610 2150 65662 2202
rect 65674 2150 65726 2202
rect 96202 2150 96254 2202
rect 96266 2150 96318 2202
rect 96330 2150 96382 2202
rect 96394 2150 96446 2202
rect 22652 2048 22704 2100
rect 23664 2048 23716 2100
rect 24768 2048 24820 2100
rect 25780 2048 25832 2100
rect 58624 2048 58676 2100
rect 59636 2048 59688 2100
rect 77668 2048 77720 2100
rect 78772 2048 78824 2100
rect 80336 2048 80388 2100
rect 81164 2048 81216 2100
rect 96712 2048 96764 2100
rect 97908 2048 97960 2100
rect 80612 1980 80664 2032
rect 81348 1980 81400 2032
rect 1124 1955 1176 1964
rect 1124 1921 1133 1955
rect 1133 1921 1167 1955
rect 1167 1921 1176 1955
rect 1124 1912 1176 1921
rect 3240 1955 3292 1964
rect 3240 1921 3249 1955
rect 3249 1921 3283 1955
rect 3283 1921 3292 1955
rect 3240 1912 3292 1921
rect 3516 1955 3568 1964
rect 3516 1921 3525 1955
rect 3525 1921 3559 1955
rect 3559 1921 3568 1955
rect 3516 1912 3568 1921
rect 3608 1912 3660 1964
rect 4620 1912 4672 1964
rect 5356 1955 5408 1964
rect 5356 1921 5365 1955
rect 5365 1921 5399 1955
rect 5399 1921 5408 1955
rect 5356 1912 5408 1921
rect 5632 1955 5684 1964
rect 5632 1921 5641 1955
rect 5641 1921 5675 1955
rect 5675 1921 5684 1955
rect 5632 1912 5684 1921
rect 7472 1955 7524 1964
rect 7472 1921 7481 1955
rect 7481 1921 7515 1955
rect 7515 1921 7524 1955
rect 7472 1912 7524 1921
rect 7748 1955 7800 1964
rect 7748 1921 7757 1955
rect 7757 1921 7791 1955
rect 7791 1921 7800 1955
rect 7748 1912 7800 1921
rect 7840 1912 7892 1964
rect 8852 1912 8904 1964
rect 9588 1955 9640 1964
rect 9588 1921 9597 1955
rect 9597 1921 9631 1955
rect 9631 1921 9640 1955
rect 9588 1912 9640 1921
rect 9864 1955 9916 1964
rect 9864 1921 9873 1955
rect 9873 1921 9907 1955
rect 9907 1921 9916 1955
rect 9864 1912 9916 1921
rect 9956 1912 10008 1964
rect 11152 1912 11204 1964
rect 11704 1955 11756 1964
rect 11704 1921 11713 1955
rect 11713 1921 11747 1955
rect 11747 1921 11756 1955
rect 11704 1912 11756 1921
rect 11888 1912 11940 1964
rect 12072 1912 12124 1964
rect 13268 1912 13320 1964
rect 13820 1955 13872 1964
rect 13820 1921 13829 1955
rect 13829 1921 13863 1955
rect 13863 1921 13872 1955
rect 13820 1912 13872 1921
rect 14096 1955 14148 1964
rect 14096 1921 14105 1955
rect 14105 1921 14139 1955
rect 14139 1921 14148 1955
rect 14096 1912 14148 1921
rect 15936 1955 15988 1964
rect 15936 1921 15945 1955
rect 15945 1921 15979 1955
rect 15979 1921 15988 1955
rect 15936 1912 15988 1921
rect 16212 1955 16264 1964
rect 16212 1921 16221 1955
rect 16221 1921 16255 1955
rect 16255 1921 16264 1955
rect 16212 1912 16264 1921
rect 18052 1955 18104 1964
rect 18052 1921 18061 1955
rect 18061 1921 18095 1955
rect 18095 1921 18104 1955
rect 18052 1912 18104 1921
rect 18328 1955 18380 1964
rect 18328 1921 18337 1955
rect 18337 1921 18371 1955
rect 18371 1921 18380 1955
rect 18328 1912 18380 1921
rect 20168 1955 20220 1964
rect 20168 1921 20177 1955
rect 20177 1921 20211 1955
rect 20211 1921 20220 1955
rect 20168 1912 20220 1921
rect 20444 1955 20496 1964
rect 20444 1921 20453 1955
rect 20453 1921 20487 1955
rect 20487 1921 20496 1955
rect 20444 1912 20496 1921
rect 22192 1912 22244 1964
rect 24400 1955 24452 1964
rect 24400 1921 24409 1955
rect 24409 1921 24443 1955
rect 24443 1921 24452 1955
rect 24400 1912 24452 1921
rect 24676 1955 24728 1964
rect 24676 1921 24685 1955
rect 24685 1921 24719 1955
rect 24719 1921 24728 1955
rect 24676 1912 24728 1921
rect 26516 1955 26568 1964
rect 26516 1921 26525 1955
rect 26525 1921 26559 1955
rect 26559 1921 26568 1955
rect 26516 1912 26568 1921
rect 26700 1912 26752 1964
rect 28632 1955 28684 1964
rect 28632 1921 28641 1955
rect 28641 1921 28675 1955
rect 28675 1921 28684 1955
rect 28632 1912 28684 1921
rect 28816 1912 28868 1964
rect 29000 1912 29052 1964
rect 30196 1912 30248 1964
rect 30748 1955 30800 1964
rect 30748 1921 30757 1955
rect 30757 1921 30791 1955
rect 30791 1921 30800 1955
rect 30748 1912 30800 1921
rect 31024 1955 31076 1964
rect 31024 1921 31033 1955
rect 31033 1921 31067 1955
rect 31067 1921 31076 1955
rect 31024 1912 31076 1921
rect 32864 1955 32916 1964
rect 32864 1921 32873 1955
rect 32873 1921 32907 1955
rect 32907 1921 32916 1955
rect 32864 1912 32916 1921
rect 33140 1955 33192 1964
rect 33140 1921 33149 1955
rect 33149 1921 33183 1955
rect 33183 1921 33192 1955
rect 33140 1912 33192 1921
rect 35256 1955 35308 1964
rect 35256 1921 35265 1955
rect 35265 1921 35299 1955
rect 35299 1921 35308 1955
rect 35256 1912 35308 1921
rect 37096 1955 37148 1964
rect 37096 1921 37105 1955
rect 37105 1921 37139 1955
rect 37139 1921 37148 1955
rect 37096 1912 37148 1921
rect 37372 1955 37424 1964
rect 37372 1921 37381 1955
rect 37381 1921 37415 1955
rect 37415 1921 37424 1955
rect 37372 1912 37424 1921
rect 39212 1955 39264 1964
rect 39212 1921 39221 1955
rect 39221 1921 39255 1955
rect 39255 1921 39264 1955
rect 39212 1912 39264 1921
rect 39396 1912 39448 1964
rect 39580 1912 39632 1964
rect 40684 1912 40736 1964
rect 41328 1955 41380 1964
rect 41328 1921 41337 1955
rect 41337 1921 41371 1955
rect 41371 1921 41380 1955
rect 41328 1912 41380 1921
rect 41604 1955 41656 1964
rect 41604 1921 41613 1955
rect 41613 1921 41647 1955
rect 41647 1921 41656 1955
rect 41604 1912 41656 1921
rect 41696 1912 41748 1964
rect 42708 1912 42760 1964
rect 43444 1955 43496 1964
rect 43444 1921 43453 1955
rect 43453 1921 43487 1955
rect 43487 1921 43496 1955
rect 43444 1912 43496 1921
rect 43720 1955 43772 1964
rect 43720 1921 43729 1955
rect 43729 1921 43763 1955
rect 43763 1921 43772 1955
rect 43720 1912 43772 1921
rect 43812 1912 43864 1964
rect 45008 1912 45060 1964
rect 45560 1955 45612 1964
rect 45560 1921 45569 1955
rect 45569 1921 45603 1955
rect 45603 1921 45612 1955
rect 45560 1912 45612 1921
rect 45836 1955 45888 1964
rect 45836 1921 45845 1955
rect 45845 1921 45879 1955
rect 45879 1921 45888 1955
rect 45836 1912 45888 1921
rect 45928 1912 45980 1964
rect 47124 1912 47176 1964
rect 47676 1955 47728 1964
rect 47676 1921 47685 1955
rect 47685 1921 47719 1955
rect 47719 1921 47728 1955
rect 47676 1912 47728 1921
rect 47860 1912 47912 1964
rect 49792 1955 49844 1964
rect 49792 1921 49801 1955
rect 49801 1921 49835 1955
rect 49835 1921 49844 1955
rect 49792 1912 49844 1921
rect 50068 1955 50120 1964
rect 50068 1921 50077 1955
rect 50077 1921 50111 1955
rect 50111 1921 50120 1955
rect 51908 1955 51960 1964
rect 50068 1912 50120 1921
rect 51908 1921 51917 1955
rect 51917 1921 51951 1955
rect 51951 1921 51960 1955
rect 51908 1912 51960 1921
rect 52184 1955 52236 1964
rect 52184 1921 52193 1955
rect 52193 1921 52227 1955
rect 52227 1921 52236 1955
rect 52184 1912 52236 1921
rect 54024 1955 54076 1964
rect 54024 1921 54033 1955
rect 54033 1921 54067 1955
rect 54067 1921 54076 1955
rect 54024 1912 54076 1921
rect 54208 1912 54260 1964
rect 54392 1912 54444 1964
rect 55404 1912 55456 1964
rect 56140 1955 56192 1964
rect 56140 1921 56149 1955
rect 56149 1921 56183 1955
rect 56183 1921 56192 1955
rect 56140 1912 56192 1921
rect 56416 1955 56468 1964
rect 56416 1921 56425 1955
rect 56425 1921 56459 1955
rect 56459 1921 56468 1955
rect 56416 1912 56468 1921
rect 58256 1955 58308 1964
rect 58256 1921 58265 1955
rect 58265 1921 58299 1955
rect 58299 1921 58308 1955
rect 58256 1912 58308 1921
rect 58440 1912 58492 1964
rect 60372 1955 60424 1964
rect 60372 1921 60381 1955
rect 60381 1921 60415 1955
rect 60415 1921 60424 1955
rect 62488 1955 62540 1964
rect 60372 1912 60424 1921
rect 62488 1921 62497 1955
rect 62497 1921 62531 1955
rect 62531 1921 62540 1955
rect 62488 1912 62540 1921
rect 62764 1955 62816 1964
rect 62764 1921 62773 1955
rect 62773 1921 62807 1955
rect 62807 1921 62816 1955
rect 62764 1912 62816 1921
rect 62856 1912 62908 1964
rect 64052 1912 64104 1964
rect 64604 1955 64656 1964
rect 64604 1921 64613 1955
rect 64613 1921 64647 1955
rect 64647 1921 64656 1955
rect 64604 1912 64656 1921
rect 64788 1912 64840 1964
rect 66720 1955 66772 1964
rect 66720 1921 66729 1955
rect 66729 1921 66763 1955
rect 66763 1921 66772 1955
rect 66720 1912 66772 1921
rect 66996 1955 67048 1964
rect 66996 1921 67005 1955
rect 67005 1921 67039 1955
rect 67039 1921 67048 1955
rect 66996 1912 67048 1921
rect 68836 1955 68888 1964
rect 68836 1921 68845 1955
rect 68845 1921 68879 1955
rect 68879 1921 68888 1955
rect 68836 1912 68888 1921
rect 69112 1955 69164 1964
rect 69112 1921 69121 1955
rect 69121 1921 69155 1955
rect 69155 1921 69164 1955
rect 69112 1912 69164 1921
rect 70952 1955 71004 1964
rect 70952 1921 70961 1955
rect 70961 1921 70995 1955
rect 70995 1921 71004 1955
rect 70952 1912 71004 1921
rect 71228 1955 71280 1964
rect 71228 1921 71237 1955
rect 71237 1921 71271 1955
rect 71271 1921 71280 1955
rect 71228 1912 71280 1921
rect 73068 1955 73120 1964
rect 73068 1921 73077 1955
rect 73077 1921 73111 1955
rect 73111 1921 73120 1955
rect 73068 1912 73120 1921
rect 73344 1955 73396 1964
rect 73344 1921 73353 1955
rect 73353 1921 73387 1955
rect 73387 1921 73396 1955
rect 73344 1912 73396 1921
rect 75184 1955 75236 1964
rect 75184 1921 75193 1955
rect 75193 1921 75227 1955
rect 75227 1921 75236 1955
rect 75184 1912 75236 1921
rect 75460 1955 75512 1964
rect 75460 1921 75469 1955
rect 75469 1921 75503 1955
rect 75503 1921 75512 1955
rect 75460 1912 75512 1921
rect 75552 1912 75604 1964
rect 76748 1912 76800 1964
rect 77576 1955 77628 1964
rect 77576 1921 77585 1955
rect 77585 1921 77619 1955
rect 77619 1921 77628 1955
rect 77576 1912 77628 1921
rect 78220 1912 78272 1964
rect 78864 1912 78916 1964
rect 79416 1955 79468 1964
rect 79416 1921 79425 1955
rect 79425 1921 79459 1955
rect 79459 1921 79468 1955
rect 79416 1912 79468 1921
rect 79600 1912 79652 1964
rect 79784 1912 79836 1964
rect 81256 1912 81308 1964
rect 81532 1955 81584 1964
rect 81532 1921 81541 1955
rect 81541 1921 81575 1955
rect 81575 1921 81584 1955
rect 81532 1912 81584 1921
rect 81716 1912 81768 1964
rect 83648 1955 83700 1964
rect 83648 1921 83657 1955
rect 83657 1921 83691 1955
rect 83691 1921 83700 1955
rect 83648 1912 83700 1921
rect 83924 1955 83976 1964
rect 83924 1921 83933 1955
rect 83933 1921 83967 1955
rect 83967 1921 83976 1955
rect 83924 1912 83976 1921
rect 85764 1955 85816 1964
rect 85764 1921 85773 1955
rect 85773 1921 85807 1955
rect 85807 1921 85816 1955
rect 85764 1912 85816 1921
rect 85948 1912 86000 1964
rect 87880 1955 87932 1964
rect 87880 1921 87889 1955
rect 87889 1921 87923 1955
rect 87923 1921 87932 1955
rect 87880 1912 87932 1921
rect 88156 1955 88208 1964
rect 88156 1921 88165 1955
rect 88165 1921 88199 1955
rect 88199 1921 88208 1955
rect 88156 1912 88208 1921
rect 88800 1912 88852 1964
rect 89260 1912 89312 1964
rect 89996 1955 90048 1964
rect 89996 1921 90005 1955
rect 90005 1921 90039 1955
rect 90039 1921 90048 1955
rect 89996 1912 90048 1921
rect 90272 1955 90324 1964
rect 90272 1921 90281 1955
rect 90281 1921 90315 1955
rect 90315 1921 90324 1955
rect 90272 1912 90324 1921
rect 90364 1912 90416 1964
rect 91376 1912 91428 1964
rect 92112 1955 92164 1964
rect 92112 1921 92121 1955
rect 92121 1921 92155 1955
rect 92155 1921 92164 1955
rect 92112 1912 92164 1921
rect 92388 1955 92440 1964
rect 92388 1921 92397 1955
rect 92397 1921 92431 1955
rect 92431 1921 92440 1955
rect 92388 1912 92440 1921
rect 92480 1912 92532 1964
rect 93492 1912 93544 1964
rect 94228 1955 94280 1964
rect 94228 1921 94237 1955
rect 94237 1921 94271 1955
rect 94271 1921 94280 1955
rect 94228 1912 94280 1921
rect 94412 1912 94464 1964
rect 95148 1912 95200 1964
rect 95792 1912 95844 1964
rect 96068 1912 96120 1964
rect 96620 1955 96672 1964
rect 96620 1921 96629 1955
rect 96629 1921 96663 1955
rect 96663 1921 96672 1955
rect 96620 1912 96672 1921
rect 97264 1912 97316 1964
rect 98000 1912 98052 1964
rect 98460 1955 98512 1964
rect 98460 1921 98469 1955
rect 98469 1921 98503 1955
rect 98503 1921 98512 1955
rect 98460 1912 98512 1921
rect 98736 1955 98788 1964
rect 98736 1921 98745 1955
rect 98745 1921 98779 1955
rect 98779 1921 98788 1955
rect 98736 1912 98788 1921
rect 100576 1955 100628 1964
rect 100576 1921 100585 1955
rect 100585 1921 100619 1955
rect 100619 1921 100628 1955
rect 100576 1912 100628 1921
rect 100852 1955 100904 1964
rect 100852 1921 100861 1955
rect 100861 1921 100895 1955
rect 100895 1921 100904 1955
rect 100852 1912 100904 1921
rect 102692 1955 102744 1964
rect 102692 1921 102701 1955
rect 102701 1921 102735 1955
rect 102735 1921 102744 1955
rect 102692 1912 102744 1921
rect 102968 1955 103020 1964
rect 102968 1921 102977 1955
rect 102977 1921 103011 1955
rect 103011 1921 103020 1955
rect 102968 1912 103020 1921
rect 104808 1955 104860 1964
rect 104808 1921 104817 1955
rect 104817 1921 104851 1955
rect 104851 1921 104860 1955
rect 104808 1912 104860 1921
rect 1216 1844 1268 1896
rect 5724 1844 5776 1896
rect 6736 1844 6788 1896
rect 10784 1844 10836 1896
rect 11244 1844 11296 1896
rect 18420 1844 18472 1896
rect 18696 1844 18748 1896
rect 20536 1844 20588 1896
rect 21548 1844 21600 1896
rect 22376 1844 22428 1896
rect 26884 1844 26936 1896
rect 28080 1844 28132 1896
rect 35072 1844 35124 1896
rect 37464 1844 37516 1896
rect 38476 1844 38528 1896
rect 56508 1844 56560 1896
rect 57520 1844 57572 1896
rect 60464 1844 60516 1896
rect 60740 1844 60792 1896
rect 61936 1844 61988 1896
rect 71320 1844 71372 1896
rect 72332 1844 72384 1896
rect 73436 1844 73488 1896
rect 74448 1844 74500 1896
rect 77300 1887 77352 1896
rect 77300 1853 77309 1887
rect 77309 1853 77343 1887
rect 77343 1853 77352 1887
rect 77300 1844 77352 1853
rect 78496 1844 78548 1896
rect 78956 1844 79008 1896
rect 88248 1844 88300 1896
rect 89444 1844 89496 1896
rect 93032 1844 93084 1896
rect 93676 1844 93728 1896
rect 94596 1844 94648 1896
rect 95700 1844 95752 1896
rect 97540 1844 97592 1896
rect 98092 1844 98144 1896
rect 104900 1844 104952 1896
rect 81164 1776 81216 1828
rect 95424 1776 95476 1828
rect 95884 1776 95936 1828
rect 2504 1751 2556 1760
rect 2504 1717 2513 1751
rect 2513 1717 2547 1751
rect 2547 1717 2556 1751
rect 2504 1708 2556 1717
rect 4160 1708 4212 1760
rect 5908 1708 5960 1760
rect 8208 1708 8260 1760
rect 11152 1751 11204 1760
rect 11152 1717 11161 1751
rect 11161 1717 11195 1751
rect 11195 1717 11204 1751
rect 11152 1708 11204 1717
rect 13268 1751 13320 1760
rect 13268 1717 13277 1751
rect 13277 1717 13311 1751
rect 13311 1717 13320 1751
rect 13268 1708 13320 1717
rect 15200 1751 15252 1760
rect 15200 1717 15209 1751
rect 15209 1717 15243 1751
rect 15243 1717 15252 1751
rect 15200 1708 15252 1717
rect 17316 1751 17368 1760
rect 17316 1717 17325 1751
rect 17325 1717 17359 1751
rect 17359 1717 17368 1751
rect 17316 1708 17368 1717
rect 18696 1708 18748 1760
rect 20720 1708 20772 1760
rect 22836 1708 22888 1760
rect 25044 1708 25096 1760
rect 28080 1751 28132 1760
rect 28080 1717 28089 1751
rect 28089 1717 28123 1751
rect 28123 1717 28132 1751
rect 28080 1708 28132 1717
rect 30196 1751 30248 1760
rect 30196 1717 30205 1751
rect 30205 1717 30239 1751
rect 30239 1717 30248 1751
rect 30196 1708 30248 1717
rect 32128 1751 32180 1760
rect 32128 1717 32137 1751
rect 32137 1717 32171 1751
rect 32171 1717 32180 1751
rect 32128 1708 32180 1717
rect 34244 1751 34296 1760
rect 34244 1717 34253 1751
rect 34253 1717 34287 1751
rect 34287 1717 34296 1751
rect 34244 1708 34296 1717
rect 35532 1708 35584 1760
rect 37648 1708 37700 1760
rect 40132 1708 40184 1760
rect 41972 1708 42024 1760
rect 45008 1751 45060 1760
rect 45008 1717 45017 1751
rect 45017 1717 45051 1751
rect 45051 1717 45060 1751
rect 45008 1708 45060 1717
rect 47124 1751 47176 1760
rect 47124 1717 47133 1751
rect 47133 1717 47167 1751
rect 47167 1717 47176 1751
rect 47124 1708 47176 1717
rect 49056 1751 49108 1760
rect 49056 1717 49065 1751
rect 49065 1717 49099 1751
rect 49099 1717 49108 1751
rect 49056 1708 49108 1717
rect 51172 1751 51224 1760
rect 51172 1717 51181 1751
rect 51181 1717 51215 1751
rect 51215 1717 51224 1751
rect 51172 1708 51224 1717
rect 52276 1708 52328 1760
rect 54760 1708 54812 1760
rect 56692 1708 56744 1760
rect 58900 1708 58952 1760
rect 61936 1751 61988 1760
rect 61936 1717 61945 1751
rect 61945 1717 61979 1751
rect 61979 1717 61988 1751
rect 61936 1708 61988 1717
rect 64052 1751 64104 1760
rect 64052 1717 64061 1751
rect 64061 1717 64095 1751
rect 64095 1717 64104 1751
rect 64052 1708 64104 1717
rect 65984 1751 66036 1760
rect 65984 1717 65993 1751
rect 65993 1717 66027 1751
rect 66027 1717 66036 1751
rect 65984 1708 66036 1717
rect 68100 1751 68152 1760
rect 68100 1717 68109 1751
rect 68109 1717 68143 1751
rect 68143 1717 68152 1751
rect 68100 1708 68152 1717
rect 69204 1708 69256 1760
rect 71504 1708 71556 1760
rect 73620 1708 73672 1760
rect 76196 1708 76248 1760
rect 78864 1751 78916 1760
rect 78864 1717 78873 1751
rect 78873 1717 78907 1751
rect 78907 1717 78916 1751
rect 78864 1708 78916 1717
rect 82912 1751 82964 1760
rect 82912 1717 82921 1751
rect 82921 1717 82955 1751
rect 82955 1717 82964 1751
rect 82912 1708 82964 1717
rect 85028 1751 85080 1760
rect 85028 1717 85037 1751
rect 85037 1717 85071 1751
rect 85071 1717 85080 1751
rect 85028 1708 85080 1717
rect 86500 1708 86552 1760
rect 88432 1708 88484 1760
rect 90732 1708 90784 1760
rect 92756 1708 92808 1760
rect 95792 1751 95844 1760
rect 95792 1717 95801 1751
rect 95801 1717 95835 1751
rect 95835 1717 95844 1751
rect 95792 1708 95844 1717
rect 97908 1751 97960 1760
rect 97908 1717 97917 1751
rect 97917 1717 97951 1751
rect 97951 1717 97960 1751
rect 97908 1708 97960 1717
rect 99840 1751 99892 1760
rect 99840 1717 99849 1751
rect 99849 1717 99883 1751
rect 99883 1717 99892 1751
rect 99840 1708 99892 1717
rect 101956 1751 102008 1760
rect 101956 1717 101965 1751
rect 101965 1717 101999 1751
rect 101999 1717 102008 1751
rect 101956 1708 102008 1717
rect 103244 1708 103296 1760
rect 105360 1708 105412 1760
rect 19402 1606 19454 1658
rect 19466 1606 19518 1658
rect 19530 1606 19582 1658
rect 19594 1606 19646 1658
rect 50122 1606 50174 1658
rect 50186 1606 50238 1658
rect 50250 1606 50302 1658
rect 50314 1606 50366 1658
rect 80842 1606 80894 1658
rect 80906 1606 80958 1658
rect 80970 1606 81022 1658
rect 81034 1606 81086 1658
rect 1032 1504 1084 1556
rect 7380 1504 7432 1556
rect 9496 1504 9548 1556
rect 13728 1504 13780 1556
rect 24308 1504 24360 1556
rect 26424 1504 26476 1556
rect 30656 1504 30708 1556
rect 41236 1504 41288 1556
rect 43352 1504 43404 1556
rect 47584 1504 47636 1556
rect 58164 1504 58216 1556
rect 64512 1504 64564 1556
rect 75092 1504 75144 1556
rect 77208 1504 77260 1556
rect 81440 1504 81492 1556
rect 92020 1504 92072 1556
rect 94136 1504 94188 1556
rect 98368 1504 98420 1556
rect 1124 1411 1176 1420
rect 1124 1377 1133 1411
rect 1133 1377 1167 1411
rect 1167 1377 1176 1411
rect 1124 1368 1176 1377
rect 2504 1368 2556 1420
rect 3240 1411 3292 1420
rect 3240 1377 3249 1411
rect 3249 1377 3283 1411
rect 3283 1377 3292 1411
rect 3240 1368 3292 1377
rect 4160 1368 4212 1420
rect 5356 1411 5408 1420
rect 5356 1377 5365 1411
rect 5365 1377 5399 1411
rect 5399 1377 5408 1411
rect 5356 1368 5408 1377
rect 5908 1368 5960 1420
rect 7472 1411 7524 1420
rect 7472 1377 7481 1411
rect 7481 1377 7515 1411
rect 7515 1377 7524 1411
rect 7472 1368 7524 1377
rect 8208 1368 8260 1420
rect 9588 1411 9640 1420
rect 9588 1377 9597 1411
rect 9597 1377 9631 1411
rect 9631 1377 9640 1411
rect 9588 1368 9640 1377
rect 11152 1368 11204 1420
rect 11704 1411 11756 1420
rect 11704 1377 11713 1411
rect 11713 1377 11747 1411
rect 11747 1377 11756 1411
rect 11704 1368 11756 1377
rect 13268 1368 13320 1420
rect 13820 1411 13872 1420
rect 13820 1377 13829 1411
rect 13829 1377 13863 1411
rect 13863 1377 13872 1411
rect 13820 1368 13872 1377
rect 15200 1368 15252 1420
rect 15936 1411 15988 1420
rect 15936 1377 15945 1411
rect 15945 1377 15979 1411
rect 15979 1377 15988 1411
rect 15936 1368 15988 1377
rect 17316 1368 17368 1420
rect 18052 1411 18104 1420
rect 18052 1377 18061 1411
rect 18061 1377 18095 1411
rect 18095 1377 18104 1411
rect 18052 1368 18104 1377
rect 18696 1368 18748 1420
rect 20168 1411 20220 1420
rect 20168 1377 20177 1411
rect 20177 1377 20211 1411
rect 20211 1377 20220 1411
rect 20168 1368 20220 1377
rect 20720 1368 20772 1420
rect 22284 1411 22336 1420
rect 22284 1377 22293 1411
rect 22293 1377 22327 1411
rect 22327 1377 22336 1411
rect 22284 1368 22336 1377
rect 22836 1368 22888 1420
rect 24400 1411 24452 1420
rect 24400 1377 24409 1411
rect 24409 1377 24443 1411
rect 24443 1377 24452 1411
rect 24400 1368 24452 1377
rect 25044 1368 25096 1420
rect 26516 1411 26568 1420
rect 26516 1377 26525 1411
rect 26525 1377 26559 1411
rect 26559 1377 26568 1411
rect 26516 1368 26568 1377
rect 28080 1368 28132 1420
rect 28632 1411 28684 1420
rect 28632 1377 28641 1411
rect 28641 1377 28675 1411
rect 28675 1377 28684 1411
rect 28632 1368 28684 1377
rect 30196 1368 30248 1420
rect 30748 1411 30800 1420
rect 30748 1377 30757 1411
rect 30757 1377 30791 1411
rect 30791 1377 30800 1411
rect 30748 1368 30800 1377
rect 32128 1368 32180 1420
rect 32864 1411 32916 1420
rect 32864 1377 32873 1411
rect 32873 1377 32907 1411
rect 32907 1377 32916 1411
rect 32864 1368 32916 1377
rect 34244 1368 34296 1420
rect 35072 1368 35124 1420
rect 35532 1368 35584 1420
rect 37096 1411 37148 1420
rect 37096 1377 37105 1411
rect 37105 1377 37139 1411
rect 37139 1377 37148 1411
rect 37096 1368 37148 1377
rect 37648 1368 37700 1420
rect 39212 1411 39264 1420
rect 39212 1377 39221 1411
rect 39221 1377 39255 1411
rect 39255 1377 39264 1411
rect 39212 1368 39264 1377
rect 40132 1368 40184 1420
rect 41328 1411 41380 1420
rect 41328 1377 41337 1411
rect 41337 1377 41371 1411
rect 41371 1377 41380 1411
rect 41328 1368 41380 1377
rect 41972 1368 42024 1420
rect 43444 1411 43496 1420
rect 43444 1377 43453 1411
rect 43453 1377 43487 1411
rect 43487 1377 43496 1411
rect 43444 1368 43496 1377
rect 45008 1368 45060 1420
rect 45560 1411 45612 1420
rect 45560 1377 45569 1411
rect 45569 1377 45603 1411
rect 45603 1377 45612 1411
rect 45560 1368 45612 1377
rect 47124 1368 47176 1420
rect 47676 1411 47728 1420
rect 47676 1377 47685 1411
rect 47685 1377 47719 1411
rect 47719 1377 47728 1411
rect 47676 1368 47728 1377
rect 49056 1368 49108 1420
rect 49792 1411 49844 1420
rect 49792 1377 49801 1411
rect 49801 1377 49835 1411
rect 49835 1377 49844 1411
rect 49792 1368 49844 1377
rect 51172 1368 51224 1420
rect 51908 1411 51960 1420
rect 51908 1377 51917 1411
rect 51917 1377 51951 1411
rect 51951 1377 51960 1411
rect 51908 1368 51960 1377
rect 52276 1368 52328 1420
rect 54024 1411 54076 1420
rect 54024 1377 54033 1411
rect 54033 1377 54067 1411
rect 54067 1377 54076 1411
rect 54024 1368 54076 1377
rect 54760 1368 54812 1420
rect 56140 1411 56192 1420
rect 56140 1377 56149 1411
rect 56149 1377 56183 1411
rect 56183 1377 56192 1411
rect 56140 1368 56192 1377
rect 56692 1368 56744 1420
rect 58256 1411 58308 1420
rect 58256 1377 58265 1411
rect 58265 1377 58299 1411
rect 58299 1377 58308 1411
rect 58256 1368 58308 1377
rect 58900 1368 58952 1420
rect 60372 1411 60424 1420
rect 60372 1377 60381 1411
rect 60381 1377 60415 1411
rect 60415 1377 60424 1411
rect 60372 1368 60424 1377
rect 61936 1368 61988 1420
rect 62488 1411 62540 1420
rect 62488 1377 62497 1411
rect 62497 1377 62531 1411
rect 62531 1377 62540 1411
rect 62488 1368 62540 1377
rect 64052 1368 64104 1420
rect 64604 1411 64656 1420
rect 64604 1377 64613 1411
rect 64613 1377 64647 1411
rect 64647 1377 64656 1411
rect 64604 1368 64656 1377
rect 65984 1368 66036 1420
rect 66720 1411 66772 1420
rect 66720 1377 66729 1411
rect 66729 1377 66763 1411
rect 66763 1377 66772 1411
rect 66720 1368 66772 1377
rect 68100 1368 68152 1420
rect 68836 1411 68888 1420
rect 68836 1377 68845 1411
rect 68845 1377 68879 1411
rect 68879 1377 68888 1411
rect 68836 1368 68888 1377
rect 69204 1368 69256 1420
rect 70952 1411 71004 1420
rect 70952 1377 70961 1411
rect 70961 1377 70995 1411
rect 70995 1377 71004 1411
rect 70952 1368 71004 1377
rect 71504 1368 71556 1420
rect 73068 1411 73120 1420
rect 73068 1377 73077 1411
rect 73077 1377 73111 1411
rect 73111 1377 73120 1411
rect 73068 1368 73120 1377
rect 73620 1368 73672 1420
rect 75184 1411 75236 1420
rect 75184 1377 75193 1411
rect 75193 1377 75227 1411
rect 75227 1377 75236 1411
rect 75184 1368 75236 1377
rect 76196 1368 76248 1420
rect 77300 1411 77352 1420
rect 77300 1377 77309 1411
rect 77309 1377 77343 1411
rect 77343 1377 77352 1411
rect 77300 1368 77352 1377
rect 78864 1368 78916 1420
rect 79416 1411 79468 1420
rect 79416 1377 79425 1411
rect 79425 1377 79459 1411
rect 79459 1377 79468 1411
rect 79416 1368 79468 1377
rect 81164 1368 81216 1420
rect 81532 1411 81584 1420
rect 81532 1377 81541 1411
rect 81541 1377 81575 1411
rect 81575 1377 81584 1411
rect 81532 1368 81584 1377
rect 82912 1368 82964 1420
rect 83648 1411 83700 1420
rect 83648 1377 83657 1411
rect 83657 1377 83691 1411
rect 83691 1377 83700 1411
rect 83648 1368 83700 1377
rect 85028 1368 85080 1420
rect 85764 1411 85816 1420
rect 85764 1377 85773 1411
rect 85773 1377 85807 1411
rect 85807 1377 85816 1411
rect 85764 1368 85816 1377
rect 86500 1368 86552 1420
rect 87880 1411 87932 1420
rect 87880 1377 87889 1411
rect 87889 1377 87923 1411
rect 87923 1377 87932 1411
rect 87880 1368 87932 1377
rect 88432 1368 88484 1420
rect 89996 1411 90048 1420
rect 89996 1377 90005 1411
rect 90005 1377 90039 1411
rect 90039 1377 90048 1411
rect 89996 1368 90048 1377
rect 90732 1368 90784 1420
rect 92112 1411 92164 1420
rect 92112 1377 92121 1411
rect 92121 1377 92155 1411
rect 92155 1377 92164 1411
rect 92112 1368 92164 1377
rect 92756 1368 92808 1420
rect 94228 1411 94280 1420
rect 94228 1377 94237 1411
rect 94237 1377 94271 1411
rect 94271 1377 94280 1411
rect 94228 1368 94280 1377
rect 95792 1368 95844 1420
rect 96068 1368 96120 1420
rect 97908 1368 97960 1420
rect 98460 1411 98512 1420
rect 98460 1377 98469 1411
rect 98469 1377 98503 1411
rect 98503 1377 98512 1411
rect 98460 1368 98512 1377
rect 99840 1368 99892 1420
rect 100576 1411 100628 1420
rect 100576 1377 100585 1411
rect 100585 1377 100619 1411
rect 100619 1377 100628 1411
rect 100576 1368 100628 1377
rect 101956 1368 102008 1420
rect 102692 1411 102744 1420
rect 102692 1377 102701 1411
rect 102701 1377 102735 1411
rect 102735 1377 102744 1411
rect 102692 1368 102744 1377
rect 103244 1368 103296 1420
rect 104808 1411 104860 1420
rect 104808 1377 104817 1411
rect 104817 1377 104851 1411
rect 104851 1377 104860 1411
rect 104808 1368 104860 1377
rect 105360 1368 105412 1420
rect 3424 1164 3476 1216
rect 5632 1164 5684 1216
rect 11612 1164 11664 1216
rect 16120 1164 16172 1216
rect 18328 1164 18380 1216
rect 20352 1164 20404 1216
rect 22560 1164 22612 1216
rect 28540 1164 28592 1216
rect 33048 1164 33100 1216
rect 35256 1164 35308 1216
rect 37280 1164 37332 1216
rect 39488 1164 39540 1216
rect 45468 1164 45520 1216
rect 49976 1164 50028 1216
rect 52184 1164 52236 1216
rect 54208 1164 54260 1216
rect 56416 1164 56468 1216
rect 60280 1164 60332 1216
rect 62396 1164 62448 1216
rect 66904 1164 66956 1216
rect 69112 1164 69164 1216
rect 71136 1164 71188 1216
rect 73344 1164 73396 1216
rect 79324 1164 79376 1216
rect 83832 1164 83884 1216
rect 86040 1164 86092 1216
rect 88064 1164 88116 1216
rect 90272 1164 90324 1216
rect 96528 1164 96580 1216
rect 100760 1164 100812 1216
rect 102968 1164 103020 1216
rect 104992 1164 105044 1216
rect 4042 1062 4094 1114
rect 4106 1062 4158 1114
rect 4170 1062 4222 1114
rect 4234 1062 4286 1114
rect 34762 1062 34814 1114
rect 34826 1062 34878 1114
rect 34890 1062 34942 1114
rect 34954 1062 35006 1114
rect 65482 1062 65534 1114
rect 65546 1062 65598 1114
rect 65610 1062 65662 1114
rect 65674 1062 65726 1114
rect 96202 1062 96254 1114
rect 96266 1062 96318 1114
rect 96330 1062 96382 1114
rect 96394 1062 96446 1114
<< metal2 >>
rect 1030 8650 1086 8704
rect 3146 8650 3202 8704
rect 1030 8648 1164 8650
rect 3146 8648 3280 8650
rect 5262 8648 5318 8704
rect 7378 8648 7434 8704
rect 9494 8648 9550 8704
rect 11610 8650 11666 8704
rect 13726 8650 13782 8704
rect 11610 8648 11744 8650
rect 13726 8648 13860 8650
rect 15842 8648 15898 8704
rect 17958 8648 18014 8704
rect 20074 8648 20130 8704
rect 22190 8648 22246 8704
rect 24306 8648 24362 8704
rect 26422 8648 26478 8704
rect 28538 8650 28594 8704
rect 30654 8650 30710 8704
rect 32770 8650 32826 8704
rect 34886 8650 34942 8704
rect 34992 8662 35112 8690
rect 34992 8650 35020 8662
rect 28538 8648 28672 8650
rect 30654 8648 30788 8650
rect 32770 8648 32904 8650
rect 34886 8648 35020 8650
rect 1044 8622 1164 8648
rect 3160 8622 3280 8648
rect 1136 7342 1164 8622
rect 3252 7342 3280 8622
rect 4016 7644 4312 7664
rect 4072 7642 4096 7644
rect 4152 7642 4176 7644
rect 4232 7642 4256 7644
rect 4094 7590 4096 7642
rect 4158 7590 4170 7642
rect 4232 7590 4234 7642
rect 4072 7588 4096 7590
rect 4152 7588 4176 7590
rect 4232 7588 4256 7590
rect 4016 7568 4312 7588
rect 5276 7342 5304 8648
rect 7392 7342 7420 8648
rect 1124 7336 1176 7342
rect 1124 7278 1176 7284
rect 3240 7336 3292 7342
rect 3240 7278 3292 7284
rect 3516 7336 3568 7342
rect 3516 7278 3568 7284
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7748 7336 7800 7342
rect 9508 7324 9536 8648
rect 11624 8622 11744 8648
rect 13740 8622 13860 8648
rect 11716 7342 11744 8622
rect 13832 7342 13860 8622
rect 15856 7426 15884 8648
rect 17972 7426 18000 8648
rect 15856 7398 15976 7426
rect 17972 7398 18092 7426
rect 15948 7342 15976 7398
rect 18064 7342 18092 7398
rect 20088 7342 20116 8648
rect 22204 7342 22232 8648
rect 24320 7426 24348 8648
rect 24320 7398 24440 7426
rect 24412 7342 24440 7398
rect 9588 7336 9640 7342
rect 9508 7296 9588 7324
rect 7748 7278 7800 7284
rect 9588 7278 9640 7284
rect 9864 7336 9916 7342
rect 9864 7278 9916 7284
rect 11704 7336 11756 7342
rect 11704 7278 11756 7284
rect 11980 7336 12032 7342
rect 11980 7278 12032 7284
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 14096 7336 14148 7342
rect 14096 7278 14148 7284
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 16212 7336 16264 7342
rect 16212 7278 16264 7284
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 18328 7336 18380 7342
rect 18328 7278 18380 7284
rect 20076 7336 20128 7342
rect 20076 7278 20128 7284
rect 20444 7336 20496 7342
rect 20444 7278 20496 7284
rect 22192 7336 22244 7342
rect 22192 7278 22244 7284
rect 22560 7336 22612 7342
rect 22560 7278 22612 7284
rect 24400 7336 24452 7342
rect 24400 7278 24452 7284
rect 24676 7336 24728 7342
rect 24676 7278 24728 7284
rect 26436 7290 26464 8648
rect 28552 8622 28672 8648
rect 30668 8622 30788 8648
rect 32784 8622 32904 8648
rect 34900 8622 35020 8648
rect 28644 7342 28672 8622
rect 30760 7342 30788 8622
rect 32876 7342 32904 8622
rect 34736 7644 35032 7664
rect 34792 7642 34816 7644
rect 34872 7642 34896 7644
rect 34952 7642 34976 7644
rect 34814 7590 34816 7642
rect 34878 7590 34890 7642
rect 34952 7590 34954 7642
rect 34792 7588 34816 7590
rect 34872 7588 34896 7590
rect 34952 7588 34976 7590
rect 34736 7568 35032 7588
rect 35084 7342 35112 8662
rect 37002 8650 37058 8704
rect 39118 8650 39174 8704
rect 37002 8648 37136 8650
rect 39118 8648 39252 8650
rect 41234 8648 41290 8704
rect 43350 8648 43406 8704
rect 45466 8650 45522 8704
rect 47582 8650 47638 8704
rect 49698 8650 49754 8704
rect 45466 8648 45600 8650
rect 47582 8648 47716 8650
rect 49698 8648 49832 8650
rect 51814 8648 51870 8704
rect 53930 8648 53986 8704
rect 56046 8648 56102 8704
rect 58162 8648 58218 8704
rect 60278 8648 60334 8704
rect 62394 8648 62450 8704
rect 64510 8648 64566 8704
rect 66626 8650 66682 8704
rect 68742 8650 68798 8704
rect 66626 8648 66760 8650
rect 68742 8648 68876 8650
rect 70858 8648 70914 8704
rect 72974 8648 73030 8704
rect 75090 8648 75146 8704
rect 77206 8648 77262 8704
rect 79322 8648 79378 8704
rect 81438 8648 81494 8704
rect 83554 8648 83610 8704
rect 85670 8648 85726 8704
rect 87786 8648 87842 8704
rect 89902 8648 89958 8704
rect 92018 8648 92074 8704
rect 94134 8648 94190 8704
rect 96080 8662 96200 8690
rect 37016 8622 37136 8648
rect 39132 8622 39252 8648
rect 37108 7342 37136 8622
rect 39224 7342 39252 8622
rect 41248 7342 41276 8648
rect 26516 7336 26568 7342
rect 26436 7284 26516 7290
rect 26436 7278 26568 7284
rect 26792 7336 26844 7342
rect 26792 7278 26844 7284
rect 28632 7336 28684 7342
rect 28632 7278 28684 7284
rect 28908 7336 28960 7342
rect 28908 7278 28960 7284
rect 30748 7336 30800 7342
rect 30748 7278 30800 7284
rect 31024 7336 31076 7342
rect 31024 7278 31076 7284
rect 32864 7336 32916 7342
rect 32864 7278 32916 7284
rect 33140 7336 33192 7342
rect 33140 7278 33192 7284
rect 35072 7336 35124 7342
rect 35072 7278 35124 7284
rect 35256 7336 35308 7342
rect 35256 7278 35308 7284
rect 37096 7336 37148 7342
rect 37096 7278 37148 7284
rect 37372 7336 37424 7342
rect 37372 7278 37424 7284
rect 39212 7336 39264 7342
rect 39212 7278 39264 7284
rect 39488 7336 39540 7342
rect 39488 7278 39540 7284
rect 41236 7336 41288 7342
rect 41236 7278 41288 7284
rect 41604 7336 41656 7342
rect 43364 7324 43392 8648
rect 45480 8622 45600 8648
rect 47596 8622 47716 8648
rect 49712 8622 49832 8648
rect 45572 7342 45600 8622
rect 47688 7342 47716 8622
rect 49804 7342 49832 8622
rect 51828 7426 51856 8648
rect 53944 7426 53972 8648
rect 51828 7398 51948 7426
rect 53944 7398 54064 7426
rect 51920 7342 51948 7398
rect 54036 7342 54064 7398
rect 56060 7342 56088 8648
rect 58176 7342 58204 8648
rect 43444 7336 43496 7342
rect 43364 7296 43444 7324
rect 41604 7278 41656 7284
rect 43444 7278 43496 7284
rect 43720 7336 43772 7342
rect 43720 7278 43772 7284
rect 45560 7336 45612 7342
rect 45560 7278 45612 7284
rect 45836 7336 45888 7342
rect 45836 7278 45888 7284
rect 47676 7336 47728 7342
rect 47676 7278 47728 7284
rect 47952 7336 48004 7342
rect 47952 7278 48004 7284
rect 49792 7336 49844 7342
rect 49792 7278 49844 7284
rect 51172 7336 51224 7342
rect 51172 7278 51224 7284
rect 51908 7336 51960 7342
rect 51908 7278 51960 7284
rect 52184 7336 52236 7342
rect 52184 7278 52236 7284
rect 54024 7336 54076 7342
rect 54024 7278 54076 7284
rect 54300 7336 54352 7342
rect 54300 7278 54352 7284
rect 56048 7336 56100 7342
rect 56048 7278 56100 7284
rect 56416 7336 56468 7342
rect 56416 7278 56468 7284
rect 58164 7336 58216 7342
rect 58164 7278 58216 7284
rect 58532 7336 58584 7342
rect 60292 7324 60320 8648
rect 62408 7426 62436 8648
rect 64524 7426 64552 8648
rect 66640 8622 66760 8648
rect 68756 8622 68876 8648
rect 65456 7644 65752 7664
rect 65512 7642 65536 7644
rect 65592 7642 65616 7644
rect 65672 7642 65696 7644
rect 65534 7590 65536 7642
rect 65598 7590 65610 7642
rect 65672 7590 65674 7642
rect 65512 7588 65536 7590
rect 65592 7588 65616 7590
rect 65672 7588 65696 7590
rect 65456 7568 65752 7588
rect 62408 7398 62528 7426
rect 64524 7398 64644 7426
rect 62500 7342 62528 7398
rect 64616 7342 64644 7398
rect 66732 7342 66760 8622
rect 68848 7342 68876 8622
rect 70872 7342 70900 8648
rect 72988 7342 73016 8648
rect 75104 7342 75132 8648
rect 77220 7342 77248 8648
rect 79336 7342 79364 8648
rect 81452 7342 81480 8648
rect 83568 7342 83596 8648
rect 85684 7342 85712 8648
rect 87800 7342 87828 8648
rect 89916 7342 89944 8648
rect 92032 7342 92060 8648
rect 60372 7336 60424 7342
rect 60292 7296 60372 7324
rect 58532 7278 58584 7284
rect 60372 7278 60424 7284
rect 60648 7336 60700 7342
rect 60648 7278 60700 7284
rect 62488 7336 62540 7342
rect 62488 7278 62540 7284
rect 62764 7336 62816 7342
rect 62764 7278 62816 7284
rect 64604 7336 64656 7342
rect 64604 7278 64656 7284
rect 64880 7336 64932 7342
rect 64880 7278 64932 7284
rect 66720 7336 66772 7342
rect 66720 7278 66772 7284
rect 66996 7336 67048 7342
rect 66996 7278 67048 7284
rect 68836 7336 68888 7342
rect 68836 7278 68888 7284
rect 69112 7336 69164 7342
rect 69112 7278 69164 7284
rect 70860 7336 70912 7342
rect 70860 7278 70912 7284
rect 71228 7336 71280 7342
rect 71228 7278 71280 7284
rect 72976 7336 73028 7342
rect 72976 7278 73028 7284
rect 73344 7336 73396 7342
rect 73344 7278 73396 7284
rect 75092 7336 75144 7342
rect 75092 7278 75144 7284
rect 75460 7336 75512 7342
rect 75460 7278 75512 7284
rect 77208 7336 77260 7342
rect 77208 7278 77260 7284
rect 77576 7336 77628 7342
rect 77576 7278 77628 7284
rect 79324 7336 79376 7342
rect 79324 7278 79376 7284
rect 79692 7336 79744 7342
rect 79692 7278 79744 7284
rect 81440 7336 81492 7342
rect 81440 7278 81492 7284
rect 81808 7336 81860 7342
rect 81808 7278 81860 7284
rect 83556 7336 83608 7342
rect 83556 7278 83608 7284
rect 83924 7336 83976 7342
rect 83924 7278 83976 7284
rect 85672 7336 85724 7342
rect 85672 7278 85724 7284
rect 86040 7336 86092 7342
rect 86040 7278 86092 7284
rect 87788 7336 87840 7342
rect 87788 7278 87840 7284
rect 88156 7336 88208 7342
rect 88156 7278 88208 7284
rect 89904 7336 89956 7342
rect 89904 7278 89956 7284
rect 90272 7336 90324 7342
rect 90272 7278 90324 7284
rect 92020 7336 92072 7342
rect 92020 7278 92072 7284
rect 92388 7336 92440 7342
rect 92388 7278 92440 7284
rect 94148 7290 94176 8648
rect 96080 7342 96108 8662
rect 96172 8650 96200 8662
rect 96250 8650 96306 8704
rect 96172 8648 96306 8650
rect 98366 8648 98422 8704
rect 100482 8648 100538 8704
rect 102598 8650 102654 8704
rect 104714 8650 104770 8704
rect 102598 8648 102732 8650
rect 104714 8648 104848 8650
rect 96172 8622 96292 8648
rect 96176 7644 96472 7664
rect 96232 7642 96256 7644
rect 96312 7642 96336 7644
rect 96392 7642 96416 7644
rect 96254 7590 96256 7642
rect 96318 7590 96330 7642
rect 96392 7590 96394 7642
rect 96232 7588 96256 7590
rect 96312 7588 96336 7590
rect 96392 7588 96416 7590
rect 96176 7568 96472 7588
rect 98380 7342 98408 8648
rect 100496 7342 100524 8648
rect 102612 8622 102732 8648
rect 104728 8622 104848 8648
rect 102704 7342 102732 8622
rect 104820 7342 104848 8622
rect 94228 7336 94280 7342
rect 94148 7284 94228 7290
rect 94148 7278 94280 7284
rect 94504 7336 94556 7342
rect 94504 7278 94556 7284
rect 96068 7336 96120 7342
rect 96068 7278 96120 7284
rect 96620 7336 96672 7342
rect 96620 7278 96672 7284
rect 98368 7336 98420 7342
rect 98368 7278 98420 7284
rect 98736 7336 98788 7342
rect 98736 7278 98788 7284
rect 100484 7336 100536 7342
rect 100484 7278 100536 7284
rect 100852 7336 100904 7342
rect 100852 7278 100904 7284
rect 102692 7336 102744 7342
rect 102692 7278 102744 7284
rect 102968 7336 103020 7342
rect 102968 7278 103020 7284
rect 104808 7336 104860 7342
rect 104808 7278 104860 7284
rect 105084 7336 105136 7342
rect 105084 7278 105136 7284
rect 1136 6866 1164 7278
rect 2596 7200 2648 7206
rect 2596 7142 2648 7148
rect 1124 6860 1176 6866
rect 1124 6802 1176 6808
rect 1136 5234 1164 6802
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 2148 6390 2176 6734
rect 2136 6384 2188 6390
rect 2136 6326 2188 6332
rect 1308 5772 1360 5778
rect 1308 5714 1360 5720
rect 1320 5234 1348 5714
rect 1124 5228 1176 5234
rect 1124 5170 1176 5176
rect 1308 5228 1360 5234
rect 1308 5170 1360 5176
rect 1136 4622 1164 5170
rect 1124 4616 1176 4622
rect 1124 4558 1176 4564
rect 1136 4146 1164 4558
rect 1124 4140 1176 4146
rect 1124 4082 1176 4088
rect 1136 3602 1164 4082
rect 1124 3596 1176 3602
rect 1124 3538 1176 3544
rect 1136 1970 1164 3538
rect 1320 3194 1348 5170
rect 2228 4480 2280 4486
rect 2228 4422 2280 4428
rect 1492 3936 1544 3942
rect 1492 3878 1544 3884
rect 1400 3528 1452 3534
rect 1400 3470 1452 3476
rect 1308 3188 1360 3194
rect 1308 3130 1360 3136
rect 1412 2990 1440 3470
rect 1400 2984 1452 2990
rect 1400 2926 1452 2932
rect 1216 2508 1268 2514
rect 1216 2450 1268 2456
rect 1228 2417 1256 2450
rect 1214 2408 1270 2417
rect 1214 2343 1270 2352
rect 1124 1964 1176 1970
rect 1124 1906 1176 1912
rect 1032 1556 1084 1562
rect 1032 1498 1084 1504
rect 1044 56 1072 1498
rect 1136 1426 1164 1906
rect 1228 1902 1256 2343
rect 1216 1896 1268 1902
rect 1216 1838 1268 1844
rect 1124 1420 1176 1426
rect 1124 1362 1176 1368
rect 1504 56 1532 3878
rect 2240 1578 2268 4422
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 2516 3738 2544 4014
rect 2504 3732 2556 3738
rect 2504 3674 2556 3680
rect 2504 1760 2556 1766
rect 2504 1702 2556 1708
rect 2148 1550 2268 1578
rect 1964 56 2084 82
rect 1030 0 1086 56
rect 1490 0 1546 56
rect 1950 54 2084 56
rect 1950 0 2006 54
rect 2056 42 2084 54
rect 2148 42 2176 1550
rect 2516 1426 2544 1702
rect 2504 1420 2556 1426
rect 2504 1362 2556 1368
rect 2332 56 2452 82
rect 2056 14 2176 42
rect 2318 54 2452 56
rect 2318 0 2374 54
rect 2424 42 2452 54
rect 2608 42 2636 7142
rect 3252 6866 3280 7278
rect 3528 7002 3556 7278
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 3516 6996 3568 7002
rect 3516 6938 3568 6944
rect 3240 6860 3292 6866
rect 3240 6802 3292 6808
rect 3252 5234 3280 6802
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 3528 6254 3556 6734
rect 4016 6556 4312 6576
rect 4072 6554 4096 6556
rect 4152 6554 4176 6556
rect 4232 6554 4256 6556
rect 4094 6502 4096 6554
rect 4158 6502 4170 6554
rect 4232 6502 4234 6554
rect 4072 6500 4096 6502
rect 4152 6500 4176 6502
rect 4232 6500 4256 6502
rect 4016 6480 4312 6500
rect 3516 6248 3568 6254
rect 3516 6190 3568 6196
rect 3516 5772 3568 5778
rect 3516 5714 3568 5720
rect 3528 5234 3556 5714
rect 4016 5468 4312 5488
rect 4072 5466 4096 5468
rect 4152 5466 4176 5468
rect 4232 5466 4256 5468
rect 4094 5414 4096 5466
rect 4158 5414 4170 5466
rect 4232 5414 4234 5466
rect 4072 5412 4096 5414
rect 4152 5412 4176 5414
rect 4232 5412 4256 5414
rect 4016 5392 4312 5412
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 3252 4690 3280 5170
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3528 4690 3556 4966
rect 3240 4684 3292 4690
rect 3240 4626 3292 4632
rect 3516 4684 3568 4690
rect 3516 4626 3568 4632
rect 3252 4146 3280 4626
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4016 4380 4312 4400
rect 4072 4378 4096 4380
rect 4152 4378 4176 4380
rect 4232 4378 4256 4380
rect 4094 4326 4096 4378
rect 4158 4326 4170 4378
rect 4232 4326 4234 4378
rect 4072 4324 4096 4326
rect 4152 4324 4176 4326
rect 4232 4324 4256 4326
rect 4016 4304 4312 4324
rect 3240 4140 3292 4146
rect 3240 4082 3292 4088
rect 3252 3602 3280 4082
rect 3884 4072 3936 4078
rect 3884 4014 3936 4020
rect 3240 3596 3292 3602
rect 3240 3538 3292 3544
rect 3252 1970 3280 3538
rect 3896 3534 3924 4014
rect 3516 3528 3568 3534
rect 3516 3470 3568 3476
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 3528 2990 3556 3470
rect 4016 3292 4312 3312
rect 4072 3290 4096 3292
rect 4152 3290 4176 3292
rect 4232 3290 4256 3292
rect 4094 3238 4096 3290
rect 4158 3238 4170 3290
rect 4232 3238 4234 3290
rect 4072 3236 4096 3238
rect 4152 3236 4176 3238
rect 4232 3236 4256 3238
rect 4016 3216 4312 3236
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3516 2508 3568 2514
rect 3516 2450 3568 2456
rect 3528 1970 3556 2450
rect 4016 2204 4312 2224
rect 4072 2202 4096 2204
rect 4152 2202 4176 2204
rect 4232 2202 4256 2204
rect 4094 2150 4096 2202
rect 4158 2150 4170 2202
rect 4232 2150 4234 2202
rect 4072 2148 4096 2150
rect 4152 2148 4176 2150
rect 4232 2148 4256 2150
rect 4016 2128 4312 2148
rect 3240 1964 3292 1970
rect 3240 1906 3292 1912
rect 3516 1964 3568 1970
rect 3516 1906 3568 1912
rect 3608 1964 3660 1970
rect 3608 1906 3660 1912
rect 3252 1426 3280 1906
rect 3240 1420 3292 1426
rect 3240 1362 3292 1368
rect 3424 1216 3476 1222
rect 3424 1158 3476 1164
rect 3160 56 3280 82
rect 2424 14 2636 42
rect 3146 54 3280 56
rect 3146 0 3202 54
rect 3252 42 3280 54
rect 3436 42 3464 1158
rect 3620 56 3648 1906
rect 4160 1760 4212 1766
rect 4160 1702 4212 1708
rect 4172 1426 4200 1702
rect 4160 1420 4212 1426
rect 4160 1362 4212 1368
rect 4016 1116 4312 1136
rect 4072 1114 4096 1116
rect 4152 1114 4176 1116
rect 4232 1114 4256 1116
rect 4094 1062 4096 1114
rect 4158 1062 4170 1114
rect 4232 1062 4234 1114
rect 4072 1060 4096 1062
rect 4152 1060 4176 1062
rect 4232 1060 4256 1062
rect 4016 1040 4312 1060
rect 4080 56 4200 82
rect 3252 14 3464 42
rect 3606 0 3662 56
rect 4066 54 4200 56
rect 4066 0 4122 54
rect 4172 42 4200 54
rect 4356 42 4384 4422
rect 4540 82 4568 7142
rect 5276 6866 5304 7278
rect 5644 7002 5672 7278
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 5632 6996 5684 7002
rect 5632 6938 5684 6944
rect 5264 6860 5316 6866
rect 5264 6802 5316 6808
rect 5276 5234 5304 6802
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5644 6254 5672 6734
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5632 5636 5684 5642
rect 5632 5578 5684 5584
rect 5644 5234 5672 5578
rect 5264 5228 5316 5234
rect 5264 5170 5316 5176
rect 5632 5228 5684 5234
rect 5632 5170 5684 5176
rect 5276 4690 5304 5170
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 5644 4690 5672 4966
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 5632 4684 5684 4690
rect 5632 4626 5684 4632
rect 5276 4146 5304 4626
rect 6276 4616 6328 4622
rect 6196 4564 6276 4570
rect 6196 4558 6328 4564
rect 6196 4542 6316 4558
rect 5264 4140 5316 4146
rect 5316 4100 5396 4128
rect 5264 4082 5316 4088
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4632 1970 4660 3878
rect 5368 3602 5396 4100
rect 6000 4072 6052 4078
rect 6000 4014 6052 4020
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5368 1970 5396 3538
rect 6012 3534 6040 4014
rect 5632 3528 5684 3534
rect 5632 3470 5684 3476
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 5644 2990 5672 3470
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 5632 2508 5684 2514
rect 5632 2450 5684 2456
rect 5644 1970 5672 2450
rect 4620 1964 4672 1970
rect 4620 1906 4672 1912
rect 5356 1964 5408 1970
rect 5356 1906 5408 1912
rect 5632 1964 5684 1970
rect 5632 1906 5684 1912
rect 5368 1426 5396 1906
rect 5724 1896 5776 1902
rect 5724 1838 5776 1844
rect 5356 1420 5408 1426
rect 5356 1362 5408 1368
rect 5632 1216 5684 1222
rect 5632 1158 5684 1164
rect 4448 56 4568 82
rect 5276 56 5396 82
rect 4172 14 4384 42
rect 4434 54 4568 56
rect 5262 54 5396 56
rect 4434 0 4490 54
rect 5262 0 5318 54
rect 5368 42 5396 54
rect 5644 42 5672 1158
rect 5736 56 5764 1838
rect 5908 1760 5960 1766
rect 5908 1702 5960 1708
rect 5920 1426 5948 1702
rect 5908 1420 5960 1426
rect 5908 1362 5960 1368
rect 6196 56 6224 4542
rect 6656 1850 6684 7142
rect 7392 6866 7420 7278
rect 7760 7002 7788 7278
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 7748 6996 7800 7002
rect 7748 6938 7800 6944
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7392 5234 7420 6802
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7760 6254 7788 6734
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 7656 5772 7708 5778
rect 7656 5714 7708 5720
rect 7668 5234 7696 5714
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7392 4690 7420 5170
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7760 4690 7788 4966
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7748 4684 7800 4690
rect 7748 4626 7800 4632
rect 7392 4146 7420 4626
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 7380 4140 7432 4146
rect 8220 4128 8248 4422
rect 7432 4100 7512 4128
rect 8220 4100 8340 4128
rect 7380 4082 7432 4088
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6748 1902 6776 3878
rect 7484 3602 7512 4100
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 7472 3596 7524 3602
rect 7472 3538 7524 3544
rect 7484 1970 7512 3538
rect 8128 3534 8156 4014
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 7760 2990 7788 3470
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7748 2576 7800 2582
rect 7748 2518 7800 2524
rect 7760 1970 7788 2518
rect 7472 1964 7524 1970
rect 7472 1906 7524 1912
rect 7748 1964 7800 1970
rect 7748 1906 7800 1912
rect 7840 1964 7892 1970
rect 7840 1906 7892 1912
rect 6564 1822 6684 1850
rect 6736 1896 6788 1902
rect 6736 1838 6788 1844
rect 6564 56 6592 1822
rect 7380 1556 7432 1562
rect 7380 1498 7432 1504
rect 7392 56 7420 1498
rect 7484 1426 7512 1906
rect 7472 1420 7524 1426
rect 7472 1362 7524 1368
rect 7852 56 7880 1906
rect 8208 1760 8260 1766
rect 8208 1702 8260 1708
rect 8220 1426 8248 1702
rect 8208 1420 8260 1426
rect 8208 1362 8260 1368
rect 8312 56 8340 4100
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8864 1970 8892 3878
rect 8852 1964 8904 1970
rect 8852 1906 8904 1912
rect 8956 1850 8984 7142
rect 9600 6866 9628 7278
rect 9876 7002 9904 7278
rect 11244 7268 11296 7274
rect 11244 7210 11296 7216
rect 9864 6996 9916 7002
rect 9864 6938 9916 6944
rect 9588 6860 9640 6866
rect 9588 6802 9640 6808
rect 9600 5234 9628 6802
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9876 6254 9904 6734
rect 9864 6248 9916 6254
rect 9864 6190 9916 6196
rect 9864 5704 9916 5710
rect 9864 5646 9916 5652
rect 9876 5234 9904 5646
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 9600 4690 9628 5170
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 9876 4690 9904 4966
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 9600 4146 9628 4626
rect 10508 4480 10560 4486
rect 10508 4422 10560 4428
rect 9588 4140 9640 4146
rect 9588 4082 9640 4088
rect 9600 3602 9628 4082
rect 9588 3596 9640 3602
rect 9588 3538 9640 3544
rect 9600 1970 9628 3538
rect 9864 3528 9916 3534
rect 9864 3470 9916 3476
rect 9876 2990 9904 3470
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 9876 1970 9904 2382
rect 9588 1964 9640 1970
rect 9588 1906 9640 1912
rect 9864 1964 9916 1970
rect 9864 1906 9916 1912
rect 9956 1964 10008 1970
rect 9956 1906 10008 1912
rect 8680 1822 8984 1850
rect 8680 56 8708 1822
rect 9496 1556 9548 1562
rect 9496 1498 9548 1504
rect 9508 56 9536 1498
rect 9600 1426 9628 1906
rect 9588 1420 9640 1426
rect 9588 1362 9640 1368
rect 9968 56 9996 1906
rect 10520 82 10548 4422
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 10980 3738 11008 4014
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 11164 1970 11192 3878
rect 11152 1964 11204 1970
rect 11152 1906 11204 1912
rect 11256 1902 11284 7210
rect 11716 6866 11744 7278
rect 11992 7002 12020 7278
rect 13360 7268 13412 7274
rect 13360 7210 13412 7216
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11716 5234 11744 6802
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 11992 6254 12020 6734
rect 11980 6248 12032 6254
rect 11980 6190 12032 6196
rect 11888 5840 11940 5846
rect 11888 5782 11940 5788
rect 11900 5234 11928 5782
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11716 4690 11744 5170
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11992 4690 12020 4966
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 11716 4146 11744 4626
rect 12624 4480 12676 4486
rect 12624 4422 12676 4428
rect 11704 4140 11756 4146
rect 11704 4082 11756 4088
rect 11716 3602 11744 4082
rect 11704 3596 11756 3602
rect 11704 3538 11756 3544
rect 11716 1970 11744 3538
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11992 2990 12020 3470
rect 11980 2984 12032 2990
rect 11980 2926 12032 2932
rect 11888 2576 11940 2582
rect 11888 2518 11940 2524
rect 11900 1970 11928 2518
rect 11704 1964 11756 1970
rect 11704 1906 11756 1912
rect 11888 1964 11940 1970
rect 11888 1906 11940 1912
rect 12072 1964 12124 1970
rect 12072 1906 12124 1912
rect 10784 1896 10836 1902
rect 10784 1838 10836 1844
rect 11244 1896 11296 1902
rect 11244 1838 11296 1844
rect 10428 56 10548 82
rect 10796 56 10824 1838
rect 11152 1760 11204 1766
rect 11152 1702 11204 1708
rect 11164 1426 11192 1702
rect 11716 1426 11744 1906
rect 11152 1420 11204 1426
rect 11152 1362 11204 1368
rect 11704 1420 11756 1426
rect 11704 1362 11756 1368
rect 11612 1216 11664 1222
rect 11612 1158 11664 1164
rect 11624 56 11652 1158
rect 12084 56 12112 1906
rect 12636 82 12664 4422
rect 13084 4072 13136 4078
rect 13084 4014 13136 4020
rect 13096 3738 13124 4014
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 13280 1970 13308 3878
rect 13268 1964 13320 1970
rect 13268 1906 13320 1912
rect 13372 1850 13400 7210
rect 13832 6866 13860 7278
rect 14108 7002 14136 7278
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 14096 6996 14148 7002
rect 14096 6938 14148 6944
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 13832 5234 13860 6802
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 14108 6254 14136 6734
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 14096 5840 14148 5846
rect 14096 5782 14148 5788
rect 14108 5234 14136 5782
rect 13820 5228 13872 5234
rect 13820 5170 13872 5176
rect 14096 5228 14148 5234
rect 14096 5170 14148 5176
rect 13832 4690 13860 5170
rect 14096 5024 14148 5030
rect 14096 4966 14148 4972
rect 14108 4690 14136 4966
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 14096 4684 14148 4690
rect 14096 4626 14148 4632
rect 13832 4146 13860 4626
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13832 3602 13860 4082
rect 14188 3936 14240 3942
rect 14188 3878 14240 3884
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 13832 1970 13860 3538
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 14108 2990 14136 3470
rect 14096 2984 14148 2990
rect 14096 2926 14148 2932
rect 14096 2576 14148 2582
rect 14096 2518 14148 2524
rect 14108 1970 14136 2518
rect 13820 1964 13872 1970
rect 13820 1906 13872 1912
rect 14096 1964 14148 1970
rect 14096 1906 14148 1912
rect 13188 1822 13400 1850
rect 12544 56 12664 82
rect 12912 56 13032 82
rect 5368 14 5672 42
rect 5722 0 5778 56
rect 6182 0 6238 56
rect 6550 0 6606 56
rect 7378 0 7434 56
rect 7838 0 7894 56
rect 8298 0 8354 56
rect 8666 0 8722 56
rect 9494 0 9550 56
rect 9954 0 10010 56
rect 10414 54 10548 56
rect 10414 0 10470 54
rect 10782 0 10838 56
rect 11610 0 11666 56
rect 12070 0 12126 56
rect 12530 54 12664 56
rect 12898 54 13032 56
rect 12530 0 12586 54
rect 12898 0 12954 54
rect 13004 42 13032 54
rect 13188 42 13216 1822
rect 13268 1760 13320 1766
rect 13268 1702 13320 1708
rect 13280 1426 13308 1702
rect 13728 1556 13780 1562
rect 13728 1498 13780 1504
rect 13268 1420 13320 1426
rect 13268 1362 13320 1368
rect 13740 56 13768 1498
rect 13832 1426 13860 1906
rect 13820 1420 13872 1426
rect 13820 1362 13872 1368
rect 14200 56 14228 3878
rect 14568 82 14596 4422
rect 15120 82 15148 7142
rect 15948 6866 15976 7278
rect 16224 7002 16252 7278
rect 17224 7200 17276 7206
rect 17224 7142 17276 7148
rect 16212 6996 16264 7002
rect 16212 6938 16264 6944
rect 15936 6860 15988 6866
rect 15936 6802 15988 6808
rect 15948 5234 15976 6802
rect 16212 6792 16264 6798
rect 16212 6734 16264 6740
rect 16224 6254 16252 6734
rect 16212 6248 16264 6254
rect 16212 6190 16264 6196
rect 16212 5772 16264 5778
rect 16212 5714 16264 5720
rect 16224 5234 16252 5714
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 16212 5228 16264 5234
rect 16212 5170 16264 5176
rect 15948 4690 15976 5170
rect 16212 5024 16264 5030
rect 16212 4966 16264 4972
rect 16224 4690 16252 4966
rect 15936 4684 15988 4690
rect 15936 4626 15988 4632
rect 16212 4684 16264 4690
rect 16212 4626 16264 4632
rect 15948 4146 15976 4626
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 15936 4140 15988 4146
rect 15936 4082 15988 4088
rect 15200 4072 15252 4078
rect 15200 4014 15252 4020
rect 15212 3738 15240 4014
rect 15200 3732 15252 3738
rect 15200 3674 15252 3680
rect 15948 3602 15976 4082
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 15936 3596 15988 3602
rect 15936 3538 15988 3544
rect 15948 1970 15976 3538
rect 16212 3528 16264 3534
rect 16212 3470 16264 3476
rect 16224 2922 16252 3470
rect 16212 2916 16264 2922
rect 16212 2858 16264 2864
rect 16212 2508 16264 2514
rect 16212 2450 16264 2456
rect 16224 1970 16252 2450
rect 15936 1964 15988 1970
rect 15936 1906 15988 1912
rect 16212 1964 16264 1970
rect 16212 1906 16264 1912
rect 15200 1760 15252 1766
rect 15200 1702 15252 1708
rect 15212 1426 15240 1702
rect 15948 1426 15976 1906
rect 15200 1420 15252 1426
rect 15200 1362 15252 1368
rect 15936 1420 15988 1426
rect 15936 1362 15988 1368
rect 16120 1216 16172 1222
rect 16120 1158 16172 1164
rect 14568 56 14688 82
rect 15028 56 15148 82
rect 15856 56 15976 82
rect 13004 14 13216 42
rect 13726 0 13782 56
rect 14186 0 14242 56
rect 14568 54 14702 56
rect 14646 0 14702 54
rect 15014 54 15148 56
rect 15842 54 15976 56
rect 15014 0 15070 54
rect 15842 0 15898 54
rect 15948 42 15976 54
rect 16132 42 16160 1158
rect 16316 56 16344 3878
rect 16868 82 16896 4422
rect 17236 82 17264 7142
rect 18064 6866 18092 7278
rect 18340 7002 18368 7278
rect 19248 7200 19300 7206
rect 19248 7142 19300 7148
rect 18328 6996 18380 7002
rect 18328 6938 18380 6944
rect 18052 6860 18104 6866
rect 18052 6802 18104 6808
rect 18064 5234 18092 6802
rect 18328 6792 18380 6798
rect 18328 6734 18380 6740
rect 18340 6254 18368 6734
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 18328 5636 18380 5642
rect 18328 5578 18380 5584
rect 18340 5234 18368 5578
rect 18052 5228 18104 5234
rect 18052 5170 18104 5176
rect 18328 5228 18380 5234
rect 18328 5170 18380 5176
rect 18064 4690 18092 5170
rect 18328 5024 18380 5030
rect 18328 4966 18380 4972
rect 18340 4690 18368 4966
rect 18052 4684 18104 4690
rect 18052 4626 18104 4632
rect 18328 4684 18380 4690
rect 18328 4626 18380 4632
rect 18064 4146 18092 4626
rect 18972 4480 19024 4486
rect 18972 4422 19024 4428
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17328 3738 17356 4014
rect 17316 3732 17368 3738
rect 17316 3674 17368 3680
rect 18064 3602 18092 4082
rect 18420 4072 18472 4078
rect 18420 4014 18472 4020
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 18064 1970 18092 3538
rect 18432 3534 18460 4014
rect 18696 3936 18748 3942
rect 18696 3878 18748 3884
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18340 2990 18368 3470
rect 18328 2984 18380 2990
rect 18328 2926 18380 2932
rect 18328 2372 18380 2378
rect 18328 2314 18380 2320
rect 18340 1970 18368 2314
rect 18052 1964 18104 1970
rect 18052 1906 18104 1912
rect 18328 1964 18380 1970
rect 18328 1906 18380 1912
rect 17316 1760 17368 1766
rect 17316 1702 17368 1708
rect 17328 1426 17356 1702
rect 18064 1426 18092 1906
rect 18708 1902 18736 3878
rect 18420 1896 18472 1902
rect 18420 1838 18472 1844
rect 18696 1896 18748 1902
rect 18696 1838 18748 1844
rect 17316 1420 17368 1426
rect 17316 1362 17368 1368
rect 18052 1420 18104 1426
rect 18052 1362 18104 1368
rect 18328 1216 18380 1222
rect 18328 1158 18380 1164
rect 16776 56 16896 82
rect 17144 56 17264 82
rect 17972 56 18092 82
rect 15948 14 16160 42
rect 16302 0 16358 56
rect 16762 54 16896 56
rect 17130 54 17264 56
rect 17958 54 18092 56
rect 16762 0 16818 54
rect 17130 0 17186 54
rect 17958 0 18014 54
rect 18064 42 18092 54
rect 18340 42 18368 1158
rect 18432 56 18460 1838
rect 18696 1760 18748 1766
rect 18696 1702 18748 1708
rect 18708 1426 18736 1702
rect 18696 1420 18748 1426
rect 18696 1362 18748 1368
rect 18984 82 19012 4422
rect 18892 56 19012 82
rect 19260 56 19288 7142
rect 19376 7100 19672 7120
rect 19432 7098 19456 7100
rect 19512 7098 19536 7100
rect 19592 7098 19616 7100
rect 19454 7046 19456 7098
rect 19518 7046 19530 7098
rect 19592 7046 19594 7098
rect 19432 7044 19456 7046
rect 19512 7044 19536 7046
rect 19592 7044 19616 7046
rect 19376 7024 19672 7044
rect 20088 6866 20116 7278
rect 20456 7002 20484 7278
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 20444 6996 20496 7002
rect 20444 6938 20496 6944
rect 20076 6860 20128 6866
rect 20076 6802 20128 6808
rect 19376 6012 19672 6032
rect 19432 6010 19456 6012
rect 19512 6010 19536 6012
rect 19592 6010 19616 6012
rect 19454 5958 19456 6010
rect 19518 5958 19530 6010
rect 19592 5958 19594 6010
rect 19432 5956 19456 5958
rect 19512 5956 19536 5958
rect 19592 5956 19616 5958
rect 19376 5936 19672 5956
rect 20088 5234 20116 6802
rect 20444 6792 20496 6798
rect 20444 6734 20496 6740
rect 20456 6254 20484 6734
rect 20444 6248 20496 6254
rect 20444 6190 20496 6196
rect 20444 5772 20496 5778
rect 20444 5714 20496 5720
rect 20456 5234 20484 5714
rect 20076 5228 20128 5234
rect 20076 5170 20128 5176
rect 20444 5228 20496 5234
rect 20444 5170 20496 5176
rect 19376 4924 19672 4944
rect 19432 4922 19456 4924
rect 19512 4922 19536 4924
rect 19592 4922 19616 4924
rect 19454 4870 19456 4922
rect 19518 4870 19530 4922
rect 19592 4870 19594 4922
rect 19432 4868 19456 4870
rect 19512 4868 19536 4870
rect 19592 4868 19616 4870
rect 19376 4848 19672 4868
rect 20088 4690 20116 5170
rect 20444 5024 20496 5030
rect 20444 4966 20496 4972
rect 20456 4690 20484 4966
rect 20076 4684 20128 4690
rect 20076 4626 20128 4632
rect 20444 4684 20496 4690
rect 20444 4626 20496 4632
rect 20088 4214 20116 4626
rect 21088 4480 21140 4486
rect 21008 4440 21088 4468
rect 20076 4208 20128 4214
rect 20128 4156 20208 4162
rect 20076 4150 20208 4156
rect 20088 4134 20208 4150
rect 19376 3836 19672 3856
rect 19432 3834 19456 3836
rect 19512 3834 19536 3836
rect 19592 3834 19616 3836
rect 19454 3782 19456 3834
rect 19518 3782 19530 3834
rect 19592 3782 19594 3834
rect 19432 3780 19456 3782
rect 19512 3780 19536 3782
rect 19592 3780 19616 3782
rect 19376 3760 19672 3780
rect 20180 3602 20208 4134
rect 20168 3596 20220 3602
rect 20168 3538 20220 3544
rect 19376 2748 19672 2768
rect 19432 2746 19456 2748
rect 19512 2746 19536 2748
rect 19592 2746 19616 2748
rect 19454 2694 19456 2746
rect 19518 2694 19530 2746
rect 19592 2694 19594 2746
rect 19432 2692 19456 2694
rect 19512 2692 19536 2694
rect 19592 2692 19616 2694
rect 19376 2672 19672 2692
rect 20180 1970 20208 3538
rect 20444 3528 20496 3534
rect 20444 3470 20496 3476
rect 20456 2990 20484 3470
rect 20444 2984 20496 2990
rect 20444 2926 20496 2932
rect 20444 2508 20496 2514
rect 20444 2450 20496 2456
rect 20456 1970 20484 2450
rect 20168 1964 20220 1970
rect 20168 1906 20220 1912
rect 20444 1964 20496 1970
rect 20444 1906 20496 1912
rect 19376 1660 19672 1680
rect 19432 1658 19456 1660
rect 19512 1658 19536 1660
rect 19592 1658 19616 1660
rect 19454 1606 19456 1658
rect 19518 1606 19530 1658
rect 19592 1606 19594 1658
rect 19432 1604 19456 1606
rect 19512 1604 19536 1606
rect 19592 1604 19616 1606
rect 19376 1584 19672 1604
rect 20180 1426 20208 1906
rect 20536 1896 20588 1902
rect 20536 1838 20588 1844
rect 20168 1420 20220 1426
rect 20168 1362 20220 1368
rect 20352 1216 20404 1222
rect 20352 1158 20404 1164
rect 20088 56 20208 82
rect 18064 14 18368 42
rect 18418 0 18474 56
rect 18878 54 19012 56
rect 18878 0 18934 54
rect 19246 0 19302 56
rect 20074 54 20208 56
rect 20074 0 20130 54
rect 20180 42 20208 54
rect 20364 42 20392 1158
rect 20548 56 20576 1838
rect 20720 1760 20772 1766
rect 20720 1702 20772 1708
rect 20732 1426 20760 1702
rect 20720 1420 20772 1426
rect 20720 1362 20772 1368
rect 21008 56 21036 4440
rect 21088 4422 21140 4428
rect 21088 4072 21140 4078
rect 21088 4014 21140 4020
rect 21100 3534 21128 4014
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 21468 82 21496 7142
rect 22204 6866 22232 7278
rect 22572 7002 22600 7278
rect 23940 7268 23992 7274
rect 23940 7210 23992 7216
rect 22560 6996 22612 7002
rect 22560 6938 22612 6944
rect 22192 6860 22244 6866
rect 22192 6802 22244 6808
rect 22204 5234 22232 6802
rect 22560 6792 22612 6798
rect 22560 6734 22612 6740
rect 22572 6254 22600 6734
rect 22560 6248 22612 6254
rect 22560 6190 22612 6196
rect 22376 5840 22428 5846
rect 22428 5788 22508 5794
rect 22376 5782 22508 5788
rect 22388 5766 22508 5782
rect 22480 5234 22508 5766
rect 23952 5234 23980 7210
rect 24412 6866 24440 7278
rect 24688 7002 24716 7278
rect 26436 7262 26556 7278
rect 25872 7200 25924 7206
rect 25872 7142 25924 7148
rect 24676 6996 24728 7002
rect 24676 6938 24728 6944
rect 24400 6860 24452 6866
rect 24400 6802 24452 6808
rect 24412 5234 24440 6802
rect 24676 6792 24728 6798
rect 24676 6734 24728 6740
rect 24688 6254 24716 6734
rect 24676 6248 24728 6254
rect 24676 6190 24728 6196
rect 24676 5840 24728 5846
rect 24676 5782 24728 5788
rect 24688 5234 24716 5782
rect 22192 5228 22244 5234
rect 22192 5170 22244 5176
rect 22468 5228 22520 5234
rect 22468 5170 22520 5176
rect 23756 5228 23808 5234
rect 23756 5170 23808 5176
rect 23940 5228 23992 5234
rect 23940 5170 23992 5176
rect 24400 5228 24452 5234
rect 24400 5170 24452 5176
rect 24676 5228 24728 5234
rect 24676 5170 24728 5176
rect 22204 4690 22232 5170
rect 22560 5024 22612 5030
rect 22560 4966 22612 4972
rect 22572 4690 22600 4966
rect 22192 4684 22244 4690
rect 22192 4626 22244 4632
rect 22560 4684 22612 4690
rect 22560 4626 22612 4632
rect 22204 4146 22232 4626
rect 23204 4480 23256 4486
rect 23204 4422 23256 4428
rect 22192 4140 22244 4146
rect 22192 4082 22244 4088
rect 21548 3936 21600 3942
rect 21548 3878 21600 3884
rect 21560 1902 21588 3878
rect 22204 3602 22232 4082
rect 22928 4072 22980 4078
rect 22928 4014 22980 4020
rect 22192 3596 22244 3602
rect 22192 3538 22244 3544
rect 22204 1970 22232 3538
rect 22940 3534 22968 4014
rect 22560 3528 22612 3534
rect 22560 3470 22612 3476
rect 22928 3528 22980 3534
rect 22928 3470 22980 3476
rect 22572 2990 22600 3470
rect 22560 2984 22612 2990
rect 22560 2926 22612 2932
rect 22376 2576 22428 2582
rect 22376 2518 22428 2524
rect 22192 1964 22244 1970
rect 22192 1906 22244 1912
rect 21548 1896 21600 1902
rect 21548 1838 21600 1844
rect 22204 1850 22232 1906
rect 22388 1902 22416 2518
rect 22652 2100 22704 2106
rect 22652 2042 22704 2048
rect 22376 1896 22428 1902
rect 22204 1822 22324 1850
rect 22376 1838 22428 1844
rect 22296 1426 22324 1822
rect 22284 1420 22336 1426
rect 22284 1362 22336 1368
rect 22560 1216 22612 1222
rect 22560 1158 22612 1164
rect 21376 56 21496 82
rect 22204 56 22324 82
rect 20180 14 20392 42
rect 20534 0 20590 56
rect 20994 0 21050 56
rect 21362 54 21496 56
rect 22190 54 22324 56
rect 21362 0 21418 54
rect 22190 0 22246 54
rect 22296 42 22324 54
rect 22572 42 22600 1158
rect 22664 56 22692 2042
rect 22836 1760 22888 1766
rect 22836 1702 22888 1708
rect 22848 1426 22876 1702
rect 22836 1420 22888 1426
rect 22836 1362 22888 1368
rect 23216 82 23244 4422
rect 23664 3936 23716 3942
rect 23664 3878 23716 3884
rect 23388 2644 23440 2650
rect 23388 2586 23440 2592
rect 23124 56 23244 82
rect 22296 14 22600 42
rect 22650 0 22706 56
rect 23110 54 23244 56
rect 23400 82 23428 2586
rect 23676 2106 23704 3878
rect 23768 2650 23796 5170
rect 24412 4690 24440 5170
rect 24676 5024 24728 5030
rect 24676 4966 24728 4972
rect 24688 4690 24716 4966
rect 24400 4684 24452 4690
rect 24400 4626 24452 4632
rect 24676 4684 24728 4690
rect 24676 4626 24728 4632
rect 24412 4146 24440 4626
rect 25320 4480 25372 4486
rect 25320 4422 25372 4428
rect 24400 4140 24452 4146
rect 24400 4082 24452 4088
rect 24412 3602 24440 4082
rect 25044 4072 25096 4078
rect 25044 4014 25096 4020
rect 24400 3596 24452 3602
rect 24400 3538 24452 3544
rect 23756 2644 23808 2650
rect 23756 2586 23808 2592
rect 23664 2100 23716 2106
rect 23664 2042 23716 2048
rect 24412 1970 24440 3538
rect 25056 3534 25084 4014
rect 24676 3528 24728 3534
rect 24676 3470 24728 3476
rect 25044 3528 25096 3534
rect 25044 3470 25096 3476
rect 24688 2990 24716 3470
rect 24676 2984 24728 2990
rect 24676 2926 24728 2932
rect 24676 2576 24728 2582
rect 24676 2518 24728 2524
rect 24688 1970 24716 2518
rect 24768 2100 24820 2106
rect 24768 2042 24820 2048
rect 24400 1964 24452 1970
rect 24400 1906 24452 1912
rect 24676 1964 24728 1970
rect 24676 1906 24728 1912
rect 24308 1556 24360 1562
rect 24308 1498 24360 1504
rect 23400 56 23520 82
rect 24320 56 24348 1498
rect 24412 1426 24440 1906
rect 24400 1420 24452 1426
rect 24400 1362 24452 1368
rect 24780 56 24808 2042
rect 25044 1760 25096 1766
rect 25044 1702 25096 1708
rect 25056 1426 25084 1702
rect 25044 1420 25096 1426
rect 25044 1362 25096 1368
rect 25332 82 25360 4422
rect 25780 3936 25832 3942
rect 25780 3878 25832 3884
rect 25792 2106 25820 3878
rect 25780 2100 25832 2106
rect 25780 2042 25832 2048
rect 25884 1986 25912 7142
rect 26528 6866 26556 7262
rect 26804 7002 26832 7278
rect 27988 7200 28040 7206
rect 27988 7142 28040 7148
rect 26792 6996 26844 7002
rect 26792 6938 26844 6944
rect 26516 6860 26568 6866
rect 26516 6802 26568 6808
rect 26528 5234 26556 6802
rect 26792 6792 26844 6798
rect 26792 6734 26844 6740
rect 26804 6254 26832 6734
rect 26792 6248 26844 6254
rect 26792 6190 26844 6196
rect 26700 5704 26752 5710
rect 26700 5646 26752 5652
rect 26712 5234 26740 5646
rect 26516 5228 26568 5234
rect 26516 5170 26568 5176
rect 26700 5228 26752 5234
rect 26700 5170 26752 5176
rect 26528 4690 26556 5170
rect 26792 5024 26844 5030
rect 26792 4966 26844 4972
rect 26804 4690 26832 4966
rect 26516 4684 26568 4690
rect 26516 4626 26568 4632
rect 26792 4684 26844 4690
rect 26792 4626 26844 4632
rect 26528 4146 26556 4626
rect 27436 4616 27488 4622
rect 27356 4576 27436 4604
rect 26516 4140 26568 4146
rect 26516 4082 26568 4088
rect 26528 3602 26556 4082
rect 26516 3596 26568 3602
rect 26516 3538 26568 3544
rect 25240 56 25360 82
rect 25608 1958 25912 1986
rect 26528 1970 26556 3538
rect 26792 3528 26844 3534
rect 26792 3470 26844 3476
rect 26804 2990 26832 3470
rect 26792 2984 26844 2990
rect 26792 2926 26844 2932
rect 26700 2440 26752 2446
rect 26700 2382 26752 2388
rect 26712 1970 26740 2382
rect 26516 1964 26568 1970
rect 25608 56 25636 1958
rect 26516 1906 26568 1912
rect 26700 1964 26752 1970
rect 26700 1906 26752 1912
rect 26424 1556 26476 1562
rect 26424 1498 26476 1504
rect 26436 56 26464 1498
rect 26528 1426 26556 1906
rect 26884 1896 26936 1902
rect 26884 1838 26936 1844
rect 26516 1420 26568 1426
rect 26516 1362 26568 1368
rect 26896 56 26924 1838
rect 27356 56 27384 4576
rect 27436 4558 27488 4564
rect 27896 4072 27948 4078
rect 27896 4014 27948 4020
rect 27908 3738 27936 4014
rect 27896 3732 27948 3738
rect 27896 3674 27948 3680
rect 28000 1578 28028 7142
rect 28644 6866 28672 7278
rect 28920 7002 28948 7278
rect 30288 7268 30340 7274
rect 30288 7210 30340 7216
rect 28908 6996 28960 7002
rect 28908 6938 28960 6944
rect 28632 6860 28684 6866
rect 28632 6802 28684 6808
rect 28644 5234 28672 6802
rect 28908 6792 28960 6798
rect 28908 6734 28960 6740
rect 28920 6254 28948 6734
rect 28908 6248 28960 6254
rect 28908 6190 28960 6196
rect 28816 5704 28868 5710
rect 28816 5646 28868 5652
rect 28828 5234 28856 5646
rect 28632 5228 28684 5234
rect 28632 5170 28684 5176
rect 28816 5228 28868 5234
rect 28816 5170 28868 5176
rect 28644 4690 28672 5170
rect 28908 5024 28960 5030
rect 28908 4966 28960 4972
rect 28920 4690 28948 4966
rect 28632 4684 28684 4690
rect 28632 4626 28684 4632
rect 28908 4684 28960 4690
rect 28908 4626 28960 4632
rect 28644 4146 28672 4626
rect 29552 4616 29604 4622
rect 29472 4564 29552 4570
rect 29472 4558 29604 4564
rect 29472 4542 29592 4558
rect 28632 4140 28684 4146
rect 28632 4082 28684 4088
rect 28080 3936 28132 3942
rect 28080 3878 28132 3884
rect 28092 1902 28120 3878
rect 28644 3602 28672 4082
rect 28632 3596 28684 3602
rect 28632 3538 28684 3544
rect 28644 1970 28672 3538
rect 28908 3528 28960 3534
rect 28908 3470 28960 3476
rect 28920 2990 28948 3470
rect 28908 2984 28960 2990
rect 28908 2926 28960 2932
rect 28816 2440 28868 2446
rect 28816 2382 28868 2388
rect 28828 1970 28856 2382
rect 28632 1964 28684 1970
rect 28632 1906 28684 1912
rect 28816 1964 28868 1970
rect 28816 1906 28868 1912
rect 29000 1964 29052 1970
rect 29000 1906 29052 1912
rect 28080 1896 28132 1902
rect 28080 1838 28132 1844
rect 28080 1760 28132 1766
rect 28080 1702 28132 1708
rect 27908 1550 28028 1578
rect 27724 56 27844 82
rect 23400 54 23534 56
rect 23110 0 23166 54
rect 23478 0 23534 54
rect 24306 0 24362 56
rect 24766 0 24822 56
rect 25226 54 25360 56
rect 25226 0 25282 54
rect 25594 0 25650 56
rect 26422 0 26478 56
rect 26882 0 26938 56
rect 27342 0 27398 56
rect 27710 54 27844 56
rect 27710 0 27766 54
rect 27816 42 27844 54
rect 27908 42 27936 1550
rect 28092 1426 28120 1702
rect 28644 1426 28672 1906
rect 28080 1420 28132 1426
rect 28080 1362 28132 1368
rect 28632 1420 28684 1426
rect 28632 1362 28684 1368
rect 28540 1216 28592 1222
rect 28540 1158 28592 1164
rect 28552 56 28580 1158
rect 29012 56 29040 1906
rect 29472 56 29500 4542
rect 30012 4072 30064 4078
rect 30012 4014 30064 4020
rect 30024 3738 30052 4014
rect 30196 3936 30248 3942
rect 30196 3878 30248 3884
rect 30012 3732 30064 3738
rect 30012 3674 30064 3680
rect 30208 1970 30236 3878
rect 30196 1964 30248 1970
rect 30196 1906 30248 1912
rect 30300 1850 30328 7210
rect 30760 6866 30788 7278
rect 31036 7002 31064 7278
rect 32036 7200 32088 7206
rect 32036 7142 32088 7148
rect 31024 6996 31076 7002
rect 31024 6938 31076 6944
rect 30748 6860 30800 6866
rect 30748 6802 30800 6808
rect 30760 5234 30788 6802
rect 31024 6792 31076 6798
rect 31024 6734 31076 6740
rect 31036 6254 31064 6734
rect 31024 6248 31076 6254
rect 31024 6190 31076 6196
rect 31024 5772 31076 5778
rect 31024 5714 31076 5720
rect 31036 5234 31064 5714
rect 30748 5228 30800 5234
rect 30748 5170 30800 5176
rect 31024 5228 31076 5234
rect 31024 5170 31076 5176
rect 30760 4690 30788 5170
rect 31024 5024 31076 5030
rect 31024 4966 31076 4972
rect 31036 4690 31064 4966
rect 30748 4684 30800 4690
rect 30748 4626 30800 4632
rect 31024 4684 31076 4690
rect 31024 4626 31076 4632
rect 30760 4146 30788 4626
rect 31484 4480 31536 4486
rect 31484 4422 31536 4428
rect 30748 4140 30800 4146
rect 30748 4082 30800 4088
rect 30760 3602 30788 4082
rect 31116 3936 31168 3942
rect 31116 3878 31168 3884
rect 30748 3596 30800 3602
rect 30748 3538 30800 3544
rect 30760 1970 30788 3538
rect 31024 3528 31076 3534
rect 31024 3470 31076 3476
rect 31036 2990 31064 3470
rect 31024 2984 31076 2990
rect 31024 2926 31076 2932
rect 31024 2508 31076 2514
rect 31024 2450 31076 2456
rect 31036 1970 31064 2450
rect 30748 1964 30800 1970
rect 30748 1906 30800 1912
rect 31024 1964 31076 1970
rect 31024 1906 31076 1912
rect 30116 1822 30328 1850
rect 29840 56 29960 82
rect 27816 14 27936 42
rect 28538 0 28594 56
rect 28998 0 29054 56
rect 29458 0 29514 56
rect 29826 54 29960 56
rect 29826 0 29882 54
rect 29932 42 29960 54
rect 30116 42 30144 1822
rect 30196 1760 30248 1766
rect 30196 1702 30248 1708
rect 30208 1426 30236 1702
rect 30656 1556 30708 1562
rect 30656 1498 30708 1504
rect 30196 1420 30248 1426
rect 30196 1362 30248 1368
rect 30668 56 30696 1498
rect 30760 1426 30788 1906
rect 30748 1420 30800 1426
rect 30748 1362 30800 1368
rect 31128 56 31156 3878
rect 31496 82 31524 4422
rect 32048 82 32076 7142
rect 32876 6866 32904 7278
rect 33152 7002 33180 7278
rect 34152 7200 34204 7206
rect 34152 7142 34204 7148
rect 33140 6996 33192 7002
rect 33140 6938 33192 6944
rect 32864 6860 32916 6866
rect 32864 6802 32916 6808
rect 32876 5234 32904 6802
rect 33140 6792 33192 6798
rect 33140 6734 33192 6740
rect 33152 6254 33180 6734
rect 33140 6248 33192 6254
rect 33140 6190 33192 6196
rect 33048 5840 33100 5846
rect 33048 5782 33100 5788
rect 33060 5234 33088 5782
rect 32864 5228 32916 5234
rect 32864 5170 32916 5176
rect 33048 5228 33100 5234
rect 33048 5170 33100 5176
rect 32876 4690 32904 5170
rect 33140 5024 33192 5030
rect 33140 4966 33192 4972
rect 33152 4690 33180 4966
rect 32864 4684 32916 4690
rect 32864 4626 32916 4632
rect 33140 4684 33192 4690
rect 33140 4626 33192 4632
rect 32876 4146 32904 4626
rect 33784 4480 33836 4486
rect 33784 4422 33836 4428
rect 32864 4140 32916 4146
rect 32864 4082 32916 4088
rect 32128 4072 32180 4078
rect 32128 4014 32180 4020
rect 32140 3738 32168 4014
rect 32128 3732 32180 3738
rect 32128 3674 32180 3680
rect 32876 3602 32904 4082
rect 33232 3936 33284 3942
rect 33232 3878 33284 3884
rect 32864 3596 32916 3602
rect 32864 3538 32916 3544
rect 32876 1970 32904 3538
rect 33140 3528 33192 3534
rect 33140 3470 33192 3476
rect 33152 2922 33180 3470
rect 33140 2916 33192 2922
rect 33140 2858 33192 2864
rect 33140 2644 33192 2650
rect 33140 2586 33192 2592
rect 33152 1970 33180 2586
rect 32864 1964 32916 1970
rect 32864 1906 32916 1912
rect 33140 1964 33192 1970
rect 33140 1906 33192 1912
rect 32128 1760 32180 1766
rect 32128 1702 32180 1708
rect 32140 1426 32168 1702
rect 32876 1426 32904 1906
rect 32128 1420 32180 1426
rect 32128 1362 32180 1368
rect 32864 1420 32916 1426
rect 32864 1362 32916 1368
rect 33048 1216 33100 1222
rect 33048 1158 33100 1164
rect 31496 56 31616 82
rect 31956 56 32076 82
rect 32784 56 32904 82
rect 29932 14 30144 42
rect 30654 0 30710 56
rect 31114 0 31170 56
rect 31496 54 31630 56
rect 31574 0 31630 54
rect 31942 54 32076 56
rect 32770 54 32904 56
rect 31942 0 31998 54
rect 32770 0 32826 54
rect 32876 42 32904 54
rect 33060 42 33088 1158
rect 33244 56 33272 3878
rect 33796 82 33824 4422
rect 34164 82 34192 7142
rect 35084 6866 35112 7278
rect 35268 7002 35296 7278
rect 36176 7200 36228 7206
rect 36176 7142 36228 7148
rect 35256 6996 35308 7002
rect 35256 6938 35308 6944
rect 35072 6860 35124 6866
rect 35072 6802 35124 6808
rect 34736 6556 35032 6576
rect 34792 6554 34816 6556
rect 34872 6554 34896 6556
rect 34952 6554 34976 6556
rect 34814 6502 34816 6554
rect 34878 6502 34890 6554
rect 34952 6502 34954 6554
rect 34792 6500 34816 6502
rect 34872 6500 34896 6502
rect 34952 6500 34976 6502
rect 34736 6480 35032 6500
rect 34736 5468 35032 5488
rect 34792 5466 34816 5468
rect 34872 5466 34896 5468
rect 34952 5466 34976 5468
rect 34814 5414 34816 5466
rect 34878 5414 34890 5466
rect 34952 5414 34954 5466
rect 34792 5412 34816 5414
rect 34872 5412 34896 5414
rect 34952 5412 34976 5414
rect 34736 5392 35032 5412
rect 35084 5166 35112 6802
rect 35256 6792 35308 6798
rect 35256 6734 35308 6740
rect 35268 6254 35296 6734
rect 35256 6248 35308 6254
rect 35256 6190 35308 6196
rect 35256 5772 35308 5778
rect 35256 5714 35308 5720
rect 35268 5234 35296 5714
rect 35256 5228 35308 5234
rect 35256 5170 35308 5176
rect 35072 5160 35124 5166
rect 35072 5102 35124 5108
rect 35084 4690 35112 5102
rect 35256 5024 35308 5030
rect 35256 4966 35308 4972
rect 35268 4690 35296 4966
rect 35072 4684 35124 4690
rect 35072 4626 35124 4632
rect 35256 4684 35308 4690
rect 35256 4626 35308 4632
rect 34736 4380 35032 4400
rect 34792 4378 34816 4380
rect 34872 4378 34896 4380
rect 34952 4378 34976 4380
rect 34814 4326 34816 4378
rect 34878 4326 34890 4378
rect 34952 4326 34954 4378
rect 34792 4324 34816 4326
rect 34872 4324 34896 4326
rect 34952 4324 34976 4326
rect 34736 4304 35032 4324
rect 35084 4078 35112 4626
rect 35900 4480 35952 4486
rect 35900 4422 35952 4428
rect 34244 4072 34296 4078
rect 34244 4014 34296 4020
rect 35072 4072 35124 4078
rect 35072 4014 35124 4020
rect 35624 4072 35676 4078
rect 35624 4014 35676 4020
rect 34256 3738 34284 4014
rect 34244 3732 34296 3738
rect 34244 3674 34296 3680
rect 35084 3602 35112 4014
rect 35348 3936 35400 3942
rect 35348 3878 35400 3884
rect 35072 3596 35124 3602
rect 35072 3538 35124 3544
rect 34736 3292 35032 3312
rect 34792 3290 34816 3292
rect 34872 3290 34896 3292
rect 34952 3290 34976 3292
rect 34814 3238 34816 3290
rect 34878 3238 34890 3290
rect 34952 3238 34954 3290
rect 34792 3236 34816 3238
rect 34872 3236 34896 3238
rect 34952 3236 34976 3238
rect 34736 3216 35032 3236
rect 34736 2204 35032 2224
rect 34792 2202 34816 2204
rect 34872 2202 34896 2204
rect 34952 2202 34976 2204
rect 34814 2150 34816 2202
rect 34878 2150 34890 2202
rect 34952 2150 34954 2202
rect 34792 2148 34816 2150
rect 34872 2148 34896 2150
rect 34952 2148 34976 2150
rect 34736 2128 35032 2148
rect 35084 1902 35112 3538
rect 35256 3528 35308 3534
rect 35256 3470 35308 3476
rect 35268 2990 35296 3470
rect 35256 2984 35308 2990
rect 35256 2926 35308 2932
rect 35256 2508 35308 2514
rect 35256 2450 35308 2456
rect 35268 1970 35296 2450
rect 35256 1964 35308 1970
rect 35256 1906 35308 1912
rect 35072 1896 35124 1902
rect 35072 1838 35124 1844
rect 34244 1760 34296 1766
rect 34244 1702 34296 1708
rect 34256 1426 34284 1702
rect 35084 1426 35112 1838
rect 34244 1420 34296 1426
rect 34244 1362 34296 1368
rect 35072 1420 35124 1426
rect 35072 1362 35124 1368
rect 35256 1216 35308 1222
rect 35256 1158 35308 1164
rect 34736 1116 35032 1136
rect 34792 1114 34816 1116
rect 34872 1114 34896 1116
rect 34952 1114 34976 1116
rect 34814 1062 34816 1114
rect 34878 1062 34890 1114
rect 34952 1062 34954 1114
rect 34792 1060 34816 1062
rect 34872 1060 34896 1062
rect 34952 1060 34976 1062
rect 34736 1040 35032 1060
rect 33704 56 33824 82
rect 34072 56 34192 82
rect 34900 56 35020 82
rect 32876 14 33088 42
rect 33230 0 33286 56
rect 33690 54 33824 56
rect 34058 54 34192 56
rect 34886 54 35020 56
rect 33690 0 33746 54
rect 34058 0 34114 54
rect 34886 0 34942 54
rect 34992 42 35020 54
rect 35268 42 35296 1158
rect 35360 56 35388 3878
rect 35636 3534 35664 4014
rect 35624 3528 35676 3534
rect 35624 3470 35676 3476
rect 35532 1760 35584 1766
rect 35532 1702 35584 1708
rect 35544 1426 35572 1702
rect 35532 1420 35584 1426
rect 35532 1362 35584 1368
rect 35912 82 35940 4422
rect 35820 56 35940 82
rect 36188 56 36216 7142
rect 37108 6866 37136 7278
rect 37384 7002 37412 7278
rect 38384 7200 38436 7206
rect 38384 7142 38436 7148
rect 37372 6996 37424 7002
rect 37372 6938 37424 6944
rect 37096 6860 37148 6866
rect 37096 6802 37148 6808
rect 37108 5234 37136 6802
rect 37372 6792 37424 6798
rect 37372 6734 37424 6740
rect 37384 6254 37412 6734
rect 37372 6248 37424 6254
rect 37372 6190 37424 6196
rect 37372 5840 37424 5846
rect 37372 5782 37424 5788
rect 37384 5234 37412 5782
rect 37096 5228 37148 5234
rect 37096 5170 37148 5176
rect 37372 5228 37424 5234
rect 37372 5170 37424 5176
rect 37108 4690 37136 5170
rect 37372 5024 37424 5030
rect 37372 4966 37424 4972
rect 37384 4690 37412 4966
rect 37096 4684 37148 4690
rect 37096 4626 37148 4632
rect 37372 4684 37424 4690
rect 37372 4626 37424 4632
rect 37108 4146 37136 4626
rect 38016 4616 38068 4622
rect 37936 4564 38016 4570
rect 37936 4558 38068 4564
rect 37936 4542 38056 4558
rect 37096 4140 37148 4146
rect 37096 4082 37148 4088
rect 37108 3602 37136 4082
rect 37740 4072 37792 4078
rect 37740 4014 37792 4020
rect 37096 3596 37148 3602
rect 37096 3538 37148 3544
rect 37108 1970 37136 3538
rect 37752 3534 37780 4014
rect 37372 3528 37424 3534
rect 37372 3470 37424 3476
rect 37740 3528 37792 3534
rect 37740 3470 37792 3476
rect 37384 2990 37412 3470
rect 37372 2984 37424 2990
rect 37372 2926 37424 2932
rect 37372 2576 37424 2582
rect 37372 2518 37424 2524
rect 37384 1970 37412 2518
rect 37096 1964 37148 1970
rect 37096 1906 37148 1912
rect 37372 1964 37424 1970
rect 37372 1906 37424 1912
rect 37108 1426 37136 1906
rect 37464 1896 37516 1902
rect 37464 1838 37516 1844
rect 37096 1420 37148 1426
rect 37096 1362 37148 1368
rect 37280 1216 37332 1222
rect 37280 1158 37332 1164
rect 37016 56 37136 82
rect 34992 14 35296 42
rect 35346 0 35402 56
rect 35806 54 35940 56
rect 35806 0 35862 54
rect 36174 0 36230 56
rect 37002 54 37136 56
rect 37002 0 37058 54
rect 37108 42 37136 54
rect 37292 42 37320 1158
rect 37476 56 37504 1838
rect 37648 1760 37700 1766
rect 37648 1702 37700 1708
rect 37660 1426 37688 1702
rect 37648 1420 37700 1426
rect 37648 1362 37700 1368
rect 37936 56 37964 4542
rect 38396 82 38424 7142
rect 39224 6866 39252 7278
rect 39500 7002 39528 7278
rect 40500 7200 40552 7206
rect 40500 7142 40552 7148
rect 39488 6996 39540 7002
rect 39488 6938 39540 6944
rect 39212 6860 39264 6866
rect 39212 6802 39264 6808
rect 39224 5234 39252 6802
rect 39396 6792 39448 6798
rect 39396 6734 39448 6740
rect 39408 6186 39436 6734
rect 39396 6180 39448 6186
rect 39396 6122 39448 6128
rect 39488 5704 39540 5710
rect 39488 5646 39540 5652
rect 39500 5234 39528 5646
rect 39212 5228 39264 5234
rect 39212 5170 39264 5176
rect 39488 5228 39540 5234
rect 39488 5170 39540 5176
rect 39224 4690 39252 5170
rect 39488 5024 39540 5030
rect 39488 4966 39540 4972
rect 39500 4690 39528 4966
rect 39212 4684 39264 4690
rect 39212 4626 39264 4632
rect 39488 4684 39540 4690
rect 39488 4626 39540 4632
rect 39224 4146 39252 4626
rect 40132 4480 40184 4486
rect 40132 4422 40184 4428
rect 39212 4140 39264 4146
rect 39212 4082 39264 4088
rect 38476 3936 38528 3942
rect 38476 3878 38528 3884
rect 38488 1902 38516 3878
rect 39224 3602 39252 4082
rect 39948 4072 40000 4078
rect 40144 4026 40172 4422
rect 39948 4014 40000 4020
rect 39212 3596 39264 3602
rect 39212 3538 39264 3544
rect 39488 3596 39540 3602
rect 39488 3538 39540 3544
rect 39224 1970 39252 3538
rect 39500 2990 39528 3538
rect 39960 3534 39988 4014
rect 40052 3998 40172 4026
rect 39948 3528 40000 3534
rect 39948 3470 40000 3476
rect 39488 2984 39540 2990
rect 39488 2926 39540 2932
rect 39396 2440 39448 2446
rect 39396 2382 39448 2388
rect 39408 1970 39436 2382
rect 39212 1964 39264 1970
rect 39212 1906 39264 1912
rect 39396 1964 39448 1970
rect 39396 1906 39448 1912
rect 39580 1964 39632 1970
rect 39580 1906 39632 1912
rect 38476 1896 38528 1902
rect 38476 1838 38528 1844
rect 39224 1426 39252 1906
rect 39212 1420 39264 1426
rect 39212 1362 39264 1368
rect 39488 1216 39540 1222
rect 39488 1158 39540 1164
rect 38304 56 38424 82
rect 39132 56 39252 82
rect 37108 14 37320 42
rect 37462 0 37518 56
rect 37922 0 37978 56
rect 38290 54 38424 56
rect 39118 54 39252 56
rect 38290 0 38346 54
rect 39118 0 39174 54
rect 39224 42 39252 54
rect 39500 42 39528 1158
rect 39592 56 39620 1906
rect 40052 56 40080 3998
rect 40408 3596 40460 3602
rect 40408 3538 40460 3544
rect 40420 3194 40448 3538
rect 40408 3188 40460 3194
rect 40408 3130 40460 3136
rect 40512 1850 40540 7142
rect 41248 6866 41276 7278
rect 41616 7002 41644 7278
rect 42892 7200 42944 7206
rect 42892 7142 42944 7148
rect 41604 6996 41656 7002
rect 41604 6938 41656 6944
rect 41236 6860 41288 6866
rect 41236 6802 41288 6808
rect 41248 5234 41276 6802
rect 41604 6792 41656 6798
rect 41604 6734 41656 6740
rect 41616 6254 41644 6734
rect 41604 6248 41656 6254
rect 41604 6190 41656 6196
rect 41604 5568 41656 5574
rect 41604 5510 41656 5516
rect 41616 5234 41644 5510
rect 41236 5228 41288 5234
rect 41236 5170 41288 5176
rect 41604 5228 41656 5234
rect 41604 5170 41656 5176
rect 41248 4690 41276 5170
rect 41604 5024 41656 5030
rect 41604 4966 41656 4972
rect 41616 4690 41644 4966
rect 41236 4684 41288 4690
rect 41236 4626 41288 4632
rect 41604 4684 41656 4690
rect 41604 4626 41656 4632
rect 41248 4146 41276 4626
rect 42248 4480 42300 4486
rect 42248 4422 42300 4428
rect 41236 4140 41288 4146
rect 41236 4082 41288 4088
rect 41248 4026 41276 4082
rect 41972 4072 42024 4078
rect 41248 3998 41368 4026
rect 41972 4014 42024 4020
rect 40592 3936 40644 3942
rect 40592 3878 40644 3884
rect 40604 3618 40632 3878
rect 40604 3590 40724 3618
rect 41340 3602 41368 3998
rect 40696 1970 40724 3590
rect 41328 3596 41380 3602
rect 41328 3538 41380 3544
rect 41340 1970 41368 3538
rect 41984 3534 42012 4014
rect 41604 3528 41656 3534
rect 41604 3470 41656 3476
rect 41972 3528 42024 3534
rect 41972 3470 42024 3476
rect 41616 2990 41644 3470
rect 41604 2984 41656 2990
rect 41604 2926 41656 2932
rect 41604 2508 41656 2514
rect 41604 2450 41656 2456
rect 41616 1970 41644 2450
rect 40684 1964 40736 1970
rect 40684 1906 40736 1912
rect 41328 1964 41380 1970
rect 41328 1906 41380 1912
rect 41604 1964 41656 1970
rect 41604 1906 41656 1912
rect 41696 1964 41748 1970
rect 41696 1906 41748 1912
rect 40420 1822 40540 1850
rect 40132 1760 40184 1766
rect 40132 1702 40184 1708
rect 40144 1426 40172 1702
rect 40132 1420 40184 1426
rect 40132 1362 40184 1368
rect 40420 56 40448 1822
rect 41236 1556 41288 1562
rect 41236 1498 41288 1504
rect 41248 56 41276 1498
rect 41340 1426 41368 1906
rect 41328 1420 41380 1426
rect 41328 1362 41380 1368
rect 41708 56 41736 1906
rect 41972 1760 42024 1766
rect 41972 1702 42024 1708
rect 41984 1426 42012 1702
rect 41972 1420 42024 1426
rect 41972 1362 42024 1368
rect 42260 82 42288 4422
rect 42708 3936 42760 3942
rect 42708 3878 42760 3884
rect 42720 1970 42748 3878
rect 42708 1964 42760 1970
rect 42708 1906 42760 1912
rect 42904 1748 42932 7142
rect 43456 6866 43484 7278
rect 43732 7002 43760 7278
rect 44916 7200 44968 7206
rect 44916 7142 44968 7148
rect 43720 6996 43772 7002
rect 43720 6938 43772 6944
rect 43444 6860 43496 6866
rect 43444 6802 43496 6808
rect 43456 5234 43484 6802
rect 43720 6792 43772 6798
rect 43720 6734 43772 6740
rect 43732 6254 43760 6734
rect 43720 6248 43772 6254
rect 43720 6190 43772 6196
rect 43720 5840 43772 5846
rect 43720 5782 43772 5788
rect 43732 5234 43760 5782
rect 43444 5228 43496 5234
rect 43444 5170 43496 5176
rect 43720 5228 43772 5234
rect 43720 5170 43772 5176
rect 43456 4690 43484 5170
rect 43720 5024 43772 5030
rect 43720 4966 43772 4972
rect 43732 4690 43760 4966
rect 43444 4684 43496 4690
rect 43444 4626 43496 4632
rect 43720 4684 43772 4690
rect 43720 4626 43772 4632
rect 43456 4146 43484 4626
rect 44364 4480 44416 4486
rect 44364 4422 44416 4428
rect 43444 4140 43496 4146
rect 43444 4082 43496 4088
rect 43456 3602 43484 4082
rect 43444 3596 43496 3602
rect 43444 3538 43496 3544
rect 43456 1970 43484 3538
rect 43720 3528 43772 3534
rect 43720 3470 43772 3476
rect 43732 2990 43760 3470
rect 43720 2984 43772 2990
rect 43720 2926 43772 2932
rect 43720 2576 43772 2582
rect 43720 2518 43772 2524
rect 43732 1970 43760 2518
rect 43444 1964 43496 1970
rect 43444 1906 43496 1912
rect 43720 1964 43772 1970
rect 43720 1906 43772 1912
rect 43812 1964 43864 1970
rect 43812 1906 43864 1912
rect 42168 56 42288 82
rect 42536 1720 42932 1748
rect 42536 56 42564 1720
rect 43352 1556 43404 1562
rect 43352 1498 43404 1504
rect 43364 56 43392 1498
rect 43456 1426 43484 1906
rect 43444 1420 43496 1426
rect 43444 1362 43496 1368
rect 43824 56 43852 1906
rect 44376 82 44404 4422
rect 44824 4072 44876 4078
rect 44824 4014 44876 4020
rect 44836 3738 44864 4014
rect 44824 3732 44876 3738
rect 44824 3674 44876 3680
rect 44928 1578 44956 7142
rect 45572 6866 45600 7278
rect 45848 7002 45876 7278
rect 47216 7268 47268 7274
rect 47216 7210 47268 7216
rect 45836 6996 45888 7002
rect 45836 6938 45888 6944
rect 45560 6860 45612 6866
rect 45560 6802 45612 6808
rect 45572 5234 45600 6802
rect 45836 6792 45888 6798
rect 45836 6734 45888 6740
rect 45848 6254 45876 6734
rect 45836 6248 45888 6254
rect 45836 6190 45888 6196
rect 45836 5704 45888 5710
rect 45836 5646 45888 5652
rect 45848 5234 45876 5646
rect 45560 5228 45612 5234
rect 45560 5170 45612 5176
rect 45836 5228 45888 5234
rect 45836 5170 45888 5176
rect 45572 4690 45600 5170
rect 45836 5024 45888 5030
rect 45836 4966 45888 4972
rect 45848 4690 45876 4966
rect 45560 4684 45612 4690
rect 45560 4626 45612 4632
rect 45836 4684 45888 4690
rect 45836 4626 45888 4632
rect 45572 4146 45600 4626
rect 46480 4480 46532 4486
rect 46480 4422 46532 4428
rect 45560 4140 45612 4146
rect 45560 4082 45612 4088
rect 45008 3936 45060 3942
rect 45008 3878 45060 3884
rect 45020 1970 45048 3878
rect 45572 3602 45600 4082
rect 45560 3596 45612 3602
rect 45560 3538 45612 3544
rect 45572 1970 45600 3538
rect 45836 3528 45888 3534
rect 45836 3470 45888 3476
rect 45848 2990 45876 3470
rect 45836 2984 45888 2990
rect 45836 2926 45888 2932
rect 45836 2440 45888 2446
rect 45836 2382 45888 2388
rect 45848 1970 45876 2382
rect 45008 1964 45060 1970
rect 45008 1906 45060 1912
rect 45560 1964 45612 1970
rect 45560 1906 45612 1912
rect 45836 1964 45888 1970
rect 45836 1906 45888 1912
rect 45928 1964 45980 1970
rect 45928 1906 45980 1912
rect 45008 1760 45060 1766
rect 45008 1702 45060 1708
rect 44836 1550 44956 1578
rect 44284 56 44404 82
rect 44652 56 44772 82
rect 39224 14 39528 42
rect 39578 0 39634 56
rect 40038 0 40094 56
rect 40406 0 40462 56
rect 41234 0 41290 56
rect 41694 0 41750 56
rect 42154 54 42288 56
rect 42154 0 42210 54
rect 42522 0 42578 56
rect 43350 0 43406 56
rect 43810 0 43866 56
rect 44270 54 44404 56
rect 44638 54 44772 56
rect 44270 0 44326 54
rect 44638 0 44694 54
rect 44744 42 44772 54
rect 44836 42 44864 1550
rect 45020 1426 45048 1702
rect 45572 1426 45600 1906
rect 45008 1420 45060 1426
rect 45008 1362 45060 1368
rect 45560 1420 45612 1426
rect 45560 1362 45612 1368
rect 45468 1216 45520 1222
rect 45468 1158 45520 1164
rect 45480 56 45508 1158
rect 45940 56 45968 1906
rect 46492 82 46520 4422
rect 46940 4072 46992 4078
rect 46940 4014 46992 4020
rect 46952 3738 46980 4014
rect 47124 3936 47176 3942
rect 47124 3878 47176 3884
rect 46940 3732 46992 3738
rect 46940 3674 46992 3680
rect 47136 1970 47164 3878
rect 47124 1964 47176 1970
rect 47124 1906 47176 1912
rect 47228 1850 47256 7210
rect 47688 6866 47716 7278
rect 47964 7002 47992 7278
rect 48964 7200 49016 7206
rect 48964 7142 49016 7148
rect 47952 6996 48004 7002
rect 47952 6938 48004 6944
rect 47676 6860 47728 6866
rect 47676 6802 47728 6808
rect 47688 5234 47716 6802
rect 47952 6792 48004 6798
rect 47952 6734 48004 6740
rect 47964 6254 47992 6734
rect 47952 6248 48004 6254
rect 47952 6190 48004 6196
rect 47860 5840 47912 5846
rect 47860 5782 47912 5788
rect 47872 5234 47900 5782
rect 47676 5228 47728 5234
rect 47676 5170 47728 5176
rect 47860 5228 47912 5234
rect 47860 5170 47912 5176
rect 47688 4690 47716 5170
rect 47952 5024 48004 5030
rect 47952 4966 48004 4972
rect 47964 4690 47992 4966
rect 47676 4684 47728 4690
rect 47676 4626 47728 4632
rect 47952 4684 48004 4690
rect 47952 4626 48004 4632
rect 47688 4146 47716 4626
rect 48412 4480 48464 4486
rect 48412 4422 48464 4428
rect 47676 4140 47728 4146
rect 47676 4082 47728 4088
rect 47688 3602 47716 4082
rect 48044 3936 48096 3942
rect 48044 3878 48096 3884
rect 47676 3596 47728 3602
rect 47676 3538 47728 3544
rect 47688 1970 47716 3538
rect 47952 3528 48004 3534
rect 47952 3470 48004 3476
rect 47964 2990 47992 3470
rect 47952 2984 48004 2990
rect 47952 2926 48004 2932
rect 47860 2576 47912 2582
rect 47860 2518 47912 2524
rect 47872 1970 47900 2518
rect 47676 1964 47728 1970
rect 47676 1906 47728 1912
rect 47860 1964 47912 1970
rect 47860 1906 47912 1912
rect 47044 1822 47256 1850
rect 46400 56 46520 82
rect 46768 56 46888 82
rect 44744 14 44864 42
rect 45466 0 45522 56
rect 45926 0 45982 56
rect 46386 54 46520 56
rect 46754 54 46888 56
rect 46386 0 46442 54
rect 46754 0 46810 54
rect 46860 42 46888 54
rect 47044 42 47072 1822
rect 47124 1760 47176 1766
rect 47124 1702 47176 1708
rect 47136 1426 47164 1702
rect 47584 1556 47636 1562
rect 47584 1498 47636 1504
rect 47124 1420 47176 1426
rect 47124 1362 47176 1368
rect 47596 56 47624 1498
rect 47688 1426 47716 1906
rect 47676 1420 47728 1426
rect 47676 1362 47728 1368
rect 48056 56 48084 3878
rect 48424 82 48452 4422
rect 48976 82 49004 7142
rect 49804 6866 49832 7278
rect 51080 7200 51132 7206
rect 51080 7142 51132 7148
rect 50096 7100 50392 7120
rect 50152 7098 50176 7100
rect 50232 7098 50256 7100
rect 50312 7098 50336 7100
rect 50174 7046 50176 7098
rect 50238 7046 50250 7098
rect 50312 7046 50314 7098
rect 50152 7044 50176 7046
rect 50232 7044 50256 7046
rect 50312 7044 50336 7046
rect 50096 7024 50392 7044
rect 49792 6860 49844 6866
rect 49792 6802 49844 6808
rect 49804 5234 49832 6802
rect 50068 6792 50120 6798
rect 50068 6734 50120 6740
rect 50080 6186 50108 6734
rect 50068 6180 50120 6186
rect 50068 6122 50120 6128
rect 50096 6012 50392 6032
rect 50152 6010 50176 6012
rect 50232 6010 50256 6012
rect 50312 6010 50336 6012
rect 50174 5958 50176 6010
rect 50238 5958 50250 6010
rect 50312 5958 50314 6010
rect 50152 5956 50176 5958
rect 50232 5956 50256 5958
rect 50312 5956 50336 5958
rect 50096 5936 50392 5956
rect 50068 5772 50120 5778
rect 50068 5714 50120 5720
rect 50080 5234 50108 5714
rect 49792 5228 49844 5234
rect 49792 5170 49844 5176
rect 50068 5228 50120 5234
rect 50068 5170 50120 5176
rect 49804 4690 49832 5170
rect 50096 4924 50392 4944
rect 50152 4922 50176 4924
rect 50232 4922 50256 4924
rect 50312 4922 50336 4924
rect 50174 4870 50176 4922
rect 50238 4870 50250 4922
rect 50312 4870 50314 4922
rect 50152 4868 50176 4870
rect 50232 4868 50256 4870
rect 50312 4868 50336 4870
rect 50096 4848 50392 4868
rect 49792 4684 49844 4690
rect 49792 4626 49844 4632
rect 49804 4146 49832 4626
rect 50712 4480 50764 4486
rect 50712 4422 50764 4428
rect 49792 4140 49844 4146
rect 49792 4082 49844 4088
rect 49056 4072 49108 4078
rect 49056 4014 49108 4020
rect 49068 3738 49096 4014
rect 49056 3732 49108 3738
rect 49056 3674 49108 3680
rect 49804 3602 49832 4082
rect 50528 3936 50580 3942
rect 50528 3878 50580 3884
rect 50096 3836 50392 3856
rect 50152 3834 50176 3836
rect 50232 3834 50256 3836
rect 50312 3834 50336 3836
rect 50174 3782 50176 3834
rect 50238 3782 50250 3834
rect 50312 3782 50314 3834
rect 50152 3780 50176 3782
rect 50232 3780 50256 3782
rect 50312 3780 50336 3782
rect 50096 3760 50392 3780
rect 49792 3596 49844 3602
rect 49792 3538 49844 3544
rect 49804 1970 49832 3538
rect 50068 3528 50120 3534
rect 50068 3470 50120 3476
rect 50080 2922 50108 3470
rect 50068 2916 50120 2922
rect 50068 2858 50120 2864
rect 50096 2748 50392 2768
rect 50152 2746 50176 2748
rect 50232 2746 50256 2748
rect 50312 2746 50336 2748
rect 50174 2694 50176 2746
rect 50238 2694 50250 2746
rect 50312 2694 50314 2746
rect 50152 2692 50176 2694
rect 50232 2692 50256 2694
rect 50312 2692 50336 2694
rect 50096 2672 50392 2692
rect 50068 2508 50120 2514
rect 50068 2450 50120 2456
rect 50080 1970 50108 2450
rect 49792 1964 49844 1970
rect 49792 1906 49844 1912
rect 50068 1964 50120 1970
rect 50068 1906 50120 1912
rect 49056 1760 49108 1766
rect 49056 1702 49108 1708
rect 49068 1426 49096 1702
rect 49804 1426 49832 1906
rect 50096 1660 50392 1680
rect 50152 1658 50176 1660
rect 50232 1658 50256 1660
rect 50312 1658 50336 1660
rect 50174 1606 50176 1658
rect 50238 1606 50250 1658
rect 50312 1606 50314 1658
rect 50152 1604 50176 1606
rect 50232 1604 50256 1606
rect 50312 1604 50336 1606
rect 50096 1584 50392 1604
rect 49056 1420 49108 1426
rect 49056 1362 49108 1368
rect 49792 1420 49844 1426
rect 49792 1362 49844 1368
rect 49976 1216 50028 1222
rect 49976 1158 50028 1164
rect 48424 56 48544 82
rect 48884 56 49004 82
rect 49712 56 49832 82
rect 46860 14 47072 42
rect 47582 0 47638 56
rect 48042 0 48098 56
rect 48424 54 48558 56
rect 48502 0 48558 54
rect 48870 54 49004 56
rect 49698 54 49832 56
rect 48870 0 48926 54
rect 49698 0 49754 54
rect 49804 42 49832 54
rect 49988 42 50016 1158
rect 50172 56 50292 82
rect 49804 14 50016 42
rect 50158 54 50292 56
rect 50158 0 50214 54
rect 50264 42 50292 54
rect 50540 42 50568 3878
rect 50724 82 50752 4422
rect 51092 82 51120 7142
rect 51184 7002 51212 7278
rect 51172 6996 51224 7002
rect 51172 6938 51224 6944
rect 51920 6866 51948 7278
rect 52196 7002 52224 7278
rect 53288 7200 53340 7206
rect 53288 7142 53340 7148
rect 52184 6996 52236 7002
rect 52184 6938 52236 6944
rect 51908 6860 51960 6866
rect 51908 6802 51960 6808
rect 51920 5234 51948 6802
rect 52184 6792 52236 6798
rect 52184 6734 52236 6740
rect 52196 6254 52224 6734
rect 52184 6248 52236 6254
rect 52184 6190 52236 6196
rect 52184 5636 52236 5642
rect 52184 5578 52236 5584
rect 52196 5234 52224 5578
rect 51908 5228 51960 5234
rect 51908 5170 51960 5176
rect 52184 5228 52236 5234
rect 52184 5170 52236 5176
rect 51172 5024 51224 5030
rect 51172 4966 51224 4972
rect 51184 4690 51212 4966
rect 51920 4690 51948 5170
rect 52184 5024 52236 5030
rect 52184 4966 52236 4972
rect 52196 4690 52224 4966
rect 51172 4684 51224 4690
rect 51172 4626 51224 4632
rect 51908 4684 51960 4690
rect 51908 4626 51960 4632
rect 52184 4684 52236 4690
rect 52184 4626 52236 4632
rect 51920 4146 51948 4626
rect 52828 4480 52880 4486
rect 52828 4422 52880 4428
rect 51908 4140 51960 4146
rect 51908 4082 51960 4088
rect 51172 4072 51224 4078
rect 51172 4014 51224 4020
rect 51184 3738 51212 4014
rect 51172 3732 51224 3738
rect 51172 3674 51224 3680
rect 51920 3602 51948 4082
rect 52276 4072 52328 4078
rect 52276 4014 52328 4020
rect 51908 3596 51960 3602
rect 51908 3538 51960 3544
rect 51920 1970 51948 3538
rect 52288 3534 52316 4014
rect 52552 3936 52604 3942
rect 52552 3878 52604 3884
rect 52184 3528 52236 3534
rect 52184 3470 52236 3476
rect 52276 3528 52328 3534
rect 52276 3470 52328 3476
rect 52196 2990 52224 3470
rect 52184 2984 52236 2990
rect 52184 2926 52236 2932
rect 52184 2372 52236 2378
rect 52184 2314 52236 2320
rect 52196 1970 52224 2314
rect 51908 1964 51960 1970
rect 51908 1906 51960 1912
rect 52184 1964 52236 1970
rect 52184 1906 52236 1912
rect 51172 1760 51224 1766
rect 51172 1702 51224 1708
rect 51184 1426 51212 1702
rect 51920 1426 51948 1906
rect 52276 1760 52328 1766
rect 52276 1702 52328 1708
rect 52288 1426 52316 1702
rect 51172 1420 51224 1426
rect 51172 1362 51224 1368
rect 51908 1420 51960 1426
rect 51908 1362 51960 1368
rect 52276 1420 52328 1426
rect 52276 1362 52328 1368
rect 52184 1216 52236 1222
rect 52184 1158 52236 1164
rect 50632 56 50752 82
rect 51000 56 51120 82
rect 51828 56 51948 82
rect 50264 14 50568 42
rect 50618 54 50752 56
rect 50986 54 51120 56
rect 51814 54 51948 56
rect 50618 0 50674 54
rect 50986 0 51042 54
rect 51814 0 51870 54
rect 51920 42 51948 54
rect 52196 42 52224 1158
rect 52288 56 52408 82
rect 51920 14 52224 42
rect 52274 54 52408 56
rect 52274 0 52330 54
rect 52380 42 52408 54
rect 52564 42 52592 3878
rect 52840 82 52868 4422
rect 52748 56 52868 82
rect 53116 56 53236 82
rect 52380 14 52592 42
rect 52734 54 52868 56
rect 53102 54 53236 56
rect 52734 0 52790 54
rect 53102 0 53158 54
rect 53208 42 53236 54
rect 53300 42 53328 7142
rect 54036 6866 54064 7278
rect 54312 7002 54340 7278
rect 55312 7200 55364 7206
rect 55312 7142 55364 7148
rect 54300 6996 54352 7002
rect 54300 6938 54352 6944
rect 54024 6860 54076 6866
rect 54024 6802 54076 6808
rect 54036 5234 54064 6802
rect 54300 6792 54352 6798
rect 54300 6734 54352 6740
rect 54312 6254 54340 6734
rect 54300 6248 54352 6254
rect 54300 6190 54352 6196
rect 54208 5772 54260 5778
rect 54208 5714 54260 5720
rect 54220 5234 54248 5714
rect 54024 5228 54076 5234
rect 54024 5170 54076 5176
rect 54208 5228 54260 5234
rect 54208 5170 54260 5176
rect 54036 4690 54064 5170
rect 54300 5024 54352 5030
rect 54300 4966 54352 4972
rect 54312 4690 54340 4966
rect 54024 4684 54076 4690
rect 54024 4626 54076 4632
rect 54300 4684 54352 4690
rect 54300 4626 54352 4632
rect 54036 4146 54064 4626
rect 54944 4480 54996 4486
rect 54944 4422 54996 4428
rect 54024 4140 54076 4146
rect 54024 4082 54076 4088
rect 54036 3602 54064 4082
rect 54668 4072 54720 4078
rect 54668 4014 54720 4020
rect 54024 3596 54076 3602
rect 54024 3538 54076 3544
rect 54036 1970 54064 3538
rect 54680 3534 54708 4014
rect 54300 3528 54352 3534
rect 54300 3470 54352 3476
rect 54668 3528 54720 3534
rect 54668 3470 54720 3476
rect 54312 2990 54340 3470
rect 54300 2984 54352 2990
rect 54300 2926 54352 2932
rect 54208 2508 54260 2514
rect 54208 2450 54260 2456
rect 54220 1970 54248 2450
rect 54024 1964 54076 1970
rect 54024 1906 54076 1912
rect 54208 1964 54260 1970
rect 54208 1906 54260 1912
rect 54392 1964 54444 1970
rect 54392 1906 54444 1912
rect 54036 1426 54064 1906
rect 54024 1420 54076 1426
rect 54024 1362 54076 1368
rect 54208 1216 54260 1222
rect 54208 1158 54260 1164
rect 53944 56 54064 82
rect 53208 14 53328 42
rect 53930 54 54064 56
rect 53930 0 53986 54
rect 54036 42 54064 54
rect 54220 42 54248 1158
rect 54404 56 54432 1906
rect 54760 1760 54812 1766
rect 54760 1702 54812 1708
rect 54772 1426 54800 1702
rect 54760 1420 54812 1426
rect 54760 1362 54812 1368
rect 54956 82 54984 4422
rect 55324 82 55352 7142
rect 56060 6866 56088 7278
rect 56428 7002 56456 7278
rect 57428 7200 57480 7206
rect 57428 7142 57480 7148
rect 56416 6996 56468 7002
rect 56416 6938 56468 6944
rect 56048 6860 56100 6866
rect 56048 6802 56100 6808
rect 56060 5234 56088 6802
rect 56416 6792 56468 6798
rect 56416 6734 56468 6740
rect 56428 6254 56456 6734
rect 56416 6248 56468 6254
rect 56416 6190 56468 6196
rect 56416 5704 56468 5710
rect 56416 5646 56468 5652
rect 56428 5234 56456 5646
rect 56048 5228 56100 5234
rect 56048 5170 56100 5176
rect 56416 5228 56468 5234
rect 56416 5170 56468 5176
rect 56060 4690 56088 5170
rect 56416 5024 56468 5030
rect 56416 4966 56468 4972
rect 56428 4690 56456 4966
rect 56048 4684 56100 4690
rect 56048 4626 56100 4632
rect 56416 4684 56468 4690
rect 56416 4626 56468 4632
rect 56060 4060 56088 4626
rect 57060 4480 57112 4486
rect 57060 4422 57112 4428
rect 56140 4072 56192 4078
rect 56060 4032 56140 4060
rect 56140 4014 56192 4020
rect 55404 3936 55456 3942
rect 55404 3878 55456 3884
rect 55416 1970 55444 3878
rect 56152 3602 56180 4014
rect 56140 3596 56192 3602
rect 56140 3538 56192 3544
rect 56152 1970 56180 3538
rect 56416 3528 56468 3534
rect 56416 3470 56468 3476
rect 56428 2990 56456 3470
rect 56416 2984 56468 2990
rect 56416 2926 56468 2932
rect 56416 2440 56468 2446
rect 56416 2382 56468 2388
rect 56428 1970 56456 2382
rect 55404 1964 55456 1970
rect 55404 1906 55456 1912
rect 56140 1964 56192 1970
rect 56140 1906 56192 1912
rect 56416 1964 56468 1970
rect 56416 1906 56468 1912
rect 56152 1426 56180 1906
rect 56508 1896 56560 1902
rect 56508 1838 56560 1844
rect 56140 1420 56192 1426
rect 56140 1362 56192 1368
rect 56416 1216 56468 1222
rect 56416 1158 56468 1164
rect 54864 56 54984 82
rect 55232 56 55352 82
rect 56060 56 56180 82
rect 54036 14 54248 42
rect 54390 0 54446 56
rect 54850 54 54984 56
rect 55218 54 55352 56
rect 56046 54 56180 56
rect 54850 0 54906 54
rect 55218 0 55274 54
rect 56046 0 56102 54
rect 56152 42 56180 54
rect 56428 42 56456 1158
rect 56520 56 56548 1838
rect 56692 1760 56744 1766
rect 56692 1702 56744 1708
rect 56704 1426 56732 1702
rect 56692 1420 56744 1426
rect 56692 1362 56744 1368
rect 57072 82 57100 4422
rect 57152 4072 57204 4078
rect 57152 4014 57204 4020
rect 57164 3534 57192 4014
rect 57152 3528 57204 3534
rect 57152 3470 57204 3476
rect 57440 1884 57468 7142
rect 58176 6866 58204 7278
rect 58544 7002 58572 7278
rect 59728 7200 59780 7206
rect 59728 7142 59780 7148
rect 58532 6996 58584 7002
rect 58532 6938 58584 6944
rect 58164 6860 58216 6866
rect 58164 6802 58216 6808
rect 58176 5234 58204 6802
rect 58532 6792 58584 6798
rect 58532 6734 58584 6740
rect 58544 6254 58572 6734
rect 58532 6248 58584 6254
rect 58532 6190 58584 6196
rect 58440 5840 58492 5846
rect 58440 5782 58492 5788
rect 58452 5234 58480 5782
rect 58164 5228 58216 5234
rect 58164 5170 58216 5176
rect 58440 5228 58492 5234
rect 58440 5170 58492 5176
rect 58176 4690 58204 5170
rect 58532 5024 58584 5030
rect 58532 4966 58584 4972
rect 58544 4690 58572 4966
rect 58164 4684 58216 4690
rect 58164 4626 58216 4632
rect 58532 4684 58584 4690
rect 58532 4626 58584 4632
rect 58176 4214 58204 4626
rect 59176 4480 59228 4486
rect 59176 4422 59228 4428
rect 58164 4208 58216 4214
rect 58216 4156 58296 4162
rect 58164 4150 58296 4156
rect 58176 4134 58296 4150
rect 57520 3936 57572 3942
rect 57520 3878 57572 3884
rect 57532 1902 57560 3878
rect 58268 3602 58296 4134
rect 58992 4072 59044 4078
rect 58992 4014 59044 4020
rect 58256 3596 58308 3602
rect 58256 3538 58308 3544
rect 58268 1970 58296 3538
rect 59004 3534 59032 4014
rect 58532 3528 58584 3534
rect 58532 3470 58584 3476
rect 58992 3528 59044 3534
rect 58992 3470 59044 3476
rect 58544 2990 58572 3470
rect 58532 2984 58584 2990
rect 58532 2926 58584 2932
rect 58440 2576 58492 2582
rect 58440 2518 58492 2524
rect 58452 1970 58480 2518
rect 58624 2100 58676 2106
rect 58624 2042 58676 2048
rect 58256 1964 58308 1970
rect 58256 1906 58308 1912
rect 58440 1964 58492 1970
rect 58440 1906 58492 1912
rect 56980 56 57100 82
rect 57348 1856 57468 1884
rect 57520 1896 57572 1902
rect 57348 56 57376 1856
rect 57520 1838 57572 1844
rect 58164 1556 58216 1562
rect 58164 1498 58216 1504
rect 58176 56 58204 1498
rect 58268 1426 58296 1906
rect 58256 1420 58308 1426
rect 58256 1362 58308 1368
rect 58636 56 58664 2042
rect 58900 1760 58952 1766
rect 58900 1702 58952 1708
rect 58912 1426 58940 1702
rect 58900 1420 58952 1426
rect 58900 1362 58952 1368
rect 59188 82 59216 4422
rect 59636 3936 59688 3942
rect 59636 3878 59688 3884
rect 59648 2106 59676 3878
rect 59636 2100 59688 2106
rect 59636 2042 59688 2048
rect 59740 1884 59768 7142
rect 60384 6798 60412 7278
rect 60660 7002 60688 7278
rect 61844 7200 61896 7206
rect 61844 7142 61896 7148
rect 60648 6996 60700 7002
rect 60648 6938 60700 6944
rect 60372 6792 60424 6798
rect 60372 6734 60424 6740
rect 60648 6792 60700 6798
rect 60648 6734 60700 6740
rect 60384 5166 60412 6734
rect 60660 6254 60688 6734
rect 60648 6248 60700 6254
rect 60648 6190 60700 6196
rect 60464 5840 60516 5846
rect 60516 5788 60596 5794
rect 60464 5782 60596 5788
rect 60476 5766 60596 5782
rect 60568 5234 60596 5766
rect 60556 5228 60608 5234
rect 60556 5170 60608 5176
rect 60372 5160 60424 5166
rect 60372 5102 60424 5108
rect 60384 4622 60412 5102
rect 60648 5024 60700 5030
rect 60648 4966 60700 4972
rect 60660 4690 60688 4966
rect 60648 4684 60700 4690
rect 60648 4626 60700 4632
rect 60372 4616 60424 4622
rect 60372 4558 60424 4564
rect 60384 4078 60412 4558
rect 61292 4480 61344 4486
rect 61292 4422 61344 4428
rect 61304 4162 61332 4422
rect 61212 4134 61332 4162
rect 60372 4072 60424 4078
rect 60372 4014 60424 4020
rect 60384 3602 60412 4014
rect 60372 3596 60424 3602
rect 60372 3538 60424 3544
rect 60384 1970 60412 3538
rect 60648 3528 60700 3534
rect 60648 3470 60700 3476
rect 60660 2990 60688 3470
rect 60648 2984 60700 2990
rect 60648 2926 60700 2932
rect 60464 2576 60516 2582
rect 60464 2518 60516 2524
rect 60372 1964 60424 1970
rect 60372 1906 60424 1912
rect 59096 56 59216 82
rect 59464 1856 59768 1884
rect 59464 56 59492 1856
rect 60384 1426 60412 1906
rect 60476 1902 60504 2518
rect 60464 1896 60516 1902
rect 60464 1838 60516 1844
rect 60740 1896 60792 1902
rect 60740 1838 60792 1844
rect 60372 1420 60424 1426
rect 60372 1362 60424 1368
rect 60280 1216 60332 1222
rect 60280 1158 60332 1164
rect 60292 56 60320 1158
rect 60752 56 60780 1838
rect 61212 56 61240 4134
rect 61292 4072 61344 4078
rect 61292 4014 61344 4020
rect 61304 3534 61332 4014
rect 61292 3528 61344 3534
rect 61292 3470 61344 3476
rect 61856 1578 61884 7142
rect 62500 6866 62528 7278
rect 62776 7002 62804 7278
rect 64144 7268 64196 7274
rect 64144 7210 64196 7216
rect 62764 6996 62816 7002
rect 62764 6938 62816 6944
rect 62488 6860 62540 6866
rect 62488 6802 62540 6808
rect 62500 5234 62528 6802
rect 62764 6792 62816 6798
rect 62764 6734 62816 6740
rect 62776 6254 62804 6734
rect 62764 6248 62816 6254
rect 62764 6190 62816 6196
rect 62764 5840 62816 5846
rect 62764 5782 62816 5788
rect 62776 5234 62804 5782
rect 62488 5228 62540 5234
rect 62488 5170 62540 5176
rect 62764 5228 62816 5234
rect 62764 5170 62816 5176
rect 62500 4690 62528 5170
rect 62764 5024 62816 5030
rect 62764 4966 62816 4972
rect 62776 4690 62804 4966
rect 62488 4684 62540 4690
rect 62488 4626 62540 4632
rect 62764 4684 62816 4690
rect 62764 4626 62816 4632
rect 62500 4146 62528 4626
rect 63408 4480 63460 4486
rect 63408 4422 63460 4428
rect 62488 4140 62540 4146
rect 62488 4082 62540 4088
rect 61936 3936 61988 3942
rect 61936 3878 61988 3884
rect 61948 1902 61976 3878
rect 62500 3602 62528 4082
rect 62488 3596 62540 3602
rect 62488 3538 62540 3544
rect 62500 1970 62528 3538
rect 62764 3528 62816 3534
rect 62764 3470 62816 3476
rect 62776 2990 62804 3470
rect 62764 2984 62816 2990
rect 62764 2926 62816 2932
rect 62764 2576 62816 2582
rect 62764 2518 62816 2524
rect 62776 1970 62804 2518
rect 62488 1964 62540 1970
rect 62488 1906 62540 1912
rect 62764 1964 62816 1970
rect 62764 1906 62816 1912
rect 62856 1964 62908 1970
rect 62856 1906 62908 1912
rect 61936 1896 61988 1902
rect 61936 1838 61988 1844
rect 61936 1760 61988 1766
rect 61936 1702 61988 1708
rect 61764 1550 61884 1578
rect 61580 56 61700 82
rect 56152 14 56456 42
rect 56506 0 56562 56
rect 56966 54 57100 56
rect 56966 0 57022 54
rect 57334 0 57390 56
rect 58162 0 58218 56
rect 58622 0 58678 56
rect 59082 54 59216 56
rect 59082 0 59138 54
rect 59450 0 59506 56
rect 60278 0 60334 56
rect 60738 0 60794 56
rect 61198 0 61254 56
rect 61566 54 61700 56
rect 61566 0 61622 54
rect 61672 42 61700 54
rect 61764 42 61792 1550
rect 61948 1426 61976 1702
rect 62500 1426 62528 1906
rect 61936 1420 61988 1426
rect 61936 1362 61988 1368
rect 62488 1420 62540 1426
rect 62488 1362 62540 1368
rect 62396 1216 62448 1222
rect 62396 1158 62448 1164
rect 62408 56 62436 1158
rect 62868 56 62896 1906
rect 63420 82 63448 4422
rect 63868 4072 63920 4078
rect 63868 4014 63920 4020
rect 63880 3738 63908 4014
rect 64052 3936 64104 3942
rect 64052 3878 64104 3884
rect 63868 3732 63920 3738
rect 63868 3674 63920 3680
rect 64064 1970 64092 3878
rect 64052 1964 64104 1970
rect 64052 1906 64104 1912
rect 64156 1850 64184 7210
rect 64616 6866 64644 7278
rect 64892 7002 64920 7278
rect 65892 7200 65944 7206
rect 65892 7142 65944 7148
rect 64880 6996 64932 7002
rect 64880 6938 64932 6944
rect 64604 6860 64656 6866
rect 64604 6802 64656 6808
rect 64616 5234 64644 6802
rect 64880 6792 64932 6798
rect 64880 6734 64932 6740
rect 64892 6254 64920 6734
rect 65456 6556 65752 6576
rect 65512 6554 65536 6556
rect 65592 6554 65616 6556
rect 65672 6554 65696 6556
rect 65534 6502 65536 6554
rect 65598 6502 65610 6554
rect 65672 6502 65674 6554
rect 65512 6500 65536 6502
rect 65592 6500 65616 6502
rect 65672 6500 65696 6502
rect 65456 6480 65752 6500
rect 64880 6248 64932 6254
rect 64880 6190 64932 6196
rect 64788 5772 64840 5778
rect 64788 5714 64840 5720
rect 64800 5234 64828 5714
rect 65456 5468 65752 5488
rect 65512 5466 65536 5468
rect 65592 5466 65616 5468
rect 65672 5466 65696 5468
rect 65534 5414 65536 5466
rect 65598 5414 65610 5466
rect 65672 5414 65674 5466
rect 65512 5412 65536 5414
rect 65592 5412 65616 5414
rect 65672 5412 65696 5414
rect 65456 5392 65752 5412
rect 64604 5228 64656 5234
rect 64604 5170 64656 5176
rect 64788 5228 64840 5234
rect 64788 5170 64840 5176
rect 64616 4690 64644 5170
rect 64880 5024 64932 5030
rect 64880 4966 64932 4972
rect 64892 4690 64920 4966
rect 64604 4684 64656 4690
rect 64604 4626 64656 4632
rect 64880 4684 64932 4690
rect 64880 4626 64932 4632
rect 64616 4146 64644 4626
rect 65340 4480 65392 4486
rect 65340 4422 65392 4428
rect 64604 4140 64656 4146
rect 64604 4082 64656 4088
rect 64616 3602 64644 4082
rect 64972 3936 65024 3942
rect 64972 3878 65024 3884
rect 64604 3596 64656 3602
rect 64604 3538 64656 3544
rect 64616 1970 64644 3538
rect 64880 3528 64932 3534
rect 64880 3470 64932 3476
rect 64892 2990 64920 3470
rect 64880 2984 64932 2990
rect 64880 2926 64932 2932
rect 64788 2508 64840 2514
rect 64788 2450 64840 2456
rect 64800 1970 64828 2450
rect 64604 1964 64656 1970
rect 64604 1906 64656 1912
rect 64788 1964 64840 1970
rect 64788 1906 64840 1912
rect 63972 1822 64184 1850
rect 63328 56 63448 82
rect 63696 56 63816 82
rect 61672 14 61792 42
rect 62394 0 62450 56
rect 62854 0 62910 56
rect 63314 54 63448 56
rect 63682 54 63816 56
rect 63314 0 63370 54
rect 63682 0 63738 54
rect 63788 42 63816 54
rect 63972 42 64000 1822
rect 64052 1760 64104 1766
rect 64052 1702 64104 1708
rect 64064 1426 64092 1702
rect 64512 1556 64564 1562
rect 64512 1498 64564 1504
rect 64052 1420 64104 1426
rect 64052 1362 64104 1368
rect 64524 56 64552 1498
rect 64616 1426 64644 1906
rect 64604 1420 64656 1426
rect 64604 1362 64656 1368
rect 64984 56 65012 3878
rect 65352 898 65380 4422
rect 65456 4380 65752 4400
rect 65512 4378 65536 4380
rect 65592 4378 65616 4380
rect 65672 4378 65696 4380
rect 65534 4326 65536 4378
rect 65598 4326 65610 4378
rect 65672 4326 65674 4378
rect 65512 4324 65536 4326
rect 65592 4324 65616 4326
rect 65672 4324 65696 4326
rect 65456 4304 65752 4324
rect 65456 3292 65752 3312
rect 65512 3290 65536 3292
rect 65592 3290 65616 3292
rect 65672 3290 65696 3292
rect 65534 3238 65536 3290
rect 65598 3238 65610 3290
rect 65672 3238 65674 3290
rect 65512 3236 65536 3238
rect 65592 3236 65616 3238
rect 65672 3236 65696 3238
rect 65456 3216 65752 3236
rect 65456 2204 65752 2224
rect 65512 2202 65536 2204
rect 65592 2202 65616 2204
rect 65672 2202 65696 2204
rect 65534 2150 65536 2202
rect 65598 2150 65610 2202
rect 65672 2150 65674 2202
rect 65512 2148 65536 2150
rect 65592 2148 65616 2150
rect 65672 2148 65696 2150
rect 65456 2128 65752 2148
rect 65456 1116 65752 1136
rect 65512 1114 65536 1116
rect 65592 1114 65616 1116
rect 65672 1114 65696 1116
rect 65534 1062 65536 1114
rect 65598 1062 65610 1114
rect 65672 1062 65674 1114
rect 65512 1060 65536 1062
rect 65592 1060 65616 1062
rect 65672 1060 65696 1062
rect 65456 1040 65752 1060
rect 65352 870 65472 898
rect 65444 56 65472 870
rect 65904 82 65932 7142
rect 66732 6866 66760 7278
rect 67008 7002 67036 7278
rect 68008 7200 68060 7206
rect 68008 7142 68060 7148
rect 66996 6996 67048 7002
rect 66996 6938 67048 6944
rect 66720 6860 66772 6866
rect 66720 6802 66772 6808
rect 66732 5234 66760 6802
rect 66996 6792 67048 6798
rect 66996 6734 67048 6740
rect 67008 6254 67036 6734
rect 66996 6248 67048 6254
rect 66996 6190 67048 6196
rect 66996 5772 67048 5778
rect 66996 5714 67048 5720
rect 67008 5234 67036 5714
rect 66720 5228 66772 5234
rect 66720 5170 66772 5176
rect 66996 5228 67048 5234
rect 66996 5170 67048 5176
rect 66732 4690 66760 5170
rect 66996 5024 67048 5030
rect 66996 4966 67048 4972
rect 67008 4690 67036 4966
rect 66720 4684 66772 4690
rect 66720 4626 66772 4632
rect 66996 4684 67048 4690
rect 66996 4626 67048 4632
rect 66732 4146 66760 4626
rect 67640 4480 67692 4486
rect 67640 4422 67692 4428
rect 66720 4140 66772 4146
rect 66720 4082 66772 4088
rect 65984 4072 66036 4078
rect 65984 4014 66036 4020
rect 65996 3738 66024 4014
rect 65984 3732 66036 3738
rect 65984 3674 66036 3680
rect 66732 3602 66760 4082
rect 67088 3936 67140 3942
rect 67088 3878 67140 3884
rect 66720 3596 66772 3602
rect 66720 3538 66772 3544
rect 66732 1970 66760 3538
rect 66996 3528 67048 3534
rect 66996 3470 67048 3476
rect 67008 2922 67036 3470
rect 66996 2916 67048 2922
rect 66996 2858 67048 2864
rect 66996 2508 67048 2514
rect 66996 2450 67048 2456
rect 67008 1970 67036 2450
rect 66720 1964 66772 1970
rect 66720 1906 66772 1912
rect 66996 1964 67048 1970
rect 66996 1906 67048 1912
rect 65984 1760 66036 1766
rect 65984 1702 66036 1708
rect 65996 1426 66024 1702
rect 66732 1426 66760 1906
rect 65984 1420 66036 1426
rect 65984 1362 66036 1368
rect 66720 1420 66772 1426
rect 66720 1362 66772 1368
rect 66904 1216 66956 1222
rect 66904 1158 66956 1164
rect 65812 56 65932 82
rect 66640 56 66760 82
rect 63788 14 64000 42
rect 64510 0 64566 56
rect 64970 0 65026 56
rect 65430 0 65486 56
rect 65798 54 65932 56
rect 66626 54 66760 56
rect 65798 0 65854 54
rect 66626 0 66682 54
rect 66732 42 66760 54
rect 66916 42 66944 1158
rect 67100 56 67128 3878
rect 67652 82 67680 4422
rect 68020 82 68048 7142
rect 68848 6866 68876 7278
rect 69124 7002 69152 7278
rect 70216 7200 70268 7206
rect 70216 7142 70268 7148
rect 69112 6996 69164 7002
rect 69112 6938 69164 6944
rect 68836 6860 68888 6866
rect 68836 6802 68888 6808
rect 68848 5234 68876 6802
rect 69112 6792 69164 6798
rect 69112 6734 69164 6740
rect 69124 6254 69152 6734
rect 69112 6248 69164 6254
rect 69112 6190 69164 6196
rect 69112 5636 69164 5642
rect 69112 5578 69164 5584
rect 69124 5234 69152 5578
rect 68836 5228 68888 5234
rect 68836 5170 68888 5176
rect 69112 5228 69164 5234
rect 69112 5170 69164 5176
rect 68848 4690 68876 5170
rect 69112 5024 69164 5030
rect 69112 4966 69164 4972
rect 69124 4690 69152 4966
rect 68836 4684 68888 4690
rect 68836 4626 68888 4632
rect 69112 4684 69164 4690
rect 69112 4626 69164 4632
rect 68848 4146 68876 4626
rect 69756 4480 69808 4486
rect 69756 4422 69808 4428
rect 68836 4140 68888 4146
rect 68836 4082 68888 4088
rect 68100 4072 68152 4078
rect 68100 4014 68152 4020
rect 68112 3738 68140 4014
rect 68100 3732 68152 3738
rect 68100 3674 68152 3680
rect 68848 3602 68876 4082
rect 69204 4072 69256 4078
rect 69204 4014 69256 4020
rect 68836 3596 68888 3602
rect 68836 3538 68888 3544
rect 68848 1970 68876 3538
rect 69216 3534 69244 4014
rect 69480 3936 69532 3942
rect 69480 3878 69532 3884
rect 69112 3528 69164 3534
rect 69112 3470 69164 3476
rect 69204 3528 69256 3534
rect 69204 3470 69256 3476
rect 69124 2990 69152 3470
rect 69112 2984 69164 2990
rect 69112 2926 69164 2932
rect 69112 2372 69164 2378
rect 69112 2314 69164 2320
rect 69124 1970 69152 2314
rect 68836 1964 68888 1970
rect 68836 1906 68888 1912
rect 69112 1964 69164 1970
rect 69112 1906 69164 1912
rect 68100 1760 68152 1766
rect 68100 1702 68152 1708
rect 68112 1426 68140 1702
rect 68848 1426 68876 1906
rect 69204 1760 69256 1766
rect 69204 1702 69256 1708
rect 69216 1426 69244 1702
rect 68100 1420 68152 1426
rect 68100 1362 68152 1368
rect 68836 1420 68888 1426
rect 68836 1362 68888 1368
rect 69204 1420 69256 1426
rect 69204 1362 69256 1368
rect 69112 1216 69164 1222
rect 69112 1158 69164 1164
rect 67560 56 67680 82
rect 67928 56 68048 82
rect 68756 56 68876 82
rect 66732 14 66944 42
rect 67086 0 67142 56
rect 67546 54 67680 56
rect 67914 54 68048 56
rect 68742 54 68876 56
rect 67546 0 67602 54
rect 67914 0 67970 54
rect 68742 0 68798 54
rect 68848 42 68876 54
rect 69124 42 69152 1158
rect 69216 56 69336 82
rect 68848 14 69152 42
rect 69202 54 69336 56
rect 69202 0 69258 54
rect 69308 42 69336 54
rect 69492 42 69520 3878
rect 69768 82 69796 4422
rect 69676 56 69796 82
rect 70044 56 70164 82
rect 69308 14 69520 42
rect 69662 54 69796 56
rect 70030 54 70164 56
rect 69662 0 69718 54
rect 70030 0 70086 54
rect 70136 42 70164 54
rect 70228 42 70256 7142
rect 70872 6866 70900 7278
rect 71240 7002 71268 7278
rect 72240 7200 72292 7206
rect 72240 7142 72292 7148
rect 71228 6996 71280 7002
rect 71228 6938 71280 6944
rect 70860 6860 70912 6866
rect 70860 6802 70912 6808
rect 70872 5234 70900 6802
rect 71228 6792 71280 6798
rect 71228 6734 71280 6740
rect 71240 6254 71268 6734
rect 71228 6248 71280 6254
rect 71228 6190 71280 6196
rect 71228 5772 71280 5778
rect 71228 5714 71280 5720
rect 71240 5234 71268 5714
rect 70860 5228 70912 5234
rect 70860 5170 70912 5176
rect 71228 5228 71280 5234
rect 71228 5170 71280 5176
rect 70872 4690 70900 5170
rect 71228 5024 71280 5030
rect 71228 4966 71280 4972
rect 71240 4690 71268 4966
rect 70860 4684 70912 4690
rect 70860 4626 70912 4632
rect 71228 4684 71280 4690
rect 71228 4626 71280 4632
rect 70872 4214 70900 4626
rect 71872 4480 71924 4486
rect 71872 4422 71924 4428
rect 70860 4208 70912 4214
rect 70912 4156 70992 4162
rect 70860 4150 70992 4156
rect 70872 4134 70992 4150
rect 70964 3602 70992 4134
rect 71688 4072 71740 4078
rect 71688 4014 71740 4020
rect 70952 3596 71004 3602
rect 70952 3538 71004 3544
rect 70964 1970 70992 3538
rect 71700 3534 71728 4014
rect 71228 3528 71280 3534
rect 71228 3470 71280 3476
rect 71688 3528 71740 3534
rect 71688 3470 71740 3476
rect 71240 2990 71268 3470
rect 71228 2984 71280 2990
rect 71228 2926 71280 2932
rect 71228 2508 71280 2514
rect 71228 2450 71280 2456
rect 71240 1970 71268 2450
rect 70952 1964 71004 1970
rect 70952 1906 71004 1912
rect 71228 1964 71280 1970
rect 71228 1906 71280 1912
rect 70964 1426 70992 1906
rect 71320 1896 71372 1902
rect 71320 1838 71372 1844
rect 70952 1420 71004 1426
rect 70952 1362 71004 1368
rect 71136 1216 71188 1222
rect 71136 1158 71188 1164
rect 70872 56 70992 82
rect 70136 14 70256 42
rect 70858 54 70992 56
rect 70858 0 70914 54
rect 70964 42 70992 54
rect 71148 42 71176 1158
rect 71332 56 71360 1838
rect 71504 1760 71556 1766
rect 71504 1702 71556 1708
rect 71516 1426 71544 1702
rect 71504 1420 71556 1426
rect 71504 1362 71556 1368
rect 71884 82 71912 4422
rect 72252 82 72280 7142
rect 72988 6866 73016 7278
rect 73356 7002 73384 7278
rect 74356 7200 74408 7206
rect 74356 7142 74408 7148
rect 73344 6996 73396 7002
rect 73344 6938 73396 6944
rect 72976 6860 73028 6866
rect 72976 6802 73028 6808
rect 72988 5234 73016 6802
rect 73344 6792 73396 6798
rect 73344 6734 73396 6740
rect 73356 6254 73384 6734
rect 73344 6248 73396 6254
rect 73344 6190 73396 6196
rect 73344 5840 73396 5846
rect 73344 5782 73396 5788
rect 73356 5234 73384 5782
rect 72976 5228 73028 5234
rect 72976 5170 73028 5176
rect 73344 5228 73396 5234
rect 73344 5170 73396 5176
rect 72988 4690 73016 5170
rect 73344 5024 73396 5030
rect 73344 4966 73396 4972
rect 73356 4690 73384 4966
rect 72976 4684 73028 4690
rect 73344 4684 73396 4690
rect 73028 4644 73108 4672
rect 72976 4626 73028 4632
rect 73080 4146 73108 4644
rect 73344 4626 73396 4632
rect 73988 4480 74040 4486
rect 73988 4422 74040 4428
rect 73068 4140 73120 4146
rect 73068 4082 73120 4088
rect 72332 3936 72384 3942
rect 72332 3878 72384 3884
rect 72344 1902 72372 3878
rect 73080 3602 73108 4082
rect 73712 4072 73764 4078
rect 73712 4014 73764 4020
rect 73068 3596 73120 3602
rect 73068 3538 73120 3544
rect 73080 1970 73108 3538
rect 73724 3534 73752 4014
rect 73344 3528 73396 3534
rect 73344 3470 73396 3476
rect 73712 3528 73764 3534
rect 73712 3470 73764 3476
rect 73356 2990 73384 3470
rect 73344 2984 73396 2990
rect 73344 2926 73396 2932
rect 73344 2576 73396 2582
rect 73344 2518 73396 2524
rect 73356 1970 73384 2518
rect 73068 1964 73120 1970
rect 73068 1906 73120 1912
rect 73344 1964 73396 1970
rect 73344 1906 73396 1912
rect 72332 1896 72384 1902
rect 72332 1838 72384 1844
rect 73080 1426 73108 1906
rect 73436 1896 73488 1902
rect 73436 1838 73488 1844
rect 73068 1420 73120 1426
rect 73068 1362 73120 1368
rect 73344 1216 73396 1222
rect 73344 1158 73396 1164
rect 71792 56 71912 82
rect 72160 56 72280 82
rect 72988 56 73108 82
rect 70964 14 71176 42
rect 71318 0 71374 56
rect 71778 54 71912 56
rect 72146 54 72280 56
rect 72974 54 73108 56
rect 71778 0 71834 54
rect 72146 0 72202 54
rect 72974 0 73030 54
rect 73080 42 73108 54
rect 73356 42 73384 1158
rect 73448 56 73476 1838
rect 73620 1760 73672 1766
rect 73620 1702 73672 1708
rect 73632 1426 73660 1702
rect 73620 1420 73672 1426
rect 73620 1362 73672 1368
rect 74000 82 74028 4422
rect 74368 1850 74396 7142
rect 75104 6866 75132 7278
rect 75472 7002 75500 7278
rect 76656 7200 76708 7206
rect 76656 7142 76708 7148
rect 75460 6996 75512 7002
rect 75460 6938 75512 6944
rect 75092 6860 75144 6866
rect 75092 6802 75144 6808
rect 75104 5234 75132 6802
rect 75368 6792 75420 6798
rect 75368 6734 75420 6740
rect 75380 6186 75408 6734
rect 75368 6180 75420 6186
rect 75368 6122 75420 6128
rect 75460 5704 75512 5710
rect 75460 5646 75512 5652
rect 75472 5234 75500 5646
rect 75092 5228 75144 5234
rect 75092 5170 75144 5176
rect 75460 5228 75512 5234
rect 75460 5170 75512 5176
rect 75104 4690 75132 5170
rect 75460 5024 75512 5030
rect 75460 4966 75512 4972
rect 75472 4690 75500 4966
rect 75092 4684 75144 4690
rect 75092 4626 75144 4632
rect 75460 4684 75512 4690
rect 75460 4626 75512 4632
rect 75104 4214 75132 4626
rect 76564 4480 76616 4486
rect 76564 4422 76616 4428
rect 75092 4208 75144 4214
rect 75144 4156 75224 4162
rect 75092 4150 75224 4156
rect 75104 4134 75224 4150
rect 74448 3936 74500 3942
rect 74448 3878 74500 3884
rect 74460 1902 74488 3878
rect 75196 3602 75224 4134
rect 75828 4072 75880 4078
rect 75828 4014 75880 4020
rect 75184 3596 75236 3602
rect 75184 3538 75236 3544
rect 75196 1970 75224 3538
rect 75840 3534 75868 4014
rect 75368 3528 75420 3534
rect 75368 3470 75420 3476
rect 75828 3528 75880 3534
rect 75828 3470 75880 3476
rect 75380 2990 75408 3470
rect 75368 2984 75420 2990
rect 75368 2926 75420 2932
rect 75460 2440 75512 2446
rect 75460 2382 75512 2388
rect 75472 1970 75500 2382
rect 75184 1964 75236 1970
rect 75184 1906 75236 1912
rect 75460 1964 75512 1970
rect 75460 1906 75512 1912
rect 75552 1964 75604 1970
rect 76576 1952 76604 4422
rect 75552 1906 75604 1912
rect 76300 1924 76604 1952
rect 73908 56 74028 82
rect 74276 1822 74396 1850
rect 74448 1896 74500 1902
rect 74448 1838 74500 1844
rect 74276 56 74304 1822
rect 75092 1556 75144 1562
rect 75092 1498 75144 1504
rect 75104 56 75132 1498
rect 75196 1426 75224 1906
rect 75184 1420 75236 1426
rect 75184 1362 75236 1368
rect 75564 56 75592 1906
rect 76196 1760 76248 1766
rect 76196 1702 76248 1708
rect 76208 1426 76236 1702
rect 76196 1420 76248 1426
rect 76196 1362 76248 1368
rect 76024 56 76144 82
rect 73080 14 73384 42
rect 73434 0 73490 56
rect 73894 54 74028 56
rect 73894 0 73950 54
rect 74262 0 74318 56
rect 75090 0 75146 56
rect 75550 0 75606 56
rect 76010 54 76144 56
rect 76010 0 76066 54
rect 76116 42 76144 54
rect 76300 42 76328 1924
rect 76668 1850 76696 7142
rect 77220 6780 77248 7278
rect 77588 7002 77616 7278
rect 78956 7268 79008 7274
rect 78956 7210 79008 7216
rect 77576 6996 77628 7002
rect 77576 6938 77628 6944
rect 77300 6792 77352 6798
rect 77220 6752 77300 6780
rect 77300 6734 77352 6740
rect 77576 6792 77628 6798
rect 77576 6734 77628 6740
rect 77312 5166 77340 6734
rect 77588 6254 77616 6734
rect 77576 6248 77628 6254
rect 77576 6190 77628 6196
rect 77576 5568 77628 5574
rect 77576 5510 77628 5516
rect 77588 5234 77616 5510
rect 77576 5228 77628 5234
rect 77576 5170 77628 5176
rect 77300 5160 77352 5166
rect 77300 5102 77352 5108
rect 77312 4622 77340 5102
rect 77576 5024 77628 5030
rect 77576 4966 77628 4972
rect 77588 4690 77616 4966
rect 77576 4684 77628 4690
rect 77576 4626 77628 4632
rect 77300 4616 77352 4622
rect 77300 4558 77352 4564
rect 77312 4078 77340 4558
rect 78864 4480 78916 4486
rect 78864 4422 78916 4428
rect 77300 4072 77352 4078
rect 77300 4014 77352 4020
rect 78680 4072 78732 4078
rect 78680 4014 78732 4020
rect 76748 3936 76800 3942
rect 76748 3878 76800 3884
rect 76760 1970 76788 3878
rect 77312 3534 77340 4014
rect 78692 3738 78720 4014
rect 78772 3936 78824 3942
rect 78772 3878 78824 3884
rect 78680 3732 78732 3738
rect 78680 3674 78732 3680
rect 77392 3596 77444 3602
rect 77392 3538 77444 3544
rect 77300 3528 77352 3534
rect 77300 3470 77352 3476
rect 76748 1964 76800 1970
rect 76748 1906 76800 1912
rect 77312 1902 77340 3470
rect 77404 3194 77432 3538
rect 77576 3528 77628 3534
rect 77576 3470 77628 3476
rect 77392 3188 77444 3194
rect 77392 3130 77444 3136
rect 77588 2990 77616 3470
rect 77576 2984 77628 2990
rect 77576 2926 77628 2932
rect 77576 2304 77628 2310
rect 77576 2246 77628 2252
rect 77588 1970 77616 2246
rect 78784 2106 78812 3878
rect 77668 2100 77720 2106
rect 77668 2042 77720 2048
rect 78772 2100 78824 2106
rect 78772 2042 78824 2048
rect 77576 1964 77628 1970
rect 77576 1906 77628 1912
rect 76392 1822 76696 1850
rect 77300 1896 77352 1902
rect 77300 1838 77352 1844
rect 76392 56 76420 1822
rect 77208 1556 77260 1562
rect 77208 1498 77260 1504
rect 77220 56 77248 1498
rect 77312 1426 77340 1838
rect 77300 1420 77352 1426
rect 77300 1362 77352 1368
rect 77680 56 77708 2042
rect 78876 1970 78904 4422
rect 78220 1964 78272 1970
rect 78140 1924 78220 1952
rect 78140 56 78168 1924
rect 78220 1906 78272 1912
rect 78864 1964 78916 1970
rect 78864 1906 78916 1912
rect 78968 1902 78996 7210
rect 79336 6866 79364 7278
rect 79704 7002 79732 7278
rect 81348 7268 81400 7274
rect 81348 7210 81400 7216
rect 80816 7100 81112 7120
rect 80872 7098 80896 7100
rect 80952 7098 80976 7100
rect 81032 7098 81056 7100
rect 80894 7046 80896 7098
rect 80958 7046 80970 7098
rect 81032 7046 81034 7098
rect 80872 7044 80896 7046
rect 80952 7044 80976 7046
rect 81032 7044 81056 7046
rect 80816 7024 81112 7044
rect 79692 6996 79744 7002
rect 79692 6938 79744 6944
rect 79324 6860 79376 6866
rect 79324 6802 79376 6808
rect 79336 5234 79364 6802
rect 79692 6792 79744 6798
rect 79692 6734 79744 6740
rect 79704 6254 79732 6734
rect 79692 6248 79744 6254
rect 79692 6190 79744 6196
rect 80816 6012 81112 6032
rect 80872 6010 80896 6012
rect 80952 6010 80976 6012
rect 81032 6010 81056 6012
rect 80894 5958 80896 6010
rect 80958 5958 80970 6010
rect 81032 5958 81034 6010
rect 80872 5956 80896 5958
rect 80952 5956 80976 5958
rect 81032 5956 81056 5958
rect 80816 5936 81112 5956
rect 79600 5840 79652 5846
rect 79600 5782 79652 5788
rect 79612 5234 79640 5782
rect 79324 5228 79376 5234
rect 79324 5170 79376 5176
rect 79600 5228 79652 5234
rect 79600 5170 79652 5176
rect 79336 4690 79364 5170
rect 79692 5024 79744 5030
rect 79692 4966 79744 4972
rect 79704 4690 79732 4966
rect 80816 4924 81112 4944
rect 80872 4922 80896 4924
rect 80952 4922 80976 4924
rect 81032 4922 81056 4924
rect 80894 4870 80896 4922
rect 80958 4870 80970 4922
rect 81032 4870 81034 4922
rect 80872 4868 80896 4870
rect 80952 4868 80976 4870
rect 81032 4868 81056 4870
rect 80816 4848 81112 4868
rect 79324 4684 79376 4690
rect 79324 4626 79376 4632
rect 79692 4684 79744 4690
rect 79692 4626 79744 4632
rect 79336 4146 79364 4626
rect 81164 4480 81216 4486
rect 81164 4422 81216 4428
rect 79324 4140 79376 4146
rect 79324 4082 79376 4088
rect 79336 4026 79364 4082
rect 80704 4072 80756 4078
rect 79336 3998 79456 4026
rect 80704 4014 80756 4020
rect 79428 3602 79456 3998
rect 80716 3738 80744 4014
rect 80816 3836 81112 3856
rect 80872 3834 80896 3836
rect 80952 3834 80976 3836
rect 81032 3834 81056 3836
rect 80894 3782 80896 3834
rect 80958 3782 80970 3834
rect 81032 3782 81034 3834
rect 80872 3780 80896 3782
rect 80952 3780 80976 3782
rect 81032 3780 81056 3782
rect 80816 3760 81112 3780
rect 80704 3732 80756 3738
rect 80704 3674 80756 3680
rect 79416 3596 79468 3602
rect 79416 3538 79468 3544
rect 79428 1970 79456 3538
rect 79692 3528 79744 3534
rect 79692 3470 79744 3476
rect 79704 2990 79732 3470
rect 79692 2984 79744 2990
rect 79692 2926 79744 2932
rect 80816 2748 81112 2768
rect 80872 2746 80896 2748
rect 80952 2746 80976 2748
rect 81032 2746 81056 2748
rect 80894 2694 80896 2746
rect 80958 2694 80970 2746
rect 81032 2694 81034 2746
rect 80872 2692 80896 2694
rect 80952 2692 80976 2694
rect 81032 2692 81056 2694
rect 80816 2672 81112 2692
rect 79600 2576 79652 2582
rect 79600 2518 79652 2524
rect 79612 1970 79640 2518
rect 81176 2106 81204 4422
rect 81256 4004 81308 4010
rect 81256 3946 81308 3952
rect 80336 2100 80388 2106
rect 80256 2060 80336 2088
rect 79416 1964 79468 1970
rect 79416 1906 79468 1912
rect 79600 1964 79652 1970
rect 79600 1906 79652 1912
rect 79784 1964 79836 1970
rect 79784 1906 79836 1912
rect 78496 1896 78548 1902
rect 78496 1838 78548 1844
rect 78956 1896 79008 1902
rect 78956 1838 79008 1844
rect 78508 56 78536 1838
rect 78864 1760 78916 1766
rect 78864 1702 78916 1708
rect 78876 1426 78904 1702
rect 79428 1426 79456 1906
rect 78864 1420 78916 1426
rect 78864 1362 78916 1368
rect 79416 1420 79468 1426
rect 79416 1362 79468 1368
rect 79324 1216 79376 1222
rect 79324 1158 79376 1164
rect 79336 56 79364 1158
rect 79796 56 79824 1906
rect 80256 56 80284 2060
rect 80336 2042 80388 2048
rect 81164 2100 81216 2106
rect 81164 2042 81216 2048
rect 80612 2032 80664 2038
rect 80612 1974 80664 1980
rect 80624 56 80652 1974
rect 81268 1970 81296 3946
rect 81360 2038 81388 7210
rect 81452 6866 81480 7278
rect 81820 7002 81848 7278
rect 82820 7200 82872 7206
rect 82820 7142 82872 7148
rect 81808 6996 81860 7002
rect 81808 6938 81860 6944
rect 81440 6860 81492 6866
rect 81440 6802 81492 6808
rect 81452 5234 81480 6802
rect 81808 6792 81860 6798
rect 81808 6734 81860 6740
rect 81820 6254 81848 6734
rect 81808 6248 81860 6254
rect 81808 6190 81860 6196
rect 81808 5772 81860 5778
rect 81808 5714 81860 5720
rect 81820 5234 81848 5714
rect 81440 5228 81492 5234
rect 81440 5170 81492 5176
rect 81808 5228 81860 5234
rect 81808 5170 81860 5176
rect 81452 4690 81480 5170
rect 81808 5024 81860 5030
rect 81808 4966 81860 4972
rect 81820 4690 81848 4966
rect 81440 4684 81492 4690
rect 81440 4626 81492 4632
rect 81808 4684 81860 4690
rect 81808 4626 81860 4632
rect 81452 4128 81480 4626
rect 82636 4480 82688 4486
rect 82636 4422 82688 4428
rect 81532 4140 81584 4146
rect 81452 4100 81532 4128
rect 81532 4082 81584 4088
rect 81544 3602 81572 4082
rect 81900 3936 81952 3942
rect 81900 3878 81952 3884
rect 81532 3596 81584 3602
rect 81532 3538 81584 3544
rect 81348 2032 81400 2038
rect 81348 1974 81400 1980
rect 81544 1970 81572 3538
rect 81808 3528 81860 3534
rect 81808 3470 81860 3476
rect 81820 2990 81848 3470
rect 81808 2984 81860 2990
rect 81808 2926 81860 2932
rect 81716 2508 81768 2514
rect 81716 2450 81768 2456
rect 81728 1970 81756 2450
rect 81256 1964 81308 1970
rect 81256 1906 81308 1912
rect 81532 1964 81584 1970
rect 81532 1906 81584 1912
rect 81716 1964 81768 1970
rect 81716 1906 81768 1912
rect 81164 1828 81216 1834
rect 81164 1770 81216 1776
rect 80816 1660 81112 1680
rect 80872 1658 80896 1660
rect 80952 1658 80976 1660
rect 81032 1658 81056 1660
rect 80894 1606 80896 1658
rect 80958 1606 80970 1658
rect 81032 1606 81034 1658
rect 80872 1604 80896 1606
rect 80952 1604 80976 1606
rect 81032 1604 81056 1606
rect 80816 1584 81112 1604
rect 81176 1426 81204 1770
rect 81440 1556 81492 1562
rect 81440 1498 81492 1504
rect 81164 1420 81216 1426
rect 81164 1362 81216 1368
rect 81452 56 81480 1498
rect 81544 1426 81572 1906
rect 81532 1420 81584 1426
rect 81532 1362 81584 1368
rect 81912 56 81940 3878
rect 82648 1748 82676 4422
rect 82372 1720 82676 1748
rect 82372 56 82400 1720
rect 82832 82 82860 7142
rect 83568 6866 83596 7278
rect 83936 7002 83964 7278
rect 85120 7200 85172 7206
rect 85120 7142 85172 7148
rect 83924 6996 83976 7002
rect 83924 6938 83976 6944
rect 83556 6860 83608 6866
rect 83556 6802 83608 6808
rect 83568 5234 83596 6802
rect 83924 6792 83976 6798
rect 83924 6734 83976 6740
rect 83936 6254 83964 6734
rect 83924 6248 83976 6254
rect 83924 6190 83976 6196
rect 83924 5840 83976 5846
rect 83924 5782 83976 5788
rect 83936 5234 83964 5782
rect 83556 5228 83608 5234
rect 83556 5170 83608 5176
rect 83924 5228 83976 5234
rect 83924 5170 83976 5176
rect 83568 4690 83596 5170
rect 83924 5024 83976 5030
rect 83924 4966 83976 4972
rect 83936 4690 83964 4966
rect 83556 4684 83608 4690
rect 83556 4626 83608 4632
rect 83924 4684 83976 4690
rect 83924 4626 83976 4632
rect 83568 4214 83596 4626
rect 84660 4480 84712 4486
rect 84660 4422 84712 4428
rect 83556 4208 83608 4214
rect 83608 4156 83688 4162
rect 83556 4150 83688 4156
rect 83568 4134 83688 4150
rect 82912 4072 82964 4078
rect 82912 4014 82964 4020
rect 82924 3738 82952 4014
rect 82912 3732 82964 3738
rect 82912 3674 82964 3680
rect 83660 3602 83688 4134
rect 84016 3936 84068 3942
rect 84016 3878 84068 3884
rect 83648 3596 83700 3602
rect 83648 3538 83700 3544
rect 83660 1970 83688 3538
rect 83924 3528 83976 3534
rect 83924 3470 83976 3476
rect 83936 2922 83964 3470
rect 83924 2916 83976 2922
rect 83924 2858 83976 2864
rect 83924 2508 83976 2514
rect 83924 2450 83976 2456
rect 83936 1970 83964 2450
rect 83648 1964 83700 1970
rect 83648 1906 83700 1912
rect 83924 1964 83976 1970
rect 83924 1906 83976 1912
rect 82912 1760 82964 1766
rect 82912 1702 82964 1708
rect 82924 1426 82952 1702
rect 83660 1426 83688 1906
rect 82912 1420 82964 1426
rect 82912 1362 82964 1368
rect 83648 1420 83700 1426
rect 83648 1362 83700 1368
rect 83832 1216 83884 1222
rect 83832 1158 83884 1164
rect 82740 56 82860 82
rect 83568 56 83688 82
rect 76116 14 76328 42
rect 76378 0 76434 56
rect 77206 0 77262 56
rect 77666 0 77722 56
rect 78126 0 78182 56
rect 78494 0 78550 56
rect 79322 0 79378 56
rect 79782 0 79838 56
rect 80242 0 80298 56
rect 80610 0 80666 56
rect 81438 0 81494 56
rect 81898 0 81954 56
rect 82358 0 82414 56
rect 82726 54 82860 56
rect 83554 54 83688 56
rect 82726 0 82782 54
rect 83554 0 83610 54
rect 83660 42 83688 54
rect 83844 42 83872 1158
rect 84028 56 84056 3878
rect 84672 1850 84700 4422
rect 85028 4072 85080 4078
rect 85028 4014 85080 4020
rect 85040 3738 85068 4014
rect 85028 3732 85080 3738
rect 85028 3674 85080 3680
rect 84488 1822 84700 1850
rect 84488 56 84516 1822
rect 85028 1760 85080 1766
rect 85028 1702 85080 1708
rect 85040 1426 85068 1702
rect 85028 1420 85080 1426
rect 85028 1362 85080 1368
rect 84856 56 84976 82
rect 83660 14 83872 42
rect 84014 0 84070 56
rect 84474 0 84530 56
rect 84842 54 84976 56
rect 84842 0 84898 54
rect 84948 42 84976 54
rect 85132 42 85160 7142
rect 85684 6866 85712 7278
rect 86052 7002 86080 7278
rect 87144 7200 87196 7206
rect 87144 7142 87196 7148
rect 86040 6996 86092 7002
rect 86040 6938 86092 6944
rect 85672 6860 85724 6866
rect 85672 6802 85724 6808
rect 85684 5234 85712 6802
rect 85948 6792 86000 6798
rect 85948 6734 86000 6740
rect 85960 6186 85988 6734
rect 85948 6180 86000 6186
rect 85948 6122 86000 6128
rect 86040 5772 86092 5778
rect 86040 5714 86092 5720
rect 86052 5234 86080 5714
rect 85672 5228 85724 5234
rect 85672 5170 85724 5176
rect 86040 5228 86092 5234
rect 86040 5170 86092 5176
rect 85684 4690 85712 5170
rect 86040 5024 86092 5030
rect 86040 4966 86092 4972
rect 86052 4690 86080 4966
rect 85672 4684 85724 4690
rect 86040 4684 86092 4690
rect 85724 4644 85804 4672
rect 85672 4626 85724 4632
rect 85776 4146 85804 4644
rect 86040 4626 86092 4632
rect 86868 4480 86920 4486
rect 86868 4422 86920 4428
rect 85764 4140 85816 4146
rect 85764 4082 85816 4088
rect 85776 3602 85804 4082
rect 86132 4072 86184 4078
rect 86132 4014 86184 4020
rect 85764 3596 85816 3602
rect 85764 3538 85816 3544
rect 85776 1970 85804 3538
rect 86144 3534 86172 4014
rect 86408 3936 86460 3942
rect 86408 3878 86460 3884
rect 85948 3528 86000 3534
rect 85948 3470 86000 3476
rect 86132 3528 86184 3534
rect 86132 3470 86184 3476
rect 85960 2990 85988 3470
rect 85948 2984 86000 2990
rect 85948 2926 86000 2932
rect 85948 2372 86000 2378
rect 85948 2314 86000 2320
rect 85960 1970 85988 2314
rect 85764 1964 85816 1970
rect 85764 1906 85816 1912
rect 85948 1964 86000 1970
rect 85948 1906 86000 1912
rect 85776 1426 85804 1906
rect 85764 1420 85816 1426
rect 85764 1362 85816 1368
rect 86040 1216 86092 1222
rect 86040 1158 86092 1164
rect 85684 56 85804 82
rect 84948 14 85160 42
rect 85670 54 85804 56
rect 85670 0 85726 54
rect 85776 42 85804 54
rect 86052 42 86080 1158
rect 86144 56 86264 82
rect 85776 14 86080 42
rect 86130 54 86264 56
rect 86130 0 86186 54
rect 86236 42 86264 54
rect 86420 42 86448 3878
rect 86500 1760 86552 1766
rect 86500 1702 86552 1708
rect 86512 1426 86540 1702
rect 86880 1578 86908 4422
rect 87052 3596 87104 3602
rect 87052 3538 87104 3544
rect 87064 3194 87092 3538
rect 87052 3188 87104 3194
rect 87052 3130 87104 3136
rect 86788 1550 86908 1578
rect 86500 1420 86552 1426
rect 86500 1362 86552 1368
rect 86604 56 86724 82
rect 86236 14 86448 42
rect 86590 54 86724 56
rect 86590 0 86646 54
rect 86696 42 86724 54
rect 86788 42 86816 1550
rect 86972 56 87092 82
rect 86696 14 86816 42
rect 86958 54 87092 56
rect 86958 0 87014 54
rect 87064 42 87092 54
rect 87156 42 87184 7142
rect 87800 6866 87828 7278
rect 88168 7002 88196 7278
rect 89168 7200 89220 7206
rect 89168 7142 89220 7148
rect 88156 6996 88208 7002
rect 88156 6938 88208 6944
rect 87788 6860 87840 6866
rect 87788 6802 87840 6808
rect 87800 5234 87828 6802
rect 88156 6792 88208 6798
rect 88156 6734 88208 6740
rect 88168 6254 88196 6734
rect 88156 6248 88208 6254
rect 88156 6190 88208 6196
rect 88156 5568 88208 5574
rect 88156 5510 88208 5516
rect 88168 5234 88196 5510
rect 87788 5228 87840 5234
rect 87788 5170 87840 5176
rect 88156 5228 88208 5234
rect 88156 5170 88208 5176
rect 87800 4690 87828 5170
rect 88156 5024 88208 5030
rect 88156 4966 88208 4972
rect 88168 4690 88196 4966
rect 87788 4684 87840 4690
rect 87788 4626 87840 4632
rect 88156 4684 88208 4690
rect 88156 4626 88208 4632
rect 87800 4214 87828 4626
rect 87788 4208 87840 4214
rect 87840 4168 87920 4196
rect 87788 4150 87840 4156
rect 87892 3602 87920 4168
rect 88524 4072 88576 4078
rect 88524 4014 88576 4020
rect 87880 3596 87932 3602
rect 87880 3538 87932 3544
rect 87892 1970 87920 3538
rect 88536 3534 88564 4014
rect 88156 3528 88208 3534
rect 88156 3470 88208 3476
rect 88524 3528 88576 3534
rect 88524 3470 88576 3476
rect 88168 2990 88196 3470
rect 88156 2984 88208 2990
rect 88156 2926 88208 2932
rect 88156 2440 88208 2446
rect 88156 2382 88208 2388
rect 88168 1970 88196 2382
rect 87880 1964 87932 1970
rect 87880 1906 87932 1912
rect 88156 1964 88208 1970
rect 88800 1964 88852 1970
rect 88156 1906 88208 1912
rect 88720 1924 88800 1952
rect 87892 1426 87920 1906
rect 88248 1896 88300 1902
rect 88248 1838 88300 1844
rect 87880 1420 87932 1426
rect 87880 1362 87932 1368
rect 88064 1216 88116 1222
rect 88064 1158 88116 1164
rect 87800 56 87920 82
rect 87064 14 87184 42
rect 87786 54 87920 56
rect 87786 0 87842 54
rect 87892 42 87920 54
rect 88076 42 88104 1158
rect 88260 56 88288 1838
rect 88432 1760 88484 1766
rect 88432 1702 88484 1708
rect 88444 1426 88472 1702
rect 88432 1420 88484 1426
rect 88432 1362 88484 1368
rect 88720 56 88748 1924
rect 88800 1906 88852 1912
rect 89180 82 89208 7142
rect 89916 6866 89944 7278
rect 90284 7002 90312 7278
rect 91468 7200 91520 7206
rect 91468 7142 91520 7148
rect 90272 6996 90324 7002
rect 90272 6938 90324 6944
rect 89904 6860 89956 6866
rect 89904 6802 89956 6808
rect 89916 5234 89944 6802
rect 90272 6792 90324 6798
rect 90272 6734 90324 6740
rect 90284 6254 90312 6734
rect 90272 6248 90324 6254
rect 90272 6190 90324 6196
rect 90272 5840 90324 5846
rect 90272 5782 90324 5788
rect 90284 5234 90312 5782
rect 89904 5228 89956 5234
rect 89904 5170 89956 5176
rect 90272 5228 90324 5234
rect 90272 5170 90324 5176
rect 89916 4690 89944 5170
rect 90272 5024 90324 5030
rect 90272 4966 90324 4972
rect 90284 4690 90312 4966
rect 89904 4684 89956 4690
rect 89904 4626 89956 4632
rect 90272 4684 90324 4690
rect 90272 4626 90324 4632
rect 89260 4480 89312 4486
rect 89260 4422 89312 4428
rect 89272 1970 89300 4422
rect 89916 4060 89944 4626
rect 91284 4480 91336 4486
rect 91284 4422 91336 4428
rect 89996 4072 90048 4078
rect 89916 4032 89996 4060
rect 89996 4014 90048 4020
rect 90640 4072 90692 4078
rect 90640 4014 90692 4020
rect 89444 3936 89496 3942
rect 89444 3878 89496 3884
rect 89260 1964 89312 1970
rect 89260 1906 89312 1912
rect 89456 1902 89484 3878
rect 90008 3602 90036 4014
rect 89996 3596 90048 3602
rect 89996 3538 90048 3544
rect 90008 1970 90036 3538
rect 90652 3534 90680 4014
rect 90272 3528 90324 3534
rect 90272 3470 90324 3476
rect 90640 3528 90692 3534
rect 90640 3470 90692 3476
rect 90284 2990 90312 3470
rect 90272 2984 90324 2990
rect 90272 2926 90324 2932
rect 90272 2576 90324 2582
rect 90272 2518 90324 2524
rect 90284 1970 90312 2518
rect 89996 1964 90048 1970
rect 89996 1906 90048 1912
rect 90272 1964 90324 1970
rect 90272 1906 90324 1912
rect 90364 1964 90416 1970
rect 90364 1906 90416 1912
rect 89444 1896 89496 1902
rect 89444 1838 89496 1844
rect 90008 1426 90036 1906
rect 89996 1420 90048 1426
rect 89996 1362 90048 1368
rect 90272 1216 90324 1222
rect 90272 1158 90324 1164
rect 89088 56 89208 82
rect 89916 56 90036 82
rect 87892 14 88104 42
rect 88246 0 88302 56
rect 88706 0 88762 56
rect 89074 54 89208 56
rect 89902 54 90036 56
rect 89074 0 89130 54
rect 89902 0 89958 54
rect 90008 42 90036 54
rect 90284 42 90312 1158
rect 90376 56 90404 1906
rect 90732 1760 90784 1766
rect 90732 1702 90784 1708
rect 90744 1426 90772 1702
rect 91296 1578 91324 4422
rect 91376 3936 91428 3942
rect 91376 3878 91428 3884
rect 91388 1970 91416 3878
rect 91376 1964 91428 1970
rect 91376 1906 91428 1912
rect 91480 1578 91508 7142
rect 92032 6866 92060 7278
rect 92400 7002 92428 7278
rect 94148 7262 94268 7278
rect 93584 7200 93636 7206
rect 93584 7142 93636 7148
rect 92388 6996 92440 7002
rect 92388 6938 92440 6944
rect 92020 6860 92072 6866
rect 92020 6802 92072 6808
rect 92032 5234 92060 6802
rect 92388 6792 92440 6798
rect 92388 6734 92440 6740
rect 92400 6254 92428 6734
rect 92388 6248 92440 6254
rect 92388 6190 92440 6196
rect 92388 5704 92440 5710
rect 92388 5646 92440 5652
rect 92400 5234 92428 5646
rect 92020 5228 92072 5234
rect 92020 5170 92072 5176
rect 92388 5228 92440 5234
rect 92388 5170 92440 5176
rect 92032 4690 92060 5170
rect 92388 5024 92440 5030
rect 92388 4966 92440 4972
rect 92400 4690 92428 4966
rect 92020 4684 92072 4690
rect 92020 4626 92072 4632
rect 92388 4684 92440 4690
rect 92388 4626 92440 4632
rect 92032 4146 92060 4626
rect 92020 4140 92072 4146
rect 92020 4082 92072 4088
rect 92032 4026 92060 4082
rect 93124 4072 93176 4078
rect 92032 3998 92152 4026
rect 93124 4014 93176 4020
rect 92124 3602 92152 3998
rect 92112 3596 92164 3602
rect 92112 3538 92164 3544
rect 92124 1970 92152 3538
rect 93136 3534 93164 4014
rect 93492 3936 93544 3942
rect 93492 3878 93544 3884
rect 92388 3528 92440 3534
rect 92388 3470 92440 3476
rect 93124 3528 93176 3534
rect 93124 3470 93176 3476
rect 92400 2990 92428 3470
rect 92388 2984 92440 2990
rect 92388 2926 92440 2932
rect 92388 2440 92440 2446
rect 92388 2382 92440 2388
rect 92400 1970 92428 2382
rect 93504 1970 93532 3878
rect 92112 1964 92164 1970
rect 92112 1906 92164 1912
rect 92388 1964 92440 1970
rect 92388 1906 92440 1912
rect 92480 1964 92532 1970
rect 92480 1906 92532 1912
rect 93492 1964 93544 1970
rect 93492 1906 93544 1912
rect 91112 1550 91324 1578
rect 91388 1550 91508 1578
rect 92020 1556 92072 1562
rect 90732 1420 90784 1426
rect 90732 1362 90784 1368
rect 90836 56 90956 82
rect 90008 14 90312 42
rect 90362 0 90418 56
rect 90822 54 90956 56
rect 90822 0 90878 54
rect 90928 42 90956 54
rect 91112 42 91140 1550
rect 91388 1442 91416 1550
rect 92020 1498 92072 1504
rect 91204 1414 91416 1442
rect 91204 56 91232 1414
rect 92032 56 92060 1498
rect 92124 1426 92152 1906
rect 92112 1420 92164 1426
rect 92112 1362 92164 1368
rect 92492 56 92520 1906
rect 93032 1896 93084 1902
rect 92952 1844 93032 1850
rect 93596 1850 93624 7142
rect 94240 6866 94268 7262
rect 94516 7002 94544 7278
rect 95884 7268 95936 7274
rect 95884 7210 95936 7216
rect 94504 6996 94556 7002
rect 94504 6938 94556 6944
rect 94228 6860 94280 6866
rect 94228 6802 94280 6808
rect 94240 5234 94268 6802
rect 94504 6792 94556 6798
rect 94504 6734 94556 6740
rect 94516 6254 94544 6734
rect 94504 6248 94556 6254
rect 94504 6190 94556 6196
rect 94412 5840 94464 5846
rect 94412 5782 94464 5788
rect 94424 5234 94452 5782
rect 94228 5228 94280 5234
rect 94228 5170 94280 5176
rect 94412 5228 94464 5234
rect 94412 5170 94464 5176
rect 94240 4690 94268 5170
rect 94504 5024 94556 5030
rect 94504 4966 94556 4972
rect 94516 4690 94544 4966
rect 94228 4684 94280 4690
rect 94228 4626 94280 4632
rect 94504 4684 94556 4690
rect 94504 4626 94556 4632
rect 93676 4480 93728 4486
rect 93676 4422 93728 4428
rect 93688 1902 93716 4422
rect 94240 4146 94268 4626
rect 95792 4480 95844 4486
rect 95792 4422 95844 4428
rect 94228 4140 94280 4146
rect 94228 4082 94280 4088
rect 94240 3602 94268 4082
rect 95608 4072 95660 4078
rect 95608 4014 95660 4020
rect 95620 3738 95648 4014
rect 95700 3936 95752 3942
rect 95700 3878 95752 3884
rect 95608 3732 95660 3738
rect 95608 3674 95660 3680
rect 94228 3596 94280 3602
rect 94228 3538 94280 3544
rect 94240 1970 94268 3538
rect 94504 3528 94556 3534
rect 94504 3470 94556 3476
rect 94516 2990 94544 3470
rect 94504 2984 94556 2990
rect 94504 2926 94556 2932
rect 94412 2576 94464 2582
rect 94412 2518 94464 2524
rect 94424 1970 94452 2518
rect 94228 1964 94280 1970
rect 94228 1906 94280 1912
rect 94412 1964 94464 1970
rect 95148 1964 95200 1970
rect 94412 1906 94464 1912
rect 95068 1924 95148 1952
rect 92952 1838 93084 1844
rect 92952 1822 93072 1838
rect 93320 1822 93624 1850
rect 93676 1896 93728 1902
rect 93676 1838 93728 1844
rect 92756 1760 92808 1766
rect 92756 1702 92808 1708
rect 92768 1426 92796 1702
rect 92756 1420 92808 1426
rect 92756 1362 92808 1368
rect 92952 56 92980 1822
rect 93320 56 93348 1822
rect 94136 1556 94188 1562
rect 94136 1498 94188 1504
rect 94148 56 94176 1498
rect 94240 1426 94268 1906
rect 94596 1896 94648 1902
rect 94596 1838 94648 1844
rect 94228 1420 94280 1426
rect 94228 1362 94280 1368
rect 94608 56 94636 1838
rect 95068 56 95096 1924
rect 95148 1906 95200 1912
rect 95712 1902 95740 3878
rect 95804 1970 95832 4422
rect 95792 1964 95844 1970
rect 95792 1906 95844 1912
rect 95700 1896 95752 1902
rect 95700 1838 95752 1844
rect 95896 1834 95924 7210
rect 96080 6866 96108 7278
rect 96632 7002 96660 7278
rect 98092 7268 98144 7274
rect 98092 7210 98144 7216
rect 96620 6996 96672 7002
rect 96620 6938 96672 6944
rect 96068 6860 96120 6866
rect 96068 6802 96120 6808
rect 96080 5234 96108 6802
rect 96620 6792 96672 6798
rect 96620 6734 96672 6740
rect 96176 6556 96472 6576
rect 96232 6554 96256 6556
rect 96312 6554 96336 6556
rect 96392 6554 96416 6556
rect 96254 6502 96256 6554
rect 96318 6502 96330 6554
rect 96392 6502 96394 6554
rect 96232 6500 96256 6502
rect 96312 6500 96336 6502
rect 96392 6500 96416 6502
rect 96176 6480 96472 6500
rect 96632 6254 96660 6734
rect 96620 6248 96672 6254
rect 96620 6190 96672 6196
rect 96436 5840 96488 5846
rect 96488 5788 96568 5794
rect 96436 5782 96568 5788
rect 96448 5766 96568 5782
rect 96176 5468 96472 5488
rect 96232 5466 96256 5468
rect 96312 5466 96336 5468
rect 96392 5466 96416 5468
rect 96254 5414 96256 5466
rect 96318 5414 96330 5466
rect 96392 5414 96394 5466
rect 96232 5412 96256 5414
rect 96312 5412 96336 5414
rect 96392 5412 96416 5414
rect 96176 5392 96472 5412
rect 96540 5234 96568 5766
rect 96068 5228 96120 5234
rect 96068 5170 96120 5176
rect 96528 5228 96580 5234
rect 96528 5170 96580 5176
rect 96080 4690 96108 5170
rect 96620 5024 96672 5030
rect 96620 4966 96672 4972
rect 96632 4690 96660 4966
rect 96068 4684 96120 4690
rect 96068 4626 96120 4632
rect 96620 4684 96672 4690
rect 96620 4626 96672 4632
rect 96080 4146 96108 4626
rect 98000 4480 98052 4486
rect 98000 4422 98052 4428
rect 96176 4380 96472 4400
rect 96232 4378 96256 4380
rect 96312 4378 96336 4380
rect 96392 4378 96416 4380
rect 96254 4326 96256 4378
rect 96318 4326 96330 4378
rect 96392 4326 96394 4378
rect 96232 4324 96256 4326
rect 96312 4324 96336 4326
rect 96392 4324 96416 4326
rect 96176 4304 96472 4324
rect 96068 4140 96120 4146
rect 96068 4082 96120 4088
rect 96080 3602 96108 4082
rect 97264 4072 97316 4078
rect 97264 4014 97316 4020
rect 96068 3596 96120 3602
rect 96068 3538 96120 3544
rect 96080 1970 96108 3538
rect 97276 3534 97304 4014
rect 97908 3936 97960 3942
rect 97908 3878 97960 3884
rect 96620 3528 96672 3534
rect 96620 3470 96672 3476
rect 97264 3528 97316 3534
rect 97264 3470 97316 3476
rect 96176 3292 96472 3312
rect 96232 3290 96256 3292
rect 96312 3290 96336 3292
rect 96392 3290 96416 3292
rect 96254 3238 96256 3290
rect 96318 3238 96330 3290
rect 96392 3238 96394 3290
rect 96232 3236 96256 3238
rect 96312 3236 96336 3238
rect 96392 3236 96416 3238
rect 96176 3216 96472 3236
rect 96632 2990 96660 3470
rect 96620 2984 96672 2990
rect 96620 2926 96672 2932
rect 96620 2576 96672 2582
rect 96620 2518 96672 2524
rect 96176 2204 96472 2224
rect 96232 2202 96256 2204
rect 96312 2202 96336 2204
rect 96392 2202 96416 2204
rect 96254 2150 96256 2202
rect 96318 2150 96330 2202
rect 96392 2150 96394 2202
rect 96232 2148 96256 2150
rect 96312 2148 96336 2150
rect 96392 2148 96416 2150
rect 96176 2128 96472 2148
rect 96632 1970 96660 2518
rect 97920 2106 97948 3878
rect 96712 2100 96764 2106
rect 96712 2042 96764 2048
rect 97908 2100 97960 2106
rect 97908 2042 97960 2048
rect 96068 1964 96120 1970
rect 96068 1906 96120 1912
rect 96620 1964 96672 1970
rect 96620 1906 96672 1912
rect 95424 1828 95476 1834
rect 95424 1770 95476 1776
rect 95884 1828 95936 1834
rect 95884 1770 95936 1776
rect 95436 56 95464 1770
rect 95792 1760 95844 1766
rect 95792 1702 95844 1708
rect 95804 1426 95832 1702
rect 96080 1426 96108 1906
rect 95792 1420 95844 1426
rect 95792 1362 95844 1368
rect 96068 1420 96120 1426
rect 96068 1362 96120 1368
rect 96528 1216 96580 1222
rect 96528 1158 96580 1164
rect 96176 1116 96472 1136
rect 96232 1114 96256 1116
rect 96312 1114 96336 1116
rect 96392 1114 96416 1116
rect 96254 1062 96256 1114
rect 96318 1062 96330 1114
rect 96392 1062 96394 1114
rect 96232 1060 96256 1062
rect 96312 1060 96336 1062
rect 96392 1060 96416 1062
rect 96176 1040 96472 1060
rect 96540 762 96568 1158
rect 96264 734 96568 762
rect 96264 56 96292 734
rect 96724 56 96752 2042
rect 98012 1970 98040 4422
rect 97264 1964 97316 1970
rect 97184 1924 97264 1952
rect 97184 56 97212 1924
rect 97264 1906 97316 1912
rect 98000 1964 98052 1970
rect 98000 1906 98052 1912
rect 98104 1902 98132 7210
rect 98380 6866 98408 7278
rect 98748 7002 98776 7278
rect 99748 7200 99800 7206
rect 99748 7142 99800 7148
rect 98736 6996 98788 7002
rect 98736 6938 98788 6944
rect 98368 6860 98420 6866
rect 98368 6802 98420 6808
rect 98380 5234 98408 6802
rect 98736 6792 98788 6798
rect 98736 6734 98788 6740
rect 98748 6254 98776 6734
rect 98736 6248 98788 6254
rect 98736 6190 98788 6196
rect 98644 5772 98696 5778
rect 98644 5714 98696 5720
rect 98656 5234 98684 5714
rect 98368 5228 98420 5234
rect 98368 5170 98420 5176
rect 98644 5228 98696 5234
rect 98644 5170 98696 5176
rect 98380 4690 98408 5170
rect 98736 5024 98788 5030
rect 98736 4966 98788 4972
rect 98748 4690 98776 4966
rect 98368 4684 98420 4690
rect 98368 4626 98420 4632
rect 98736 4684 98788 4690
rect 98736 4626 98788 4632
rect 98380 4146 98408 4626
rect 99380 4480 99432 4486
rect 99380 4422 99432 4428
rect 98368 4140 98420 4146
rect 98420 4100 98500 4128
rect 98368 4082 98420 4088
rect 98472 3602 98500 4100
rect 98828 3936 98880 3942
rect 98828 3878 98880 3884
rect 98460 3596 98512 3602
rect 98460 3538 98512 3544
rect 98472 1970 98500 3538
rect 98736 3528 98788 3534
rect 98736 3470 98788 3476
rect 98748 2990 98776 3470
rect 98736 2984 98788 2990
rect 98736 2926 98788 2932
rect 98736 2576 98788 2582
rect 98736 2518 98788 2524
rect 98748 1970 98776 2518
rect 98460 1964 98512 1970
rect 98460 1906 98512 1912
rect 98736 1964 98788 1970
rect 98736 1906 98788 1912
rect 97540 1896 97592 1902
rect 97540 1838 97592 1844
rect 98092 1896 98144 1902
rect 98092 1838 98144 1844
rect 97552 56 97580 1838
rect 97908 1760 97960 1766
rect 97908 1702 97960 1708
rect 97920 1426 97948 1702
rect 98368 1556 98420 1562
rect 98368 1498 98420 1504
rect 97908 1420 97960 1426
rect 97908 1362 97960 1368
rect 98380 56 98408 1498
rect 98472 1426 98500 1906
rect 98460 1420 98512 1426
rect 98460 1362 98512 1368
rect 98840 56 98868 3878
rect 99392 1850 99420 4422
rect 99300 1822 99420 1850
rect 99300 56 99328 1822
rect 99760 82 99788 7142
rect 100496 6866 100524 7278
rect 100864 7002 100892 7278
rect 101864 7200 101916 7206
rect 101864 7142 101916 7148
rect 100852 6996 100904 7002
rect 100852 6938 100904 6944
rect 100484 6860 100536 6866
rect 100484 6802 100536 6808
rect 100496 5234 100524 6802
rect 100852 6792 100904 6798
rect 100852 6734 100904 6740
rect 100864 6254 100892 6734
rect 100852 6248 100904 6254
rect 100852 6190 100904 6196
rect 100760 5772 100812 5778
rect 100760 5714 100812 5720
rect 100772 5234 100800 5714
rect 100484 5228 100536 5234
rect 100484 5170 100536 5176
rect 100760 5228 100812 5234
rect 100760 5170 100812 5176
rect 100496 4690 100524 5170
rect 100852 5024 100904 5030
rect 100852 4966 100904 4972
rect 100864 4690 100892 4966
rect 100484 4684 100536 4690
rect 100484 4626 100536 4632
rect 100852 4684 100904 4690
rect 100852 4626 100904 4632
rect 100496 4146 100524 4626
rect 101588 4480 101640 4486
rect 101588 4422 101640 4428
rect 100484 4140 100536 4146
rect 100536 4100 100616 4128
rect 100484 4082 100536 4088
rect 99840 4072 99892 4078
rect 99840 4014 99892 4020
rect 99852 3738 99880 4014
rect 99840 3732 99892 3738
rect 99840 3674 99892 3680
rect 100588 3602 100616 4100
rect 100944 3936 100996 3942
rect 100944 3878 100996 3884
rect 100576 3596 100628 3602
rect 100576 3538 100628 3544
rect 100588 1970 100616 3538
rect 100852 3528 100904 3534
rect 100852 3470 100904 3476
rect 100864 2990 100892 3470
rect 100852 2984 100904 2990
rect 100852 2926 100904 2932
rect 100852 2508 100904 2514
rect 100852 2450 100904 2456
rect 100864 1970 100892 2450
rect 100576 1964 100628 1970
rect 100576 1906 100628 1912
rect 100852 1964 100904 1970
rect 100852 1906 100904 1912
rect 99840 1760 99892 1766
rect 99840 1702 99892 1708
rect 99852 1426 99880 1702
rect 100588 1426 100616 1906
rect 99840 1420 99892 1426
rect 99840 1362 99892 1368
rect 100576 1420 100628 1426
rect 100576 1362 100628 1368
rect 100760 1216 100812 1222
rect 100760 1158 100812 1164
rect 99668 56 99788 82
rect 100496 56 100616 82
rect 90928 14 91140 42
rect 91190 0 91246 56
rect 92018 0 92074 56
rect 92478 0 92534 56
rect 92938 0 92994 56
rect 93306 0 93362 56
rect 94134 0 94190 56
rect 94594 0 94650 56
rect 95054 0 95110 56
rect 95422 0 95478 56
rect 96250 0 96306 56
rect 96710 0 96766 56
rect 97170 0 97226 56
rect 97538 0 97594 56
rect 98366 0 98422 56
rect 98826 0 98882 56
rect 99286 0 99342 56
rect 99654 54 99788 56
rect 100482 54 100616 56
rect 99654 0 99710 54
rect 100482 0 100538 54
rect 100588 42 100616 54
rect 100772 42 100800 1158
rect 100956 56 100984 3878
rect 101600 2122 101628 4422
rect 101416 2094 101628 2122
rect 101416 56 101444 2094
rect 101876 82 101904 7142
rect 102704 6866 102732 7278
rect 102980 7002 103008 7278
rect 103888 7200 103940 7206
rect 103888 7142 103940 7148
rect 102968 6996 103020 7002
rect 102968 6938 103020 6944
rect 102692 6860 102744 6866
rect 102692 6802 102744 6808
rect 102704 5234 102732 6802
rect 102968 6792 103020 6798
rect 102968 6734 103020 6740
rect 102980 6254 103008 6734
rect 102968 6248 103020 6254
rect 102968 6190 103020 6196
rect 102968 5772 103020 5778
rect 102968 5714 103020 5720
rect 102980 5234 103008 5714
rect 102692 5228 102744 5234
rect 102692 5170 102744 5176
rect 102968 5228 103020 5234
rect 102968 5170 103020 5176
rect 102704 4690 102732 5170
rect 102968 5024 103020 5030
rect 102968 4966 103020 4972
rect 102980 4690 103008 4966
rect 102692 4684 102744 4690
rect 102692 4626 102744 4632
rect 102968 4684 103020 4690
rect 102968 4626 103020 4632
rect 102704 4146 102732 4626
rect 103796 4480 103848 4486
rect 103796 4422 103848 4428
rect 102692 4140 102744 4146
rect 102692 4082 102744 4088
rect 101956 4072 102008 4078
rect 101956 4014 102008 4020
rect 101968 3738 101996 4014
rect 101956 3732 102008 3738
rect 101956 3674 102008 3680
rect 102704 3602 102732 4082
rect 103612 4072 103664 4078
rect 103612 4014 103664 4020
rect 103060 3936 103112 3942
rect 103060 3878 103112 3884
rect 102692 3596 102744 3602
rect 102692 3538 102744 3544
rect 102704 1970 102732 3538
rect 102968 3528 103020 3534
rect 102968 3470 103020 3476
rect 102980 2990 103008 3470
rect 102968 2984 103020 2990
rect 102968 2926 103020 2932
rect 102968 2372 103020 2378
rect 102968 2314 103020 2320
rect 102980 1970 103008 2314
rect 102692 1964 102744 1970
rect 102692 1906 102744 1912
rect 102968 1964 103020 1970
rect 102968 1906 103020 1912
rect 101956 1760 102008 1766
rect 101956 1702 102008 1708
rect 101968 1426 101996 1702
rect 102704 1426 102732 1906
rect 101956 1420 102008 1426
rect 101956 1362 102008 1368
rect 102692 1420 102744 1426
rect 102692 1362 102744 1368
rect 102968 1216 103020 1222
rect 102968 1158 103020 1164
rect 101784 56 101904 82
rect 102612 56 102732 82
rect 100588 14 100800 42
rect 100942 0 100998 56
rect 101402 0 101458 56
rect 101770 54 101904 56
rect 102598 54 102732 56
rect 101770 0 101826 54
rect 102598 0 102654 54
rect 102704 42 102732 54
rect 102980 42 103008 1158
rect 103072 56 103100 3878
rect 103624 3534 103652 4014
rect 103612 3528 103664 3534
rect 103612 3470 103664 3476
rect 103244 1760 103296 1766
rect 103244 1702 103296 1708
rect 103256 1426 103284 1702
rect 103808 1578 103836 4422
rect 103716 1550 103836 1578
rect 103244 1420 103296 1426
rect 103244 1362 103296 1368
rect 103532 56 103652 82
rect 102704 14 103008 42
rect 103058 0 103114 56
rect 103518 54 103652 56
rect 103518 0 103574 54
rect 103624 42 103652 54
rect 103716 42 103744 1550
rect 103900 56 103928 7142
rect 104820 6866 104848 7278
rect 105096 7002 105124 7278
rect 106188 7200 106240 7206
rect 106188 7142 106240 7148
rect 105084 6996 105136 7002
rect 105084 6938 105136 6944
rect 104808 6860 104860 6866
rect 104808 6802 104860 6808
rect 104820 5234 104848 6802
rect 105084 6792 105136 6798
rect 105084 6734 105136 6740
rect 105096 6254 105124 6734
rect 105084 6248 105136 6254
rect 105084 6190 105136 6196
rect 105096 5846 105124 6190
rect 105084 5840 105136 5846
rect 105084 5782 105136 5788
rect 104992 5772 105044 5778
rect 104992 5714 105044 5720
rect 105004 5234 105032 5714
rect 104808 5228 104860 5234
rect 104808 5170 104860 5176
rect 104992 5228 105044 5234
rect 104992 5170 105044 5176
rect 104820 4690 104848 5170
rect 105084 5024 105136 5030
rect 105084 4966 105136 4972
rect 105096 4690 105124 4966
rect 104808 4684 104860 4690
rect 104808 4626 104860 4632
rect 105084 4684 105136 4690
rect 105084 4626 105136 4632
rect 104820 4146 104848 4626
rect 106004 4480 106056 4486
rect 106004 4422 106056 4428
rect 104808 4140 104860 4146
rect 104808 4082 104860 4088
rect 104820 3602 104848 4082
rect 105452 4072 105504 4078
rect 105452 4014 105504 4020
rect 105176 3936 105228 3942
rect 105176 3878 105228 3884
rect 104808 3596 104860 3602
rect 104808 3538 104860 3544
rect 104820 1970 104848 3538
rect 105084 3528 105136 3534
rect 105084 3470 105136 3476
rect 105096 2990 105124 3470
rect 105084 2984 105136 2990
rect 105084 2926 105136 2932
rect 105096 2582 105124 2926
rect 104900 2576 104952 2582
rect 104900 2518 104952 2524
rect 105084 2576 105136 2582
rect 105084 2518 105136 2524
rect 104808 1964 104860 1970
rect 104808 1906 104860 1912
rect 104820 1426 104848 1906
rect 104912 1902 104940 2518
rect 104900 1896 104952 1902
rect 104900 1838 104952 1844
rect 104808 1420 104860 1426
rect 104808 1362 104860 1368
rect 104992 1216 105044 1222
rect 104992 1158 105044 1164
rect 104728 56 104848 82
rect 103624 14 103744 42
rect 103886 0 103942 56
rect 104714 54 104848 56
rect 104714 0 104770 54
rect 104820 42 104848 54
rect 105004 42 105032 1158
rect 105188 56 105216 3878
rect 105464 3534 105492 4014
rect 105452 3528 105504 3534
rect 105452 3470 105504 3476
rect 105360 1760 105412 1766
rect 105360 1702 105412 1708
rect 105372 1426 105400 1702
rect 106016 1578 106044 4422
rect 105924 1550 106044 1578
rect 105360 1420 105412 1426
rect 105360 1362 105412 1368
rect 105648 56 105768 82
rect 104820 14 105032 42
rect 105174 0 105230 56
rect 105634 54 105768 56
rect 105634 0 105690 54
rect 105740 42 105768 54
rect 105924 42 105952 1550
rect 106016 56 106136 82
rect 105740 14 105952 42
rect 106002 54 106136 56
rect 106002 0 106058 54
rect 106108 42 106136 54
rect 106200 42 106228 7142
rect 106108 14 106228 42
<< via2 >>
rect 4016 7642 4072 7644
rect 4096 7642 4152 7644
rect 4176 7642 4232 7644
rect 4256 7642 4312 7644
rect 4016 7590 4042 7642
rect 4042 7590 4072 7642
rect 4096 7590 4106 7642
rect 4106 7590 4152 7642
rect 4176 7590 4222 7642
rect 4222 7590 4232 7642
rect 4256 7590 4286 7642
rect 4286 7590 4312 7642
rect 4016 7588 4072 7590
rect 4096 7588 4152 7590
rect 4176 7588 4232 7590
rect 4256 7588 4312 7590
rect 34736 7642 34792 7644
rect 34816 7642 34872 7644
rect 34896 7642 34952 7644
rect 34976 7642 35032 7644
rect 34736 7590 34762 7642
rect 34762 7590 34792 7642
rect 34816 7590 34826 7642
rect 34826 7590 34872 7642
rect 34896 7590 34942 7642
rect 34942 7590 34952 7642
rect 34976 7590 35006 7642
rect 35006 7590 35032 7642
rect 34736 7588 34792 7590
rect 34816 7588 34872 7590
rect 34896 7588 34952 7590
rect 34976 7588 35032 7590
rect 65456 7642 65512 7644
rect 65536 7642 65592 7644
rect 65616 7642 65672 7644
rect 65696 7642 65752 7644
rect 65456 7590 65482 7642
rect 65482 7590 65512 7642
rect 65536 7590 65546 7642
rect 65546 7590 65592 7642
rect 65616 7590 65662 7642
rect 65662 7590 65672 7642
rect 65696 7590 65726 7642
rect 65726 7590 65752 7642
rect 65456 7588 65512 7590
rect 65536 7588 65592 7590
rect 65616 7588 65672 7590
rect 65696 7588 65752 7590
rect 96176 7642 96232 7644
rect 96256 7642 96312 7644
rect 96336 7642 96392 7644
rect 96416 7642 96472 7644
rect 96176 7590 96202 7642
rect 96202 7590 96232 7642
rect 96256 7590 96266 7642
rect 96266 7590 96312 7642
rect 96336 7590 96382 7642
rect 96382 7590 96392 7642
rect 96416 7590 96446 7642
rect 96446 7590 96472 7642
rect 96176 7588 96232 7590
rect 96256 7588 96312 7590
rect 96336 7588 96392 7590
rect 96416 7588 96472 7590
rect 1214 2352 1270 2408
rect 4016 6554 4072 6556
rect 4096 6554 4152 6556
rect 4176 6554 4232 6556
rect 4256 6554 4312 6556
rect 4016 6502 4042 6554
rect 4042 6502 4072 6554
rect 4096 6502 4106 6554
rect 4106 6502 4152 6554
rect 4176 6502 4222 6554
rect 4222 6502 4232 6554
rect 4256 6502 4286 6554
rect 4286 6502 4312 6554
rect 4016 6500 4072 6502
rect 4096 6500 4152 6502
rect 4176 6500 4232 6502
rect 4256 6500 4312 6502
rect 4016 5466 4072 5468
rect 4096 5466 4152 5468
rect 4176 5466 4232 5468
rect 4256 5466 4312 5468
rect 4016 5414 4042 5466
rect 4042 5414 4072 5466
rect 4096 5414 4106 5466
rect 4106 5414 4152 5466
rect 4176 5414 4222 5466
rect 4222 5414 4232 5466
rect 4256 5414 4286 5466
rect 4286 5414 4312 5466
rect 4016 5412 4072 5414
rect 4096 5412 4152 5414
rect 4176 5412 4232 5414
rect 4256 5412 4312 5414
rect 4016 4378 4072 4380
rect 4096 4378 4152 4380
rect 4176 4378 4232 4380
rect 4256 4378 4312 4380
rect 4016 4326 4042 4378
rect 4042 4326 4072 4378
rect 4096 4326 4106 4378
rect 4106 4326 4152 4378
rect 4176 4326 4222 4378
rect 4222 4326 4232 4378
rect 4256 4326 4286 4378
rect 4286 4326 4312 4378
rect 4016 4324 4072 4326
rect 4096 4324 4152 4326
rect 4176 4324 4232 4326
rect 4256 4324 4312 4326
rect 4016 3290 4072 3292
rect 4096 3290 4152 3292
rect 4176 3290 4232 3292
rect 4256 3290 4312 3292
rect 4016 3238 4042 3290
rect 4042 3238 4072 3290
rect 4096 3238 4106 3290
rect 4106 3238 4152 3290
rect 4176 3238 4222 3290
rect 4222 3238 4232 3290
rect 4256 3238 4286 3290
rect 4286 3238 4312 3290
rect 4016 3236 4072 3238
rect 4096 3236 4152 3238
rect 4176 3236 4232 3238
rect 4256 3236 4312 3238
rect 4016 2202 4072 2204
rect 4096 2202 4152 2204
rect 4176 2202 4232 2204
rect 4256 2202 4312 2204
rect 4016 2150 4042 2202
rect 4042 2150 4072 2202
rect 4096 2150 4106 2202
rect 4106 2150 4152 2202
rect 4176 2150 4222 2202
rect 4222 2150 4232 2202
rect 4256 2150 4286 2202
rect 4286 2150 4312 2202
rect 4016 2148 4072 2150
rect 4096 2148 4152 2150
rect 4176 2148 4232 2150
rect 4256 2148 4312 2150
rect 4016 1114 4072 1116
rect 4096 1114 4152 1116
rect 4176 1114 4232 1116
rect 4256 1114 4312 1116
rect 4016 1062 4042 1114
rect 4042 1062 4072 1114
rect 4096 1062 4106 1114
rect 4106 1062 4152 1114
rect 4176 1062 4222 1114
rect 4222 1062 4232 1114
rect 4256 1062 4286 1114
rect 4286 1062 4312 1114
rect 4016 1060 4072 1062
rect 4096 1060 4152 1062
rect 4176 1060 4232 1062
rect 4256 1060 4312 1062
rect 19376 7098 19432 7100
rect 19456 7098 19512 7100
rect 19536 7098 19592 7100
rect 19616 7098 19672 7100
rect 19376 7046 19402 7098
rect 19402 7046 19432 7098
rect 19456 7046 19466 7098
rect 19466 7046 19512 7098
rect 19536 7046 19582 7098
rect 19582 7046 19592 7098
rect 19616 7046 19646 7098
rect 19646 7046 19672 7098
rect 19376 7044 19432 7046
rect 19456 7044 19512 7046
rect 19536 7044 19592 7046
rect 19616 7044 19672 7046
rect 19376 6010 19432 6012
rect 19456 6010 19512 6012
rect 19536 6010 19592 6012
rect 19616 6010 19672 6012
rect 19376 5958 19402 6010
rect 19402 5958 19432 6010
rect 19456 5958 19466 6010
rect 19466 5958 19512 6010
rect 19536 5958 19582 6010
rect 19582 5958 19592 6010
rect 19616 5958 19646 6010
rect 19646 5958 19672 6010
rect 19376 5956 19432 5958
rect 19456 5956 19512 5958
rect 19536 5956 19592 5958
rect 19616 5956 19672 5958
rect 19376 4922 19432 4924
rect 19456 4922 19512 4924
rect 19536 4922 19592 4924
rect 19616 4922 19672 4924
rect 19376 4870 19402 4922
rect 19402 4870 19432 4922
rect 19456 4870 19466 4922
rect 19466 4870 19512 4922
rect 19536 4870 19582 4922
rect 19582 4870 19592 4922
rect 19616 4870 19646 4922
rect 19646 4870 19672 4922
rect 19376 4868 19432 4870
rect 19456 4868 19512 4870
rect 19536 4868 19592 4870
rect 19616 4868 19672 4870
rect 19376 3834 19432 3836
rect 19456 3834 19512 3836
rect 19536 3834 19592 3836
rect 19616 3834 19672 3836
rect 19376 3782 19402 3834
rect 19402 3782 19432 3834
rect 19456 3782 19466 3834
rect 19466 3782 19512 3834
rect 19536 3782 19582 3834
rect 19582 3782 19592 3834
rect 19616 3782 19646 3834
rect 19646 3782 19672 3834
rect 19376 3780 19432 3782
rect 19456 3780 19512 3782
rect 19536 3780 19592 3782
rect 19616 3780 19672 3782
rect 19376 2746 19432 2748
rect 19456 2746 19512 2748
rect 19536 2746 19592 2748
rect 19616 2746 19672 2748
rect 19376 2694 19402 2746
rect 19402 2694 19432 2746
rect 19456 2694 19466 2746
rect 19466 2694 19512 2746
rect 19536 2694 19582 2746
rect 19582 2694 19592 2746
rect 19616 2694 19646 2746
rect 19646 2694 19672 2746
rect 19376 2692 19432 2694
rect 19456 2692 19512 2694
rect 19536 2692 19592 2694
rect 19616 2692 19672 2694
rect 19376 1658 19432 1660
rect 19456 1658 19512 1660
rect 19536 1658 19592 1660
rect 19616 1658 19672 1660
rect 19376 1606 19402 1658
rect 19402 1606 19432 1658
rect 19456 1606 19466 1658
rect 19466 1606 19512 1658
rect 19536 1606 19582 1658
rect 19582 1606 19592 1658
rect 19616 1606 19646 1658
rect 19646 1606 19672 1658
rect 19376 1604 19432 1606
rect 19456 1604 19512 1606
rect 19536 1604 19592 1606
rect 19616 1604 19672 1606
rect 34736 6554 34792 6556
rect 34816 6554 34872 6556
rect 34896 6554 34952 6556
rect 34976 6554 35032 6556
rect 34736 6502 34762 6554
rect 34762 6502 34792 6554
rect 34816 6502 34826 6554
rect 34826 6502 34872 6554
rect 34896 6502 34942 6554
rect 34942 6502 34952 6554
rect 34976 6502 35006 6554
rect 35006 6502 35032 6554
rect 34736 6500 34792 6502
rect 34816 6500 34872 6502
rect 34896 6500 34952 6502
rect 34976 6500 35032 6502
rect 34736 5466 34792 5468
rect 34816 5466 34872 5468
rect 34896 5466 34952 5468
rect 34976 5466 35032 5468
rect 34736 5414 34762 5466
rect 34762 5414 34792 5466
rect 34816 5414 34826 5466
rect 34826 5414 34872 5466
rect 34896 5414 34942 5466
rect 34942 5414 34952 5466
rect 34976 5414 35006 5466
rect 35006 5414 35032 5466
rect 34736 5412 34792 5414
rect 34816 5412 34872 5414
rect 34896 5412 34952 5414
rect 34976 5412 35032 5414
rect 34736 4378 34792 4380
rect 34816 4378 34872 4380
rect 34896 4378 34952 4380
rect 34976 4378 35032 4380
rect 34736 4326 34762 4378
rect 34762 4326 34792 4378
rect 34816 4326 34826 4378
rect 34826 4326 34872 4378
rect 34896 4326 34942 4378
rect 34942 4326 34952 4378
rect 34976 4326 35006 4378
rect 35006 4326 35032 4378
rect 34736 4324 34792 4326
rect 34816 4324 34872 4326
rect 34896 4324 34952 4326
rect 34976 4324 35032 4326
rect 34736 3290 34792 3292
rect 34816 3290 34872 3292
rect 34896 3290 34952 3292
rect 34976 3290 35032 3292
rect 34736 3238 34762 3290
rect 34762 3238 34792 3290
rect 34816 3238 34826 3290
rect 34826 3238 34872 3290
rect 34896 3238 34942 3290
rect 34942 3238 34952 3290
rect 34976 3238 35006 3290
rect 35006 3238 35032 3290
rect 34736 3236 34792 3238
rect 34816 3236 34872 3238
rect 34896 3236 34952 3238
rect 34976 3236 35032 3238
rect 34736 2202 34792 2204
rect 34816 2202 34872 2204
rect 34896 2202 34952 2204
rect 34976 2202 35032 2204
rect 34736 2150 34762 2202
rect 34762 2150 34792 2202
rect 34816 2150 34826 2202
rect 34826 2150 34872 2202
rect 34896 2150 34942 2202
rect 34942 2150 34952 2202
rect 34976 2150 35006 2202
rect 35006 2150 35032 2202
rect 34736 2148 34792 2150
rect 34816 2148 34872 2150
rect 34896 2148 34952 2150
rect 34976 2148 35032 2150
rect 34736 1114 34792 1116
rect 34816 1114 34872 1116
rect 34896 1114 34952 1116
rect 34976 1114 35032 1116
rect 34736 1062 34762 1114
rect 34762 1062 34792 1114
rect 34816 1062 34826 1114
rect 34826 1062 34872 1114
rect 34896 1062 34942 1114
rect 34942 1062 34952 1114
rect 34976 1062 35006 1114
rect 35006 1062 35032 1114
rect 34736 1060 34792 1062
rect 34816 1060 34872 1062
rect 34896 1060 34952 1062
rect 34976 1060 35032 1062
rect 50096 7098 50152 7100
rect 50176 7098 50232 7100
rect 50256 7098 50312 7100
rect 50336 7098 50392 7100
rect 50096 7046 50122 7098
rect 50122 7046 50152 7098
rect 50176 7046 50186 7098
rect 50186 7046 50232 7098
rect 50256 7046 50302 7098
rect 50302 7046 50312 7098
rect 50336 7046 50366 7098
rect 50366 7046 50392 7098
rect 50096 7044 50152 7046
rect 50176 7044 50232 7046
rect 50256 7044 50312 7046
rect 50336 7044 50392 7046
rect 50096 6010 50152 6012
rect 50176 6010 50232 6012
rect 50256 6010 50312 6012
rect 50336 6010 50392 6012
rect 50096 5958 50122 6010
rect 50122 5958 50152 6010
rect 50176 5958 50186 6010
rect 50186 5958 50232 6010
rect 50256 5958 50302 6010
rect 50302 5958 50312 6010
rect 50336 5958 50366 6010
rect 50366 5958 50392 6010
rect 50096 5956 50152 5958
rect 50176 5956 50232 5958
rect 50256 5956 50312 5958
rect 50336 5956 50392 5958
rect 50096 4922 50152 4924
rect 50176 4922 50232 4924
rect 50256 4922 50312 4924
rect 50336 4922 50392 4924
rect 50096 4870 50122 4922
rect 50122 4870 50152 4922
rect 50176 4870 50186 4922
rect 50186 4870 50232 4922
rect 50256 4870 50302 4922
rect 50302 4870 50312 4922
rect 50336 4870 50366 4922
rect 50366 4870 50392 4922
rect 50096 4868 50152 4870
rect 50176 4868 50232 4870
rect 50256 4868 50312 4870
rect 50336 4868 50392 4870
rect 50096 3834 50152 3836
rect 50176 3834 50232 3836
rect 50256 3834 50312 3836
rect 50336 3834 50392 3836
rect 50096 3782 50122 3834
rect 50122 3782 50152 3834
rect 50176 3782 50186 3834
rect 50186 3782 50232 3834
rect 50256 3782 50302 3834
rect 50302 3782 50312 3834
rect 50336 3782 50366 3834
rect 50366 3782 50392 3834
rect 50096 3780 50152 3782
rect 50176 3780 50232 3782
rect 50256 3780 50312 3782
rect 50336 3780 50392 3782
rect 50096 2746 50152 2748
rect 50176 2746 50232 2748
rect 50256 2746 50312 2748
rect 50336 2746 50392 2748
rect 50096 2694 50122 2746
rect 50122 2694 50152 2746
rect 50176 2694 50186 2746
rect 50186 2694 50232 2746
rect 50256 2694 50302 2746
rect 50302 2694 50312 2746
rect 50336 2694 50366 2746
rect 50366 2694 50392 2746
rect 50096 2692 50152 2694
rect 50176 2692 50232 2694
rect 50256 2692 50312 2694
rect 50336 2692 50392 2694
rect 50096 1658 50152 1660
rect 50176 1658 50232 1660
rect 50256 1658 50312 1660
rect 50336 1658 50392 1660
rect 50096 1606 50122 1658
rect 50122 1606 50152 1658
rect 50176 1606 50186 1658
rect 50186 1606 50232 1658
rect 50256 1606 50302 1658
rect 50302 1606 50312 1658
rect 50336 1606 50366 1658
rect 50366 1606 50392 1658
rect 50096 1604 50152 1606
rect 50176 1604 50232 1606
rect 50256 1604 50312 1606
rect 50336 1604 50392 1606
rect 65456 6554 65512 6556
rect 65536 6554 65592 6556
rect 65616 6554 65672 6556
rect 65696 6554 65752 6556
rect 65456 6502 65482 6554
rect 65482 6502 65512 6554
rect 65536 6502 65546 6554
rect 65546 6502 65592 6554
rect 65616 6502 65662 6554
rect 65662 6502 65672 6554
rect 65696 6502 65726 6554
rect 65726 6502 65752 6554
rect 65456 6500 65512 6502
rect 65536 6500 65592 6502
rect 65616 6500 65672 6502
rect 65696 6500 65752 6502
rect 65456 5466 65512 5468
rect 65536 5466 65592 5468
rect 65616 5466 65672 5468
rect 65696 5466 65752 5468
rect 65456 5414 65482 5466
rect 65482 5414 65512 5466
rect 65536 5414 65546 5466
rect 65546 5414 65592 5466
rect 65616 5414 65662 5466
rect 65662 5414 65672 5466
rect 65696 5414 65726 5466
rect 65726 5414 65752 5466
rect 65456 5412 65512 5414
rect 65536 5412 65592 5414
rect 65616 5412 65672 5414
rect 65696 5412 65752 5414
rect 65456 4378 65512 4380
rect 65536 4378 65592 4380
rect 65616 4378 65672 4380
rect 65696 4378 65752 4380
rect 65456 4326 65482 4378
rect 65482 4326 65512 4378
rect 65536 4326 65546 4378
rect 65546 4326 65592 4378
rect 65616 4326 65662 4378
rect 65662 4326 65672 4378
rect 65696 4326 65726 4378
rect 65726 4326 65752 4378
rect 65456 4324 65512 4326
rect 65536 4324 65592 4326
rect 65616 4324 65672 4326
rect 65696 4324 65752 4326
rect 65456 3290 65512 3292
rect 65536 3290 65592 3292
rect 65616 3290 65672 3292
rect 65696 3290 65752 3292
rect 65456 3238 65482 3290
rect 65482 3238 65512 3290
rect 65536 3238 65546 3290
rect 65546 3238 65592 3290
rect 65616 3238 65662 3290
rect 65662 3238 65672 3290
rect 65696 3238 65726 3290
rect 65726 3238 65752 3290
rect 65456 3236 65512 3238
rect 65536 3236 65592 3238
rect 65616 3236 65672 3238
rect 65696 3236 65752 3238
rect 65456 2202 65512 2204
rect 65536 2202 65592 2204
rect 65616 2202 65672 2204
rect 65696 2202 65752 2204
rect 65456 2150 65482 2202
rect 65482 2150 65512 2202
rect 65536 2150 65546 2202
rect 65546 2150 65592 2202
rect 65616 2150 65662 2202
rect 65662 2150 65672 2202
rect 65696 2150 65726 2202
rect 65726 2150 65752 2202
rect 65456 2148 65512 2150
rect 65536 2148 65592 2150
rect 65616 2148 65672 2150
rect 65696 2148 65752 2150
rect 65456 1114 65512 1116
rect 65536 1114 65592 1116
rect 65616 1114 65672 1116
rect 65696 1114 65752 1116
rect 65456 1062 65482 1114
rect 65482 1062 65512 1114
rect 65536 1062 65546 1114
rect 65546 1062 65592 1114
rect 65616 1062 65662 1114
rect 65662 1062 65672 1114
rect 65696 1062 65726 1114
rect 65726 1062 65752 1114
rect 65456 1060 65512 1062
rect 65536 1060 65592 1062
rect 65616 1060 65672 1062
rect 65696 1060 65752 1062
rect 80816 7098 80872 7100
rect 80896 7098 80952 7100
rect 80976 7098 81032 7100
rect 81056 7098 81112 7100
rect 80816 7046 80842 7098
rect 80842 7046 80872 7098
rect 80896 7046 80906 7098
rect 80906 7046 80952 7098
rect 80976 7046 81022 7098
rect 81022 7046 81032 7098
rect 81056 7046 81086 7098
rect 81086 7046 81112 7098
rect 80816 7044 80872 7046
rect 80896 7044 80952 7046
rect 80976 7044 81032 7046
rect 81056 7044 81112 7046
rect 80816 6010 80872 6012
rect 80896 6010 80952 6012
rect 80976 6010 81032 6012
rect 81056 6010 81112 6012
rect 80816 5958 80842 6010
rect 80842 5958 80872 6010
rect 80896 5958 80906 6010
rect 80906 5958 80952 6010
rect 80976 5958 81022 6010
rect 81022 5958 81032 6010
rect 81056 5958 81086 6010
rect 81086 5958 81112 6010
rect 80816 5956 80872 5958
rect 80896 5956 80952 5958
rect 80976 5956 81032 5958
rect 81056 5956 81112 5958
rect 80816 4922 80872 4924
rect 80896 4922 80952 4924
rect 80976 4922 81032 4924
rect 81056 4922 81112 4924
rect 80816 4870 80842 4922
rect 80842 4870 80872 4922
rect 80896 4870 80906 4922
rect 80906 4870 80952 4922
rect 80976 4870 81022 4922
rect 81022 4870 81032 4922
rect 81056 4870 81086 4922
rect 81086 4870 81112 4922
rect 80816 4868 80872 4870
rect 80896 4868 80952 4870
rect 80976 4868 81032 4870
rect 81056 4868 81112 4870
rect 80816 3834 80872 3836
rect 80896 3834 80952 3836
rect 80976 3834 81032 3836
rect 81056 3834 81112 3836
rect 80816 3782 80842 3834
rect 80842 3782 80872 3834
rect 80896 3782 80906 3834
rect 80906 3782 80952 3834
rect 80976 3782 81022 3834
rect 81022 3782 81032 3834
rect 81056 3782 81086 3834
rect 81086 3782 81112 3834
rect 80816 3780 80872 3782
rect 80896 3780 80952 3782
rect 80976 3780 81032 3782
rect 81056 3780 81112 3782
rect 80816 2746 80872 2748
rect 80896 2746 80952 2748
rect 80976 2746 81032 2748
rect 81056 2746 81112 2748
rect 80816 2694 80842 2746
rect 80842 2694 80872 2746
rect 80896 2694 80906 2746
rect 80906 2694 80952 2746
rect 80976 2694 81022 2746
rect 81022 2694 81032 2746
rect 81056 2694 81086 2746
rect 81086 2694 81112 2746
rect 80816 2692 80872 2694
rect 80896 2692 80952 2694
rect 80976 2692 81032 2694
rect 81056 2692 81112 2694
rect 80816 1658 80872 1660
rect 80896 1658 80952 1660
rect 80976 1658 81032 1660
rect 81056 1658 81112 1660
rect 80816 1606 80842 1658
rect 80842 1606 80872 1658
rect 80896 1606 80906 1658
rect 80906 1606 80952 1658
rect 80976 1606 81022 1658
rect 81022 1606 81032 1658
rect 81056 1606 81086 1658
rect 81086 1606 81112 1658
rect 80816 1604 80872 1606
rect 80896 1604 80952 1606
rect 80976 1604 81032 1606
rect 81056 1604 81112 1606
rect 96176 6554 96232 6556
rect 96256 6554 96312 6556
rect 96336 6554 96392 6556
rect 96416 6554 96472 6556
rect 96176 6502 96202 6554
rect 96202 6502 96232 6554
rect 96256 6502 96266 6554
rect 96266 6502 96312 6554
rect 96336 6502 96382 6554
rect 96382 6502 96392 6554
rect 96416 6502 96446 6554
rect 96446 6502 96472 6554
rect 96176 6500 96232 6502
rect 96256 6500 96312 6502
rect 96336 6500 96392 6502
rect 96416 6500 96472 6502
rect 96176 5466 96232 5468
rect 96256 5466 96312 5468
rect 96336 5466 96392 5468
rect 96416 5466 96472 5468
rect 96176 5414 96202 5466
rect 96202 5414 96232 5466
rect 96256 5414 96266 5466
rect 96266 5414 96312 5466
rect 96336 5414 96382 5466
rect 96382 5414 96392 5466
rect 96416 5414 96446 5466
rect 96446 5414 96472 5466
rect 96176 5412 96232 5414
rect 96256 5412 96312 5414
rect 96336 5412 96392 5414
rect 96416 5412 96472 5414
rect 96176 4378 96232 4380
rect 96256 4378 96312 4380
rect 96336 4378 96392 4380
rect 96416 4378 96472 4380
rect 96176 4326 96202 4378
rect 96202 4326 96232 4378
rect 96256 4326 96266 4378
rect 96266 4326 96312 4378
rect 96336 4326 96382 4378
rect 96382 4326 96392 4378
rect 96416 4326 96446 4378
rect 96446 4326 96472 4378
rect 96176 4324 96232 4326
rect 96256 4324 96312 4326
rect 96336 4324 96392 4326
rect 96416 4324 96472 4326
rect 96176 3290 96232 3292
rect 96256 3290 96312 3292
rect 96336 3290 96392 3292
rect 96416 3290 96472 3292
rect 96176 3238 96202 3290
rect 96202 3238 96232 3290
rect 96256 3238 96266 3290
rect 96266 3238 96312 3290
rect 96336 3238 96382 3290
rect 96382 3238 96392 3290
rect 96416 3238 96446 3290
rect 96446 3238 96472 3290
rect 96176 3236 96232 3238
rect 96256 3236 96312 3238
rect 96336 3236 96392 3238
rect 96416 3236 96472 3238
rect 96176 2202 96232 2204
rect 96256 2202 96312 2204
rect 96336 2202 96392 2204
rect 96416 2202 96472 2204
rect 96176 2150 96202 2202
rect 96202 2150 96232 2202
rect 96256 2150 96266 2202
rect 96266 2150 96312 2202
rect 96336 2150 96382 2202
rect 96382 2150 96392 2202
rect 96416 2150 96446 2202
rect 96446 2150 96472 2202
rect 96176 2148 96232 2150
rect 96256 2148 96312 2150
rect 96336 2148 96392 2150
rect 96416 2148 96472 2150
rect 96176 1114 96232 1116
rect 96256 1114 96312 1116
rect 96336 1114 96392 1116
rect 96416 1114 96472 1116
rect 96176 1062 96202 1114
rect 96202 1062 96232 1114
rect 96256 1062 96266 1114
rect 96266 1062 96312 1114
rect 96336 1062 96382 1114
rect 96382 1062 96392 1114
rect 96416 1062 96446 1114
rect 96446 1062 96472 1114
rect 96176 1060 96232 1062
rect 96256 1060 96312 1062
rect 96336 1060 96392 1062
rect 96416 1060 96472 1062
<< metal3 >>
rect 4004 7648 4324 7649
rect 4004 7584 4012 7648
rect 4076 7584 4092 7648
rect 4156 7584 4172 7648
rect 4236 7584 4252 7648
rect 4316 7584 4324 7648
rect 4004 7583 4324 7584
rect 34724 7648 35044 7649
rect 34724 7584 34732 7648
rect 34796 7584 34812 7648
rect 34876 7584 34892 7648
rect 34956 7584 34972 7648
rect 35036 7584 35044 7648
rect 34724 7583 35044 7584
rect 65444 7648 65764 7649
rect 65444 7584 65452 7648
rect 65516 7584 65532 7648
rect 65596 7584 65612 7648
rect 65676 7584 65692 7648
rect 65756 7584 65764 7648
rect 65444 7583 65764 7584
rect 96164 7648 96484 7649
rect 96164 7584 96172 7648
rect 96236 7584 96252 7648
rect 96316 7584 96332 7648
rect 96396 7584 96412 7648
rect 96476 7584 96484 7648
rect 96164 7583 96484 7584
rect 19364 7104 19684 7105
rect 19364 7040 19372 7104
rect 19436 7040 19452 7104
rect 19516 7040 19532 7104
rect 19596 7040 19612 7104
rect 19676 7040 19684 7104
rect 19364 7039 19684 7040
rect 50084 7104 50404 7105
rect 50084 7040 50092 7104
rect 50156 7040 50172 7104
rect 50236 7040 50252 7104
rect 50316 7040 50332 7104
rect 50396 7040 50404 7104
rect 50084 7039 50404 7040
rect 80804 7104 81124 7105
rect 80804 7040 80812 7104
rect 80876 7040 80892 7104
rect 80956 7040 80972 7104
rect 81036 7040 81052 7104
rect 81116 7040 81124 7104
rect 80804 7039 81124 7040
rect 4004 6560 4324 6561
rect 4004 6496 4012 6560
rect 4076 6496 4092 6560
rect 4156 6496 4172 6560
rect 4236 6496 4252 6560
rect 4316 6496 4324 6560
rect 4004 6495 4324 6496
rect 34724 6560 35044 6561
rect 34724 6496 34732 6560
rect 34796 6496 34812 6560
rect 34876 6496 34892 6560
rect 34956 6496 34972 6560
rect 35036 6496 35044 6560
rect 34724 6495 35044 6496
rect 65444 6560 65764 6561
rect 65444 6496 65452 6560
rect 65516 6496 65532 6560
rect 65596 6496 65612 6560
rect 65676 6496 65692 6560
rect 65756 6496 65764 6560
rect 65444 6495 65764 6496
rect 96164 6560 96484 6561
rect 96164 6496 96172 6560
rect 96236 6496 96252 6560
rect 96316 6496 96332 6560
rect 96396 6496 96412 6560
rect 96476 6496 96484 6560
rect 96164 6495 96484 6496
rect 19364 6016 19684 6017
rect 19364 5952 19372 6016
rect 19436 5952 19452 6016
rect 19516 5952 19532 6016
rect 19596 5952 19612 6016
rect 19676 5952 19684 6016
rect 19364 5951 19684 5952
rect 50084 6016 50404 6017
rect 50084 5952 50092 6016
rect 50156 5952 50172 6016
rect 50236 5952 50252 6016
rect 50316 5952 50332 6016
rect 50396 5952 50404 6016
rect 50084 5951 50404 5952
rect 80804 6016 81124 6017
rect 80804 5952 80812 6016
rect 80876 5952 80892 6016
rect 80956 5952 80972 6016
rect 81036 5952 81052 6016
rect 81116 5952 81124 6016
rect 80804 5951 81124 5952
rect 4004 5472 4324 5473
rect 4004 5408 4012 5472
rect 4076 5408 4092 5472
rect 4156 5408 4172 5472
rect 4236 5408 4252 5472
rect 4316 5408 4324 5472
rect 4004 5407 4324 5408
rect 34724 5472 35044 5473
rect 34724 5408 34732 5472
rect 34796 5408 34812 5472
rect 34876 5408 34892 5472
rect 34956 5408 34972 5472
rect 35036 5408 35044 5472
rect 34724 5407 35044 5408
rect 65444 5472 65764 5473
rect 65444 5408 65452 5472
rect 65516 5408 65532 5472
rect 65596 5408 65612 5472
rect 65676 5408 65692 5472
rect 65756 5408 65764 5472
rect 65444 5407 65764 5408
rect 96164 5472 96484 5473
rect 96164 5408 96172 5472
rect 96236 5408 96252 5472
rect 96316 5408 96332 5472
rect 96396 5408 96412 5472
rect 96476 5408 96484 5472
rect 96164 5407 96484 5408
rect 19364 4928 19684 4929
rect 19364 4864 19372 4928
rect 19436 4864 19452 4928
rect 19516 4864 19532 4928
rect 19596 4864 19612 4928
rect 19676 4864 19684 4928
rect 19364 4863 19684 4864
rect 50084 4928 50404 4929
rect 50084 4864 50092 4928
rect 50156 4864 50172 4928
rect 50236 4864 50252 4928
rect 50316 4864 50332 4928
rect 50396 4864 50404 4928
rect 50084 4863 50404 4864
rect 80804 4928 81124 4929
rect 80804 4864 80812 4928
rect 80876 4864 80892 4928
rect 80956 4864 80972 4928
rect 81036 4864 81052 4928
rect 81116 4864 81124 4928
rect 80804 4863 81124 4864
rect 4004 4384 4324 4385
rect 4004 4320 4012 4384
rect 4076 4320 4092 4384
rect 4156 4320 4172 4384
rect 4236 4320 4252 4384
rect 4316 4320 4324 4384
rect 4004 4319 4324 4320
rect 34724 4384 35044 4385
rect 34724 4320 34732 4384
rect 34796 4320 34812 4384
rect 34876 4320 34892 4384
rect 34956 4320 34972 4384
rect 35036 4320 35044 4384
rect 34724 4319 35044 4320
rect 65444 4384 65764 4385
rect 65444 4320 65452 4384
rect 65516 4320 65532 4384
rect 65596 4320 65612 4384
rect 65676 4320 65692 4384
rect 65756 4320 65764 4384
rect 65444 4319 65764 4320
rect 96164 4384 96484 4385
rect 96164 4320 96172 4384
rect 96236 4320 96252 4384
rect 96316 4320 96332 4384
rect 96396 4320 96412 4384
rect 96476 4320 96484 4384
rect 96164 4319 96484 4320
rect 19364 3840 19684 3841
rect 19364 3776 19372 3840
rect 19436 3776 19452 3840
rect 19516 3776 19532 3840
rect 19596 3776 19612 3840
rect 19676 3776 19684 3840
rect 19364 3775 19684 3776
rect 50084 3840 50404 3841
rect 50084 3776 50092 3840
rect 50156 3776 50172 3840
rect 50236 3776 50252 3840
rect 50316 3776 50332 3840
rect 50396 3776 50404 3840
rect 50084 3775 50404 3776
rect 80804 3840 81124 3841
rect 80804 3776 80812 3840
rect 80876 3776 80892 3840
rect 80956 3776 80972 3840
rect 81036 3776 81052 3840
rect 81116 3776 81124 3840
rect 80804 3775 81124 3776
rect 4004 3296 4324 3297
rect 4004 3232 4012 3296
rect 4076 3232 4092 3296
rect 4156 3232 4172 3296
rect 4236 3232 4252 3296
rect 4316 3232 4324 3296
rect 4004 3231 4324 3232
rect 34724 3296 35044 3297
rect 34724 3232 34732 3296
rect 34796 3232 34812 3296
rect 34876 3232 34892 3296
rect 34956 3232 34972 3296
rect 35036 3232 35044 3296
rect 34724 3231 35044 3232
rect 65444 3296 65764 3297
rect 65444 3232 65452 3296
rect 65516 3232 65532 3296
rect 65596 3232 65612 3296
rect 65676 3232 65692 3296
rect 65756 3232 65764 3296
rect 65444 3231 65764 3232
rect 96164 3296 96484 3297
rect 96164 3232 96172 3296
rect 96236 3232 96252 3296
rect 96316 3232 96332 3296
rect 96396 3232 96412 3296
rect 96476 3232 96484 3296
rect 96164 3231 96484 3232
rect 19364 2752 19684 2753
rect 19364 2688 19372 2752
rect 19436 2688 19452 2752
rect 19516 2688 19532 2752
rect 19596 2688 19612 2752
rect 19676 2688 19684 2752
rect 19364 2687 19684 2688
rect 50084 2752 50404 2753
rect 50084 2688 50092 2752
rect 50156 2688 50172 2752
rect 50236 2688 50252 2752
rect 50316 2688 50332 2752
rect 50396 2688 50404 2752
rect 50084 2687 50404 2688
rect 80804 2752 81124 2753
rect 80804 2688 80812 2752
rect 80876 2688 80892 2752
rect 80956 2688 80972 2752
rect 81036 2688 81052 2752
rect 81116 2688 81124 2752
rect 80804 2687 81124 2688
rect 1209 2410 1275 2413
rect 30 2408 1275 2410
rect 30 2352 1214 2408
rect 1270 2352 1275 2408
rect 30 2350 1275 2352
rect 30 2168 90 2350
rect 1209 2347 1275 2350
rect 4004 2208 4324 2209
rect 0 2048 120 2168
rect 4004 2144 4012 2208
rect 4076 2144 4092 2208
rect 4156 2144 4172 2208
rect 4236 2144 4252 2208
rect 4316 2144 4324 2208
rect 4004 2143 4324 2144
rect 34724 2208 35044 2209
rect 34724 2144 34732 2208
rect 34796 2144 34812 2208
rect 34876 2144 34892 2208
rect 34956 2144 34972 2208
rect 35036 2144 35044 2208
rect 34724 2143 35044 2144
rect 65444 2208 65764 2209
rect 65444 2144 65452 2208
rect 65516 2144 65532 2208
rect 65596 2144 65612 2208
rect 65676 2144 65692 2208
rect 65756 2144 65764 2208
rect 65444 2143 65764 2144
rect 96164 2208 96484 2209
rect 96164 2144 96172 2208
rect 96236 2144 96252 2208
rect 96316 2144 96332 2208
rect 96396 2144 96412 2208
rect 96476 2144 96484 2208
rect 96164 2143 96484 2144
rect 19364 1664 19684 1665
rect 19364 1600 19372 1664
rect 19436 1600 19452 1664
rect 19516 1600 19532 1664
rect 19596 1600 19612 1664
rect 19676 1600 19684 1664
rect 19364 1599 19684 1600
rect 50084 1664 50404 1665
rect 50084 1600 50092 1664
rect 50156 1600 50172 1664
rect 50236 1600 50252 1664
rect 50316 1600 50332 1664
rect 50396 1600 50404 1664
rect 50084 1599 50404 1600
rect 80804 1664 81124 1665
rect 80804 1600 80812 1664
rect 80876 1600 80892 1664
rect 80956 1600 80972 1664
rect 81036 1600 81052 1664
rect 81116 1600 81124 1664
rect 80804 1599 81124 1600
rect 4004 1120 4324 1121
rect 4004 1056 4012 1120
rect 4076 1056 4092 1120
rect 4156 1056 4172 1120
rect 4236 1056 4252 1120
rect 4316 1056 4324 1120
rect 4004 1055 4324 1056
rect 34724 1120 35044 1121
rect 34724 1056 34732 1120
rect 34796 1056 34812 1120
rect 34876 1056 34892 1120
rect 34956 1056 34972 1120
rect 35036 1056 35044 1120
rect 34724 1055 35044 1056
rect 65444 1120 65764 1121
rect 65444 1056 65452 1120
rect 65516 1056 65532 1120
rect 65596 1056 65612 1120
rect 65676 1056 65692 1120
rect 65756 1056 65764 1120
rect 65444 1055 65764 1056
rect 96164 1120 96484 1121
rect 96164 1056 96172 1120
rect 96236 1056 96252 1120
rect 96316 1056 96332 1120
rect 96396 1056 96412 1120
rect 96476 1056 96484 1120
rect 96164 1055 96484 1056
<< via3 >>
rect 4012 7644 4076 7648
rect 4012 7588 4016 7644
rect 4016 7588 4072 7644
rect 4072 7588 4076 7644
rect 4012 7584 4076 7588
rect 4092 7644 4156 7648
rect 4092 7588 4096 7644
rect 4096 7588 4152 7644
rect 4152 7588 4156 7644
rect 4092 7584 4156 7588
rect 4172 7644 4236 7648
rect 4172 7588 4176 7644
rect 4176 7588 4232 7644
rect 4232 7588 4236 7644
rect 4172 7584 4236 7588
rect 4252 7644 4316 7648
rect 4252 7588 4256 7644
rect 4256 7588 4312 7644
rect 4312 7588 4316 7644
rect 4252 7584 4316 7588
rect 34732 7644 34796 7648
rect 34732 7588 34736 7644
rect 34736 7588 34792 7644
rect 34792 7588 34796 7644
rect 34732 7584 34796 7588
rect 34812 7644 34876 7648
rect 34812 7588 34816 7644
rect 34816 7588 34872 7644
rect 34872 7588 34876 7644
rect 34812 7584 34876 7588
rect 34892 7644 34956 7648
rect 34892 7588 34896 7644
rect 34896 7588 34952 7644
rect 34952 7588 34956 7644
rect 34892 7584 34956 7588
rect 34972 7644 35036 7648
rect 34972 7588 34976 7644
rect 34976 7588 35032 7644
rect 35032 7588 35036 7644
rect 34972 7584 35036 7588
rect 65452 7644 65516 7648
rect 65452 7588 65456 7644
rect 65456 7588 65512 7644
rect 65512 7588 65516 7644
rect 65452 7584 65516 7588
rect 65532 7644 65596 7648
rect 65532 7588 65536 7644
rect 65536 7588 65592 7644
rect 65592 7588 65596 7644
rect 65532 7584 65596 7588
rect 65612 7644 65676 7648
rect 65612 7588 65616 7644
rect 65616 7588 65672 7644
rect 65672 7588 65676 7644
rect 65612 7584 65676 7588
rect 65692 7644 65756 7648
rect 65692 7588 65696 7644
rect 65696 7588 65752 7644
rect 65752 7588 65756 7644
rect 65692 7584 65756 7588
rect 96172 7644 96236 7648
rect 96172 7588 96176 7644
rect 96176 7588 96232 7644
rect 96232 7588 96236 7644
rect 96172 7584 96236 7588
rect 96252 7644 96316 7648
rect 96252 7588 96256 7644
rect 96256 7588 96312 7644
rect 96312 7588 96316 7644
rect 96252 7584 96316 7588
rect 96332 7644 96396 7648
rect 96332 7588 96336 7644
rect 96336 7588 96392 7644
rect 96392 7588 96396 7644
rect 96332 7584 96396 7588
rect 96412 7644 96476 7648
rect 96412 7588 96416 7644
rect 96416 7588 96472 7644
rect 96472 7588 96476 7644
rect 96412 7584 96476 7588
rect 19372 7100 19436 7104
rect 19372 7044 19376 7100
rect 19376 7044 19432 7100
rect 19432 7044 19436 7100
rect 19372 7040 19436 7044
rect 19452 7100 19516 7104
rect 19452 7044 19456 7100
rect 19456 7044 19512 7100
rect 19512 7044 19516 7100
rect 19452 7040 19516 7044
rect 19532 7100 19596 7104
rect 19532 7044 19536 7100
rect 19536 7044 19592 7100
rect 19592 7044 19596 7100
rect 19532 7040 19596 7044
rect 19612 7100 19676 7104
rect 19612 7044 19616 7100
rect 19616 7044 19672 7100
rect 19672 7044 19676 7100
rect 19612 7040 19676 7044
rect 50092 7100 50156 7104
rect 50092 7044 50096 7100
rect 50096 7044 50152 7100
rect 50152 7044 50156 7100
rect 50092 7040 50156 7044
rect 50172 7100 50236 7104
rect 50172 7044 50176 7100
rect 50176 7044 50232 7100
rect 50232 7044 50236 7100
rect 50172 7040 50236 7044
rect 50252 7100 50316 7104
rect 50252 7044 50256 7100
rect 50256 7044 50312 7100
rect 50312 7044 50316 7100
rect 50252 7040 50316 7044
rect 50332 7100 50396 7104
rect 50332 7044 50336 7100
rect 50336 7044 50392 7100
rect 50392 7044 50396 7100
rect 50332 7040 50396 7044
rect 80812 7100 80876 7104
rect 80812 7044 80816 7100
rect 80816 7044 80872 7100
rect 80872 7044 80876 7100
rect 80812 7040 80876 7044
rect 80892 7100 80956 7104
rect 80892 7044 80896 7100
rect 80896 7044 80952 7100
rect 80952 7044 80956 7100
rect 80892 7040 80956 7044
rect 80972 7100 81036 7104
rect 80972 7044 80976 7100
rect 80976 7044 81032 7100
rect 81032 7044 81036 7100
rect 80972 7040 81036 7044
rect 81052 7100 81116 7104
rect 81052 7044 81056 7100
rect 81056 7044 81112 7100
rect 81112 7044 81116 7100
rect 81052 7040 81116 7044
rect 4012 6556 4076 6560
rect 4012 6500 4016 6556
rect 4016 6500 4072 6556
rect 4072 6500 4076 6556
rect 4012 6496 4076 6500
rect 4092 6556 4156 6560
rect 4092 6500 4096 6556
rect 4096 6500 4152 6556
rect 4152 6500 4156 6556
rect 4092 6496 4156 6500
rect 4172 6556 4236 6560
rect 4172 6500 4176 6556
rect 4176 6500 4232 6556
rect 4232 6500 4236 6556
rect 4172 6496 4236 6500
rect 4252 6556 4316 6560
rect 4252 6500 4256 6556
rect 4256 6500 4312 6556
rect 4312 6500 4316 6556
rect 4252 6496 4316 6500
rect 34732 6556 34796 6560
rect 34732 6500 34736 6556
rect 34736 6500 34792 6556
rect 34792 6500 34796 6556
rect 34732 6496 34796 6500
rect 34812 6556 34876 6560
rect 34812 6500 34816 6556
rect 34816 6500 34872 6556
rect 34872 6500 34876 6556
rect 34812 6496 34876 6500
rect 34892 6556 34956 6560
rect 34892 6500 34896 6556
rect 34896 6500 34952 6556
rect 34952 6500 34956 6556
rect 34892 6496 34956 6500
rect 34972 6556 35036 6560
rect 34972 6500 34976 6556
rect 34976 6500 35032 6556
rect 35032 6500 35036 6556
rect 34972 6496 35036 6500
rect 65452 6556 65516 6560
rect 65452 6500 65456 6556
rect 65456 6500 65512 6556
rect 65512 6500 65516 6556
rect 65452 6496 65516 6500
rect 65532 6556 65596 6560
rect 65532 6500 65536 6556
rect 65536 6500 65592 6556
rect 65592 6500 65596 6556
rect 65532 6496 65596 6500
rect 65612 6556 65676 6560
rect 65612 6500 65616 6556
rect 65616 6500 65672 6556
rect 65672 6500 65676 6556
rect 65612 6496 65676 6500
rect 65692 6556 65756 6560
rect 65692 6500 65696 6556
rect 65696 6500 65752 6556
rect 65752 6500 65756 6556
rect 65692 6496 65756 6500
rect 96172 6556 96236 6560
rect 96172 6500 96176 6556
rect 96176 6500 96232 6556
rect 96232 6500 96236 6556
rect 96172 6496 96236 6500
rect 96252 6556 96316 6560
rect 96252 6500 96256 6556
rect 96256 6500 96312 6556
rect 96312 6500 96316 6556
rect 96252 6496 96316 6500
rect 96332 6556 96396 6560
rect 96332 6500 96336 6556
rect 96336 6500 96392 6556
rect 96392 6500 96396 6556
rect 96332 6496 96396 6500
rect 96412 6556 96476 6560
rect 96412 6500 96416 6556
rect 96416 6500 96472 6556
rect 96472 6500 96476 6556
rect 96412 6496 96476 6500
rect 19372 6012 19436 6016
rect 19372 5956 19376 6012
rect 19376 5956 19432 6012
rect 19432 5956 19436 6012
rect 19372 5952 19436 5956
rect 19452 6012 19516 6016
rect 19452 5956 19456 6012
rect 19456 5956 19512 6012
rect 19512 5956 19516 6012
rect 19452 5952 19516 5956
rect 19532 6012 19596 6016
rect 19532 5956 19536 6012
rect 19536 5956 19592 6012
rect 19592 5956 19596 6012
rect 19532 5952 19596 5956
rect 19612 6012 19676 6016
rect 19612 5956 19616 6012
rect 19616 5956 19672 6012
rect 19672 5956 19676 6012
rect 19612 5952 19676 5956
rect 50092 6012 50156 6016
rect 50092 5956 50096 6012
rect 50096 5956 50152 6012
rect 50152 5956 50156 6012
rect 50092 5952 50156 5956
rect 50172 6012 50236 6016
rect 50172 5956 50176 6012
rect 50176 5956 50232 6012
rect 50232 5956 50236 6012
rect 50172 5952 50236 5956
rect 50252 6012 50316 6016
rect 50252 5956 50256 6012
rect 50256 5956 50312 6012
rect 50312 5956 50316 6012
rect 50252 5952 50316 5956
rect 50332 6012 50396 6016
rect 50332 5956 50336 6012
rect 50336 5956 50392 6012
rect 50392 5956 50396 6012
rect 50332 5952 50396 5956
rect 80812 6012 80876 6016
rect 80812 5956 80816 6012
rect 80816 5956 80872 6012
rect 80872 5956 80876 6012
rect 80812 5952 80876 5956
rect 80892 6012 80956 6016
rect 80892 5956 80896 6012
rect 80896 5956 80952 6012
rect 80952 5956 80956 6012
rect 80892 5952 80956 5956
rect 80972 6012 81036 6016
rect 80972 5956 80976 6012
rect 80976 5956 81032 6012
rect 81032 5956 81036 6012
rect 80972 5952 81036 5956
rect 81052 6012 81116 6016
rect 81052 5956 81056 6012
rect 81056 5956 81112 6012
rect 81112 5956 81116 6012
rect 81052 5952 81116 5956
rect 4012 5468 4076 5472
rect 4012 5412 4016 5468
rect 4016 5412 4072 5468
rect 4072 5412 4076 5468
rect 4012 5408 4076 5412
rect 4092 5468 4156 5472
rect 4092 5412 4096 5468
rect 4096 5412 4152 5468
rect 4152 5412 4156 5468
rect 4092 5408 4156 5412
rect 4172 5468 4236 5472
rect 4172 5412 4176 5468
rect 4176 5412 4232 5468
rect 4232 5412 4236 5468
rect 4172 5408 4236 5412
rect 4252 5468 4316 5472
rect 4252 5412 4256 5468
rect 4256 5412 4312 5468
rect 4312 5412 4316 5468
rect 4252 5408 4316 5412
rect 34732 5468 34796 5472
rect 34732 5412 34736 5468
rect 34736 5412 34792 5468
rect 34792 5412 34796 5468
rect 34732 5408 34796 5412
rect 34812 5468 34876 5472
rect 34812 5412 34816 5468
rect 34816 5412 34872 5468
rect 34872 5412 34876 5468
rect 34812 5408 34876 5412
rect 34892 5468 34956 5472
rect 34892 5412 34896 5468
rect 34896 5412 34952 5468
rect 34952 5412 34956 5468
rect 34892 5408 34956 5412
rect 34972 5468 35036 5472
rect 34972 5412 34976 5468
rect 34976 5412 35032 5468
rect 35032 5412 35036 5468
rect 34972 5408 35036 5412
rect 65452 5468 65516 5472
rect 65452 5412 65456 5468
rect 65456 5412 65512 5468
rect 65512 5412 65516 5468
rect 65452 5408 65516 5412
rect 65532 5468 65596 5472
rect 65532 5412 65536 5468
rect 65536 5412 65592 5468
rect 65592 5412 65596 5468
rect 65532 5408 65596 5412
rect 65612 5468 65676 5472
rect 65612 5412 65616 5468
rect 65616 5412 65672 5468
rect 65672 5412 65676 5468
rect 65612 5408 65676 5412
rect 65692 5468 65756 5472
rect 65692 5412 65696 5468
rect 65696 5412 65752 5468
rect 65752 5412 65756 5468
rect 65692 5408 65756 5412
rect 96172 5468 96236 5472
rect 96172 5412 96176 5468
rect 96176 5412 96232 5468
rect 96232 5412 96236 5468
rect 96172 5408 96236 5412
rect 96252 5468 96316 5472
rect 96252 5412 96256 5468
rect 96256 5412 96312 5468
rect 96312 5412 96316 5468
rect 96252 5408 96316 5412
rect 96332 5468 96396 5472
rect 96332 5412 96336 5468
rect 96336 5412 96392 5468
rect 96392 5412 96396 5468
rect 96332 5408 96396 5412
rect 96412 5468 96476 5472
rect 96412 5412 96416 5468
rect 96416 5412 96472 5468
rect 96472 5412 96476 5468
rect 96412 5408 96476 5412
rect 19372 4924 19436 4928
rect 19372 4868 19376 4924
rect 19376 4868 19432 4924
rect 19432 4868 19436 4924
rect 19372 4864 19436 4868
rect 19452 4924 19516 4928
rect 19452 4868 19456 4924
rect 19456 4868 19512 4924
rect 19512 4868 19516 4924
rect 19452 4864 19516 4868
rect 19532 4924 19596 4928
rect 19532 4868 19536 4924
rect 19536 4868 19592 4924
rect 19592 4868 19596 4924
rect 19532 4864 19596 4868
rect 19612 4924 19676 4928
rect 19612 4868 19616 4924
rect 19616 4868 19672 4924
rect 19672 4868 19676 4924
rect 19612 4864 19676 4868
rect 50092 4924 50156 4928
rect 50092 4868 50096 4924
rect 50096 4868 50152 4924
rect 50152 4868 50156 4924
rect 50092 4864 50156 4868
rect 50172 4924 50236 4928
rect 50172 4868 50176 4924
rect 50176 4868 50232 4924
rect 50232 4868 50236 4924
rect 50172 4864 50236 4868
rect 50252 4924 50316 4928
rect 50252 4868 50256 4924
rect 50256 4868 50312 4924
rect 50312 4868 50316 4924
rect 50252 4864 50316 4868
rect 50332 4924 50396 4928
rect 50332 4868 50336 4924
rect 50336 4868 50392 4924
rect 50392 4868 50396 4924
rect 50332 4864 50396 4868
rect 80812 4924 80876 4928
rect 80812 4868 80816 4924
rect 80816 4868 80872 4924
rect 80872 4868 80876 4924
rect 80812 4864 80876 4868
rect 80892 4924 80956 4928
rect 80892 4868 80896 4924
rect 80896 4868 80952 4924
rect 80952 4868 80956 4924
rect 80892 4864 80956 4868
rect 80972 4924 81036 4928
rect 80972 4868 80976 4924
rect 80976 4868 81032 4924
rect 81032 4868 81036 4924
rect 80972 4864 81036 4868
rect 81052 4924 81116 4928
rect 81052 4868 81056 4924
rect 81056 4868 81112 4924
rect 81112 4868 81116 4924
rect 81052 4864 81116 4868
rect 4012 4380 4076 4384
rect 4012 4324 4016 4380
rect 4016 4324 4072 4380
rect 4072 4324 4076 4380
rect 4012 4320 4076 4324
rect 4092 4380 4156 4384
rect 4092 4324 4096 4380
rect 4096 4324 4152 4380
rect 4152 4324 4156 4380
rect 4092 4320 4156 4324
rect 4172 4380 4236 4384
rect 4172 4324 4176 4380
rect 4176 4324 4232 4380
rect 4232 4324 4236 4380
rect 4172 4320 4236 4324
rect 4252 4380 4316 4384
rect 4252 4324 4256 4380
rect 4256 4324 4312 4380
rect 4312 4324 4316 4380
rect 4252 4320 4316 4324
rect 34732 4380 34796 4384
rect 34732 4324 34736 4380
rect 34736 4324 34792 4380
rect 34792 4324 34796 4380
rect 34732 4320 34796 4324
rect 34812 4380 34876 4384
rect 34812 4324 34816 4380
rect 34816 4324 34872 4380
rect 34872 4324 34876 4380
rect 34812 4320 34876 4324
rect 34892 4380 34956 4384
rect 34892 4324 34896 4380
rect 34896 4324 34952 4380
rect 34952 4324 34956 4380
rect 34892 4320 34956 4324
rect 34972 4380 35036 4384
rect 34972 4324 34976 4380
rect 34976 4324 35032 4380
rect 35032 4324 35036 4380
rect 34972 4320 35036 4324
rect 65452 4380 65516 4384
rect 65452 4324 65456 4380
rect 65456 4324 65512 4380
rect 65512 4324 65516 4380
rect 65452 4320 65516 4324
rect 65532 4380 65596 4384
rect 65532 4324 65536 4380
rect 65536 4324 65592 4380
rect 65592 4324 65596 4380
rect 65532 4320 65596 4324
rect 65612 4380 65676 4384
rect 65612 4324 65616 4380
rect 65616 4324 65672 4380
rect 65672 4324 65676 4380
rect 65612 4320 65676 4324
rect 65692 4380 65756 4384
rect 65692 4324 65696 4380
rect 65696 4324 65752 4380
rect 65752 4324 65756 4380
rect 65692 4320 65756 4324
rect 96172 4380 96236 4384
rect 96172 4324 96176 4380
rect 96176 4324 96232 4380
rect 96232 4324 96236 4380
rect 96172 4320 96236 4324
rect 96252 4380 96316 4384
rect 96252 4324 96256 4380
rect 96256 4324 96312 4380
rect 96312 4324 96316 4380
rect 96252 4320 96316 4324
rect 96332 4380 96396 4384
rect 96332 4324 96336 4380
rect 96336 4324 96392 4380
rect 96392 4324 96396 4380
rect 96332 4320 96396 4324
rect 96412 4380 96476 4384
rect 96412 4324 96416 4380
rect 96416 4324 96472 4380
rect 96472 4324 96476 4380
rect 96412 4320 96476 4324
rect 19372 3836 19436 3840
rect 19372 3780 19376 3836
rect 19376 3780 19432 3836
rect 19432 3780 19436 3836
rect 19372 3776 19436 3780
rect 19452 3836 19516 3840
rect 19452 3780 19456 3836
rect 19456 3780 19512 3836
rect 19512 3780 19516 3836
rect 19452 3776 19516 3780
rect 19532 3836 19596 3840
rect 19532 3780 19536 3836
rect 19536 3780 19592 3836
rect 19592 3780 19596 3836
rect 19532 3776 19596 3780
rect 19612 3836 19676 3840
rect 19612 3780 19616 3836
rect 19616 3780 19672 3836
rect 19672 3780 19676 3836
rect 19612 3776 19676 3780
rect 50092 3836 50156 3840
rect 50092 3780 50096 3836
rect 50096 3780 50152 3836
rect 50152 3780 50156 3836
rect 50092 3776 50156 3780
rect 50172 3836 50236 3840
rect 50172 3780 50176 3836
rect 50176 3780 50232 3836
rect 50232 3780 50236 3836
rect 50172 3776 50236 3780
rect 50252 3836 50316 3840
rect 50252 3780 50256 3836
rect 50256 3780 50312 3836
rect 50312 3780 50316 3836
rect 50252 3776 50316 3780
rect 50332 3836 50396 3840
rect 50332 3780 50336 3836
rect 50336 3780 50392 3836
rect 50392 3780 50396 3836
rect 50332 3776 50396 3780
rect 80812 3836 80876 3840
rect 80812 3780 80816 3836
rect 80816 3780 80872 3836
rect 80872 3780 80876 3836
rect 80812 3776 80876 3780
rect 80892 3836 80956 3840
rect 80892 3780 80896 3836
rect 80896 3780 80952 3836
rect 80952 3780 80956 3836
rect 80892 3776 80956 3780
rect 80972 3836 81036 3840
rect 80972 3780 80976 3836
rect 80976 3780 81032 3836
rect 81032 3780 81036 3836
rect 80972 3776 81036 3780
rect 81052 3836 81116 3840
rect 81052 3780 81056 3836
rect 81056 3780 81112 3836
rect 81112 3780 81116 3836
rect 81052 3776 81116 3780
rect 4012 3292 4076 3296
rect 4012 3236 4016 3292
rect 4016 3236 4072 3292
rect 4072 3236 4076 3292
rect 4012 3232 4076 3236
rect 4092 3292 4156 3296
rect 4092 3236 4096 3292
rect 4096 3236 4152 3292
rect 4152 3236 4156 3292
rect 4092 3232 4156 3236
rect 4172 3292 4236 3296
rect 4172 3236 4176 3292
rect 4176 3236 4232 3292
rect 4232 3236 4236 3292
rect 4172 3232 4236 3236
rect 4252 3292 4316 3296
rect 4252 3236 4256 3292
rect 4256 3236 4312 3292
rect 4312 3236 4316 3292
rect 4252 3232 4316 3236
rect 34732 3292 34796 3296
rect 34732 3236 34736 3292
rect 34736 3236 34792 3292
rect 34792 3236 34796 3292
rect 34732 3232 34796 3236
rect 34812 3292 34876 3296
rect 34812 3236 34816 3292
rect 34816 3236 34872 3292
rect 34872 3236 34876 3292
rect 34812 3232 34876 3236
rect 34892 3292 34956 3296
rect 34892 3236 34896 3292
rect 34896 3236 34952 3292
rect 34952 3236 34956 3292
rect 34892 3232 34956 3236
rect 34972 3292 35036 3296
rect 34972 3236 34976 3292
rect 34976 3236 35032 3292
rect 35032 3236 35036 3292
rect 34972 3232 35036 3236
rect 65452 3292 65516 3296
rect 65452 3236 65456 3292
rect 65456 3236 65512 3292
rect 65512 3236 65516 3292
rect 65452 3232 65516 3236
rect 65532 3292 65596 3296
rect 65532 3236 65536 3292
rect 65536 3236 65592 3292
rect 65592 3236 65596 3292
rect 65532 3232 65596 3236
rect 65612 3292 65676 3296
rect 65612 3236 65616 3292
rect 65616 3236 65672 3292
rect 65672 3236 65676 3292
rect 65612 3232 65676 3236
rect 65692 3292 65756 3296
rect 65692 3236 65696 3292
rect 65696 3236 65752 3292
rect 65752 3236 65756 3292
rect 65692 3232 65756 3236
rect 96172 3292 96236 3296
rect 96172 3236 96176 3292
rect 96176 3236 96232 3292
rect 96232 3236 96236 3292
rect 96172 3232 96236 3236
rect 96252 3292 96316 3296
rect 96252 3236 96256 3292
rect 96256 3236 96312 3292
rect 96312 3236 96316 3292
rect 96252 3232 96316 3236
rect 96332 3292 96396 3296
rect 96332 3236 96336 3292
rect 96336 3236 96392 3292
rect 96392 3236 96396 3292
rect 96332 3232 96396 3236
rect 96412 3292 96476 3296
rect 96412 3236 96416 3292
rect 96416 3236 96472 3292
rect 96472 3236 96476 3292
rect 96412 3232 96476 3236
rect 19372 2748 19436 2752
rect 19372 2692 19376 2748
rect 19376 2692 19432 2748
rect 19432 2692 19436 2748
rect 19372 2688 19436 2692
rect 19452 2748 19516 2752
rect 19452 2692 19456 2748
rect 19456 2692 19512 2748
rect 19512 2692 19516 2748
rect 19452 2688 19516 2692
rect 19532 2748 19596 2752
rect 19532 2692 19536 2748
rect 19536 2692 19592 2748
rect 19592 2692 19596 2748
rect 19532 2688 19596 2692
rect 19612 2748 19676 2752
rect 19612 2692 19616 2748
rect 19616 2692 19672 2748
rect 19672 2692 19676 2748
rect 19612 2688 19676 2692
rect 50092 2748 50156 2752
rect 50092 2692 50096 2748
rect 50096 2692 50152 2748
rect 50152 2692 50156 2748
rect 50092 2688 50156 2692
rect 50172 2748 50236 2752
rect 50172 2692 50176 2748
rect 50176 2692 50232 2748
rect 50232 2692 50236 2748
rect 50172 2688 50236 2692
rect 50252 2748 50316 2752
rect 50252 2692 50256 2748
rect 50256 2692 50312 2748
rect 50312 2692 50316 2748
rect 50252 2688 50316 2692
rect 50332 2748 50396 2752
rect 50332 2692 50336 2748
rect 50336 2692 50392 2748
rect 50392 2692 50396 2748
rect 50332 2688 50396 2692
rect 80812 2748 80876 2752
rect 80812 2692 80816 2748
rect 80816 2692 80872 2748
rect 80872 2692 80876 2748
rect 80812 2688 80876 2692
rect 80892 2748 80956 2752
rect 80892 2692 80896 2748
rect 80896 2692 80952 2748
rect 80952 2692 80956 2748
rect 80892 2688 80956 2692
rect 80972 2748 81036 2752
rect 80972 2692 80976 2748
rect 80976 2692 81032 2748
rect 81032 2692 81036 2748
rect 80972 2688 81036 2692
rect 81052 2748 81116 2752
rect 81052 2692 81056 2748
rect 81056 2692 81112 2748
rect 81112 2692 81116 2748
rect 81052 2688 81116 2692
rect 4012 2204 4076 2208
rect 4012 2148 4016 2204
rect 4016 2148 4072 2204
rect 4072 2148 4076 2204
rect 4012 2144 4076 2148
rect 4092 2204 4156 2208
rect 4092 2148 4096 2204
rect 4096 2148 4152 2204
rect 4152 2148 4156 2204
rect 4092 2144 4156 2148
rect 4172 2204 4236 2208
rect 4172 2148 4176 2204
rect 4176 2148 4232 2204
rect 4232 2148 4236 2204
rect 4172 2144 4236 2148
rect 4252 2204 4316 2208
rect 4252 2148 4256 2204
rect 4256 2148 4312 2204
rect 4312 2148 4316 2204
rect 4252 2144 4316 2148
rect 34732 2204 34796 2208
rect 34732 2148 34736 2204
rect 34736 2148 34792 2204
rect 34792 2148 34796 2204
rect 34732 2144 34796 2148
rect 34812 2204 34876 2208
rect 34812 2148 34816 2204
rect 34816 2148 34872 2204
rect 34872 2148 34876 2204
rect 34812 2144 34876 2148
rect 34892 2204 34956 2208
rect 34892 2148 34896 2204
rect 34896 2148 34952 2204
rect 34952 2148 34956 2204
rect 34892 2144 34956 2148
rect 34972 2204 35036 2208
rect 34972 2148 34976 2204
rect 34976 2148 35032 2204
rect 35032 2148 35036 2204
rect 34972 2144 35036 2148
rect 65452 2204 65516 2208
rect 65452 2148 65456 2204
rect 65456 2148 65512 2204
rect 65512 2148 65516 2204
rect 65452 2144 65516 2148
rect 65532 2204 65596 2208
rect 65532 2148 65536 2204
rect 65536 2148 65592 2204
rect 65592 2148 65596 2204
rect 65532 2144 65596 2148
rect 65612 2204 65676 2208
rect 65612 2148 65616 2204
rect 65616 2148 65672 2204
rect 65672 2148 65676 2204
rect 65612 2144 65676 2148
rect 65692 2204 65756 2208
rect 65692 2148 65696 2204
rect 65696 2148 65752 2204
rect 65752 2148 65756 2204
rect 65692 2144 65756 2148
rect 96172 2204 96236 2208
rect 96172 2148 96176 2204
rect 96176 2148 96232 2204
rect 96232 2148 96236 2204
rect 96172 2144 96236 2148
rect 96252 2204 96316 2208
rect 96252 2148 96256 2204
rect 96256 2148 96312 2204
rect 96312 2148 96316 2204
rect 96252 2144 96316 2148
rect 96332 2204 96396 2208
rect 96332 2148 96336 2204
rect 96336 2148 96392 2204
rect 96392 2148 96396 2204
rect 96332 2144 96396 2148
rect 96412 2204 96476 2208
rect 96412 2148 96416 2204
rect 96416 2148 96472 2204
rect 96472 2148 96476 2204
rect 96412 2144 96476 2148
rect 19372 1660 19436 1664
rect 19372 1604 19376 1660
rect 19376 1604 19432 1660
rect 19432 1604 19436 1660
rect 19372 1600 19436 1604
rect 19452 1660 19516 1664
rect 19452 1604 19456 1660
rect 19456 1604 19512 1660
rect 19512 1604 19516 1660
rect 19452 1600 19516 1604
rect 19532 1660 19596 1664
rect 19532 1604 19536 1660
rect 19536 1604 19592 1660
rect 19592 1604 19596 1660
rect 19532 1600 19596 1604
rect 19612 1660 19676 1664
rect 19612 1604 19616 1660
rect 19616 1604 19672 1660
rect 19672 1604 19676 1660
rect 19612 1600 19676 1604
rect 50092 1660 50156 1664
rect 50092 1604 50096 1660
rect 50096 1604 50152 1660
rect 50152 1604 50156 1660
rect 50092 1600 50156 1604
rect 50172 1660 50236 1664
rect 50172 1604 50176 1660
rect 50176 1604 50232 1660
rect 50232 1604 50236 1660
rect 50172 1600 50236 1604
rect 50252 1660 50316 1664
rect 50252 1604 50256 1660
rect 50256 1604 50312 1660
rect 50312 1604 50316 1660
rect 50252 1600 50316 1604
rect 50332 1660 50396 1664
rect 50332 1604 50336 1660
rect 50336 1604 50392 1660
rect 50392 1604 50396 1660
rect 50332 1600 50396 1604
rect 80812 1660 80876 1664
rect 80812 1604 80816 1660
rect 80816 1604 80872 1660
rect 80872 1604 80876 1660
rect 80812 1600 80876 1604
rect 80892 1660 80956 1664
rect 80892 1604 80896 1660
rect 80896 1604 80952 1660
rect 80952 1604 80956 1660
rect 80892 1600 80956 1604
rect 80972 1660 81036 1664
rect 80972 1604 80976 1660
rect 80976 1604 81032 1660
rect 81032 1604 81036 1660
rect 80972 1600 81036 1604
rect 81052 1660 81116 1664
rect 81052 1604 81056 1660
rect 81056 1604 81112 1660
rect 81112 1604 81116 1660
rect 81052 1600 81116 1604
rect 4012 1116 4076 1120
rect 4012 1060 4016 1116
rect 4016 1060 4072 1116
rect 4072 1060 4076 1116
rect 4012 1056 4076 1060
rect 4092 1116 4156 1120
rect 4092 1060 4096 1116
rect 4096 1060 4152 1116
rect 4152 1060 4156 1116
rect 4092 1056 4156 1060
rect 4172 1116 4236 1120
rect 4172 1060 4176 1116
rect 4176 1060 4232 1116
rect 4232 1060 4236 1116
rect 4172 1056 4236 1060
rect 4252 1116 4316 1120
rect 4252 1060 4256 1116
rect 4256 1060 4312 1116
rect 4312 1060 4316 1116
rect 4252 1056 4316 1060
rect 34732 1116 34796 1120
rect 34732 1060 34736 1116
rect 34736 1060 34792 1116
rect 34792 1060 34796 1116
rect 34732 1056 34796 1060
rect 34812 1116 34876 1120
rect 34812 1060 34816 1116
rect 34816 1060 34872 1116
rect 34872 1060 34876 1116
rect 34812 1056 34876 1060
rect 34892 1116 34956 1120
rect 34892 1060 34896 1116
rect 34896 1060 34952 1116
rect 34952 1060 34956 1116
rect 34892 1056 34956 1060
rect 34972 1116 35036 1120
rect 34972 1060 34976 1116
rect 34976 1060 35032 1116
rect 35032 1060 35036 1116
rect 34972 1056 35036 1060
rect 65452 1116 65516 1120
rect 65452 1060 65456 1116
rect 65456 1060 65512 1116
rect 65512 1060 65516 1116
rect 65452 1056 65516 1060
rect 65532 1116 65596 1120
rect 65532 1060 65536 1116
rect 65536 1060 65592 1116
rect 65592 1060 65596 1116
rect 65532 1056 65596 1060
rect 65612 1116 65676 1120
rect 65612 1060 65616 1116
rect 65616 1060 65672 1116
rect 65672 1060 65676 1116
rect 65612 1056 65676 1060
rect 65692 1116 65756 1120
rect 65692 1060 65696 1116
rect 65696 1060 65752 1116
rect 65752 1060 65756 1116
rect 65692 1056 65756 1060
rect 96172 1116 96236 1120
rect 96172 1060 96176 1116
rect 96176 1060 96232 1116
rect 96232 1060 96236 1116
rect 96172 1056 96236 1060
rect 96252 1116 96316 1120
rect 96252 1060 96256 1116
rect 96256 1060 96312 1116
rect 96312 1060 96316 1116
rect 96252 1056 96316 1060
rect 96332 1116 96396 1120
rect 96332 1060 96336 1116
rect 96336 1060 96392 1116
rect 96392 1060 96396 1116
rect 96332 1056 96396 1060
rect 96412 1116 96476 1120
rect 96412 1060 96416 1116
rect 96416 1060 96472 1116
rect 96472 1060 96476 1116
rect 96412 1056 96476 1060
<< metal4 >>
rect 4004 7648 4324 7664
rect 4004 7584 4012 7648
rect 4076 7584 4092 7648
rect 4156 7584 4172 7648
rect 4236 7584 4252 7648
rect 4316 7584 4324 7648
rect 4004 6560 4324 7584
rect 4004 6496 4012 6560
rect 4076 6496 4092 6560
rect 4156 6496 4172 6560
rect 4236 6496 4252 6560
rect 4316 6496 4324 6560
rect 4004 5472 4324 6496
rect 4004 5408 4012 5472
rect 4076 5408 4092 5472
rect 4156 5408 4172 5472
rect 4236 5408 4252 5472
rect 4316 5408 4324 5472
rect 4004 4384 4324 5408
rect 4004 4320 4012 4384
rect 4076 4320 4092 4384
rect 4156 4320 4172 4384
rect 4236 4320 4252 4384
rect 4316 4320 4324 4384
rect 4004 3296 4324 4320
rect 4004 3232 4012 3296
rect 4076 3232 4092 3296
rect 4156 3232 4172 3296
rect 4236 3232 4252 3296
rect 4316 3232 4324 3296
rect 4004 2208 4324 3232
rect 4004 2144 4012 2208
rect 4076 2144 4092 2208
rect 4156 2144 4172 2208
rect 4236 2144 4252 2208
rect 4316 2144 4324 2208
rect 4004 1120 4324 2144
rect 4004 1056 4012 1120
rect 4076 1056 4092 1120
rect 4156 1056 4172 1120
rect 4236 1056 4252 1120
rect 4316 1056 4324 1120
rect 4004 1040 4324 1056
rect 19364 7104 19684 7664
rect 19364 7040 19372 7104
rect 19436 7040 19452 7104
rect 19516 7040 19532 7104
rect 19596 7040 19612 7104
rect 19676 7040 19684 7104
rect 19364 6016 19684 7040
rect 19364 5952 19372 6016
rect 19436 5952 19452 6016
rect 19516 5952 19532 6016
rect 19596 5952 19612 6016
rect 19676 5952 19684 6016
rect 19364 4928 19684 5952
rect 19364 4864 19372 4928
rect 19436 4864 19452 4928
rect 19516 4864 19532 4928
rect 19596 4864 19612 4928
rect 19676 4864 19684 4928
rect 19364 3840 19684 4864
rect 19364 3776 19372 3840
rect 19436 3776 19452 3840
rect 19516 3776 19532 3840
rect 19596 3776 19612 3840
rect 19676 3776 19684 3840
rect 19364 2752 19684 3776
rect 19364 2688 19372 2752
rect 19436 2688 19452 2752
rect 19516 2688 19532 2752
rect 19596 2688 19612 2752
rect 19676 2688 19684 2752
rect 19364 1664 19684 2688
rect 19364 1600 19372 1664
rect 19436 1600 19452 1664
rect 19516 1600 19532 1664
rect 19596 1600 19612 1664
rect 19676 1600 19684 1664
rect 19364 1040 19684 1600
rect 34724 7648 35044 7664
rect 34724 7584 34732 7648
rect 34796 7584 34812 7648
rect 34876 7584 34892 7648
rect 34956 7584 34972 7648
rect 35036 7584 35044 7648
rect 34724 6560 35044 7584
rect 34724 6496 34732 6560
rect 34796 6496 34812 6560
rect 34876 6496 34892 6560
rect 34956 6496 34972 6560
rect 35036 6496 35044 6560
rect 34724 5472 35044 6496
rect 34724 5408 34732 5472
rect 34796 5408 34812 5472
rect 34876 5408 34892 5472
rect 34956 5408 34972 5472
rect 35036 5408 35044 5472
rect 34724 4384 35044 5408
rect 34724 4320 34732 4384
rect 34796 4320 34812 4384
rect 34876 4320 34892 4384
rect 34956 4320 34972 4384
rect 35036 4320 35044 4384
rect 34724 3296 35044 4320
rect 34724 3232 34732 3296
rect 34796 3232 34812 3296
rect 34876 3232 34892 3296
rect 34956 3232 34972 3296
rect 35036 3232 35044 3296
rect 34724 2208 35044 3232
rect 34724 2144 34732 2208
rect 34796 2144 34812 2208
rect 34876 2144 34892 2208
rect 34956 2144 34972 2208
rect 35036 2144 35044 2208
rect 34724 1120 35044 2144
rect 34724 1056 34732 1120
rect 34796 1056 34812 1120
rect 34876 1056 34892 1120
rect 34956 1056 34972 1120
rect 35036 1056 35044 1120
rect 34724 1040 35044 1056
rect 50084 7104 50404 7664
rect 50084 7040 50092 7104
rect 50156 7040 50172 7104
rect 50236 7040 50252 7104
rect 50316 7040 50332 7104
rect 50396 7040 50404 7104
rect 50084 6016 50404 7040
rect 50084 5952 50092 6016
rect 50156 5952 50172 6016
rect 50236 5952 50252 6016
rect 50316 5952 50332 6016
rect 50396 5952 50404 6016
rect 50084 4928 50404 5952
rect 50084 4864 50092 4928
rect 50156 4864 50172 4928
rect 50236 4864 50252 4928
rect 50316 4864 50332 4928
rect 50396 4864 50404 4928
rect 50084 3840 50404 4864
rect 50084 3776 50092 3840
rect 50156 3776 50172 3840
rect 50236 3776 50252 3840
rect 50316 3776 50332 3840
rect 50396 3776 50404 3840
rect 50084 2752 50404 3776
rect 50084 2688 50092 2752
rect 50156 2688 50172 2752
rect 50236 2688 50252 2752
rect 50316 2688 50332 2752
rect 50396 2688 50404 2752
rect 50084 1664 50404 2688
rect 50084 1600 50092 1664
rect 50156 1600 50172 1664
rect 50236 1600 50252 1664
rect 50316 1600 50332 1664
rect 50396 1600 50404 1664
rect 50084 1040 50404 1600
rect 65444 7648 65764 7664
rect 65444 7584 65452 7648
rect 65516 7584 65532 7648
rect 65596 7584 65612 7648
rect 65676 7584 65692 7648
rect 65756 7584 65764 7648
rect 65444 6560 65764 7584
rect 65444 6496 65452 6560
rect 65516 6496 65532 6560
rect 65596 6496 65612 6560
rect 65676 6496 65692 6560
rect 65756 6496 65764 6560
rect 65444 5472 65764 6496
rect 65444 5408 65452 5472
rect 65516 5408 65532 5472
rect 65596 5408 65612 5472
rect 65676 5408 65692 5472
rect 65756 5408 65764 5472
rect 65444 4384 65764 5408
rect 65444 4320 65452 4384
rect 65516 4320 65532 4384
rect 65596 4320 65612 4384
rect 65676 4320 65692 4384
rect 65756 4320 65764 4384
rect 65444 3296 65764 4320
rect 65444 3232 65452 3296
rect 65516 3232 65532 3296
rect 65596 3232 65612 3296
rect 65676 3232 65692 3296
rect 65756 3232 65764 3296
rect 65444 2208 65764 3232
rect 65444 2144 65452 2208
rect 65516 2144 65532 2208
rect 65596 2144 65612 2208
rect 65676 2144 65692 2208
rect 65756 2144 65764 2208
rect 65444 1120 65764 2144
rect 65444 1056 65452 1120
rect 65516 1056 65532 1120
rect 65596 1056 65612 1120
rect 65676 1056 65692 1120
rect 65756 1056 65764 1120
rect 65444 1040 65764 1056
rect 80804 7104 81124 7664
rect 80804 7040 80812 7104
rect 80876 7040 80892 7104
rect 80956 7040 80972 7104
rect 81036 7040 81052 7104
rect 81116 7040 81124 7104
rect 80804 6016 81124 7040
rect 80804 5952 80812 6016
rect 80876 5952 80892 6016
rect 80956 5952 80972 6016
rect 81036 5952 81052 6016
rect 81116 5952 81124 6016
rect 80804 4928 81124 5952
rect 80804 4864 80812 4928
rect 80876 4864 80892 4928
rect 80956 4864 80972 4928
rect 81036 4864 81052 4928
rect 81116 4864 81124 4928
rect 80804 3840 81124 4864
rect 80804 3776 80812 3840
rect 80876 3776 80892 3840
rect 80956 3776 80972 3840
rect 81036 3776 81052 3840
rect 81116 3776 81124 3840
rect 80804 2752 81124 3776
rect 80804 2688 80812 2752
rect 80876 2688 80892 2752
rect 80956 2688 80972 2752
rect 81036 2688 81052 2752
rect 81116 2688 81124 2752
rect 80804 1664 81124 2688
rect 80804 1600 80812 1664
rect 80876 1600 80892 1664
rect 80956 1600 80972 1664
rect 81036 1600 81052 1664
rect 81116 1600 81124 1664
rect 80804 1040 81124 1600
rect 96164 7648 96484 7664
rect 96164 7584 96172 7648
rect 96236 7584 96252 7648
rect 96316 7584 96332 7648
rect 96396 7584 96412 7648
rect 96476 7584 96484 7648
rect 96164 6560 96484 7584
rect 96164 6496 96172 6560
rect 96236 6496 96252 6560
rect 96316 6496 96332 6560
rect 96396 6496 96412 6560
rect 96476 6496 96484 6560
rect 96164 5472 96484 6496
rect 96164 5408 96172 5472
rect 96236 5408 96252 5472
rect 96316 5408 96332 5472
rect 96396 5408 96412 5472
rect 96476 5408 96484 5472
rect 96164 4384 96484 5408
rect 96164 4320 96172 4384
rect 96236 4320 96252 4384
rect 96316 4320 96332 4384
rect 96396 4320 96412 4384
rect 96476 4320 96484 4384
rect 96164 3296 96484 4320
rect 96164 3232 96172 3296
rect 96236 3232 96252 3296
rect 96316 3232 96332 3296
rect 96396 3232 96412 3296
rect 96476 3232 96484 3296
rect 96164 2208 96484 3232
rect 96164 2144 96172 2208
rect 96236 2144 96252 2208
rect 96316 2144 96332 2208
rect 96396 2144 96412 2208
rect 96476 2144 96484 2208
rect 96164 1120 96484 2144
rect 96164 1056 96172 1120
rect 96236 1056 96252 1120
rect 96316 1056 96332 1120
rect 96396 1056 96412 1120
rect 96476 1056 96484 1120
rect 96164 1040 96484 1056
use sky130_fd_sc_hd__dfxtp_4  dff2_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 1104 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 2852 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  dff1_0
timestamp 1607194113
transform 1 0 1104 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_0
timestamp 1607194113
transform 1 0 2852 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 2944 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_1
timestamp 1607194113
transform 1 0 3220 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  decap1_0
timestamp 1607194113
transform 1 0 2944 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_1
timestamp 1607194113
transform 1 0 3220 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_1
timestamp 1607194113
transform 1 0 4968 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_1
timestamp 1607194113
transform 1 0 5060 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_2
timestamp 1607194113
transform 1 0 5336 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_1
timestamp 1607194113
transform 1 0 4968 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_1
timestamp 1607194113
transform 1 0 5060 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_2
timestamp 1607194113
transform 1 0 5336 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_2
timestamp 1607194113
transform 1 0 7084 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_2
timestamp 1607194113
transform 1 0 7176 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_3
timestamp 1607194113
transform 1 0 7452 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_2
timestamp 1607194113
transform 1 0 7084 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_2
timestamp 1607194113
transform 1 0 7176 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_3
timestamp 1607194113
transform 1 0 7452 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_3
timestamp 1607194113
transform 1 0 9200 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_3
timestamp 1607194113
transform 1 0 9292 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_4
timestamp 1607194113
transform 1 0 9568 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_3
timestamp 1607194113
transform 1 0 9200 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_3
timestamp 1607194113
transform 1 0 9292 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_4
timestamp 1607194113
transform 1 0 9568 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_4
timestamp 1607194113
transform 1 0 11316 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_4
timestamp 1607194113
transform 1 0 11408 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_5
timestamp 1607194113
transform 1 0 11684 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_4
timestamp 1607194113
transform 1 0 11316 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_4
timestamp 1607194113
transform 1 0 11408 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_5
timestamp 1607194113
transform 1 0 11684 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_5
timestamp 1607194113
transform 1 0 13432 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_5
timestamp 1607194113
transform 1 0 13524 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_6
timestamp 1607194113
transform 1 0 13800 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_5
timestamp 1607194113
transform 1 0 13432 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_5
timestamp 1607194113
transform 1 0 13524 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_6
timestamp 1607194113
transform 1 0 13800 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_6
timestamp 1607194113
transform 1 0 15548 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_6
timestamp 1607194113
transform 1 0 15640 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_6
timestamp 1607194113
transform 1 0 15548 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_6
timestamp 1607194113
transform 1 0 15640 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_7
timestamp 1607194113
transform 1 0 15916 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  dff1_7
timestamp 1607194113
transform 1 0 15916 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_7
timestamp 1607194113
transform 1 0 17664 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_7
timestamp 1607194113
transform 1 0 17756 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_8
timestamp 1607194113
transform 1 0 18032 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_7
timestamp 1607194113
transform 1 0 17664 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_7
timestamp 1607194113
transform 1 0 17756 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_8
timestamp 1607194113
transform 1 0 18032 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_8
timestamp 1607194113
transform 1 0 19780 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_8
timestamp 1607194113
transform 1 0 19872 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_9
timestamp 1607194113
transform 1 0 20148 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_8
timestamp 1607194113
transform 1 0 19780 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_8
timestamp 1607194113
transform 1 0 19872 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_9
timestamp 1607194113
transform 1 0 20148 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_9
timestamp 1607194113
transform 1 0 21896 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_9
timestamp 1607194113
transform 1 0 21988 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_10
timestamp 1607194113
transform 1 0 22264 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_9
timestamp 1607194113
transform 1 0 21896 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_9
timestamp 1607194113
transform 1 0 21988 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_10
timestamp 1607194113
transform 1 0 22264 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_10
timestamp 1607194113
transform 1 0 24012 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_10
timestamp 1607194113
transform 1 0 24104 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_11
timestamp 1607194113
transform 1 0 24380 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_10
timestamp 1607194113
transform 1 0 24012 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_10
timestamp 1607194113
transform 1 0 24104 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_11
timestamp 1607194113
transform 1 0 24380 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_11
timestamp 1607194113
transform 1 0 26128 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_11
timestamp 1607194113
transform 1 0 26220 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_12
timestamp 1607194113
transform 1 0 26496 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_11
timestamp 1607194113
transform 1 0 26128 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_11
timestamp 1607194113
transform 1 0 26220 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_12
timestamp 1607194113
transform 1 0 26496 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_12
timestamp 1607194113
transform 1 0 28244 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_12
timestamp 1607194113
transform 1 0 28336 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_12
timestamp 1607194113
transform 1 0 28244 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_12
timestamp 1607194113
transform 1 0 28336 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_13
timestamp 1607194113
transform 1 0 28612 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  dff1_13
timestamp 1607194113
transform 1 0 28612 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_13
timestamp 1607194113
transform 1 0 30360 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_13
timestamp 1607194113
transform 1 0 30452 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_14
timestamp 1607194113
transform 1 0 30728 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_13
timestamp 1607194113
transform 1 0 30360 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_13
timestamp 1607194113
transform 1 0 30452 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_14
timestamp 1607194113
transform 1 0 30728 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_14
timestamp 1607194113
transform 1 0 32476 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_14
timestamp 1607194113
transform 1 0 32568 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_15
timestamp 1607194113
transform 1 0 32844 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_14
timestamp 1607194113
transform 1 0 32476 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_14
timestamp 1607194113
transform 1 0 32568 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_15
timestamp 1607194113
transform 1 0 32844 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_15
timestamp 1607194113
transform 1 0 34592 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_15
timestamp 1607194113
transform 1 0 34684 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_16
timestamp 1607194113
transform 1 0 34960 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_15
timestamp 1607194113
transform 1 0 34592 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_15
timestamp 1607194113
transform 1 0 34684 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_16
timestamp 1607194113
transform 1 0 34960 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_16
timestamp 1607194113
transform 1 0 36708 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_16
timestamp 1607194113
transform 1 0 36800 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_17
timestamp 1607194113
transform 1 0 37076 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_16
timestamp 1607194113
transform 1 0 36708 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_16
timestamp 1607194113
transform 1 0 36800 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_17
timestamp 1607194113
transform 1 0 37076 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_17
timestamp 1607194113
transform 1 0 38824 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_17
timestamp 1607194113
transform 1 0 38916 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_18
timestamp 1607194113
transform 1 0 39192 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_17
timestamp 1607194113
transform 1 0 38824 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_17
timestamp 1607194113
transform 1 0 38916 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_18
timestamp 1607194113
transform 1 0 39192 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_18
timestamp 1607194113
transform 1 0 40940 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_18
timestamp 1607194113
transform 1 0 41032 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_18
timestamp 1607194113
transform 1 0 40940 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_18
timestamp 1607194113
transform 1 0 41032 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_19
timestamp 1607194113
transform 1 0 41308 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_19
timestamp 1607194113
transform 1 0 43056 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  dff1_19
timestamp 1607194113
transform 1 0 41308 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_19
timestamp 1607194113
transform 1 0 43056 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_19
timestamp 1607194113
transform 1 0 43148 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_20
timestamp 1607194113
transform 1 0 43424 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  decap1_19
timestamp 1607194113
transform 1 0 43148 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_20
timestamp 1607194113
transform 1 0 43424 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_20
timestamp 1607194113
transform 1 0 45172 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_20
timestamp 1607194113
transform 1 0 45264 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_21
timestamp 1607194113
transform 1 0 45540 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_20
timestamp 1607194113
transform 1 0 45172 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_20
timestamp 1607194113
transform 1 0 45264 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_21
timestamp 1607194113
transform 1 0 45540 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_21
timestamp 1607194113
transform 1 0 47288 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_21
timestamp 1607194113
transform 1 0 47380 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_22
timestamp 1607194113
transform 1 0 47656 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_21
timestamp 1607194113
transform 1 0 47288 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_21
timestamp 1607194113
transform 1 0 47380 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_22
timestamp 1607194113
transform 1 0 47656 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_22
timestamp 1607194113
transform 1 0 49404 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_22
timestamp 1607194113
transform 1 0 49496 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_23
timestamp 1607194113
transform 1 0 49772 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_22
timestamp 1607194113
transform 1 0 49404 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_22
timestamp 1607194113
transform 1 0 49496 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_23
timestamp 1607194113
transform 1 0 49772 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_23
timestamp 1607194113
transform 1 0 51520 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_23
timestamp 1607194113
transform 1 0 51612 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_24
timestamp 1607194113
transform 1 0 51888 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_23
timestamp 1607194113
transform 1 0 51520 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_23
timestamp 1607194113
transform 1 0 51612 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_24
timestamp 1607194113
transform 1 0 51888 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_24
timestamp 1607194113
transform 1 0 53636 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_24
timestamp 1607194113
transform 1 0 53728 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_25
timestamp 1607194113
transform 1 0 54004 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_24
timestamp 1607194113
transform 1 0 53636 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_24
timestamp 1607194113
transform 1 0 53728 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_25
timestamp 1607194113
transform 1 0 54004 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_25
timestamp 1607194113
transform 1 0 55752 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_25
timestamp 1607194113
transform 1 0 55844 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_25
timestamp 1607194113
transform 1 0 55752 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_25
timestamp 1607194113
transform 1 0 55844 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_26
timestamp 1607194113
transform 1 0 56120 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  dff1_26
timestamp 1607194113
transform 1 0 56120 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_26
timestamp 1607194113
transform 1 0 57868 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_26
timestamp 1607194113
transform 1 0 57960 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_27
timestamp 1607194113
transform 1 0 58236 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_26
timestamp 1607194113
transform 1 0 57868 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_26
timestamp 1607194113
transform 1 0 57960 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_27
timestamp 1607194113
transform 1 0 58236 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_27
timestamp 1607194113
transform 1 0 59984 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_27
timestamp 1607194113
transform 1 0 60076 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_28
timestamp 1607194113
transform 1 0 60352 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_27
timestamp 1607194113
transform 1 0 59984 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_27
timestamp 1607194113
transform 1 0 60076 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_28
timestamp 1607194113
transform 1 0 60352 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_28
timestamp 1607194113
transform 1 0 62100 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_28
timestamp 1607194113
transform 1 0 62192 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_29
timestamp 1607194113
transform 1 0 62468 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_28
timestamp 1607194113
transform 1 0 62100 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_28
timestamp 1607194113
transform 1 0 62192 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_29
timestamp 1607194113
transform 1 0 62468 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_29
timestamp 1607194113
transform 1 0 64216 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_29
timestamp 1607194113
transform 1 0 64308 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_30
timestamp 1607194113
transform 1 0 64584 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_29
timestamp 1607194113
transform 1 0 64216 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_29
timestamp 1607194113
transform 1 0 64308 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_30
timestamp 1607194113
transform 1 0 64584 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_30
timestamp 1607194113
transform 1 0 66332 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_30
timestamp 1607194113
transform 1 0 66424 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_31
timestamp 1607194113
transform 1 0 66700 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_30
timestamp 1607194113
transform 1 0 66332 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_30
timestamp 1607194113
transform 1 0 66424 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_31
timestamp 1607194113
transform 1 0 66700 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_31
timestamp 1607194113
transform 1 0 68448 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_31
timestamp 1607194113
transform 1 0 68540 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_31
timestamp 1607194113
transform 1 0 68448 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_31
timestamp 1607194113
transform 1 0 68540 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_32
timestamp 1607194113
transform 1 0 68816 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  dff1_32
timestamp 1607194113
transform 1 0 68816 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_32
timestamp 1607194113
transform 1 0 70564 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_32
timestamp 1607194113
transform 1 0 70656 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_33
timestamp 1607194113
transform 1 0 70932 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_32
timestamp 1607194113
transform 1 0 70564 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_32
timestamp 1607194113
transform 1 0 70656 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_33
timestamp 1607194113
transform 1 0 70932 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_33
timestamp 1607194113
transform 1 0 72680 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_33
timestamp 1607194113
transform 1 0 72772 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_34
timestamp 1607194113
transform 1 0 73048 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_33
timestamp 1607194113
transform 1 0 72680 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_33
timestamp 1607194113
transform 1 0 72772 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_34
timestamp 1607194113
transform 1 0 73048 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_34
timestamp 1607194113
transform 1 0 74796 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_34
timestamp 1607194113
transform 1 0 74888 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_35
timestamp 1607194113
transform 1 0 75164 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_34
timestamp 1607194113
transform 1 0 74796 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_34
timestamp 1607194113
transform 1 0 74888 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_35
timestamp 1607194113
transform 1 0 75164 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_35
timestamp 1607194113
transform 1 0 76912 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_35
timestamp 1607194113
transform 1 0 77004 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_36
timestamp 1607194113
transform 1 0 77280 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_35
timestamp 1607194113
transform 1 0 76912 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_35
timestamp 1607194113
transform 1 0 77004 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_36
timestamp 1607194113
transform 1 0 77280 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_36
timestamp 1607194113
transform 1 0 79028 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_36
timestamp 1607194113
transform 1 0 79120 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_37
timestamp 1607194113
transform 1 0 79396 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_36
timestamp 1607194113
transform 1 0 79028 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_36
timestamp 1607194113
transform 1 0 79120 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_37
timestamp 1607194113
transform 1 0 79396 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_37
timestamp 1607194113
transform 1 0 81144 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_37
timestamp 1607194113
transform 1 0 81236 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_37
timestamp 1607194113
transform 1 0 81144 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_37
timestamp 1607194113
transform 1 0 81236 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_38
timestamp 1607194113
transform 1 0 81512 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  dff1_38
timestamp 1607194113
transform 1 0 81512 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_38
timestamp 1607194113
transform 1 0 83260 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_38
timestamp 1607194113
transform 1 0 83352 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_39
timestamp 1607194113
transform 1 0 83628 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_38
timestamp 1607194113
transform 1 0 83260 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_38
timestamp 1607194113
transform 1 0 83352 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_39
timestamp 1607194113
transform 1 0 83628 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_39
timestamp 1607194113
transform 1 0 85376 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_39
timestamp 1607194113
transform 1 0 85468 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_40
timestamp 1607194113
transform 1 0 85744 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_39
timestamp 1607194113
transform 1 0 85376 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_39
timestamp 1607194113
transform 1 0 85468 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_40
timestamp 1607194113
transform 1 0 85744 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_40
timestamp 1607194113
transform 1 0 87492 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_40
timestamp 1607194113
transform 1 0 87584 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_41
timestamp 1607194113
transform 1 0 87860 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_40
timestamp 1607194113
transform 1 0 87492 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_40
timestamp 1607194113
transform 1 0 87584 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_41
timestamp 1607194113
transform 1 0 87860 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_41
timestamp 1607194113
transform 1 0 89608 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_41
timestamp 1607194113
transform 1 0 89700 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_42
timestamp 1607194113
transform 1 0 89976 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_41
timestamp 1607194113
transform 1 0 89608 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_41
timestamp 1607194113
transform 1 0 89700 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_42
timestamp 1607194113
transform 1 0 89976 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_42
timestamp 1607194113
transform 1 0 91724 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_42
timestamp 1607194113
transform 1 0 91816 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_43
timestamp 1607194113
transform 1 0 92092 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_42
timestamp 1607194113
transform 1 0 91724 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_42
timestamp 1607194113
transform 1 0 91816 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_43
timestamp 1607194113
transform 1 0 92092 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_43
timestamp 1607194113
transform 1 0 93840 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_43
timestamp 1607194113
transform 1 0 93932 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_43
timestamp 1607194113
transform 1 0 93840 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_43
timestamp 1607194113
transform 1 0 93932 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_44
timestamp 1607194113
transform 1 0 94208 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_44
timestamp 1607194113
transform 1 0 95956 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  dff1_44
timestamp 1607194113
transform 1 0 94208 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_44
timestamp 1607194113
transform 1 0 95956 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_44
timestamp 1607194113
transform 1 0 96048 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_45
timestamp 1607194113
transform 1 0 96324 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  decap1_44
timestamp 1607194113
transform 1 0 96048 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_45
timestamp 1607194113
transform 1 0 96324 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_45
timestamp 1607194113
transform 1 0 98072 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_45
timestamp 1607194113
transform 1 0 98164 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_46
timestamp 1607194113
transform 1 0 98440 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_45
timestamp 1607194113
transform 1 0 98072 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_45
timestamp 1607194113
transform 1 0 98164 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_46
timestamp 1607194113
transform 1 0 98440 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_46
timestamp 1607194113
transform 1 0 100188 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_46
timestamp 1607194113
transform 1 0 100280 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_47
timestamp 1607194113
transform 1 0 100556 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_46
timestamp 1607194113
transform 1 0 100188 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_46
timestamp 1607194113
transform 1 0 100280 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_47
timestamp 1607194113
transform 1 0 100556 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_47
timestamp 1607194113
transform 1 0 102304 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_47
timestamp 1607194113
transform 1 0 102396 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_48
timestamp 1607194113
transform 1 0 102672 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_47
timestamp 1607194113
transform 1 0 102304 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_47
timestamp 1607194113
transform 1 0 102396 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_48
timestamp 1607194113
transform 1 0 102672 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_48
timestamp 1607194113
transform 1 0 104420 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_48
timestamp 1607194113
transform 1 0 104512 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_49
timestamp 1607194113
transform 1 0 104788 0 -1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_48
timestamp 1607194113
transform 1 0 104420 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_48
timestamp 1607194113
transform 1 0 104512 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_49
timestamp 1607194113
transform 1 0 104788 0 1 1632
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap0_49
timestamp 1607194113
transform 1 0 106536 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap0_49
timestamp 1607194113
transform 1 0 106628 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap1_49
timestamp 1607194113
transform 1 0 106536 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap1_49
timestamp 1607194113
transform 1 0 106628 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  delay_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 1104 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_0
timestamp 1607194113
transform 1 0 1472 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_0
timestamp 1607194113
transform 1 0 1564 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_0
timestamp 1607194113
transform 1 0 1840 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 1932 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 2668 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 3036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_1
timestamp 1607194113
transform 1 0 3220 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_1
timestamp 1607194113
transform 1 0 3588 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_1
timestamp 1607194113
transform 1 0 3680 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_17
timestamp 1607194113
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_18
timestamp 1607194113
transform 1 0 4048 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_19
timestamp 1607194113
transform 1 0 4784 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_20
timestamp 1607194113
transform 1 0 5152 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_2
timestamp 1607194113
transform 1 0 5336 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_2
timestamp 1607194113
transform 1 0 5704 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_2
timestamp 1607194113
transform 1 0 5796 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_33
timestamp 1607194113
transform 1 0 6072 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_34
timestamp 1607194113
transform 1 0 6164 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_35
timestamp 1607194113
transform 1 0 6900 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_36
timestamp 1607194113
transform 1 0 7268 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_3
timestamp 1607194113
transform 1 0 7452 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_3
timestamp 1607194113
transform 1 0 7820 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_3
timestamp 1607194113
transform 1 0 7912 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_49
timestamp 1607194113
transform 1 0 8188 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_50
timestamp 1607194113
transform 1 0 8280 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_51
timestamp 1607194113
transform 1 0 9016 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_52
timestamp 1607194113
transform 1 0 9384 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_4
timestamp 1607194113
transform 1 0 9568 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_4
timestamp 1607194113
transform 1 0 9936 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_4
timestamp 1607194113
transform 1 0 10028 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_65
timestamp 1607194113
transform 1 0 10304 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_66
timestamp 1607194113
transform 1 0 10396 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_67
timestamp 1607194113
transform 1 0 11132 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_68
timestamp 1607194113
transform 1 0 11500 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_5
timestamp 1607194113
transform 1 0 11684 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_5
timestamp 1607194113
transform 1 0 12052 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_5
timestamp 1607194113
transform 1 0 12144 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_81
timestamp 1607194113
transform 1 0 12420 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_82
timestamp 1607194113
transform 1 0 12512 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_83
timestamp 1607194113
transform 1 0 13248 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_84
timestamp 1607194113
transform 1 0 13616 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_6
timestamp 1607194113
transform 1 0 13800 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_6
timestamp 1607194113
transform 1 0 14168 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_6
timestamp 1607194113
transform 1 0 14260 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_97
timestamp 1607194113
transform 1 0 14536 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_98
timestamp 1607194113
transform 1 0 14628 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_99
timestamp 1607194113
transform 1 0 15364 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_100
timestamp 1607194113
transform 1 0 15732 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_7
timestamp 1607194113
transform 1 0 15916 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_7
timestamp 1607194113
transform 1 0 16284 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_7
timestamp 1607194113
transform 1 0 16376 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_113
timestamp 1607194113
transform 1 0 16652 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_114
timestamp 1607194113
transform 1 0 16744 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_115
timestamp 1607194113
transform 1 0 17480 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_116
timestamp 1607194113
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_8
timestamp 1607194113
transform 1 0 18032 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_8
timestamp 1607194113
transform 1 0 18400 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_8
timestamp 1607194113
transform 1 0 18492 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_129
timestamp 1607194113
transform 1 0 18768 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_130
timestamp 1607194113
transform 1 0 18860 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_131
timestamp 1607194113
transform 1 0 19596 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_132
timestamp 1607194113
transform 1 0 19964 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_9
timestamp 1607194113
transform 1 0 20148 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_9
timestamp 1607194113
transform 1 0 20516 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_9
timestamp 1607194113
transform 1 0 20608 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_145
timestamp 1607194113
transform 1 0 20884 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_146
timestamp 1607194113
transform 1 0 20976 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_147
timestamp 1607194113
transform 1 0 21712 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_148
timestamp 1607194113
transform 1 0 22080 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_10
timestamp 1607194113
transform 1 0 22264 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_10
timestamp 1607194113
transform 1 0 22632 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_10
timestamp 1607194113
transform 1 0 22724 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_161
timestamp 1607194113
transform 1 0 23000 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_162
timestamp 1607194113
transform 1 0 23092 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_163
timestamp 1607194113
transform 1 0 23828 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_164
timestamp 1607194113
transform 1 0 24196 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_11
timestamp 1607194113
transform 1 0 24380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_11
timestamp 1607194113
transform 1 0 24748 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_11
timestamp 1607194113
transform 1 0 24840 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_177
timestamp 1607194113
transform 1 0 25116 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_178
timestamp 1607194113
transform 1 0 25208 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_179
timestamp 1607194113
transform 1 0 25944 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_180
timestamp 1607194113
transform 1 0 26312 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_12
timestamp 1607194113
transform 1 0 26496 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_12
timestamp 1607194113
transform 1 0 26864 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_12
timestamp 1607194113
transform 1 0 26956 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_193
timestamp 1607194113
transform 1 0 27232 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_194
timestamp 1607194113
transform 1 0 27324 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_195
timestamp 1607194113
transform 1 0 28060 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_196
timestamp 1607194113
transform 1 0 28428 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_13
timestamp 1607194113
transform 1 0 28612 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_13
timestamp 1607194113
transform 1 0 28980 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_13
timestamp 1607194113
transform 1 0 29072 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_209
timestamp 1607194113
transform 1 0 29348 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_210
timestamp 1607194113
transform 1 0 29440 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_211
timestamp 1607194113
transform 1 0 30176 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_212
timestamp 1607194113
transform 1 0 30544 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_14
timestamp 1607194113
transform 1 0 30728 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_14
timestamp 1607194113
transform 1 0 31096 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_14
timestamp 1607194113
transform 1 0 31188 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_225
timestamp 1607194113
transform 1 0 31464 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_226
timestamp 1607194113
transform 1 0 31556 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_227
timestamp 1607194113
transform 1 0 32292 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_228
timestamp 1607194113
transform 1 0 32660 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_15
timestamp 1607194113
transform 1 0 32844 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_15
timestamp 1607194113
transform 1 0 33212 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_15
timestamp 1607194113
transform 1 0 33304 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_241
timestamp 1607194113
transform 1 0 33580 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_242
timestamp 1607194113
transform 1 0 33672 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_243
timestamp 1607194113
transform 1 0 34408 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_244
timestamp 1607194113
transform 1 0 34776 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_16
timestamp 1607194113
transform 1 0 34960 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_16
timestamp 1607194113
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_16
timestamp 1607194113
transform 1 0 35420 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_257
timestamp 1607194113
transform 1 0 35696 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_258
timestamp 1607194113
transform 1 0 35788 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_259
timestamp 1607194113
transform 1 0 36524 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_260
timestamp 1607194113
transform 1 0 36892 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_17
timestamp 1607194113
transform 1 0 37076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_17
timestamp 1607194113
transform 1 0 37444 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_17
timestamp 1607194113
transform 1 0 37536 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_273
timestamp 1607194113
transform 1 0 37812 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_274
timestamp 1607194113
transform 1 0 37904 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_275
timestamp 1607194113
transform 1 0 38640 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_276
timestamp 1607194113
transform 1 0 39008 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_18
timestamp 1607194113
transform 1 0 39192 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_18
timestamp 1607194113
transform 1 0 39560 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_18
timestamp 1607194113
transform 1 0 39652 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_289
timestamp 1607194113
transform 1 0 39928 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_290
timestamp 1607194113
transform 1 0 40020 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_291
timestamp 1607194113
transform 1 0 40756 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_292
timestamp 1607194113
transform 1 0 41124 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_19
timestamp 1607194113
transform 1 0 41308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_19
timestamp 1607194113
transform 1 0 41676 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_19
timestamp 1607194113
transform 1 0 41768 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_305
timestamp 1607194113
transform 1 0 42044 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_306
timestamp 1607194113
transform 1 0 42136 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_307
timestamp 1607194113
transform 1 0 42872 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_308
timestamp 1607194113
transform 1 0 43240 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_20
timestamp 1607194113
transform 1 0 43424 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_20
timestamp 1607194113
transform 1 0 43792 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_20
timestamp 1607194113
transform 1 0 43884 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_321
timestamp 1607194113
transform 1 0 44160 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_322
timestamp 1607194113
transform 1 0 44252 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_323
timestamp 1607194113
transform 1 0 44988 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_324
timestamp 1607194113
transform 1 0 45356 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_21
timestamp 1607194113
transform 1 0 45540 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_21
timestamp 1607194113
transform 1 0 45908 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_21
timestamp 1607194113
transform 1 0 46000 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_337
timestamp 1607194113
transform 1 0 46276 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_338
timestamp 1607194113
transform 1 0 46368 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_339
timestamp 1607194113
transform 1 0 47104 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_340
timestamp 1607194113
transform 1 0 47472 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_22
timestamp 1607194113
transform 1 0 47656 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_22
timestamp 1607194113
transform 1 0 48024 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_22
timestamp 1607194113
transform 1 0 48116 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_353
timestamp 1607194113
transform 1 0 48392 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_354
timestamp 1607194113
transform 1 0 48484 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_355
timestamp 1607194113
transform 1 0 49220 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_356
timestamp 1607194113
transform 1 0 49588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_23
timestamp 1607194113
transform 1 0 49772 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_23
timestamp 1607194113
transform 1 0 50140 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_23
timestamp 1607194113
transform 1 0 50232 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_369
timestamp 1607194113
transform 1 0 50508 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_370
timestamp 1607194113
transform 1 0 50600 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_371
timestamp 1607194113
transform 1 0 51336 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_372
timestamp 1607194113
transform 1 0 51704 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_24
timestamp 1607194113
transform 1 0 51888 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_24
timestamp 1607194113
transform 1 0 52256 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_24
timestamp 1607194113
transform 1 0 52348 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_385
timestamp 1607194113
transform 1 0 52624 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_386
timestamp 1607194113
transform 1 0 52716 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_387
timestamp 1607194113
transform 1 0 53452 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_388
timestamp 1607194113
transform 1 0 53820 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_25
timestamp 1607194113
transform 1 0 54004 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_25
timestamp 1607194113
transform 1 0 54372 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_25
timestamp 1607194113
transform 1 0 54464 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_401
timestamp 1607194113
transform 1 0 54740 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_402
timestamp 1607194113
transform 1 0 54832 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_403
timestamp 1607194113
transform 1 0 55568 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_404
timestamp 1607194113
transform 1 0 55936 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_26
timestamp 1607194113
transform 1 0 56120 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_26
timestamp 1607194113
transform 1 0 56488 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_26
timestamp 1607194113
transform 1 0 56580 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_417
timestamp 1607194113
transform 1 0 56856 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_418
timestamp 1607194113
transform 1 0 56948 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_419
timestamp 1607194113
transform 1 0 57684 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_420
timestamp 1607194113
transform 1 0 58052 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_27
timestamp 1607194113
transform 1 0 58236 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_27
timestamp 1607194113
transform 1 0 58604 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_27
timestamp 1607194113
transform 1 0 58696 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_433
timestamp 1607194113
transform 1 0 58972 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_434
timestamp 1607194113
transform 1 0 59064 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_435
timestamp 1607194113
transform 1 0 59800 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_436
timestamp 1607194113
transform 1 0 60168 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_28
timestamp 1607194113
transform 1 0 60352 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_28
timestamp 1607194113
transform 1 0 60720 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_28
timestamp 1607194113
transform 1 0 60812 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_449
timestamp 1607194113
transform 1 0 61088 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_450
timestamp 1607194113
transform 1 0 61180 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_451
timestamp 1607194113
transform 1 0 61916 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_452
timestamp 1607194113
transform 1 0 62284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_29
timestamp 1607194113
transform 1 0 62468 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_29
timestamp 1607194113
transform 1 0 62836 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_29
timestamp 1607194113
transform 1 0 62928 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_465
timestamp 1607194113
transform 1 0 63204 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_466
timestamp 1607194113
transform 1 0 63296 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_467
timestamp 1607194113
transform 1 0 64032 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_468
timestamp 1607194113
transform 1 0 64400 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_30
timestamp 1607194113
transform 1 0 64584 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_30
timestamp 1607194113
transform 1 0 64952 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_30
timestamp 1607194113
transform 1 0 65044 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_481
timestamp 1607194113
transform 1 0 65320 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_482
timestamp 1607194113
transform 1 0 65412 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_483
timestamp 1607194113
transform 1 0 66148 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_484
timestamp 1607194113
transform 1 0 66516 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_31
timestamp 1607194113
transform 1 0 66700 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_31
timestamp 1607194113
transform 1 0 67068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_31
timestamp 1607194113
transform 1 0 67160 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_497
timestamp 1607194113
transform 1 0 67436 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_498
timestamp 1607194113
transform 1 0 67528 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_499
timestamp 1607194113
transform 1 0 68264 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_500
timestamp 1607194113
transform 1 0 68632 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_32
timestamp 1607194113
transform 1 0 68816 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_32
timestamp 1607194113
transform 1 0 69184 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_32
timestamp 1607194113
transform 1 0 69276 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_513
timestamp 1607194113
transform 1 0 69552 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_514
timestamp 1607194113
transform 1 0 69644 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_515
timestamp 1607194113
transform 1 0 70380 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_516
timestamp 1607194113
transform 1 0 70748 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_33
timestamp 1607194113
transform 1 0 70932 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_33
timestamp 1607194113
transform 1 0 71300 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_33
timestamp 1607194113
transform 1 0 71392 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_529
timestamp 1607194113
transform 1 0 71668 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_530
timestamp 1607194113
transform 1 0 71760 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_531
timestamp 1607194113
transform 1 0 72496 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_532
timestamp 1607194113
transform 1 0 72864 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_34
timestamp 1607194113
transform 1 0 73048 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_34
timestamp 1607194113
transform 1 0 73416 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_34
timestamp 1607194113
transform 1 0 73508 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_545
timestamp 1607194113
transform 1 0 73784 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_546
timestamp 1607194113
transform 1 0 73876 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_547
timestamp 1607194113
transform 1 0 74612 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_548
timestamp 1607194113
transform 1 0 74980 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_35
timestamp 1607194113
transform 1 0 75164 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_35
timestamp 1607194113
transform 1 0 75532 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_35
timestamp 1607194113
transform 1 0 75624 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_561
timestamp 1607194113
transform 1 0 75900 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_562
timestamp 1607194113
transform 1 0 75992 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_563
timestamp 1607194113
transform 1 0 76728 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_564
timestamp 1607194113
transform 1 0 77096 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_36
timestamp 1607194113
transform 1 0 77280 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_36
timestamp 1607194113
transform 1 0 77648 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_36
timestamp 1607194113
transform 1 0 77740 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_577
timestamp 1607194113
transform 1 0 78016 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_578
timestamp 1607194113
transform 1 0 78108 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_579
timestamp 1607194113
transform 1 0 78844 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_580
timestamp 1607194113
transform 1 0 79212 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_37
timestamp 1607194113
transform 1 0 79396 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_37
timestamp 1607194113
transform 1 0 79764 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_37
timestamp 1607194113
transform 1 0 79856 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_593
timestamp 1607194113
transform 1 0 80132 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_594
timestamp 1607194113
transform 1 0 80224 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_595
timestamp 1607194113
transform 1 0 80960 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_596
timestamp 1607194113
transform 1 0 81328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_38
timestamp 1607194113
transform 1 0 81512 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_38
timestamp 1607194113
transform 1 0 81880 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_38
timestamp 1607194113
transform 1 0 81972 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_609
timestamp 1607194113
transform 1 0 82248 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_610
timestamp 1607194113
transform 1 0 82340 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_611
timestamp 1607194113
transform 1 0 83076 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_612
timestamp 1607194113
transform 1 0 83444 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_39
timestamp 1607194113
transform 1 0 83628 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_39
timestamp 1607194113
transform 1 0 83996 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_39
timestamp 1607194113
transform 1 0 84088 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_625
timestamp 1607194113
transform 1 0 84364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_626
timestamp 1607194113
transform 1 0 84456 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_627
timestamp 1607194113
transform 1 0 85192 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_628
timestamp 1607194113
transform 1 0 85560 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_40
timestamp 1607194113
transform 1 0 85744 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_40
timestamp 1607194113
transform 1 0 86112 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_40
timestamp 1607194113
transform 1 0 86204 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_641
timestamp 1607194113
transform 1 0 86480 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_642
timestamp 1607194113
transform 1 0 86572 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_643
timestamp 1607194113
transform 1 0 87308 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_644
timestamp 1607194113
transform 1 0 87676 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_41
timestamp 1607194113
transform 1 0 87860 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_41
timestamp 1607194113
transform 1 0 88228 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_41
timestamp 1607194113
transform 1 0 88320 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_657
timestamp 1607194113
transform 1 0 88596 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_658
timestamp 1607194113
transform 1 0 88688 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_659
timestamp 1607194113
transform 1 0 89424 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_660
timestamp 1607194113
transform 1 0 89792 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_42
timestamp 1607194113
transform 1 0 89976 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_42
timestamp 1607194113
transform 1 0 90344 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_42
timestamp 1607194113
transform 1 0 90436 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_673
timestamp 1607194113
transform 1 0 90712 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_674
timestamp 1607194113
transform 1 0 90804 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_675
timestamp 1607194113
transform 1 0 91540 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_676
timestamp 1607194113
transform 1 0 91908 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_43
timestamp 1607194113
transform 1 0 92092 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_43
timestamp 1607194113
transform 1 0 92460 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_43
timestamp 1607194113
transform 1 0 92552 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_689
timestamp 1607194113
transform 1 0 92828 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_690
timestamp 1607194113
transform 1 0 92920 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_691
timestamp 1607194113
transform 1 0 93656 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_692
timestamp 1607194113
transform 1 0 94024 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_44
timestamp 1607194113
transform 1 0 94208 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_44
timestamp 1607194113
transform 1 0 94576 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_44
timestamp 1607194113
transform 1 0 94668 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_705
timestamp 1607194113
transform 1 0 94944 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_706
timestamp 1607194113
transform 1 0 95036 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_707
timestamp 1607194113
transform 1 0 95772 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_708
timestamp 1607194113
transform 1 0 96140 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_45
timestamp 1607194113
transform 1 0 96324 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_45
timestamp 1607194113
transform 1 0 96692 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_45
timestamp 1607194113
transform 1 0 96784 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_721
timestamp 1607194113
transform 1 0 97060 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_722
timestamp 1607194113
transform 1 0 97152 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_723
timestamp 1607194113
transform 1 0 97888 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_724
timestamp 1607194113
transform 1 0 98256 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_46
timestamp 1607194113
transform 1 0 98440 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_46
timestamp 1607194113
transform 1 0 98808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_46
timestamp 1607194113
transform 1 0 98900 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_737
timestamp 1607194113
transform 1 0 99176 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_738
timestamp 1607194113
transform 1 0 99268 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_739
timestamp 1607194113
transform 1 0 100004 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_740
timestamp 1607194113
transform 1 0 100372 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_47
timestamp 1607194113
transform 1 0 100556 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_47
timestamp 1607194113
transform 1 0 100924 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_47
timestamp 1607194113
transform 1 0 101016 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_753
timestamp 1607194113
transform 1 0 101292 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_754
timestamp 1607194113
transform 1 0 101384 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_755
timestamp 1607194113
transform 1 0 102120 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_756
timestamp 1607194113
transform 1 0 102488 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_48
timestamp 1607194113
transform 1 0 102672 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_48
timestamp 1607194113
transform 1 0 103040 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_48
timestamp 1607194113
transform 1 0 103132 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_769
timestamp 1607194113
transform 1 0 103408 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_770
timestamp 1607194113
transform 1 0 103500 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_771
timestamp 1607194113
transform 1 0 104236 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_772
timestamp 1607194113
transform 1 0 104604 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_49
timestamp 1607194113
transform 1 0 104788 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap2_49
timestamp 1607194113
transform 1 0 105156 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap2_49
timestamp 1607194113
transform 1 0 105248 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_785
timestamp 1607194113
transform 1 0 105524 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_786
timestamp 1607194113
transform 1 0 105616 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_787
timestamp 1607194113
transform 1 0 106352 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_788
timestamp 1607194113
transform 1 0 106720 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_99
timestamp 1607194113
transform -1 0 1472 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_0
timestamp 1607194113
transform 1 0 1472 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_0
timestamp 1607194113
transform 1 0 1564 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_4
timestamp 1607194113
transform 1 0 1840 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_5
timestamp 1607194113
transform 1 0 1932 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_6
timestamp 1607194113
transform 1 0 2668 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_7
timestamp 1607194113
transform 1 0 3036 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_98
timestamp 1607194113
transform -1 0 3588 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_1
timestamp 1607194113
transform 1 0 3588 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_1
timestamp 1607194113
transform 1 0 3680 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_21
timestamp 1607194113
transform 1 0 3956 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_22
timestamp 1607194113
transform 1 0 4048 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_23
timestamp 1607194113
transform 1 0 4784 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_24
timestamp 1607194113
transform 1 0 5152 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_97
timestamp 1607194113
transform -1 0 5704 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_2
timestamp 1607194113
transform 1 0 5704 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_2
timestamp 1607194113
transform 1 0 5796 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_37
timestamp 1607194113
transform 1 0 6072 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_38
timestamp 1607194113
transform 1 0 6164 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_39
timestamp 1607194113
transform 1 0 6900 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_40
timestamp 1607194113
transform 1 0 7268 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_96
timestamp 1607194113
transform -1 0 7820 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_3
timestamp 1607194113
transform 1 0 7820 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_3
timestamp 1607194113
transform 1 0 7912 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_53
timestamp 1607194113
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_54
timestamp 1607194113
transform 1 0 8280 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_55
timestamp 1607194113
transform 1 0 9016 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_56
timestamp 1607194113
transform 1 0 9384 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_95
timestamp 1607194113
transform -1 0 9936 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_4
timestamp 1607194113
transform 1 0 9936 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_4
timestamp 1607194113
transform 1 0 10028 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_69
timestamp 1607194113
transform 1 0 10304 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_70
timestamp 1607194113
transform 1 0 10396 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_71
timestamp 1607194113
transform 1 0 11132 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_72
timestamp 1607194113
transform 1 0 11500 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_94
timestamp 1607194113
transform -1 0 12052 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_5
timestamp 1607194113
transform 1 0 12052 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_5
timestamp 1607194113
transform 1 0 12144 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_85
timestamp 1607194113
transform 1 0 12420 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_86
timestamp 1607194113
transform 1 0 12512 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_87
timestamp 1607194113
transform 1 0 13248 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_88
timestamp 1607194113
transform 1 0 13616 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_93
timestamp 1607194113
transform -1 0 14168 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_6
timestamp 1607194113
transform 1 0 14168 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_6
timestamp 1607194113
transform 1 0 14260 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_101
timestamp 1607194113
transform 1 0 14536 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_102
timestamp 1607194113
transform 1 0 14628 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_103
timestamp 1607194113
transform 1 0 15364 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_104
timestamp 1607194113
transform 1 0 15732 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_92
timestamp 1607194113
transform -1 0 16284 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_7
timestamp 1607194113
transform 1 0 16284 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_7
timestamp 1607194113
transform 1 0 16376 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_117
timestamp 1607194113
transform 1 0 16652 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_118
timestamp 1607194113
transform 1 0 16744 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_119
timestamp 1607194113
transform 1 0 17480 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_120
timestamp 1607194113
transform 1 0 17848 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_91
timestamp 1607194113
transform -1 0 18400 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_8
timestamp 1607194113
transform 1 0 18400 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_8
timestamp 1607194113
transform 1 0 18492 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_133
timestamp 1607194113
transform 1 0 18768 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_134
timestamp 1607194113
transform 1 0 18860 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_135
timestamp 1607194113
transform 1 0 19596 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_136
timestamp 1607194113
transform 1 0 19964 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_90
timestamp 1607194113
transform -1 0 20516 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_9
timestamp 1607194113
transform 1 0 20516 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_9
timestamp 1607194113
transform 1 0 20608 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_149
timestamp 1607194113
transform 1 0 20884 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_150
timestamp 1607194113
transform 1 0 20976 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_151
timestamp 1607194113
transform 1 0 21712 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_152
timestamp 1607194113
transform 1 0 22080 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_89
timestamp 1607194113
transform -1 0 22632 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_10
timestamp 1607194113
transform 1 0 22632 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_10
timestamp 1607194113
transform 1 0 22724 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_165
timestamp 1607194113
transform 1 0 23000 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_166
timestamp 1607194113
transform 1 0 23092 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_167
timestamp 1607194113
transform 1 0 23828 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_168
timestamp 1607194113
transform 1 0 24196 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_88
timestamp 1607194113
transform -1 0 24748 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_11
timestamp 1607194113
transform 1 0 24748 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_11
timestamp 1607194113
transform 1 0 24840 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_181
timestamp 1607194113
transform 1 0 25116 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_182
timestamp 1607194113
transform 1 0 25208 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_183
timestamp 1607194113
transform 1 0 25944 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_184
timestamp 1607194113
transform 1 0 26312 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_87
timestamp 1607194113
transform -1 0 26864 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_12
timestamp 1607194113
transform 1 0 26864 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_12
timestamp 1607194113
transform 1 0 26956 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_197
timestamp 1607194113
transform 1 0 27232 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_198
timestamp 1607194113
transform 1 0 27324 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_199
timestamp 1607194113
transform 1 0 28060 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_200
timestamp 1607194113
transform 1 0 28428 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_86
timestamp 1607194113
transform -1 0 28980 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_13
timestamp 1607194113
transform 1 0 28980 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_13
timestamp 1607194113
transform 1 0 29072 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_213
timestamp 1607194113
transform 1 0 29348 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_214
timestamp 1607194113
transform 1 0 29440 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_215
timestamp 1607194113
transform 1 0 30176 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_216
timestamp 1607194113
transform 1 0 30544 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_85
timestamp 1607194113
transform -1 0 31096 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_14
timestamp 1607194113
transform 1 0 31096 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_14
timestamp 1607194113
transform 1 0 31188 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_229
timestamp 1607194113
transform 1 0 31464 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_230
timestamp 1607194113
transform 1 0 31556 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_231
timestamp 1607194113
transform 1 0 32292 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_232
timestamp 1607194113
transform 1 0 32660 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_84
timestamp 1607194113
transform -1 0 33212 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_15
timestamp 1607194113
transform 1 0 33212 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_15
timestamp 1607194113
transform 1 0 33304 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_245
timestamp 1607194113
transform 1 0 33580 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_246
timestamp 1607194113
transform 1 0 33672 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_247
timestamp 1607194113
transform 1 0 34408 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_248
timestamp 1607194113
transform 1 0 34776 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_83
timestamp 1607194113
transform -1 0 35328 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_16
timestamp 1607194113
transform 1 0 35328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_16
timestamp 1607194113
transform 1 0 35420 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_261
timestamp 1607194113
transform 1 0 35696 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_262
timestamp 1607194113
transform 1 0 35788 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_263
timestamp 1607194113
transform 1 0 36524 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_264
timestamp 1607194113
transform 1 0 36892 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_82
timestamp 1607194113
transform -1 0 37444 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_17
timestamp 1607194113
transform 1 0 37444 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_17
timestamp 1607194113
transform 1 0 37536 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_277
timestamp 1607194113
transform 1 0 37812 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_278
timestamp 1607194113
transform 1 0 37904 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_279
timestamp 1607194113
transform 1 0 38640 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_280
timestamp 1607194113
transform 1 0 39008 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_81
timestamp 1607194113
transform -1 0 39560 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_18
timestamp 1607194113
transform 1 0 39560 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_18
timestamp 1607194113
transform 1 0 39652 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_293
timestamp 1607194113
transform 1 0 39928 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_294
timestamp 1607194113
transform 1 0 40020 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_295
timestamp 1607194113
transform 1 0 40756 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_296
timestamp 1607194113
transform 1 0 41124 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_80
timestamp 1607194113
transform -1 0 41676 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_19
timestamp 1607194113
transform 1 0 41676 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_19
timestamp 1607194113
transform 1 0 41768 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_309
timestamp 1607194113
transform 1 0 42044 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_310
timestamp 1607194113
transform 1 0 42136 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_311
timestamp 1607194113
transform 1 0 42872 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_312
timestamp 1607194113
transform 1 0 43240 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_79
timestamp 1607194113
transform -1 0 43792 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_20
timestamp 1607194113
transform 1 0 43792 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_20
timestamp 1607194113
transform 1 0 43884 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_325
timestamp 1607194113
transform 1 0 44160 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_326
timestamp 1607194113
transform 1 0 44252 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_327
timestamp 1607194113
transform 1 0 44988 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_328
timestamp 1607194113
transform 1 0 45356 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_78
timestamp 1607194113
transform -1 0 45908 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_21
timestamp 1607194113
transform 1 0 45908 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_21
timestamp 1607194113
transform 1 0 46000 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_341
timestamp 1607194113
transform 1 0 46276 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_342
timestamp 1607194113
transform 1 0 46368 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_343
timestamp 1607194113
transform 1 0 47104 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_344
timestamp 1607194113
transform 1 0 47472 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_77
timestamp 1607194113
transform -1 0 48024 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_22
timestamp 1607194113
transform 1 0 48024 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_22
timestamp 1607194113
transform 1 0 48116 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_357
timestamp 1607194113
transform 1 0 48392 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_358
timestamp 1607194113
transform 1 0 48484 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_359
timestamp 1607194113
transform 1 0 49220 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_360
timestamp 1607194113
transform 1 0 49588 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_76
timestamp 1607194113
transform -1 0 50140 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_23
timestamp 1607194113
transform 1 0 50140 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_23
timestamp 1607194113
transform 1 0 50232 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_373
timestamp 1607194113
transform 1 0 50508 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_374
timestamp 1607194113
transform 1 0 50600 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_375
timestamp 1607194113
transform 1 0 51336 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_376
timestamp 1607194113
transform 1 0 51704 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_75
timestamp 1607194113
transform -1 0 52256 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_24
timestamp 1607194113
transform 1 0 52256 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_24
timestamp 1607194113
transform 1 0 52348 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_389
timestamp 1607194113
transform 1 0 52624 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_390
timestamp 1607194113
transform 1 0 52716 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_391
timestamp 1607194113
transform 1 0 53452 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_392
timestamp 1607194113
transform 1 0 53820 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_74
timestamp 1607194113
transform -1 0 54372 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_25
timestamp 1607194113
transform 1 0 54372 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_25
timestamp 1607194113
transform 1 0 54464 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_405
timestamp 1607194113
transform 1 0 54740 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_406
timestamp 1607194113
transform 1 0 54832 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_407
timestamp 1607194113
transform 1 0 55568 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_408
timestamp 1607194113
transform 1 0 55936 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_73
timestamp 1607194113
transform -1 0 56488 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_26
timestamp 1607194113
transform 1 0 56488 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_26
timestamp 1607194113
transform 1 0 56580 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_421
timestamp 1607194113
transform 1 0 56856 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_422
timestamp 1607194113
transform 1 0 56948 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_423
timestamp 1607194113
transform 1 0 57684 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_424
timestamp 1607194113
transform 1 0 58052 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_72
timestamp 1607194113
transform -1 0 58604 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_27
timestamp 1607194113
transform 1 0 58604 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_27
timestamp 1607194113
transform 1 0 58696 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_437
timestamp 1607194113
transform 1 0 58972 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_438
timestamp 1607194113
transform 1 0 59064 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_439
timestamp 1607194113
transform 1 0 59800 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_440
timestamp 1607194113
transform 1 0 60168 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_71
timestamp 1607194113
transform -1 0 60720 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_28
timestamp 1607194113
transform 1 0 60720 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_28
timestamp 1607194113
transform 1 0 60812 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_453
timestamp 1607194113
transform 1 0 61088 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_454
timestamp 1607194113
transform 1 0 61180 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_455
timestamp 1607194113
transform 1 0 61916 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_456
timestamp 1607194113
transform 1 0 62284 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_70
timestamp 1607194113
transform -1 0 62836 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_29
timestamp 1607194113
transform 1 0 62836 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_29
timestamp 1607194113
transform 1 0 62928 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_469
timestamp 1607194113
transform 1 0 63204 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_470
timestamp 1607194113
transform 1 0 63296 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_471
timestamp 1607194113
transform 1 0 64032 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_472
timestamp 1607194113
transform 1 0 64400 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_69
timestamp 1607194113
transform -1 0 64952 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_30
timestamp 1607194113
transform 1 0 64952 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_30
timestamp 1607194113
transform 1 0 65044 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_485
timestamp 1607194113
transform 1 0 65320 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_486
timestamp 1607194113
transform 1 0 65412 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_487
timestamp 1607194113
transform 1 0 66148 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_488
timestamp 1607194113
transform 1 0 66516 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_68
timestamp 1607194113
transform -1 0 67068 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_31
timestamp 1607194113
transform 1 0 67068 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_31
timestamp 1607194113
transform 1 0 67160 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_501
timestamp 1607194113
transform 1 0 67436 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_502
timestamp 1607194113
transform 1 0 67528 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_503
timestamp 1607194113
transform 1 0 68264 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_504
timestamp 1607194113
transform 1 0 68632 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_67
timestamp 1607194113
transform -1 0 69184 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_32
timestamp 1607194113
transform 1 0 69184 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_32
timestamp 1607194113
transform 1 0 69276 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_517
timestamp 1607194113
transform 1 0 69552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_518
timestamp 1607194113
transform 1 0 69644 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_519
timestamp 1607194113
transform 1 0 70380 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_520
timestamp 1607194113
transform 1 0 70748 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_66
timestamp 1607194113
transform -1 0 71300 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_33
timestamp 1607194113
transform 1 0 71300 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_33
timestamp 1607194113
transform 1 0 71392 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_533
timestamp 1607194113
transform 1 0 71668 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_534
timestamp 1607194113
transform 1 0 71760 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_535
timestamp 1607194113
transform 1 0 72496 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_536
timestamp 1607194113
transform 1 0 72864 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_65
timestamp 1607194113
transform -1 0 73416 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_34
timestamp 1607194113
transform 1 0 73416 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_34
timestamp 1607194113
transform 1 0 73508 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_549
timestamp 1607194113
transform 1 0 73784 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_550
timestamp 1607194113
transform 1 0 73876 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_551
timestamp 1607194113
transform 1 0 74612 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_552
timestamp 1607194113
transform 1 0 74980 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_64
timestamp 1607194113
transform -1 0 75532 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_35
timestamp 1607194113
transform 1 0 75532 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_35
timestamp 1607194113
transform 1 0 75624 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_565
timestamp 1607194113
transform 1 0 75900 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_566
timestamp 1607194113
transform 1 0 75992 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_567
timestamp 1607194113
transform 1 0 76728 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_568
timestamp 1607194113
transform 1 0 77096 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_63
timestamp 1607194113
transform -1 0 77648 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_36
timestamp 1607194113
transform 1 0 77648 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_36
timestamp 1607194113
transform 1 0 77740 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_581
timestamp 1607194113
transform 1 0 78016 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_582
timestamp 1607194113
transform 1 0 78108 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_583
timestamp 1607194113
transform 1 0 78844 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_584
timestamp 1607194113
transform 1 0 79212 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_62
timestamp 1607194113
transform -1 0 79764 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_37
timestamp 1607194113
transform 1 0 79764 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_37
timestamp 1607194113
transform 1 0 79856 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_597
timestamp 1607194113
transform 1 0 80132 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_598
timestamp 1607194113
transform 1 0 80224 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_599
timestamp 1607194113
transform 1 0 80960 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_600
timestamp 1607194113
transform 1 0 81328 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_61
timestamp 1607194113
transform -1 0 81880 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_38
timestamp 1607194113
transform 1 0 81880 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_38
timestamp 1607194113
transform 1 0 81972 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_613
timestamp 1607194113
transform 1 0 82248 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_614
timestamp 1607194113
transform 1 0 82340 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_615
timestamp 1607194113
transform 1 0 83076 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_616
timestamp 1607194113
transform 1 0 83444 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_60
timestamp 1607194113
transform -1 0 83996 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_39
timestamp 1607194113
transform 1 0 83996 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_39
timestamp 1607194113
transform 1 0 84088 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_629
timestamp 1607194113
transform 1 0 84364 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_630
timestamp 1607194113
transform 1 0 84456 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_631
timestamp 1607194113
transform 1 0 85192 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_632
timestamp 1607194113
transform 1 0 85560 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_59
timestamp 1607194113
transform -1 0 86112 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_40
timestamp 1607194113
transform 1 0 86112 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_40
timestamp 1607194113
transform 1 0 86204 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_645
timestamp 1607194113
transform 1 0 86480 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_646
timestamp 1607194113
transform 1 0 86572 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_647
timestamp 1607194113
transform 1 0 87308 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_648
timestamp 1607194113
transform 1 0 87676 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_58
timestamp 1607194113
transform -1 0 88228 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_41
timestamp 1607194113
transform 1 0 88228 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_41
timestamp 1607194113
transform 1 0 88320 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_661
timestamp 1607194113
transform 1 0 88596 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_662
timestamp 1607194113
transform 1 0 88688 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_663
timestamp 1607194113
transform 1 0 89424 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_664
timestamp 1607194113
transform 1 0 89792 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_57
timestamp 1607194113
transform -1 0 90344 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_42
timestamp 1607194113
transform 1 0 90344 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_42
timestamp 1607194113
transform 1 0 90436 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_677
timestamp 1607194113
transform 1 0 90712 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_678
timestamp 1607194113
transform 1 0 90804 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_679
timestamp 1607194113
transform 1 0 91540 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_680
timestamp 1607194113
transform 1 0 91908 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_56
timestamp 1607194113
transform -1 0 92460 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_43
timestamp 1607194113
transform 1 0 92460 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_43
timestamp 1607194113
transform 1 0 92552 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_693
timestamp 1607194113
transform 1 0 92828 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_694
timestamp 1607194113
transform 1 0 92920 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_695
timestamp 1607194113
transform 1 0 93656 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_696
timestamp 1607194113
transform 1 0 94024 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_55
timestamp 1607194113
transform -1 0 94576 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_44
timestamp 1607194113
transform 1 0 94576 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_44
timestamp 1607194113
transform 1 0 94668 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_709
timestamp 1607194113
transform 1 0 94944 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_710
timestamp 1607194113
transform 1 0 95036 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_711
timestamp 1607194113
transform 1 0 95772 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_712
timestamp 1607194113
transform 1 0 96140 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_54
timestamp 1607194113
transform -1 0 96692 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_45
timestamp 1607194113
transform 1 0 96692 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_45
timestamp 1607194113
transform 1 0 96784 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_725
timestamp 1607194113
transform 1 0 97060 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_726
timestamp 1607194113
transform 1 0 97152 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_727
timestamp 1607194113
transform 1 0 97888 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_728
timestamp 1607194113
transform 1 0 98256 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_53
timestamp 1607194113
transform -1 0 98808 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_46
timestamp 1607194113
transform 1 0 98808 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_46
timestamp 1607194113
transform 1 0 98900 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_741
timestamp 1607194113
transform 1 0 99176 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_742
timestamp 1607194113
transform 1 0 99268 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_743
timestamp 1607194113
transform 1 0 100004 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_744
timestamp 1607194113
transform 1 0 100372 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_52
timestamp 1607194113
transform -1 0 100924 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_47
timestamp 1607194113
transform 1 0 100924 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_47
timestamp 1607194113
transform 1 0 101016 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_757
timestamp 1607194113
transform 1 0 101292 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_758
timestamp 1607194113
transform 1 0 101384 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_759
timestamp 1607194113
transform 1 0 102120 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_760
timestamp 1607194113
transform 1 0 102488 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_51
timestamp 1607194113
transform -1 0 103040 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_48
timestamp 1607194113
transform 1 0 103040 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_48
timestamp 1607194113
transform 1 0 103132 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_773
timestamp 1607194113
transform 1 0 103408 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_774
timestamp 1607194113
transform 1 0 103500 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_775
timestamp 1607194113
transform 1 0 104236 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_776
timestamp 1607194113
transform 1 0 104604 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_50
timestamp 1607194113
transform -1 0 105156 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap3_49
timestamp 1607194113
transform 1 0 105156 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap3_49
timestamp 1607194113
transform 1 0 105248 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_789
timestamp 1607194113
transform 1 0 105524 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_790
timestamp 1607194113
transform 1 0 105616 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_791
timestamp 1607194113
transform 1 0 106352 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_792
timestamp 1607194113
transform 1 0 106720 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  dff1_99
timestamp 1607194113
transform 1 0 1104 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_0
timestamp 1607194113
transform 1 0 2852 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_0
timestamp 1607194113
transform 1 0 2944 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_98
timestamp 1607194113
transform 1 0 3220 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_1
timestamp 1607194113
transform 1 0 4968 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_1
timestamp 1607194113
transform 1 0 5060 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_97
timestamp 1607194113
transform 1 0 5336 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_2
timestamp 1607194113
transform 1 0 7084 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_2
timestamp 1607194113
transform 1 0 7176 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_96
timestamp 1607194113
transform 1 0 7452 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_3
timestamp 1607194113
transform 1 0 9200 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_3
timestamp 1607194113
transform 1 0 9292 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_95
timestamp 1607194113
transform 1 0 9568 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_4
timestamp 1607194113
transform 1 0 11316 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_4
timestamp 1607194113
transform 1 0 11408 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_94
timestamp 1607194113
transform 1 0 11684 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_5
timestamp 1607194113
transform 1 0 13432 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_5
timestamp 1607194113
transform 1 0 13524 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_93
timestamp 1607194113
transform 1 0 13800 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_6
timestamp 1607194113
transform 1 0 15548 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_6
timestamp 1607194113
transform 1 0 15640 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_92
timestamp 1607194113
transform 1 0 15916 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_7
timestamp 1607194113
transform 1 0 17664 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_7
timestamp 1607194113
transform 1 0 17756 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_91
timestamp 1607194113
transform 1 0 18032 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_8
timestamp 1607194113
transform 1 0 19780 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_8
timestamp 1607194113
transform 1 0 19872 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_90
timestamp 1607194113
transform 1 0 20148 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_9
timestamp 1607194113
transform 1 0 21896 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_9
timestamp 1607194113
transform 1 0 21988 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_89
timestamp 1607194113
transform 1 0 22264 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_10
timestamp 1607194113
transform 1 0 24012 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_10
timestamp 1607194113
transform 1 0 24104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_88
timestamp 1607194113
transform 1 0 24380 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_11
timestamp 1607194113
transform 1 0 26128 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_11
timestamp 1607194113
transform 1 0 26220 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_87
timestamp 1607194113
transform 1 0 26496 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_12
timestamp 1607194113
transform 1 0 28244 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_12
timestamp 1607194113
transform 1 0 28336 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_86
timestamp 1607194113
transform 1 0 28612 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_13
timestamp 1607194113
transform 1 0 30360 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_13
timestamp 1607194113
transform 1 0 30452 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_85
timestamp 1607194113
transform 1 0 30728 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_14
timestamp 1607194113
transform 1 0 32476 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_14
timestamp 1607194113
transform 1 0 32568 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_84
timestamp 1607194113
transform 1 0 32844 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_15
timestamp 1607194113
transform 1 0 34592 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_15
timestamp 1607194113
transform 1 0 34684 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_83
timestamp 1607194113
transform 1 0 34960 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_16
timestamp 1607194113
transform 1 0 36708 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_16
timestamp 1607194113
transform 1 0 36800 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_82
timestamp 1607194113
transform 1 0 37076 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_17
timestamp 1607194113
transform 1 0 38824 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_17
timestamp 1607194113
transform 1 0 38916 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_81
timestamp 1607194113
transform 1 0 39192 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_18
timestamp 1607194113
transform 1 0 40940 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_18
timestamp 1607194113
transform 1 0 41032 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_80
timestamp 1607194113
transform 1 0 41308 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_19
timestamp 1607194113
transform 1 0 43056 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_19
timestamp 1607194113
transform 1 0 43148 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_79
timestamp 1607194113
transform 1 0 43424 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_20
timestamp 1607194113
transform 1 0 45172 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_20
timestamp 1607194113
transform 1 0 45264 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_78
timestamp 1607194113
transform 1 0 45540 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_21
timestamp 1607194113
transform 1 0 47288 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_21
timestamp 1607194113
transform 1 0 47380 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_77
timestamp 1607194113
transform 1 0 47656 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_22
timestamp 1607194113
transform 1 0 49404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_22
timestamp 1607194113
transform 1 0 49496 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_76
timestamp 1607194113
transform 1 0 49772 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_23
timestamp 1607194113
transform 1 0 51520 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_23
timestamp 1607194113
transform 1 0 51612 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_75
timestamp 1607194113
transform 1 0 51888 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_24
timestamp 1607194113
transform 1 0 53636 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_24
timestamp 1607194113
transform 1 0 53728 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_74
timestamp 1607194113
transform 1 0 54004 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_25
timestamp 1607194113
transform 1 0 55752 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_25
timestamp 1607194113
transform 1 0 55844 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_73
timestamp 1607194113
transform 1 0 56120 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_26
timestamp 1607194113
transform 1 0 57868 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_26
timestamp 1607194113
transform 1 0 57960 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_72
timestamp 1607194113
transform 1 0 58236 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_27
timestamp 1607194113
transform 1 0 59984 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_27
timestamp 1607194113
transform 1 0 60076 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_71
timestamp 1607194113
transform 1 0 60352 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_28
timestamp 1607194113
transform 1 0 62100 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_28
timestamp 1607194113
transform 1 0 62192 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_70
timestamp 1607194113
transform 1 0 62468 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_29
timestamp 1607194113
transform 1 0 64216 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_29
timestamp 1607194113
transform 1 0 64308 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_69
timestamp 1607194113
transform 1 0 64584 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_30
timestamp 1607194113
transform 1 0 66332 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_30
timestamp 1607194113
transform 1 0 66424 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_68
timestamp 1607194113
transform 1 0 66700 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_31
timestamp 1607194113
transform 1 0 68448 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_31
timestamp 1607194113
transform 1 0 68540 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_67
timestamp 1607194113
transform 1 0 68816 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_32
timestamp 1607194113
transform 1 0 70564 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_32
timestamp 1607194113
transform 1 0 70656 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_66
timestamp 1607194113
transform 1 0 70932 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_33
timestamp 1607194113
transform 1 0 72680 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_33
timestamp 1607194113
transform 1 0 72772 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_65
timestamp 1607194113
transform 1 0 73048 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_34
timestamp 1607194113
transform 1 0 74796 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_34
timestamp 1607194113
transform 1 0 74888 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_64
timestamp 1607194113
transform 1 0 75164 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_35
timestamp 1607194113
transform 1 0 76912 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_35
timestamp 1607194113
transform 1 0 77004 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_63
timestamp 1607194113
transform 1 0 77280 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_36
timestamp 1607194113
transform 1 0 79028 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_36
timestamp 1607194113
transform 1 0 79120 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_62
timestamp 1607194113
transform 1 0 79396 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_37
timestamp 1607194113
transform 1 0 81144 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_37
timestamp 1607194113
transform 1 0 81236 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_61
timestamp 1607194113
transform 1 0 81512 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_38
timestamp 1607194113
transform 1 0 83260 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_38
timestamp 1607194113
transform 1 0 83352 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_60
timestamp 1607194113
transform 1 0 83628 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_39
timestamp 1607194113
transform 1 0 85376 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_39
timestamp 1607194113
transform 1 0 85468 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_59
timestamp 1607194113
transform 1 0 85744 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_40
timestamp 1607194113
transform 1 0 87492 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_40
timestamp 1607194113
transform 1 0 87584 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_58
timestamp 1607194113
transform 1 0 87860 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_41
timestamp 1607194113
transform 1 0 89608 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_41
timestamp 1607194113
transform 1 0 89700 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_57
timestamp 1607194113
transform 1 0 89976 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_42
timestamp 1607194113
transform 1 0 91724 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_42
timestamp 1607194113
transform 1 0 91816 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_56
timestamp 1607194113
transform 1 0 92092 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_43
timestamp 1607194113
transform 1 0 93840 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_43
timestamp 1607194113
transform 1 0 93932 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_55
timestamp 1607194113
transform 1 0 94208 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_44
timestamp 1607194113
transform 1 0 95956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_44
timestamp 1607194113
transform 1 0 96048 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_54
timestamp 1607194113
transform 1 0 96324 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_45
timestamp 1607194113
transform 1 0 98072 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_45
timestamp 1607194113
transform 1 0 98164 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_53
timestamp 1607194113
transform 1 0 98440 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_46
timestamp 1607194113
transform 1 0 100188 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_46
timestamp 1607194113
transform 1 0 100280 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_52
timestamp 1607194113
transform 1 0 100556 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_47
timestamp 1607194113
transform 1 0 102304 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_47
timestamp 1607194113
transform 1 0 102396 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_51
timestamp 1607194113
transform 1 0 102672 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_48
timestamp 1607194113
transform 1 0 104420 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_48
timestamp 1607194113
transform 1 0 104512 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_50
timestamp 1607194113
transform 1 0 104788 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap4_49
timestamp 1607194113
transform 1 0 106536 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap4_49
timestamp 1607194113
transform 1 0 106628 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_99
timestamp 1607194113
transform 1 0 1104 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_0
timestamp 1607194113
transform 1 0 2852 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_0
timestamp 1607194113
transform 1 0 2944 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_98
timestamp 1607194113
transform 1 0 3220 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_1
timestamp 1607194113
transform 1 0 4968 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_1
timestamp 1607194113
transform 1 0 5060 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_97
timestamp 1607194113
transform 1 0 5336 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_2
timestamp 1607194113
transform 1 0 7084 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_2
timestamp 1607194113
transform 1 0 7176 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_96
timestamp 1607194113
transform 1 0 7452 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_3
timestamp 1607194113
transform 1 0 9200 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_3
timestamp 1607194113
transform 1 0 9292 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_95
timestamp 1607194113
transform 1 0 9568 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_4
timestamp 1607194113
transform 1 0 11316 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_4
timestamp 1607194113
transform 1 0 11408 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_94
timestamp 1607194113
transform 1 0 11684 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_5
timestamp 1607194113
transform 1 0 13432 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_5
timestamp 1607194113
transform 1 0 13524 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_93
timestamp 1607194113
transform 1 0 13800 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_6
timestamp 1607194113
transform 1 0 15548 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_6
timestamp 1607194113
transform 1 0 15640 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_92
timestamp 1607194113
transform 1 0 15916 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_7
timestamp 1607194113
transform 1 0 17664 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_7
timestamp 1607194113
transform 1 0 17756 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_91
timestamp 1607194113
transform 1 0 18032 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_8
timestamp 1607194113
transform 1 0 19780 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_8
timestamp 1607194113
transform 1 0 19872 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_90
timestamp 1607194113
transform 1 0 20148 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_9
timestamp 1607194113
transform 1 0 21896 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_9
timestamp 1607194113
transform 1 0 21988 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_89
timestamp 1607194113
transform 1 0 22264 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_10
timestamp 1607194113
transform 1 0 24012 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_10
timestamp 1607194113
transform 1 0 24104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_88
timestamp 1607194113
transform 1 0 24380 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_11
timestamp 1607194113
transform 1 0 26128 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_11
timestamp 1607194113
transform 1 0 26220 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_87
timestamp 1607194113
transform 1 0 26496 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_12
timestamp 1607194113
transform 1 0 28244 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_12
timestamp 1607194113
transform 1 0 28336 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_86
timestamp 1607194113
transform 1 0 28612 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_13
timestamp 1607194113
transform 1 0 30360 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_13
timestamp 1607194113
transform 1 0 30452 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_85
timestamp 1607194113
transform 1 0 30728 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_14
timestamp 1607194113
transform 1 0 32476 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_14
timestamp 1607194113
transform 1 0 32568 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_84
timestamp 1607194113
transform 1 0 32844 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_15
timestamp 1607194113
transform 1 0 34592 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_15
timestamp 1607194113
transform 1 0 34684 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_83
timestamp 1607194113
transform 1 0 34960 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_16
timestamp 1607194113
transform 1 0 36708 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_16
timestamp 1607194113
transform 1 0 36800 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_82
timestamp 1607194113
transform 1 0 37076 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_17
timestamp 1607194113
transform 1 0 38824 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_17
timestamp 1607194113
transform 1 0 38916 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_81
timestamp 1607194113
transform 1 0 39192 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_18
timestamp 1607194113
transform 1 0 40940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_18
timestamp 1607194113
transform 1 0 41032 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_80
timestamp 1607194113
transform 1 0 41308 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_19
timestamp 1607194113
transform 1 0 43056 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_19
timestamp 1607194113
transform 1 0 43148 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_79
timestamp 1607194113
transform 1 0 43424 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_20
timestamp 1607194113
transform 1 0 45172 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_20
timestamp 1607194113
transform 1 0 45264 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_78
timestamp 1607194113
transform 1 0 45540 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_21
timestamp 1607194113
transform 1 0 47288 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_21
timestamp 1607194113
transform 1 0 47380 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_77
timestamp 1607194113
transform 1 0 47656 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_22
timestamp 1607194113
transform 1 0 49404 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_22
timestamp 1607194113
transform 1 0 49496 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_76
timestamp 1607194113
transform 1 0 49772 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_23
timestamp 1607194113
transform 1 0 51520 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_23
timestamp 1607194113
transform 1 0 51612 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_75
timestamp 1607194113
transform 1 0 51888 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_24
timestamp 1607194113
transform 1 0 53636 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_24
timestamp 1607194113
transform 1 0 53728 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_74
timestamp 1607194113
transform 1 0 54004 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_25
timestamp 1607194113
transform 1 0 55752 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_25
timestamp 1607194113
transform 1 0 55844 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_73
timestamp 1607194113
transform 1 0 56120 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_26
timestamp 1607194113
transform 1 0 57868 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_26
timestamp 1607194113
transform 1 0 57960 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_72
timestamp 1607194113
transform 1 0 58236 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_27
timestamp 1607194113
transform 1 0 59984 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_27
timestamp 1607194113
transform 1 0 60076 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_71
timestamp 1607194113
transform 1 0 60352 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_28
timestamp 1607194113
transform 1 0 62100 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_28
timestamp 1607194113
transform 1 0 62192 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_70
timestamp 1607194113
transform 1 0 62468 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_29
timestamp 1607194113
transform 1 0 64216 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_29
timestamp 1607194113
transform 1 0 64308 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_69
timestamp 1607194113
transform 1 0 64584 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_30
timestamp 1607194113
transform 1 0 66332 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_30
timestamp 1607194113
transform 1 0 66424 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_68
timestamp 1607194113
transform 1 0 66700 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_31
timestamp 1607194113
transform 1 0 68448 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_31
timestamp 1607194113
transform 1 0 68540 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_67
timestamp 1607194113
transform 1 0 68816 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_32
timestamp 1607194113
transform 1 0 70564 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_32
timestamp 1607194113
transform 1 0 70656 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_66
timestamp 1607194113
transform 1 0 70932 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_33
timestamp 1607194113
transform 1 0 72680 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_33
timestamp 1607194113
transform 1 0 72772 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_65
timestamp 1607194113
transform 1 0 73048 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_34
timestamp 1607194113
transform 1 0 74796 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_34
timestamp 1607194113
transform 1 0 74888 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_64
timestamp 1607194113
transform 1 0 75164 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_35
timestamp 1607194113
transform 1 0 76912 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_35
timestamp 1607194113
transform 1 0 77004 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_63
timestamp 1607194113
transform 1 0 77280 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_36
timestamp 1607194113
transform 1 0 79028 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_36
timestamp 1607194113
transform 1 0 79120 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_62
timestamp 1607194113
transform 1 0 79396 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_37
timestamp 1607194113
transform 1 0 81144 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_37
timestamp 1607194113
transform 1 0 81236 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_61
timestamp 1607194113
transform 1 0 81512 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_38
timestamp 1607194113
transform 1 0 83260 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_38
timestamp 1607194113
transform 1 0 83352 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_60
timestamp 1607194113
transform 1 0 83628 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_39
timestamp 1607194113
transform 1 0 85376 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_39
timestamp 1607194113
transform 1 0 85468 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_59
timestamp 1607194113
transform 1 0 85744 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_40
timestamp 1607194113
transform 1 0 87492 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_40
timestamp 1607194113
transform 1 0 87584 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_58
timestamp 1607194113
transform 1 0 87860 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_41
timestamp 1607194113
transform 1 0 89608 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_41
timestamp 1607194113
transform 1 0 89700 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_57
timestamp 1607194113
transform 1 0 89976 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_42
timestamp 1607194113
transform 1 0 91724 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_42
timestamp 1607194113
transform 1 0 91816 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_56
timestamp 1607194113
transform 1 0 92092 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_43
timestamp 1607194113
transform 1 0 93840 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_43
timestamp 1607194113
transform 1 0 93932 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_55
timestamp 1607194113
transform 1 0 94208 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_44
timestamp 1607194113
transform 1 0 95956 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_44
timestamp 1607194113
transform 1 0 96048 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_54
timestamp 1607194113
transform 1 0 96324 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_45
timestamp 1607194113
transform 1 0 98072 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_45
timestamp 1607194113
transform 1 0 98164 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_53
timestamp 1607194113
transform 1 0 98440 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_46
timestamp 1607194113
transform 1 0 100188 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_46
timestamp 1607194113
transform 1 0 100280 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_52
timestamp 1607194113
transform 1 0 100556 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_47
timestamp 1607194113
transform 1 0 102304 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_47
timestamp 1607194113
transform 1 0 102396 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_51
timestamp 1607194113
transform 1 0 102672 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_48
timestamp 1607194113
transform 1 0 104420 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_48
timestamp 1607194113
transform 1 0 104512 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_50
timestamp 1607194113
transform 1 0 104788 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap5_49
timestamp 1607194113
transform 1 0 106536 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap5_49
timestamp 1607194113
transform 1 0 106628 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_100
timestamp 1607194113
transform 1 0 1104 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_0
timestamp 1607194113
transform 1 0 2852 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  dff1_100
timestamp 1607194113
transform 1 0 1104 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_0
timestamp 1607194113
transform 1 0 2852 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_0
timestamp 1607194113
transform 1 0 2944 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_101
timestamp 1607194113
transform 1 0 3220 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  decap7_0
timestamp 1607194113
transform 1 0 2944 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_101
timestamp 1607194113
transform 1 0 3220 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_1
timestamp 1607194113
transform 1 0 4968 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_1
timestamp 1607194113
transform 1 0 5060 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_102
timestamp 1607194113
transform 1 0 5336 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_1
timestamp 1607194113
transform 1 0 4968 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_1
timestamp 1607194113
transform 1 0 5060 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_102
timestamp 1607194113
transform 1 0 5336 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_2
timestamp 1607194113
transform 1 0 7084 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_2
timestamp 1607194113
transform 1 0 7176 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_103
timestamp 1607194113
transform 1 0 7452 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_2
timestamp 1607194113
transform 1 0 7084 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_2
timestamp 1607194113
transform 1 0 7176 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_103
timestamp 1607194113
transform 1 0 7452 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_3
timestamp 1607194113
transform 1 0 9200 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_3
timestamp 1607194113
transform 1 0 9292 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_104
timestamp 1607194113
transform 1 0 9568 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_3
timestamp 1607194113
transform 1 0 9200 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_3
timestamp 1607194113
transform 1 0 9292 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_104
timestamp 1607194113
transform 1 0 9568 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_4
timestamp 1607194113
transform 1 0 11316 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_4
timestamp 1607194113
transform 1 0 11408 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_105
timestamp 1607194113
transform 1 0 11684 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_4
timestamp 1607194113
transform 1 0 11316 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_4
timestamp 1607194113
transform 1 0 11408 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_105
timestamp 1607194113
transform 1 0 11684 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_5
timestamp 1607194113
transform 1 0 13432 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_5
timestamp 1607194113
transform 1 0 13524 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_106
timestamp 1607194113
transform 1 0 13800 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_5
timestamp 1607194113
transform 1 0 13432 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_5
timestamp 1607194113
transform 1 0 13524 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_106
timestamp 1607194113
transform 1 0 13800 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_6
timestamp 1607194113
transform 1 0 15548 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_6
timestamp 1607194113
transform 1 0 15640 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_6
timestamp 1607194113
transform 1 0 15548 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_6
timestamp 1607194113
transform 1 0 15640 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_107
timestamp 1607194113
transform 1 0 15916 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  dff1_107
timestamp 1607194113
transform 1 0 15916 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_7
timestamp 1607194113
transform 1 0 17664 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_7
timestamp 1607194113
transform 1 0 17756 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_108
timestamp 1607194113
transform 1 0 18032 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_7
timestamp 1607194113
transform 1 0 17664 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_7
timestamp 1607194113
transform 1 0 17756 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_108
timestamp 1607194113
transform 1 0 18032 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_8
timestamp 1607194113
transform 1 0 19780 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_8
timestamp 1607194113
transform 1 0 19872 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_109
timestamp 1607194113
transform 1 0 20148 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_8
timestamp 1607194113
transform 1 0 19780 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_8
timestamp 1607194113
transform 1 0 19872 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_109
timestamp 1607194113
transform 1 0 20148 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_9
timestamp 1607194113
transform 1 0 21896 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_9
timestamp 1607194113
transform 1 0 21988 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_110
timestamp 1607194113
transform 1 0 22264 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_9
timestamp 1607194113
transform 1 0 21896 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_9
timestamp 1607194113
transform 1 0 21988 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_110
timestamp 1607194113
transform 1 0 22264 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_10
timestamp 1607194113
transform 1 0 24012 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_10
timestamp 1607194113
transform 1 0 24104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_111
timestamp 1607194113
transform 1 0 24380 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_10
timestamp 1607194113
transform 1 0 24012 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_10
timestamp 1607194113
transform 1 0 24104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_111
timestamp 1607194113
transform 1 0 24380 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_11
timestamp 1607194113
transform 1 0 26128 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_11
timestamp 1607194113
transform 1 0 26220 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_112
timestamp 1607194113
transform 1 0 26496 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_11
timestamp 1607194113
transform 1 0 26128 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_11
timestamp 1607194113
transform 1 0 26220 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_112
timestamp 1607194113
transform 1 0 26496 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_12
timestamp 1607194113
transform 1 0 28244 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_12
timestamp 1607194113
transform 1 0 28336 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_12
timestamp 1607194113
transform 1 0 28244 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_12
timestamp 1607194113
transform 1 0 28336 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_113
timestamp 1607194113
transform 1 0 28612 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  dff1_113
timestamp 1607194113
transform 1 0 28612 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_13
timestamp 1607194113
transform 1 0 30360 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_13
timestamp 1607194113
transform 1 0 30452 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_114
timestamp 1607194113
transform 1 0 30728 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_13
timestamp 1607194113
transform 1 0 30360 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_13
timestamp 1607194113
transform 1 0 30452 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_114
timestamp 1607194113
transform 1 0 30728 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_14
timestamp 1607194113
transform 1 0 32476 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_14
timestamp 1607194113
transform 1 0 32568 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_115
timestamp 1607194113
transform 1 0 32844 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_14
timestamp 1607194113
transform 1 0 32476 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_14
timestamp 1607194113
transform 1 0 32568 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_115
timestamp 1607194113
transform 1 0 32844 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_15
timestamp 1607194113
transform 1 0 34592 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_15
timestamp 1607194113
transform 1 0 34684 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_116
timestamp 1607194113
transform 1 0 34960 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_15
timestamp 1607194113
transform 1 0 34592 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_15
timestamp 1607194113
transform 1 0 34684 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_116
timestamp 1607194113
transform 1 0 34960 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_16
timestamp 1607194113
transform 1 0 36708 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_16
timestamp 1607194113
transform 1 0 36800 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_117
timestamp 1607194113
transform 1 0 37076 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_16
timestamp 1607194113
transform 1 0 36708 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_16
timestamp 1607194113
transform 1 0 36800 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_117
timestamp 1607194113
transform 1 0 37076 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_17
timestamp 1607194113
transform 1 0 38824 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_17
timestamp 1607194113
transform 1 0 38916 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_118
timestamp 1607194113
transform 1 0 39192 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_17
timestamp 1607194113
transform 1 0 38824 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_17
timestamp 1607194113
transform 1 0 38916 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_118
timestamp 1607194113
transform 1 0 39192 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_18
timestamp 1607194113
transform 1 0 40940 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_18
timestamp 1607194113
transform 1 0 41032 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_18
timestamp 1607194113
transform 1 0 40940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_18
timestamp 1607194113
transform 1 0 41032 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_119
timestamp 1607194113
transform 1 0 41308 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_19
timestamp 1607194113
transform 1 0 43056 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  dff1_119
timestamp 1607194113
transform 1 0 41308 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_19
timestamp 1607194113
transform 1 0 43056 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_19
timestamp 1607194113
transform 1 0 43148 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_120
timestamp 1607194113
transform 1 0 43424 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  decap7_19
timestamp 1607194113
transform 1 0 43148 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_120
timestamp 1607194113
transform 1 0 43424 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_20
timestamp 1607194113
transform 1 0 45172 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_20
timestamp 1607194113
transform 1 0 45264 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_121
timestamp 1607194113
transform 1 0 45540 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_20
timestamp 1607194113
transform 1 0 45172 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_20
timestamp 1607194113
transform 1 0 45264 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_121
timestamp 1607194113
transform 1 0 45540 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_21
timestamp 1607194113
transform 1 0 47288 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_21
timestamp 1607194113
transform 1 0 47380 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_122
timestamp 1607194113
transform 1 0 47656 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_21
timestamp 1607194113
transform 1 0 47288 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_21
timestamp 1607194113
transform 1 0 47380 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_122
timestamp 1607194113
transform 1 0 47656 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_22
timestamp 1607194113
transform 1 0 49404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_22
timestamp 1607194113
transform 1 0 49496 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_123
timestamp 1607194113
transform 1 0 49772 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_22
timestamp 1607194113
transform 1 0 49404 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_22
timestamp 1607194113
transform 1 0 49496 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_123
timestamp 1607194113
transform 1 0 49772 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_23
timestamp 1607194113
transform 1 0 51520 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_23
timestamp 1607194113
transform 1 0 51612 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_124
timestamp 1607194113
transform 1 0 51888 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_23
timestamp 1607194113
transform 1 0 51520 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_23
timestamp 1607194113
transform 1 0 51612 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_124
timestamp 1607194113
transform 1 0 51888 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_24
timestamp 1607194113
transform 1 0 53636 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_24
timestamp 1607194113
transform 1 0 53728 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_125
timestamp 1607194113
transform 1 0 54004 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_24
timestamp 1607194113
transform 1 0 53636 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_24
timestamp 1607194113
transform 1 0 53728 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_125
timestamp 1607194113
transform 1 0 54004 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_25
timestamp 1607194113
transform 1 0 55752 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_25
timestamp 1607194113
transform 1 0 55844 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_25
timestamp 1607194113
transform 1 0 55752 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_25
timestamp 1607194113
transform 1 0 55844 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_126
timestamp 1607194113
transform 1 0 56120 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  dff1_126
timestamp 1607194113
transform 1 0 56120 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_26
timestamp 1607194113
transform 1 0 57868 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_26
timestamp 1607194113
transform 1 0 57960 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_127
timestamp 1607194113
transform 1 0 58236 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_26
timestamp 1607194113
transform 1 0 57868 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_26
timestamp 1607194113
transform 1 0 57960 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_127
timestamp 1607194113
transform 1 0 58236 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_27
timestamp 1607194113
transform 1 0 59984 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_27
timestamp 1607194113
transform 1 0 60076 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_128
timestamp 1607194113
transform 1 0 60352 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_27
timestamp 1607194113
transform 1 0 59984 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_27
timestamp 1607194113
transform 1 0 60076 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_128
timestamp 1607194113
transform 1 0 60352 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_28
timestamp 1607194113
transform 1 0 62100 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_28
timestamp 1607194113
transform 1 0 62192 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_129
timestamp 1607194113
transform 1 0 62468 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_28
timestamp 1607194113
transform 1 0 62100 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_28
timestamp 1607194113
transform 1 0 62192 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_129
timestamp 1607194113
transform 1 0 62468 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_29
timestamp 1607194113
transform 1 0 64216 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_29
timestamp 1607194113
transform 1 0 64308 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_130
timestamp 1607194113
transform 1 0 64584 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_29
timestamp 1607194113
transform 1 0 64216 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_29
timestamp 1607194113
transform 1 0 64308 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_130
timestamp 1607194113
transform 1 0 64584 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_30
timestamp 1607194113
transform 1 0 66332 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_30
timestamp 1607194113
transform 1 0 66424 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_131
timestamp 1607194113
transform 1 0 66700 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_30
timestamp 1607194113
transform 1 0 66332 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_30
timestamp 1607194113
transform 1 0 66424 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_131
timestamp 1607194113
transform 1 0 66700 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_31
timestamp 1607194113
transform 1 0 68448 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_31
timestamp 1607194113
transform 1 0 68540 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_31
timestamp 1607194113
transform 1 0 68448 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_31
timestamp 1607194113
transform 1 0 68540 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_132
timestamp 1607194113
transform 1 0 68816 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  dff1_132
timestamp 1607194113
transform 1 0 68816 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_32
timestamp 1607194113
transform 1 0 70564 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_32
timestamp 1607194113
transform 1 0 70656 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_133
timestamp 1607194113
transform 1 0 70932 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_32
timestamp 1607194113
transform 1 0 70564 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_32
timestamp 1607194113
transform 1 0 70656 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_133
timestamp 1607194113
transform 1 0 70932 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_33
timestamp 1607194113
transform 1 0 72680 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_33
timestamp 1607194113
transform 1 0 72772 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_134
timestamp 1607194113
transform 1 0 73048 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_33
timestamp 1607194113
transform 1 0 72680 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_33
timestamp 1607194113
transform 1 0 72772 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_134
timestamp 1607194113
transform 1 0 73048 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_34
timestamp 1607194113
transform 1 0 74796 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_34
timestamp 1607194113
transform 1 0 74888 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_135
timestamp 1607194113
transform 1 0 75164 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_34
timestamp 1607194113
transform 1 0 74796 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_34
timestamp 1607194113
transform 1 0 74888 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_135
timestamp 1607194113
transform 1 0 75164 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_35
timestamp 1607194113
transform 1 0 76912 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_35
timestamp 1607194113
transform 1 0 77004 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_136
timestamp 1607194113
transform 1 0 77280 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_35
timestamp 1607194113
transform 1 0 76912 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_35
timestamp 1607194113
transform 1 0 77004 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_136
timestamp 1607194113
transform 1 0 77280 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_36
timestamp 1607194113
transform 1 0 79028 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_36
timestamp 1607194113
transform 1 0 79120 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_137
timestamp 1607194113
transform 1 0 79396 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_36
timestamp 1607194113
transform 1 0 79028 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_36
timestamp 1607194113
transform 1 0 79120 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_137
timestamp 1607194113
transform 1 0 79396 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_37
timestamp 1607194113
transform 1 0 81144 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_37
timestamp 1607194113
transform 1 0 81236 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_37
timestamp 1607194113
transform 1 0 81144 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_37
timestamp 1607194113
transform 1 0 81236 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_138
timestamp 1607194113
transform 1 0 81512 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  dff1_138
timestamp 1607194113
transform 1 0 81512 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_38
timestamp 1607194113
transform 1 0 83260 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_38
timestamp 1607194113
transform 1 0 83352 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_139
timestamp 1607194113
transform 1 0 83628 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_38
timestamp 1607194113
transform 1 0 83260 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_38
timestamp 1607194113
transform 1 0 83352 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_139
timestamp 1607194113
transform 1 0 83628 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_39
timestamp 1607194113
transform 1 0 85376 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_39
timestamp 1607194113
transform 1 0 85468 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_140
timestamp 1607194113
transform 1 0 85744 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_39
timestamp 1607194113
transform 1 0 85376 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_39
timestamp 1607194113
transform 1 0 85468 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_140
timestamp 1607194113
transform 1 0 85744 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_40
timestamp 1607194113
transform 1 0 87492 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_40
timestamp 1607194113
transform 1 0 87584 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_141
timestamp 1607194113
transform 1 0 87860 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_40
timestamp 1607194113
transform 1 0 87492 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_40
timestamp 1607194113
transform 1 0 87584 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_141
timestamp 1607194113
transform 1 0 87860 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_41
timestamp 1607194113
transform 1 0 89608 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_41
timestamp 1607194113
transform 1 0 89700 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_142
timestamp 1607194113
transform 1 0 89976 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_41
timestamp 1607194113
transform 1 0 89608 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_41
timestamp 1607194113
transform 1 0 89700 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_142
timestamp 1607194113
transform 1 0 89976 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_42
timestamp 1607194113
transform 1 0 91724 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_42
timestamp 1607194113
transform 1 0 91816 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_143
timestamp 1607194113
transform 1 0 92092 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_42
timestamp 1607194113
transform 1 0 91724 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_42
timestamp 1607194113
transform 1 0 91816 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_143
timestamp 1607194113
transform 1 0 92092 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_43
timestamp 1607194113
transform 1 0 93840 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_43
timestamp 1607194113
transform 1 0 93932 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_43
timestamp 1607194113
transform 1 0 93840 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_43
timestamp 1607194113
transform 1 0 93932 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_144
timestamp 1607194113
transform 1 0 94208 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_44
timestamp 1607194113
transform 1 0 95956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  dff1_144
timestamp 1607194113
transform 1 0 94208 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_44
timestamp 1607194113
transform 1 0 95956 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_44
timestamp 1607194113
transform 1 0 96048 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_145
timestamp 1607194113
transform 1 0 96324 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  decap7_44
timestamp 1607194113
transform 1 0 96048 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_145
timestamp 1607194113
transform 1 0 96324 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_45
timestamp 1607194113
transform 1 0 98072 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_45
timestamp 1607194113
transform 1 0 98164 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_146
timestamp 1607194113
transform 1 0 98440 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_45
timestamp 1607194113
transform 1 0 98072 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_45
timestamp 1607194113
transform 1 0 98164 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_146
timestamp 1607194113
transform 1 0 98440 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_46
timestamp 1607194113
transform 1 0 100188 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_46
timestamp 1607194113
transform 1 0 100280 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_147
timestamp 1607194113
transform 1 0 100556 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_46
timestamp 1607194113
transform 1 0 100188 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_46
timestamp 1607194113
transform 1 0 100280 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_147
timestamp 1607194113
transform 1 0 100556 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_47
timestamp 1607194113
transform 1 0 102304 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_47
timestamp 1607194113
transform 1 0 102396 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_148
timestamp 1607194113
transform 1 0 102672 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_47
timestamp 1607194113
transform 1 0 102304 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_47
timestamp 1607194113
transform 1 0 102396 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_148
timestamp 1607194113
transform 1 0 102672 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_48
timestamp 1607194113
transform 1 0 104420 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_48
timestamp 1607194113
transform 1 0 104512 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_149
timestamp 1607194113
transform 1 0 104788 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_48
timestamp 1607194113
transform 1 0 104420 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_48
timestamp 1607194113
transform 1 0 104512 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_149
timestamp 1607194113
transform 1 0 104788 0 1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap6_49
timestamp 1607194113
transform 1 0 106536 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap6_49
timestamp 1607194113
transform 1 0 106628 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap7_49
timestamp 1607194113
transform 1 0 106536 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap7_49
timestamp 1607194113
transform 1 0 106628 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  delay_100
timestamp 1607194113
transform 1 0 1104 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_0
timestamp 1607194113
transform 1 0 1472 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_0
timestamp 1607194113
transform 1 0 1564 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_8
timestamp 1607194113
transform 1 0 1840 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_9
timestamp 1607194113
transform 1 0 1932 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_10
timestamp 1607194113
transform 1 0 2668 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_11
timestamp 1607194113
transform 1 0 3036 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_101
timestamp 1607194113
transform 1 0 3220 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_1
timestamp 1607194113
transform 1 0 3588 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_1
timestamp 1607194113
transform 1 0 3680 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_25
timestamp 1607194113
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_26
timestamp 1607194113
transform 1 0 4048 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_27
timestamp 1607194113
transform 1 0 4784 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_28
timestamp 1607194113
transform 1 0 5152 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_102
timestamp 1607194113
transform 1 0 5336 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_2
timestamp 1607194113
transform 1 0 5704 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_2
timestamp 1607194113
transform 1 0 5796 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_41
timestamp 1607194113
transform 1 0 6072 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_42
timestamp 1607194113
transform 1 0 6164 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_43
timestamp 1607194113
transform 1 0 6900 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_44
timestamp 1607194113
transform 1 0 7268 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_103
timestamp 1607194113
transform 1 0 7452 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_3
timestamp 1607194113
transform 1 0 7820 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_3
timestamp 1607194113
transform 1 0 7912 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_57
timestamp 1607194113
transform 1 0 8188 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_58
timestamp 1607194113
transform 1 0 8280 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_59
timestamp 1607194113
transform 1 0 9016 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_60
timestamp 1607194113
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_104
timestamp 1607194113
transform 1 0 9568 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_4
timestamp 1607194113
transform 1 0 9936 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_4
timestamp 1607194113
transform 1 0 10028 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_73
timestamp 1607194113
transform 1 0 10304 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_74
timestamp 1607194113
transform 1 0 10396 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_75
timestamp 1607194113
transform 1 0 11132 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_76
timestamp 1607194113
transform 1 0 11500 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_105
timestamp 1607194113
transform 1 0 11684 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_5
timestamp 1607194113
transform 1 0 12052 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_5
timestamp 1607194113
transform 1 0 12144 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_89
timestamp 1607194113
transform 1 0 12420 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_90
timestamp 1607194113
transform 1 0 12512 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_91
timestamp 1607194113
transform 1 0 13248 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_92
timestamp 1607194113
transform 1 0 13616 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_106
timestamp 1607194113
transform 1 0 13800 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_6
timestamp 1607194113
transform 1 0 14168 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_6
timestamp 1607194113
transform 1 0 14260 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_105
timestamp 1607194113
transform 1 0 14536 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_106
timestamp 1607194113
transform 1 0 14628 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_107
timestamp 1607194113
transform 1 0 15364 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_108
timestamp 1607194113
transform 1 0 15732 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_107
timestamp 1607194113
transform 1 0 15916 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_7
timestamp 1607194113
transform 1 0 16284 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_7
timestamp 1607194113
transform 1 0 16376 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_121
timestamp 1607194113
transform 1 0 16652 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_122
timestamp 1607194113
transform 1 0 16744 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_123
timestamp 1607194113
transform 1 0 17480 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_124
timestamp 1607194113
transform 1 0 17848 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_108
timestamp 1607194113
transform 1 0 18032 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_8
timestamp 1607194113
transform 1 0 18400 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_8
timestamp 1607194113
transform 1 0 18492 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_137
timestamp 1607194113
transform 1 0 18768 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_138
timestamp 1607194113
transform 1 0 18860 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_139
timestamp 1607194113
transform 1 0 19596 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_140
timestamp 1607194113
transform 1 0 19964 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_109
timestamp 1607194113
transform 1 0 20148 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_9
timestamp 1607194113
transform 1 0 20516 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_9
timestamp 1607194113
transform 1 0 20608 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_153
timestamp 1607194113
transform 1 0 20884 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_154
timestamp 1607194113
transform 1 0 20976 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_155
timestamp 1607194113
transform 1 0 21712 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_156
timestamp 1607194113
transform 1 0 22080 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_110
timestamp 1607194113
transform 1 0 22264 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_10
timestamp 1607194113
transform 1 0 22632 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_10
timestamp 1607194113
transform 1 0 22724 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_169
timestamp 1607194113
transform 1 0 23000 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_170
timestamp 1607194113
transform 1 0 23092 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_171
timestamp 1607194113
transform 1 0 23828 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_172
timestamp 1607194113
transform 1 0 24196 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_111
timestamp 1607194113
transform 1 0 24380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_11
timestamp 1607194113
transform 1 0 24748 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_11
timestamp 1607194113
transform 1 0 24840 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_185
timestamp 1607194113
transform 1 0 25116 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_186
timestamp 1607194113
transform 1 0 25208 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_187
timestamp 1607194113
transform 1 0 25944 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_188
timestamp 1607194113
transform 1 0 26312 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_112
timestamp 1607194113
transform 1 0 26496 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_12
timestamp 1607194113
transform 1 0 26864 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_12
timestamp 1607194113
transform 1 0 26956 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_201
timestamp 1607194113
transform 1 0 27232 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_202
timestamp 1607194113
transform 1 0 27324 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_203
timestamp 1607194113
transform 1 0 28060 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_204
timestamp 1607194113
transform 1 0 28428 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_113
timestamp 1607194113
transform 1 0 28612 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_13
timestamp 1607194113
transform 1 0 28980 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_13
timestamp 1607194113
transform 1 0 29072 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_217
timestamp 1607194113
transform 1 0 29348 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_218
timestamp 1607194113
transform 1 0 29440 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_219
timestamp 1607194113
transform 1 0 30176 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_220
timestamp 1607194113
transform 1 0 30544 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_114
timestamp 1607194113
transform 1 0 30728 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_14
timestamp 1607194113
transform 1 0 31096 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_14
timestamp 1607194113
transform 1 0 31188 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_233
timestamp 1607194113
transform 1 0 31464 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_234
timestamp 1607194113
transform 1 0 31556 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_235
timestamp 1607194113
transform 1 0 32292 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_236
timestamp 1607194113
transform 1 0 32660 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_115
timestamp 1607194113
transform 1 0 32844 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_15
timestamp 1607194113
transform 1 0 33212 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_15
timestamp 1607194113
transform 1 0 33304 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_249
timestamp 1607194113
transform 1 0 33580 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_250
timestamp 1607194113
transform 1 0 33672 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_251
timestamp 1607194113
transform 1 0 34408 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_252
timestamp 1607194113
transform 1 0 34776 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_116
timestamp 1607194113
transform 1 0 34960 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_16
timestamp 1607194113
transform 1 0 35328 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_16
timestamp 1607194113
transform 1 0 35420 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_265
timestamp 1607194113
transform 1 0 35696 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_266
timestamp 1607194113
transform 1 0 35788 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_267
timestamp 1607194113
transform 1 0 36524 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_268
timestamp 1607194113
transform 1 0 36892 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_117
timestamp 1607194113
transform 1 0 37076 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_17
timestamp 1607194113
transform 1 0 37444 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_17
timestamp 1607194113
transform 1 0 37536 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_281
timestamp 1607194113
transform 1 0 37812 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_282
timestamp 1607194113
transform 1 0 37904 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_283
timestamp 1607194113
transform 1 0 38640 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_284
timestamp 1607194113
transform 1 0 39008 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_118
timestamp 1607194113
transform 1 0 39192 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_18
timestamp 1607194113
transform 1 0 39560 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_18
timestamp 1607194113
transform 1 0 39652 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_297
timestamp 1607194113
transform 1 0 39928 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_298
timestamp 1607194113
transform 1 0 40020 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_299
timestamp 1607194113
transform 1 0 40756 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_300
timestamp 1607194113
transform 1 0 41124 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_119
timestamp 1607194113
transform 1 0 41308 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_19
timestamp 1607194113
transform 1 0 41676 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_19
timestamp 1607194113
transform 1 0 41768 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_313
timestamp 1607194113
transform 1 0 42044 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_314
timestamp 1607194113
transform 1 0 42136 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_315
timestamp 1607194113
transform 1 0 42872 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_316
timestamp 1607194113
transform 1 0 43240 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_120
timestamp 1607194113
transform 1 0 43424 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_20
timestamp 1607194113
transform 1 0 43792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_20
timestamp 1607194113
transform 1 0 43884 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_329
timestamp 1607194113
transform 1 0 44160 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_330
timestamp 1607194113
transform 1 0 44252 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_331
timestamp 1607194113
transform 1 0 44988 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_332
timestamp 1607194113
transform 1 0 45356 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_121
timestamp 1607194113
transform 1 0 45540 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_21
timestamp 1607194113
transform 1 0 45908 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_21
timestamp 1607194113
transform 1 0 46000 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_345
timestamp 1607194113
transform 1 0 46276 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_346
timestamp 1607194113
transform 1 0 46368 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_347
timestamp 1607194113
transform 1 0 47104 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_348
timestamp 1607194113
transform 1 0 47472 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_122
timestamp 1607194113
transform 1 0 47656 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_22
timestamp 1607194113
transform 1 0 48024 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_22
timestamp 1607194113
transform 1 0 48116 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_361
timestamp 1607194113
transform 1 0 48392 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_362
timestamp 1607194113
transform 1 0 48484 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_363
timestamp 1607194113
transform 1 0 49220 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_364
timestamp 1607194113
transform 1 0 49588 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_123
timestamp 1607194113
transform 1 0 49772 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_23
timestamp 1607194113
transform 1 0 50140 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_23
timestamp 1607194113
transform 1 0 50232 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_377
timestamp 1607194113
transform 1 0 50508 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_378
timestamp 1607194113
transform 1 0 50600 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_379
timestamp 1607194113
transform 1 0 51336 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_380
timestamp 1607194113
transform 1 0 51704 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_124
timestamp 1607194113
transform 1 0 51888 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_24
timestamp 1607194113
transform 1 0 52256 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_24
timestamp 1607194113
transform 1 0 52348 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_393
timestamp 1607194113
transform 1 0 52624 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_394
timestamp 1607194113
transform 1 0 52716 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_395
timestamp 1607194113
transform 1 0 53452 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_396
timestamp 1607194113
transform 1 0 53820 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_125
timestamp 1607194113
transform 1 0 54004 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_25
timestamp 1607194113
transform 1 0 54372 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_25
timestamp 1607194113
transform 1 0 54464 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_409
timestamp 1607194113
transform 1 0 54740 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_410
timestamp 1607194113
transform 1 0 54832 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_411
timestamp 1607194113
transform 1 0 55568 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_412
timestamp 1607194113
transform 1 0 55936 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_126
timestamp 1607194113
transform 1 0 56120 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_26
timestamp 1607194113
transform 1 0 56488 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_26
timestamp 1607194113
transform 1 0 56580 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_425
timestamp 1607194113
transform 1 0 56856 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_426
timestamp 1607194113
transform 1 0 56948 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_427
timestamp 1607194113
transform 1 0 57684 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_428
timestamp 1607194113
transform 1 0 58052 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_127
timestamp 1607194113
transform 1 0 58236 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_27
timestamp 1607194113
transform 1 0 58604 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_27
timestamp 1607194113
transform 1 0 58696 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_441
timestamp 1607194113
transform 1 0 58972 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_442
timestamp 1607194113
transform 1 0 59064 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_443
timestamp 1607194113
transform 1 0 59800 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_444
timestamp 1607194113
transform 1 0 60168 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_128
timestamp 1607194113
transform 1 0 60352 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_28
timestamp 1607194113
transform 1 0 60720 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_28
timestamp 1607194113
transform 1 0 60812 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_457
timestamp 1607194113
transform 1 0 61088 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_458
timestamp 1607194113
transform 1 0 61180 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_459
timestamp 1607194113
transform 1 0 61916 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_460
timestamp 1607194113
transform 1 0 62284 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_129
timestamp 1607194113
transform 1 0 62468 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_29
timestamp 1607194113
transform 1 0 62836 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_29
timestamp 1607194113
transform 1 0 62928 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_473
timestamp 1607194113
transform 1 0 63204 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_474
timestamp 1607194113
transform 1 0 63296 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_475
timestamp 1607194113
transform 1 0 64032 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_476
timestamp 1607194113
transform 1 0 64400 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_130
timestamp 1607194113
transform 1 0 64584 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_30
timestamp 1607194113
transform 1 0 64952 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_30
timestamp 1607194113
transform 1 0 65044 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_489
timestamp 1607194113
transform 1 0 65320 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_490
timestamp 1607194113
transform 1 0 65412 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_491
timestamp 1607194113
transform 1 0 66148 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_492
timestamp 1607194113
transform 1 0 66516 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_131
timestamp 1607194113
transform 1 0 66700 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_31
timestamp 1607194113
transform 1 0 67068 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_31
timestamp 1607194113
transform 1 0 67160 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_505
timestamp 1607194113
transform 1 0 67436 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_506
timestamp 1607194113
transform 1 0 67528 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_507
timestamp 1607194113
transform 1 0 68264 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_508
timestamp 1607194113
transform 1 0 68632 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_132
timestamp 1607194113
transform 1 0 68816 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_32
timestamp 1607194113
transform 1 0 69184 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_32
timestamp 1607194113
transform 1 0 69276 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_521
timestamp 1607194113
transform 1 0 69552 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_522
timestamp 1607194113
transform 1 0 69644 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_523
timestamp 1607194113
transform 1 0 70380 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_524
timestamp 1607194113
transform 1 0 70748 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_133
timestamp 1607194113
transform 1 0 70932 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_33
timestamp 1607194113
transform 1 0 71300 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_33
timestamp 1607194113
transform 1 0 71392 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_537
timestamp 1607194113
transform 1 0 71668 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_538
timestamp 1607194113
transform 1 0 71760 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_539
timestamp 1607194113
transform 1 0 72496 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_540
timestamp 1607194113
transform 1 0 72864 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_134
timestamp 1607194113
transform 1 0 73048 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_34
timestamp 1607194113
transform 1 0 73416 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_34
timestamp 1607194113
transform 1 0 73508 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_553
timestamp 1607194113
transform 1 0 73784 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_554
timestamp 1607194113
transform 1 0 73876 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_555
timestamp 1607194113
transform 1 0 74612 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_556
timestamp 1607194113
transform 1 0 74980 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_135
timestamp 1607194113
transform 1 0 75164 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_35
timestamp 1607194113
transform 1 0 75532 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_35
timestamp 1607194113
transform 1 0 75624 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_569
timestamp 1607194113
transform 1 0 75900 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_570
timestamp 1607194113
transform 1 0 75992 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_571
timestamp 1607194113
transform 1 0 76728 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_572
timestamp 1607194113
transform 1 0 77096 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_136
timestamp 1607194113
transform 1 0 77280 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_36
timestamp 1607194113
transform 1 0 77648 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_36
timestamp 1607194113
transform 1 0 77740 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_585
timestamp 1607194113
transform 1 0 78016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_586
timestamp 1607194113
transform 1 0 78108 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_587
timestamp 1607194113
transform 1 0 78844 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_588
timestamp 1607194113
transform 1 0 79212 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_137
timestamp 1607194113
transform 1 0 79396 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_37
timestamp 1607194113
transform 1 0 79764 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_37
timestamp 1607194113
transform 1 0 79856 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_601
timestamp 1607194113
transform 1 0 80132 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_602
timestamp 1607194113
transform 1 0 80224 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_603
timestamp 1607194113
transform 1 0 80960 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_604
timestamp 1607194113
transform 1 0 81328 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_138
timestamp 1607194113
transform 1 0 81512 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_38
timestamp 1607194113
transform 1 0 81880 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_38
timestamp 1607194113
transform 1 0 81972 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_617
timestamp 1607194113
transform 1 0 82248 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_618
timestamp 1607194113
transform 1 0 82340 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_619
timestamp 1607194113
transform 1 0 83076 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_620
timestamp 1607194113
transform 1 0 83444 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_139
timestamp 1607194113
transform 1 0 83628 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_39
timestamp 1607194113
transform 1 0 83996 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_39
timestamp 1607194113
transform 1 0 84088 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_633
timestamp 1607194113
transform 1 0 84364 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_634
timestamp 1607194113
transform 1 0 84456 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_635
timestamp 1607194113
transform 1 0 85192 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_636
timestamp 1607194113
transform 1 0 85560 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_140
timestamp 1607194113
transform 1 0 85744 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_40
timestamp 1607194113
transform 1 0 86112 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_40
timestamp 1607194113
transform 1 0 86204 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_649
timestamp 1607194113
transform 1 0 86480 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_650
timestamp 1607194113
transform 1 0 86572 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_651
timestamp 1607194113
transform 1 0 87308 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_652
timestamp 1607194113
transform 1 0 87676 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_141
timestamp 1607194113
transform 1 0 87860 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_41
timestamp 1607194113
transform 1 0 88228 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_41
timestamp 1607194113
transform 1 0 88320 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_665
timestamp 1607194113
transform 1 0 88596 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_666
timestamp 1607194113
transform 1 0 88688 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_667
timestamp 1607194113
transform 1 0 89424 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_668
timestamp 1607194113
transform 1 0 89792 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_142
timestamp 1607194113
transform 1 0 89976 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_42
timestamp 1607194113
transform 1 0 90344 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_42
timestamp 1607194113
transform 1 0 90436 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_681
timestamp 1607194113
transform 1 0 90712 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_682
timestamp 1607194113
transform 1 0 90804 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_683
timestamp 1607194113
transform 1 0 91540 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_684
timestamp 1607194113
transform 1 0 91908 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_143
timestamp 1607194113
transform 1 0 92092 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_43
timestamp 1607194113
transform 1 0 92460 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_43
timestamp 1607194113
transform 1 0 92552 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_697
timestamp 1607194113
transform 1 0 92828 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_698
timestamp 1607194113
transform 1 0 92920 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_699
timestamp 1607194113
transform 1 0 93656 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_700
timestamp 1607194113
transform 1 0 94024 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_144
timestamp 1607194113
transform 1 0 94208 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_44
timestamp 1607194113
transform 1 0 94576 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_44
timestamp 1607194113
transform 1 0 94668 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_713
timestamp 1607194113
transform 1 0 94944 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_714
timestamp 1607194113
transform 1 0 95036 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_715
timestamp 1607194113
transform 1 0 95772 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_716
timestamp 1607194113
transform 1 0 96140 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_145
timestamp 1607194113
transform 1 0 96324 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_45
timestamp 1607194113
transform 1 0 96692 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_45
timestamp 1607194113
transform 1 0 96784 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_729
timestamp 1607194113
transform 1 0 97060 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_730
timestamp 1607194113
transform 1 0 97152 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_731
timestamp 1607194113
transform 1 0 97888 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_732
timestamp 1607194113
transform 1 0 98256 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_146
timestamp 1607194113
transform 1 0 98440 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_46
timestamp 1607194113
transform 1 0 98808 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_46
timestamp 1607194113
transform 1 0 98900 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_745
timestamp 1607194113
transform 1 0 99176 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_746
timestamp 1607194113
transform 1 0 99268 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_747
timestamp 1607194113
transform 1 0 100004 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_748
timestamp 1607194113
transform 1 0 100372 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_147
timestamp 1607194113
transform 1 0 100556 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_47
timestamp 1607194113
transform 1 0 100924 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_47
timestamp 1607194113
transform 1 0 101016 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_761
timestamp 1607194113
transform 1 0 101292 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_762
timestamp 1607194113
transform 1 0 101384 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_763
timestamp 1607194113
transform 1 0 102120 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_764
timestamp 1607194113
transform 1 0 102488 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_148
timestamp 1607194113
transform 1 0 102672 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_48
timestamp 1607194113
transform 1 0 103040 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_48
timestamp 1607194113
transform 1 0 103132 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_777
timestamp 1607194113
transform 1 0 103408 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_778
timestamp 1607194113
transform 1 0 103500 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_779
timestamp 1607194113
transform 1 0 104236 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_780
timestamp 1607194113
transform 1 0 104604 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_149
timestamp 1607194113
transform 1 0 104788 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap8_49
timestamp 1607194113
transform 1 0 105156 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap8_49
timestamp 1607194113
transform 1 0 105248 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_793
timestamp 1607194113
transform 1 0 105524 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_794
timestamp 1607194113
transform 1 0 105616 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_795
timestamp 1607194113
transform 1 0 106352 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_796
timestamp 1607194113
transform 1 0 106720 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_0
timestamp 1607194113
transform 1 0 1104 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_0
timestamp 1607194113
transform 1 0 1196 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_12
timestamp 1607194113
transform 1 0 1472 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_13
timestamp 1607194113
transform 1 0 1564 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_14
timestamp 1607194113
transform 1 0 2300 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_15
timestamp 1607194113
transform 1 0 2392 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILL_16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607194113
transform 1 0 3128 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  delay_198
timestamp 1607194113
transform -1 0 3588 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_1
timestamp 1607194113
transform 1 0 3588 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_1
timestamp 1607194113
transform 1 0 3680 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_29
timestamp 1607194113
transform 1 0 3956 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_30
timestamp 1607194113
transform 1 0 4048 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_31
timestamp 1607194113
transform 1 0 4784 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_32
timestamp 1607194113
transform 1 0 5152 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_197
timestamp 1607194113
transform -1 0 5704 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_2
timestamp 1607194113
transform 1 0 5704 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_2
timestamp 1607194113
transform 1 0 5796 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_45
timestamp 1607194113
transform 1 0 6072 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_46
timestamp 1607194113
transform 1 0 6164 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_47
timestamp 1607194113
transform 1 0 6900 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_48
timestamp 1607194113
transform 1 0 7268 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_196
timestamp 1607194113
transform -1 0 7820 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_3
timestamp 1607194113
transform 1 0 7820 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_3
timestamp 1607194113
transform 1 0 7912 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_61
timestamp 1607194113
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_62
timestamp 1607194113
transform 1 0 8280 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_63
timestamp 1607194113
transform 1 0 9016 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_64
timestamp 1607194113
transform 1 0 9384 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_195
timestamp 1607194113
transform -1 0 9936 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_4
timestamp 1607194113
transform 1 0 9936 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_4
timestamp 1607194113
transform 1 0 10028 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_77
timestamp 1607194113
transform 1 0 10304 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_78
timestamp 1607194113
transform 1 0 10396 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_79
timestamp 1607194113
transform 1 0 11132 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_80
timestamp 1607194113
transform 1 0 11500 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_194
timestamp 1607194113
transform -1 0 12052 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_5
timestamp 1607194113
transform 1 0 12052 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_5
timestamp 1607194113
transform 1 0 12144 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_93
timestamp 1607194113
transform 1 0 12420 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_94
timestamp 1607194113
transform 1 0 12512 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_95
timestamp 1607194113
transform 1 0 13248 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_96
timestamp 1607194113
transform 1 0 13616 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_193
timestamp 1607194113
transform -1 0 14168 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_6
timestamp 1607194113
transform 1 0 14168 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_6
timestamp 1607194113
transform 1 0 14260 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_109
timestamp 1607194113
transform 1 0 14536 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_110
timestamp 1607194113
transform 1 0 14628 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_111
timestamp 1607194113
transform 1 0 15364 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_112
timestamp 1607194113
transform 1 0 15732 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_192
timestamp 1607194113
transform -1 0 16284 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_7
timestamp 1607194113
transform 1 0 16284 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_7
timestamp 1607194113
transform 1 0 16376 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_125
timestamp 1607194113
transform 1 0 16652 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_126
timestamp 1607194113
transform 1 0 16744 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_127
timestamp 1607194113
transform 1 0 17480 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_128
timestamp 1607194113
transform 1 0 17848 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_191
timestamp 1607194113
transform -1 0 18400 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_8
timestamp 1607194113
transform 1 0 18400 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_8
timestamp 1607194113
transform 1 0 18492 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_141
timestamp 1607194113
transform 1 0 18768 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_142
timestamp 1607194113
transform 1 0 18860 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_143
timestamp 1607194113
transform 1 0 19596 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_144
timestamp 1607194113
transform 1 0 19964 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_190
timestamp 1607194113
transform -1 0 20516 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_9
timestamp 1607194113
transform 1 0 20516 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_9
timestamp 1607194113
transform 1 0 20608 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_157
timestamp 1607194113
transform 1 0 20884 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_158
timestamp 1607194113
transform 1 0 20976 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_159
timestamp 1607194113
transform 1 0 21712 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_160
timestamp 1607194113
transform 1 0 22080 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_189
timestamp 1607194113
transform -1 0 22632 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_10
timestamp 1607194113
transform 1 0 22632 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_10
timestamp 1607194113
transform 1 0 22724 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_173
timestamp 1607194113
transform 1 0 23000 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_174
timestamp 1607194113
transform 1 0 23092 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_175
timestamp 1607194113
transform 1 0 23828 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_176
timestamp 1607194113
transform 1 0 24196 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_188
timestamp 1607194113
transform -1 0 24748 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_11
timestamp 1607194113
transform 1 0 24748 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_11
timestamp 1607194113
transform 1 0 24840 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_189
timestamp 1607194113
transform 1 0 25116 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_190
timestamp 1607194113
transform 1 0 25208 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_191
timestamp 1607194113
transform 1 0 25944 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_192
timestamp 1607194113
transform 1 0 26312 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_187
timestamp 1607194113
transform -1 0 26864 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_12
timestamp 1607194113
transform 1 0 26864 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_12
timestamp 1607194113
transform 1 0 26956 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_205
timestamp 1607194113
transform 1 0 27232 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_206
timestamp 1607194113
transform 1 0 27324 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_207
timestamp 1607194113
transform 1 0 28060 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_208
timestamp 1607194113
transform 1 0 28428 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_186
timestamp 1607194113
transform -1 0 28980 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_13
timestamp 1607194113
transform 1 0 28980 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_13
timestamp 1607194113
transform 1 0 29072 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_221
timestamp 1607194113
transform 1 0 29348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_222
timestamp 1607194113
transform 1 0 29440 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_223
timestamp 1607194113
transform 1 0 30176 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_224
timestamp 1607194113
transform 1 0 30544 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_185
timestamp 1607194113
transform -1 0 31096 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_14
timestamp 1607194113
transform 1 0 31096 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_14
timestamp 1607194113
transform 1 0 31188 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_237
timestamp 1607194113
transform 1 0 31464 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_238
timestamp 1607194113
transform 1 0 31556 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_239
timestamp 1607194113
transform 1 0 32292 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_240
timestamp 1607194113
transform 1 0 32660 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_184
timestamp 1607194113
transform -1 0 33212 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_15
timestamp 1607194113
transform 1 0 33212 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_15
timestamp 1607194113
transform 1 0 33304 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_253
timestamp 1607194113
transform 1 0 33580 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_254
timestamp 1607194113
transform 1 0 33672 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_255
timestamp 1607194113
transform 1 0 34408 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_256
timestamp 1607194113
transform 1 0 34776 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_183
timestamp 1607194113
transform -1 0 35328 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_16
timestamp 1607194113
transform 1 0 35328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_16
timestamp 1607194113
transform 1 0 35420 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_269
timestamp 1607194113
transform 1 0 35696 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_270
timestamp 1607194113
transform 1 0 35788 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_271
timestamp 1607194113
transform 1 0 36524 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_272
timestamp 1607194113
transform 1 0 36892 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_182
timestamp 1607194113
transform -1 0 37444 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_17
timestamp 1607194113
transform 1 0 37444 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_17
timestamp 1607194113
transform 1 0 37536 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_285
timestamp 1607194113
transform 1 0 37812 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_286
timestamp 1607194113
transform 1 0 37904 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_287
timestamp 1607194113
transform 1 0 38640 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_288
timestamp 1607194113
transform 1 0 39008 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_181
timestamp 1607194113
transform -1 0 39560 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_18
timestamp 1607194113
transform 1 0 39560 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_18
timestamp 1607194113
transform 1 0 39652 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_301
timestamp 1607194113
transform 1 0 39928 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_302
timestamp 1607194113
transform 1 0 40020 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_303
timestamp 1607194113
transform 1 0 40756 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_304
timestamp 1607194113
transform 1 0 41124 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_180
timestamp 1607194113
transform -1 0 41676 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_19
timestamp 1607194113
transform 1 0 41676 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_19
timestamp 1607194113
transform 1 0 41768 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_317
timestamp 1607194113
transform 1 0 42044 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_318
timestamp 1607194113
transform 1 0 42136 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_319
timestamp 1607194113
transform 1 0 42872 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_320
timestamp 1607194113
transform 1 0 43240 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_179
timestamp 1607194113
transform -1 0 43792 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_20
timestamp 1607194113
transform 1 0 43792 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_20
timestamp 1607194113
transform 1 0 43884 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_333
timestamp 1607194113
transform 1 0 44160 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_334
timestamp 1607194113
transform 1 0 44252 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_335
timestamp 1607194113
transform 1 0 44988 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_336
timestamp 1607194113
transform 1 0 45356 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_178
timestamp 1607194113
transform -1 0 45908 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_21
timestamp 1607194113
transform 1 0 45908 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_21
timestamp 1607194113
transform 1 0 46000 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_349
timestamp 1607194113
transform 1 0 46276 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_350
timestamp 1607194113
transform 1 0 46368 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_351
timestamp 1607194113
transform 1 0 47104 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_352
timestamp 1607194113
transform 1 0 47472 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_177
timestamp 1607194113
transform -1 0 48024 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_22
timestamp 1607194113
transform 1 0 48024 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_22
timestamp 1607194113
transform 1 0 48116 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_365
timestamp 1607194113
transform 1 0 48392 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_366
timestamp 1607194113
transform 1 0 48484 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_367
timestamp 1607194113
transform 1 0 49220 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_368
timestamp 1607194113
transform 1 0 49588 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_176
timestamp 1607194113
transform -1 0 50140 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_23
timestamp 1607194113
transform 1 0 50140 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_23
timestamp 1607194113
transform 1 0 50232 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_381
timestamp 1607194113
transform 1 0 50508 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_382
timestamp 1607194113
transform 1 0 50600 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_383
timestamp 1607194113
transform 1 0 51336 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_384
timestamp 1607194113
transform 1 0 51704 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_175
timestamp 1607194113
transform -1 0 52256 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_24
timestamp 1607194113
transform 1 0 52256 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_24
timestamp 1607194113
transform 1 0 52348 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_397
timestamp 1607194113
transform 1 0 52624 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_398
timestamp 1607194113
transform 1 0 52716 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_399
timestamp 1607194113
transform 1 0 53452 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_400
timestamp 1607194113
transform 1 0 53820 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_174
timestamp 1607194113
transform -1 0 54372 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_25
timestamp 1607194113
transform 1 0 54372 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_25
timestamp 1607194113
transform 1 0 54464 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_413
timestamp 1607194113
transform 1 0 54740 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_414
timestamp 1607194113
transform 1 0 54832 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_415
timestamp 1607194113
transform 1 0 55568 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_416
timestamp 1607194113
transform 1 0 55936 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_173
timestamp 1607194113
transform -1 0 56488 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_26
timestamp 1607194113
transform 1 0 56488 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_26
timestamp 1607194113
transform 1 0 56580 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_429
timestamp 1607194113
transform 1 0 56856 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_430
timestamp 1607194113
transform 1 0 56948 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_431
timestamp 1607194113
transform 1 0 57684 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_432
timestamp 1607194113
transform 1 0 58052 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_172
timestamp 1607194113
transform -1 0 58604 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_27
timestamp 1607194113
transform 1 0 58604 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_27
timestamp 1607194113
transform 1 0 58696 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_445
timestamp 1607194113
transform 1 0 58972 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_446
timestamp 1607194113
transform 1 0 59064 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_447
timestamp 1607194113
transform 1 0 59800 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_448
timestamp 1607194113
transform 1 0 60168 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_171
timestamp 1607194113
transform -1 0 60720 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_28
timestamp 1607194113
transform 1 0 60720 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_28
timestamp 1607194113
transform 1 0 60812 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_461
timestamp 1607194113
transform 1 0 61088 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_462
timestamp 1607194113
transform 1 0 61180 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_463
timestamp 1607194113
transform 1 0 61916 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_464
timestamp 1607194113
transform 1 0 62284 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_170
timestamp 1607194113
transform -1 0 62836 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_29
timestamp 1607194113
transform 1 0 62836 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_29
timestamp 1607194113
transform 1 0 62928 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_477
timestamp 1607194113
transform 1 0 63204 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_478
timestamp 1607194113
transform 1 0 63296 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_479
timestamp 1607194113
transform 1 0 64032 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_480
timestamp 1607194113
transform 1 0 64400 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_169
timestamp 1607194113
transform -1 0 64952 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_30
timestamp 1607194113
transform 1 0 64952 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_30
timestamp 1607194113
transform 1 0 65044 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_493
timestamp 1607194113
transform 1 0 65320 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_494
timestamp 1607194113
transform 1 0 65412 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_495
timestamp 1607194113
transform 1 0 66148 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_496
timestamp 1607194113
transform 1 0 66516 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_168
timestamp 1607194113
transform -1 0 67068 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_31
timestamp 1607194113
transform 1 0 67068 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_31
timestamp 1607194113
transform 1 0 67160 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_509
timestamp 1607194113
transform 1 0 67436 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_510
timestamp 1607194113
transform 1 0 67528 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_511
timestamp 1607194113
transform 1 0 68264 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_512
timestamp 1607194113
transform 1 0 68632 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_167
timestamp 1607194113
transform -1 0 69184 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_32
timestamp 1607194113
transform 1 0 69184 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_32
timestamp 1607194113
transform 1 0 69276 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_525
timestamp 1607194113
transform 1 0 69552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_526
timestamp 1607194113
transform 1 0 69644 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_527
timestamp 1607194113
transform 1 0 70380 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_528
timestamp 1607194113
transform 1 0 70748 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_166
timestamp 1607194113
transform -1 0 71300 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_33
timestamp 1607194113
transform 1 0 71300 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_33
timestamp 1607194113
transform 1 0 71392 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_541
timestamp 1607194113
transform 1 0 71668 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_542
timestamp 1607194113
transform 1 0 71760 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_543
timestamp 1607194113
transform 1 0 72496 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_544
timestamp 1607194113
transform 1 0 72864 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_165
timestamp 1607194113
transform -1 0 73416 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_34
timestamp 1607194113
transform 1 0 73416 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_34
timestamp 1607194113
transform 1 0 73508 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_557
timestamp 1607194113
transform 1 0 73784 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_558
timestamp 1607194113
transform 1 0 73876 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_559
timestamp 1607194113
transform 1 0 74612 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_560
timestamp 1607194113
transform 1 0 74980 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_164
timestamp 1607194113
transform -1 0 75532 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_35
timestamp 1607194113
transform 1 0 75532 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_35
timestamp 1607194113
transform 1 0 75624 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_573
timestamp 1607194113
transform 1 0 75900 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_574
timestamp 1607194113
transform 1 0 75992 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_575
timestamp 1607194113
transform 1 0 76728 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_576
timestamp 1607194113
transform 1 0 77096 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_163
timestamp 1607194113
transform -1 0 77648 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_36
timestamp 1607194113
transform 1 0 77648 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_36
timestamp 1607194113
transform 1 0 77740 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_589
timestamp 1607194113
transform 1 0 78016 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_590
timestamp 1607194113
transform 1 0 78108 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_591
timestamp 1607194113
transform 1 0 78844 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_592
timestamp 1607194113
transform 1 0 79212 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_162
timestamp 1607194113
transform -1 0 79764 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_37
timestamp 1607194113
transform 1 0 79764 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_37
timestamp 1607194113
transform 1 0 79856 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_605
timestamp 1607194113
transform 1 0 80132 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_606
timestamp 1607194113
transform 1 0 80224 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_607
timestamp 1607194113
transform 1 0 80960 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_608
timestamp 1607194113
transform 1 0 81328 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_161
timestamp 1607194113
transform -1 0 81880 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_38
timestamp 1607194113
transform 1 0 81880 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_38
timestamp 1607194113
transform 1 0 81972 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_621
timestamp 1607194113
transform 1 0 82248 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_622
timestamp 1607194113
transform 1 0 82340 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_623
timestamp 1607194113
transform 1 0 83076 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_624
timestamp 1607194113
transform 1 0 83444 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_160
timestamp 1607194113
transform -1 0 83996 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_39
timestamp 1607194113
transform 1 0 83996 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_39
timestamp 1607194113
transform 1 0 84088 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_637
timestamp 1607194113
transform 1 0 84364 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_638
timestamp 1607194113
transform 1 0 84456 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_639
timestamp 1607194113
transform 1 0 85192 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_640
timestamp 1607194113
transform 1 0 85560 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_159
timestamp 1607194113
transform -1 0 86112 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_40
timestamp 1607194113
transform 1 0 86112 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_40
timestamp 1607194113
transform 1 0 86204 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_653
timestamp 1607194113
transform 1 0 86480 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_654
timestamp 1607194113
transform 1 0 86572 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_655
timestamp 1607194113
transform 1 0 87308 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_656
timestamp 1607194113
transform 1 0 87676 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_158
timestamp 1607194113
transform -1 0 88228 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_41
timestamp 1607194113
transform 1 0 88228 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_41
timestamp 1607194113
transform 1 0 88320 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_669
timestamp 1607194113
transform 1 0 88596 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_670
timestamp 1607194113
transform 1 0 88688 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_671
timestamp 1607194113
transform 1 0 89424 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_672
timestamp 1607194113
transform 1 0 89792 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_157
timestamp 1607194113
transform -1 0 90344 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_42
timestamp 1607194113
transform 1 0 90344 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_42
timestamp 1607194113
transform 1 0 90436 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_685
timestamp 1607194113
transform 1 0 90712 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_686
timestamp 1607194113
transform 1 0 90804 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_687
timestamp 1607194113
transform 1 0 91540 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_688
timestamp 1607194113
transform 1 0 91908 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_156
timestamp 1607194113
transform -1 0 92460 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_43
timestamp 1607194113
transform 1 0 92460 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_43
timestamp 1607194113
transform 1 0 92552 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_701
timestamp 1607194113
transform 1 0 92828 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_702
timestamp 1607194113
transform 1 0 92920 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_703
timestamp 1607194113
transform 1 0 93656 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_704
timestamp 1607194113
transform 1 0 94024 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_155
timestamp 1607194113
transform -1 0 94576 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_44
timestamp 1607194113
transform 1 0 94576 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_44
timestamp 1607194113
transform 1 0 94668 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_717
timestamp 1607194113
transform 1 0 94944 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_718
timestamp 1607194113
transform 1 0 95036 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_719
timestamp 1607194113
transform 1 0 95772 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_720
timestamp 1607194113
transform 1 0 96140 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_154
timestamp 1607194113
transform -1 0 96692 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_45
timestamp 1607194113
transform 1 0 96692 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_45
timestamp 1607194113
transform 1 0 96784 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_733
timestamp 1607194113
transform 1 0 97060 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_734
timestamp 1607194113
transform 1 0 97152 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_735
timestamp 1607194113
transform 1 0 97888 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_736
timestamp 1607194113
transform 1 0 98256 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_153
timestamp 1607194113
transform -1 0 98808 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_46
timestamp 1607194113
transform 1 0 98808 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_46
timestamp 1607194113
transform 1 0 98900 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_749
timestamp 1607194113
transform 1 0 99176 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_750
timestamp 1607194113
transform 1 0 99268 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_751
timestamp 1607194113
transform 1 0 100004 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_752
timestamp 1607194113
transform 1 0 100372 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_152
timestamp 1607194113
transform -1 0 100924 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_47
timestamp 1607194113
transform 1 0 100924 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_47
timestamp 1607194113
transform 1 0 101016 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_765
timestamp 1607194113
transform 1 0 101292 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_766
timestamp 1607194113
transform 1 0 101384 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_767
timestamp 1607194113
transform 1 0 102120 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_768
timestamp 1607194113
transform 1 0 102488 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_151
timestamp 1607194113
transform -1 0 103040 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_48
timestamp 1607194113
transform 1 0 103040 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_48
timestamp 1607194113
transform 1 0 103132 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_781
timestamp 1607194113
transform 1 0 103408 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_782
timestamp 1607194113
transform 1 0 103500 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_783
timestamp 1607194113
transform 1 0 104236 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_784
timestamp 1607194113
transform 1 0 104604 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  delay_150
timestamp 1607194113
transform -1 0 105156 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap9_49
timestamp 1607194113
transform 1 0 105156 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap9_49
timestamp 1607194113
transform 1 0 105248 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  FILL_797
timestamp 1607194113
transform 1 0 105524 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_8  FILL_798
timestamp 1607194113
transform 1 0 105616 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_4  FILL_799
timestamp 1607194113
transform 1 0 106352 0 1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILL_800
timestamp 1607194113
transform 1 0 106720 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  dff1_199
timestamp 1607194113
transform 1 0 1104 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_0
timestamp 1607194113
transform 1 0 2852 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_0
timestamp 1607194113
transform 1 0 2944 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_198
timestamp 1607194113
transform 1 0 3220 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_1
timestamp 1607194113
transform 1 0 4968 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_1
timestamp 1607194113
transform 1 0 5060 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_197
timestamp 1607194113
transform 1 0 5336 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_2
timestamp 1607194113
transform 1 0 7084 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_2
timestamp 1607194113
transform 1 0 7176 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_196
timestamp 1607194113
transform 1 0 7452 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_3
timestamp 1607194113
transform 1 0 9200 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_3
timestamp 1607194113
transform 1 0 9292 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_195
timestamp 1607194113
transform 1 0 9568 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_4
timestamp 1607194113
transform 1 0 11316 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_4
timestamp 1607194113
transform 1 0 11408 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_194
timestamp 1607194113
transform 1 0 11684 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_5
timestamp 1607194113
transform 1 0 13432 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_5
timestamp 1607194113
transform 1 0 13524 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_193
timestamp 1607194113
transform 1 0 13800 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_6
timestamp 1607194113
transform 1 0 15548 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_6
timestamp 1607194113
transform 1 0 15640 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_192
timestamp 1607194113
transform 1 0 15916 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_7
timestamp 1607194113
transform 1 0 17664 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_7
timestamp 1607194113
transform 1 0 17756 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_191
timestamp 1607194113
transform 1 0 18032 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_8
timestamp 1607194113
transform 1 0 19780 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_8
timestamp 1607194113
transform 1 0 19872 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_190
timestamp 1607194113
transform 1 0 20148 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_9
timestamp 1607194113
transform 1 0 21896 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_9
timestamp 1607194113
transform 1 0 21988 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_189
timestamp 1607194113
transform 1 0 22264 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_10
timestamp 1607194113
transform 1 0 24012 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_10
timestamp 1607194113
transform 1 0 24104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_188
timestamp 1607194113
transform 1 0 24380 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_11
timestamp 1607194113
transform 1 0 26128 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_11
timestamp 1607194113
transform 1 0 26220 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_187
timestamp 1607194113
transform 1 0 26496 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_12
timestamp 1607194113
transform 1 0 28244 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_12
timestamp 1607194113
transform 1 0 28336 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_186
timestamp 1607194113
transform 1 0 28612 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_13
timestamp 1607194113
transform 1 0 30360 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_13
timestamp 1607194113
transform 1 0 30452 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_185
timestamp 1607194113
transform 1 0 30728 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_14
timestamp 1607194113
transform 1 0 32476 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_14
timestamp 1607194113
transform 1 0 32568 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_184
timestamp 1607194113
transform 1 0 32844 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_15
timestamp 1607194113
transform 1 0 34592 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_15
timestamp 1607194113
transform 1 0 34684 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_183
timestamp 1607194113
transform 1 0 34960 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_16
timestamp 1607194113
transform 1 0 36708 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_16
timestamp 1607194113
transform 1 0 36800 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_182
timestamp 1607194113
transform 1 0 37076 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_17
timestamp 1607194113
transform 1 0 38824 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_17
timestamp 1607194113
transform 1 0 38916 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_181
timestamp 1607194113
transform 1 0 39192 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_18
timestamp 1607194113
transform 1 0 40940 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_18
timestamp 1607194113
transform 1 0 41032 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_180
timestamp 1607194113
transform 1 0 41308 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_19
timestamp 1607194113
transform 1 0 43056 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_19
timestamp 1607194113
transform 1 0 43148 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_179
timestamp 1607194113
transform 1 0 43424 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_20
timestamp 1607194113
transform 1 0 45172 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_20
timestamp 1607194113
transform 1 0 45264 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_178
timestamp 1607194113
transform 1 0 45540 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_21
timestamp 1607194113
transform 1 0 47288 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_21
timestamp 1607194113
transform 1 0 47380 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_177
timestamp 1607194113
transform 1 0 47656 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_22
timestamp 1607194113
transform 1 0 49404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_22
timestamp 1607194113
transform 1 0 49496 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_176
timestamp 1607194113
transform 1 0 49772 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_23
timestamp 1607194113
transform 1 0 51520 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_23
timestamp 1607194113
transform 1 0 51612 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_175
timestamp 1607194113
transform 1 0 51888 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_24
timestamp 1607194113
transform 1 0 53636 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_24
timestamp 1607194113
transform 1 0 53728 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_174
timestamp 1607194113
transform 1 0 54004 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_25
timestamp 1607194113
transform 1 0 55752 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_25
timestamp 1607194113
transform 1 0 55844 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_173
timestamp 1607194113
transform 1 0 56120 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_26
timestamp 1607194113
transform 1 0 57868 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_26
timestamp 1607194113
transform 1 0 57960 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_172
timestamp 1607194113
transform 1 0 58236 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_27
timestamp 1607194113
transform 1 0 59984 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_27
timestamp 1607194113
transform 1 0 60076 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_171
timestamp 1607194113
transform 1 0 60352 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_28
timestamp 1607194113
transform 1 0 62100 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_28
timestamp 1607194113
transform 1 0 62192 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_170
timestamp 1607194113
transform 1 0 62468 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_29
timestamp 1607194113
transform 1 0 64216 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_29
timestamp 1607194113
transform 1 0 64308 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_169
timestamp 1607194113
transform 1 0 64584 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_30
timestamp 1607194113
transform 1 0 66332 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_30
timestamp 1607194113
transform 1 0 66424 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_168
timestamp 1607194113
transform 1 0 66700 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_31
timestamp 1607194113
transform 1 0 68448 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_31
timestamp 1607194113
transform 1 0 68540 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_167
timestamp 1607194113
transform 1 0 68816 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_32
timestamp 1607194113
transform 1 0 70564 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_32
timestamp 1607194113
transform 1 0 70656 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_166
timestamp 1607194113
transform 1 0 70932 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_33
timestamp 1607194113
transform 1 0 72680 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_33
timestamp 1607194113
transform 1 0 72772 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_165
timestamp 1607194113
transform 1 0 73048 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_34
timestamp 1607194113
transform 1 0 74796 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_34
timestamp 1607194113
transform 1 0 74888 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_164
timestamp 1607194113
transform 1 0 75164 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_35
timestamp 1607194113
transform 1 0 76912 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_35
timestamp 1607194113
transform 1 0 77004 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_163
timestamp 1607194113
transform 1 0 77280 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_36
timestamp 1607194113
transform 1 0 79028 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_36
timestamp 1607194113
transform 1 0 79120 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_162
timestamp 1607194113
transform 1 0 79396 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_37
timestamp 1607194113
transform 1 0 81144 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_37
timestamp 1607194113
transform 1 0 81236 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_161
timestamp 1607194113
transform 1 0 81512 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_38
timestamp 1607194113
transform 1 0 83260 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_38
timestamp 1607194113
transform 1 0 83352 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_160
timestamp 1607194113
transform 1 0 83628 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_39
timestamp 1607194113
transform 1 0 85376 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_39
timestamp 1607194113
transform 1 0 85468 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_159
timestamp 1607194113
transform 1 0 85744 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_40
timestamp 1607194113
transform 1 0 87492 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_40
timestamp 1607194113
transform 1 0 87584 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_158
timestamp 1607194113
transform 1 0 87860 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_41
timestamp 1607194113
transform 1 0 89608 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_41
timestamp 1607194113
transform 1 0 89700 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_157
timestamp 1607194113
transform 1 0 89976 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_42
timestamp 1607194113
transform 1 0 91724 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_42
timestamp 1607194113
transform 1 0 91816 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_156
timestamp 1607194113
transform 1 0 92092 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_43
timestamp 1607194113
transform 1 0 93840 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_43
timestamp 1607194113
transform 1 0 93932 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_155
timestamp 1607194113
transform 1 0 94208 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_44
timestamp 1607194113
transform 1 0 95956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_44
timestamp 1607194113
transform 1 0 96048 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_154
timestamp 1607194113
transform 1 0 96324 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_45
timestamp 1607194113
transform 1 0 98072 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_45
timestamp 1607194113
transform 1 0 98164 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_153
timestamp 1607194113
transform 1 0 98440 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_46
timestamp 1607194113
transform 1 0 100188 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_46
timestamp 1607194113
transform 1 0 100280 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_152
timestamp 1607194113
transform 1 0 100556 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_47
timestamp 1607194113
transform 1 0 102304 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_47
timestamp 1607194113
transform 1 0 102396 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_151
timestamp 1607194113
transform 1 0 102672 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_48
timestamp 1607194113
transform 1 0 104420 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_48
timestamp 1607194113
transform 1 0 104512 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff1_150
timestamp 1607194113
transform 1 0 104788 0 -1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap10_49
timestamp 1607194113
transform 1 0 106536 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap10_49
timestamp 1607194113
transform 1 0 106628 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_199
timestamp 1607194113
transform 1 0 1104 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_0
timestamp 1607194113
transform 1 0 2852 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_0
timestamp 1607194113
transform 1 0 2944 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_198
timestamp 1607194113
transform 1 0 3220 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_1
timestamp 1607194113
transform 1 0 4968 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_1
timestamp 1607194113
transform 1 0 5060 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_197
timestamp 1607194113
transform 1 0 5336 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_2
timestamp 1607194113
transform 1 0 7084 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_2
timestamp 1607194113
transform 1 0 7176 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_196
timestamp 1607194113
transform 1 0 7452 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_3
timestamp 1607194113
transform 1 0 9200 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_3
timestamp 1607194113
transform 1 0 9292 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_195
timestamp 1607194113
transform 1 0 9568 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_4
timestamp 1607194113
transform 1 0 11316 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_4
timestamp 1607194113
transform 1 0 11408 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_194
timestamp 1607194113
transform 1 0 11684 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_5
timestamp 1607194113
transform 1 0 13432 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_5
timestamp 1607194113
transform 1 0 13524 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_193
timestamp 1607194113
transform 1 0 13800 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_6
timestamp 1607194113
transform 1 0 15548 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_6
timestamp 1607194113
transform 1 0 15640 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_192
timestamp 1607194113
transform 1 0 15916 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_7
timestamp 1607194113
transform 1 0 17664 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_7
timestamp 1607194113
transform 1 0 17756 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_191
timestamp 1607194113
transform 1 0 18032 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_8
timestamp 1607194113
transform 1 0 19780 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_8
timestamp 1607194113
transform 1 0 19872 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_190
timestamp 1607194113
transform 1 0 20148 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_9
timestamp 1607194113
transform 1 0 21896 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_9
timestamp 1607194113
transform 1 0 21988 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_189
timestamp 1607194113
transform 1 0 22264 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_10
timestamp 1607194113
transform 1 0 24012 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_10
timestamp 1607194113
transform 1 0 24104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_188
timestamp 1607194113
transform 1 0 24380 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_11
timestamp 1607194113
transform 1 0 26128 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_11
timestamp 1607194113
transform 1 0 26220 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_187
timestamp 1607194113
transform 1 0 26496 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_12
timestamp 1607194113
transform 1 0 28244 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_12
timestamp 1607194113
transform 1 0 28336 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_186
timestamp 1607194113
transform 1 0 28612 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_13
timestamp 1607194113
transform 1 0 30360 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_13
timestamp 1607194113
transform 1 0 30452 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_185
timestamp 1607194113
transform 1 0 30728 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_14
timestamp 1607194113
transform 1 0 32476 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_14
timestamp 1607194113
transform 1 0 32568 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_184
timestamp 1607194113
transform 1 0 32844 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_15
timestamp 1607194113
transform 1 0 34592 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_15
timestamp 1607194113
transform 1 0 34684 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_183
timestamp 1607194113
transform 1 0 34960 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_16
timestamp 1607194113
transform 1 0 36708 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_16
timestamp 1607194113
transform 1 0 36800 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_182
timestamp 1607194113
transform 1 0 37076 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_17
timestamp 1607194113
transform 1 0 38824 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_17
timestamp 1607194113
transform 1 0 38916 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_181
timestamp 1607194113
transform 1 0 39192 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_18
timestamp 1607194113
transform 1 0 40940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_18
timestamp 1607194113
transform 1 0 41032 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_180
timestamp 1607194113
transform 1 0 41308 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_19
timestamp 1607194113
transform 1 0 43056 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_19
timestamp 1607194113
transform 1 0 43148 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_179
timestamp 1607194113
transform 1 0 43424 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_20
timestamp 1607194113
transform 1 0 45172 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_20
timestamp 1607194113
transform 1 0 45264 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_178
timestamp 1607194113
transform 1 0 45540 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_21
timestamp 1607194113
transform 1 0 47288 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_21
timestamp 1607194113
transform 1 0 47380 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_177
timestamp 1607194113
transform 1 0 47656 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_22
timestamp 1607194113
transform 1 0 49404 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_22
timestamp 1607194113
transform 1 0 49496 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_176
timestamp 1607194113
transform 1 0 49772 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_23
timestamp 1607194113
transform 1 0 51520 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_23
timestamp 1607194113
transform 1 0 51612 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_175
timestamp 1607194113
transform 1 0 51888 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_24
timestamp 1607194113
transform 1 0 53636 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_24
timestamp 1607194113
transform 1 0 53728 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_174
timestamp 1607194113
transform 1 0 54004 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_25
timestamp 1607194113
transform 1 0 55752 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_25
timestamp 1607194113
transform 1 0 55844 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_173
timestamp 1607194113
transform 1 0 56120 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_26
timestamp 1607194113
transform 1 0 57868 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_26
timestamp 1607194113
transform 1 0 57960 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_172
timestamp 1607194113
transform 1 0 58236 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_27
timestamp 1607194113
transform 1 0 59984 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_27
timestamp 1607194113
transform 1 0 60076 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_171
timestamp 1607194113
transform 1 0 60352 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_28
timestamp 1607194113
transform 1 0 62100 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_28
timestamp 1607194113
transform 1 0 62192 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_170
timestamp 1607194113
transform 1 0 62468 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_29
timestamp 1607194113
transform 1 0 64216 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_29
timestamp 1607194113
transform 1 0 64308 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_169
timestamp 1607194113
transform 1 0 64584 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_30
timestamp 1607194113
transform 1 0 66332 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_30
timestamp 1607194113
transform 1 0 66424 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_168
timestamp 1607194113
transform 1 0 66700 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_31
timestamp 1607194113
transform 1 0 68448 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_31
timestamp 1607194113
transform 1 0 68540 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_167
timestamp 1607194113
transform 1 0 68816 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_32
timestamp 1607194113
transform 1 0 70564 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_32
timestamp 1607194113
transform 1 0 70656 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_166
timestamp 1607194113
transform 1 0 70932 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_33
timestamp 1607194113
transform 1 0 72680 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_33
timestamp 1607194113
transform 1 0 72772 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_165
timestamp 1607194113
transform 1 0 73048 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_34
timestamp 1607194113
transform 1 0 74796 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_34
timestamp 1607194113
transform 1 0 74888 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_164
timestamp 1607194113
transform 1 0 75164 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_35
timestamp 1607194113
transform 1 0 76912 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_35
timestamp 1607194113
transform 1 0 77004 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_163
timestamp 1607194113
transform 1 0 77280 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_36
timestamp 1607194113
transform 1 0 79028 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_36
timestamp 1607194113
transform 1 0 79120 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_162
timestamp 1607194113
transform 1 0 79396 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_37
timestamp 1607194113
transform 1 0 81144 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_37
timestamp 1607194113
transform 1 0 81236 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_161
timestamp 1607194113
transform 1 0 81512 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_38
timestamp 1607194113
transform 1 0 83260 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_38
timestamp 1607194113
transform 1 0 83352 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_160
timestamp 1607194113
transform 1 0 83628 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_39
timestamp 1607194113
transform 1 0 85376 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_39
timestamp 1607194113
transform 1 0 85468 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_159
timestamp 1607194113
transform 1 0 85744 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_40
timestamp 1607194113
transform 1 0 87492 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_40
timestamp 1607194113
transform 1 0 87584 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_158
timestamp 1607194113
transform 1 0 87860 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_41
timestamp 1607194113
transform 1 0 89608 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_41
timestamp 1607194113
transform 1 0 89700 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_157
timestamp 1607194113
transform 1 0 89976 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_42
timestamp 1607194113
transform 1 0 91724 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_42
timestamp 1607194113
transform 1 0 91816 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_156
timestamp 1607194113
transform 1 0 92092 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_43
timestamp 1607194113
transform 1 0 93840 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_43
timestamp 1607194113
transform 1 0 93932 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_155
timestamp 1607194113
transform 1 0 94208 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_44
timestamp 1607194113
transform 1 0 95956 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_44
timestamp 1607194113
transform 1 0 96048 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_154
timestamp 1607194113
transform 1 0 96324 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_45
timestamp 1607194113
transform 1 0 98072 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_45
timestamp 1607194113
transform 1 0 98164 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_153
timestamp 1607194113
transform 1 0 98440 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_46
timestamp 1607194113
transform 1 0 100188 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_46
timestamp 1607194113
transform 1 0 100280 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_152
timestamp 1607194113
transform 1 0 100556 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_47
timestamp 1607194113
transform 1 0 102304 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_47
timestamp 1607194113
transform 1 0 102396 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_151
timestamp 1607194113
transform 1 0 102672 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_48
timestamp 1607194113
transform 1 0 104420 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_48
timestamp 1607194113
transform 1 0 104512 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  dff2_150
timestamp 1607194113
transform 1 0 104788 0 1 7072
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  tap11_49
timestamp 1607194113
transform 1 0 106536 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  decap11_49
timestamp 1607194113
transform 1 0 106628 0 1 7072
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 2048 120 2168 6 inp_i
port 0 nsew default input
rlabel metal2 s 1030 0 1086 56 6 tap_o[0]
port 1 nsew default tristate
rlabel metal2 s 3146 0 3202 56 6 tap_o[1]
port 2 nsew default tristate
rlabel metal2 s 5262 0 5318 56 6 tap_o[2]
port 3 nsew default tristate
rlabel metal2 s 7378 0 7434 56 6 tap_o[3]
port 4 nsew default tristate
rlabel metal2 s 9494 0 9550 56 6 tap_o[4]
port 5 nsew default tristate
rlabel metal2 s 11610 0 11666 56 6 tap_o[5]
port 6 nsew default tristate
rlabel metal2 s 13726 0 13782 56 6 tap_o[6]
port 7 nsew default tristate
rlabel metal2 s 15842 0 15898 56 6 tap_o[7]
port 8 nsew default tristate
rlabel metal2 s 17958 0 18014 56 6 tap_o[8]
port 9 nsew default tristate
rlabel metal2 s 20074 0 20130 56 6 tap_o[9]
port 10 nsew default tristate
rlabel metal2 s 22190 0 22246 56 6 tap_o[10]
port 11 nsew default tristate
rlabel metal2 s 24306 0 24362 56 6 tap_o[11]
port 12 nsew default tristate
rlabel metal2 s 26422 0 26478 56 6 tap_o[12]
port 13 nsew default tristate
rlabel metal2 s 28538 0 28594 56 6 tap_o[13]
port 14 nsew default tristate
rlabel metal2 s 30654 0 30710 56 6 tap_o[14]
port 15 nsew default tristate
rlabel metal2 s 32770 0 32826 56 6 tap_o[15]
port 16 nsew default tristate
rlabel metal2 s 34886 0 34942 56 6 tap_o[16]
port 17 nsew default tristate
rlabel metal2 s 37002 0 37058 56 6 tap_o[17]
port 18 nsew default tristate
rlabel metal2 s 39118 0 39174 56 6 tap_o[18]
port 19 nsew default tristate
rlabel metal2 s 41234 0 41290 56 6 tap_o[19]
port 20 nsew default tristate
rlabel metal2 s 43350 0 43406 56 6 tap_o[20]
port 21 nsew default tristate
rlabel metal2 s 45466 0 45522 56 6 tap_o[21]
port 22 nsew default tristate
rlabel metal2 s 47582 0 47638 56 6 tap_o[22]
port 23 nsew default tristate
rlabel metal2 s 49698 0 49754 56 6 tap_o[23]
port 24 nsew default tristate
rlabel metal2 s 51814 0 51870 56 6 tap_o[24]
port 25 nsew default tristate
rlabel metal2 s 53930 0 53986 56 6 tap_o[25]
port 26 nsew default tristate
rlabel metal2 s 56046 0 56102 56 6 tap_o[26]
port 27 nsew default tristate
rlabel metal2 s 58162 0 58218 56 6 tap_o[27]
port 28 nsew default tristate
rlabel metal2 s 60278 0 60334 56 6 tap_o[28]
port 29 nsew default tristate
rlabel metal2 s 62394 0 62450 56 6 tap_o[29]
port 30 nsew default tristate
rlabel metal2 s 64510 0 64566 56 6 tap_o[30]
port 31 nsew default tristate
rlabel metal2 s 66626 0 66682 56 6 tap_o[31]
port 32 nsew default tristate
rlabel metal2 s 68742 0 68798 56 6 tap_o[32]
port 33 nsew default tristate
rlabel metal2 s 70858 0 70914 56 6 tap_o[33]
port 34 nsew default tristate
rlabel metal2 s 72974 0 73030 56 6 tap_o[34]
port 35 nsew default tristate
rlabel metal2 s 75090 0 75146 56 6 tap_o[35]
port 36 nsew default tristate
rlabel metal2 s 77206 0 77262 56 6 tap_o[36]
port 37 nsew default tristate
rlabel metal2 s 79322 0 79378 56 6 tap_o[37]
port 38 nsew default tristate
rlabel metal2 s 81438 0 81494 56 6 tap_o[38]
port 39 nsew default tristate
rlabel metal2 s 83554 0 83610 56 6 tap_o[39]
port 40 nsew default tristate
rlabel metal2 s 85670 0 85726 56 6 tap_o[40]
port 41 nsew default tristate
rlabel metal2 s 87786 0 87842 56 6 tap_o[41]
port 42 nsew default tristate
rlabel metal2 s 89902 0 89958 56 6 tap_o[42]
port 43 nsew default tristate
rlabel metal2 s 92018 0 92074 56 6 tap_o[43]
port 44 nsew default tristate
rlabel metal2 s 94134 0 94190 56 6 tap_o[44]
port 45 nsew default tristate
rlabel metal2 s 96250 0 96306 56 6 tap_o[45]
port 46 nsew default tristate
rlabel metal2 s 98366 0 98422 56 6 tap_o[46]
port 47 nsew default tristate
rlabel metal2 s 100482 0 100538 56 6 tap_o[47]
port 48 nsew default tristate
rlabel metal2 s 102598 0 102654 56 6 tap_o[48]
port 49 nsew default tristate
rlabel metal2 s 104714 0 104770 56 6 tap_o[49]
port 50 nsew default tristate
rlabel metal2 s 105174 0 105230 56 6 tap_o[50]
port 51 nsew default tristate
rlabel metal2 s 103058 0 103114 56 6 tap_o[51]
port 52 nsew default tristate
rlabel metal2 s 100942 0 100998 56 6 tap_o[52]
port 53 nsew default tristate
rlabel metal2 s 98826 0 98882 56 6 tap_o[53]
port 54 nsew default tristate
rlabel metal2 s 96710 0 96766 56 6 tap_o[54]
port 55 nsew default tristate
rlabel metal2 s 94594 0 94650 56 6 tap_o[55]
port 56 nsew default tristate
rlabel metal2 s 92478 0 92534 56 6 tap_o[56]
port 57 nsew default tristate
rlabel metal2 s 90362 0 90418 56 6 tap_o[57]
port 58 nsew default tristate
rlabel metal2 s 88246 0 88302 56 6 tap_o[58]
port 59 nsew default tristate
rlabel metal2 s 86130 0 86186 56 6 tap_o[59]
port 60 nsew default tristate
rlabel metal2 s 84014 0 84070 56 6 tap_o[60]
port 61 nsew default tristate
rlabel metal2 s 81898 0 81954 56 6 tap_o[61]
port 62 nsew default tristate
rlabel metal2 s 79782 0 79838 56 6 tap_o[62]
port 63 nsew default tristate
rlabel metal2 s 77666 0 77722 56 6 tap_o[63]
port 64 nsew default tristate
rlabel metal2 s 75550 0 75606 56 6 tap_o[64]
port 65 nsew default tristate
rlabel metal2 s 73434 0 73490 56 6 tap_o[65]
port 66 nsew default tristate
rlabel metal2 s 71318 0 71374 56 6 tap_o[66]
port 67 nsew default tristate
rlabel metal2 s 69202 0 69258 56 6 tap_o[67]
port 68 nsew default tristate
rlabel metal2 s 67086 0 67142 56 6 tap_o[68]
port 69 nsew default tristate
rlabel metal2 s 64970 0 65026 56 6 tap_o[69]
port 70 nsew default tristate
rlabel metal2 s 62854 0 62910 56 6 tap_o[70]
port 71 nsew default tristate
rlabel metal2 s 60738 0 60794 56 6 tap_o[71]
port 72 nsew default tristate
rlabel metal2 s 58622 0 58678 56 6 tap_o[72]
port 73 nsew default tristate
rlabel metal2 s 56506 0 56562 56 6 tap_o[73]
port 74 nsew default tristate
rlabel metal2 s 54390 0 54446 56 6 tap_o[74]
port 75 nsew default tristate
rlabel metal2 s 52274 0 52330 56 6 tap_o[75]
port 76 nsew default tristate
rlabel metal2 s 50158 0 50214 56 6 tap_o[76]
port 77 nsew default tristate
rlabel metal2 s 48042 0 48098 56 6 tap_o[77]
port 78 nsew default tristate
rlabel metal2 s 45926 0 45982 56 6 tap_o[78]
port 79 nsew default tristate
rlabel metal2 s 43810 0 43866 56 6 tap_o[79]
port 80 nsew default tristate
rlabel metal2 s 41694 0 41750 56 6 tap_o[80]
port 81 nsew default tristate
rlabel metal2 s 39578 0 39634 56 6 tap_o[81]
port 82 nsew default tristate
rlabel metal2 s 37462 0 37518 56 6 tap_o[82]
port 83 nsew default tristate
rlabel metal2 s 35346 0 35402 56 6 tap_o[83]
port 84 nsew default tristate
rlabel metal2 s 33230 0 33286 56 6 tap_o[84]
port 85 nsew default tristate
rlabel metal2 s 31114 0 31170 56 6 tap_o[85]
port 86 nsew default tristate
rlabel metal2 s 28998 0 29054 56 6 tap_o[86]
port 87 nsew default tristate
rlabel metal2 s 26882 0 26938 56 6 tap_o[87]
port 88 nsew default tristate
rlabel metal2 s 24766 0 24822 56 6 tap_o[88]
port 89 nsew default tristate
rlabel metal2 s 22650 0 22706 56 6 tap_o[89]
port 90 nsew default tristate
rlabel metal2 s 20534 0 20590 56 6 tap_o[90]
port 91 nsew default tristate
rlabel metal2 s 18418 0 18474 56 6 tap_o[91]
port 92 nsew default tristate
rlabel metal2 s 16302 0 16358 56 6 tap_o[92]
port 93 nsew default tristate
rlabel metal2 s 14186 0 14242 56 6 tap_o[93]
port 94 nsew default tristate
rlabel metal2 s 12070 0 12126 56 6 tap_o[94]
port 95 nsew default tristate
rlabel metal2 s 9954 0 10010 56 6 tap_o[95]
port 96 nsew default tristate
rlabel metal2 s 7838 0 7894 56 6 tap_o[96]
port 97 nsew default tristate
rlabel metal2 s 5722 0 5778 56 6 tap_o[97]
port 98 nsew default tristate
rlabel metal2 s 3606 0 3662 56 6 tap_o[98]
port 99 nsew default tristate
rlabel metal2 s 1490 0 1546 56 6 tap_o[99]
port 100 nsew default tristate
rlabel metal2 s 1950 0 2006 56 6 tap_o[100]
port 101 nsew default tristate
rlabel metal2 s 4066 0 4122 56 6 tap_o[101]
port 102 nsew default tristate
rlabel metal2 s 6182 0 6238 56 6 tap_o[102]
port 103 nsew default tristate
rlabel metal2 s 8298 0 8354 56 6 tap_o[103]
port 104 nsew default tristate
rlabel metal2 s 10414 0 10470 56 6 tap_o[104]
port 105 nsew default tristate
rlabel metal2 s 12530 0 12586 56 6 tap_o[105]
port 106 nsew default tristate
rlabel metal2 s 14646 0 14702 56 6 tap_o[106]
port 107 nsew default tristate
rlabel metal2 s 16762 0 16818 56 6 tap_o[107]
port 108 nsew default tristate
rlabel metal2 s 18878 0 18934 56 6 tap_o[108]
port 109 nsew default tristate
rlabel metal2 s 20994 0 21050 56 6 tap_o[109]
port 110 nsew default tristate
rlabel metal2 s 23110 0 23166 56 6 tap_o[110]
port 111 nsew default tristate
rlabel metal2 s 25226 0 25282 56 6 tap_o[111]
port 112 nsew default tristate
rlabel metal2 s 27342 0 27398 56 6 tap_o[112]
port 113 nsew default tristate
rlabel metal2 s 29458 0 29514 56 6 tap_o[113]
port 114 nsew default tristate
rlabel metal2 s 31574 0 31630 56 6 tap_o[114]
port 115 nsew default tristate
rlabel metal2 s 33690 0 33746 56 6 tap_o[115]
port 116 nsew default tristate
rlabel metal2 s 35806 0 35862 56 6 tap_o[116]
port 117 nsew default tristate
rlabel metal2 s 37922 0 37978 56 6 tap_o[117]
port 118 nsew default tristate
rlabel metal2 s 40038 0 40094 56 6 tap_o[118]
port 119 nsew default tristate
rlabel metal2 s 42154 0 42210 56 6 tap_o[119]
port 120 nsew default tristate
rlabel metal2 s 44270 0 44326 56 6 tap_o[120]
port 121 nsew default tristate
rlabel metal2 s 46386 0 46442 56 6 tap_o[121]
port 122 nsew default tristate
rlabel metal2 s 48502 0 48558 56 6 tap_o[122]
port 123 nsew default tristate
rlabel metal2 s 50618 0 50674 56 6 tap_o[123]
port 124 nsew default tristate
rlabel metal2 s 52734 0 52790 56 6 tap_o[124]
port 125 nsew default tristate
rlabel metal2 s 54850 0 54906 56 6 tap_o[125]
port 126 nsew default tristate
rlabel metal2 s 56966 0 57022 56 6 tap_o[126]
port 127 nsew default tristate
rlabel metal2 s 59082 0 59138 56 6 tap_o[127]
port 128 nsew default tristate
rlabel metal2 s 61198 0 61254 56 6 tap_o[128]
port 129 nsew default tristate
rlabel metal2 s 63314 0 63370 56 6 tap_o[129]
port 130 nsew default tristate
rlabel metal2 s 65430 0 65486 56 6 tap_o[130]
port 131 nsew default tristate
rlabel metal2 s 67546 0 67602 56 6 tap_o[131]
port 132 nsew default tristate
rlabel metal2 s 69662 0 69718 56 6 tap_o[132]
port 133 nsew default tristate
rlabel metal2 s 71778 0 71834 56 6 tap_o[133]
port 134 nsew default tristate
rlabel metal2 s 73894 0 73950 56 6 tap_o[134]
port 135 nsew default tristate
rlabel metal2 s 76010 0 76066 56 6 tap_o[135]
port 136 nsew default tristate
rlabel metal2 s 78126 0 78182 56 6 tap_o[136]
port 137 nsew default tristate
rlabel metal2 s 80242 0 80298 56 6 tap_o[137]
port 138 nsew default tristate
rlabel metal2 s 82358 0 82414 56 6 tap_o[138]
port 139 nsew default tristate
rlabel metal2 s 84474 0 84530 56 6 tap_o[139]
port 140 nsew default tristate
rlabel metal2 s 86590 0 86646 56 6 tap_o[140]
port 141 nsew default tristate
rlabel metal2 s 88706 0 88762 56 6 tap_o[141]
port 142 nsew default tristate
rlabel metal2 s 90822 0 90878 56 6 tap_o[142]
port 143 nsew default tristate
rlabel metal2 s 92938 0 92994 56 6 tap_o[143]
port 144 nsew default tristate
rlabel metal2 s 95054 0 95110 56 6 tap_o[144]
port 145 nsew default tristate
rlabel metal2 s 97170 0 97226 56 6 tap_o[145]
port 146 nsew default tristate
rlabel metal2 s 99286 0 99342 56 6 tap_o[146]
port 147 nsew default tristate
rlabel metal2 s 101402 0 101458 56 6 tap_o[147]
port 148 nsew default tristate
rlabel metal2 s 103518 0 103574 56 6 tap_o[148]
port 149 nsew default tristate
rlabel metal2 s 105634 0 105690 56 6 tap_o[149]
port 150 nsew default tristate
rlabel metal2 s 106002 0 106058 56 6 tap_o[150]
port 151 nsew default tristate
rlabel metal2 s 103886 0 103942 56 6 tap_o[151]
port 152 nsew default tristate
rlabel metal2 s 101770 0 101826 56 6 tap_o[152]
port 153 nsew default tristate
rlabel metal2 s 99654 0 99710 56 6 tap_o[153]
port 154 nsew default tristate
rlabel metal2 s 97538 0 97594 56 6 tap_o[154]
port 155 nsew default tristate
rlabel metal2 s 95422 0 95478 56 6 tap_o[155]
port 156 nsew default tristate
rlabel metal2 s 93306 0 93362 56 6 tap_o[156]
port 157 nsew default tristate
rlabel metal2 s 91190 0 91246 56 6 tap_o[157]
port 158 nsew default tristate
rlabel metal2 s 89074 0 89130 56 6 tap_o[158]
port 159 nsew default tristate
rlabel metal2 s 86958 0 87014 56 6 tap_o[159]
port 160 nsew default tristate
rlabel metal2 s 84842 0 84898 56 6 tap_o[160]
port 161 nsew default tristate
rlabel metal2 s 82726 0 82782 56 6 tap_o[161]
port 162 nsew default tristate
rlabel metal2 s 80610 0 80666 56 6 tap_o[162]
port 163 nsew default tristate
rlabel metal2 s 78494 0 78550 56 6 tap_o[163]
port 164 nsew default tristate
rlabel metal2 s 76378 0 76434 56 6 tap_o[164]
port 165 nsew default tristate
rlabel metal2 s 74262 0 74318 56 6 tap_o[165]
port 166 nsew default tristate
rlabel metal2 s 72146 0 72202 56 6 tap_o[166]
port 167 nsew default tristate
rlabel metal2 s 70030 0 70086 56 6 tap_o[167]
port 168 nsew default tristate
rlabel metal2 s 67914 0 67970 56 6 tap_o[168]
port 169 nsew default tristate
rlabel metal2 s 65798 0 65854 56 6 tap_o[169]
port 170 nsew default tristate
rlabel metal2 s 63682 0 63738 56 6 tap_o[170]
port 171 nsew default tristate
rlabel metal2 s 61566 0 61622 56 6 tap_o[171]
port 172 nsew default tristate
rlabel metal2 s 59450 0 59506 56 6 tap_o[172]
port 173 nsew default tristate
rlabel metal2 s 57334 0 57390 56 6 tap_o[173]
port 174 nsew default tristate
rlabel metal2 s 55218 0 55274 56 6 tap_o[174]
port 175 nsew default tristate
rlabel metal2 s 53102 0 53158 56 6 tap_o[175]
port 176 nsew default tristate
rlabel metal2 s 50986 0 51042 56 6 tap_o[176]
port 177 nsew default tristate
rlabel metal2 s 48870 0 48926 56 6 tap_o[177]
port 178 nsew default tristate
rlabel metal2 s 46754 0 46810 56 6 tap_o[178]
port 179 nsew default tristate
rlabel metal2 s 44638 0 44694 56 6 tap_o[179]
port 180 nsew default tristate
rlabel metal2 s 42522 0 42578 56 6 tap_o[180]
port 181 nsew default tristate
rlabel metal2 s 40406 0 40462 56 6 tap_o[181]
port 182 nsew default tristate
rlabel metal2 s 38290 0 38346 56 6 tap_o[182]
port 183 nsew default tristate
rlabel metal2 s 36174 0 36230 56 6 tap_o[183]
port 184 nsew default tristate
rlabel metal2 s 34058 0 34114 56 6 tap_o[184]
port 185 nsew default tristate
rlabel metal2 s 31942 0 31998 56 6 tap_o[185]
port 186 nsew default tristate
rlabel metal2 s 29826 0 29882 56 6 tap_o[186]
port 187 nsew default tristate
rlabel metal2 s 27710 0 27766 56 6 tap_o[187]
port 188 nsew default tristate
rlabel metal2 s 25594 0 25650 56 6 tap_o[188]
port 189 nsew default tristate
rlabel metal2 s 23478 0 23534 56 6 tap_o[189]
port 190 nsew default tristate
rlabel metal2 s 21362 0 21418 56 6 tap_o[190]
port 191 nsew default tristate
rlabel metal2 s 19246 0 19302 56 6 tap_o[191]
port 192 nsew default tristate
rlabel metal2 s 17130 0 17186 56 6 tap_o[192]
port 193 nsew default tristate
rlabel metal2 s 15014 0 15070 56 6 tap_o[193]
port 194 nsew default tristate
rlabel metal2 s 12898 0 12954 56 6 tap_o[194]
port 195 nsew default tristate
rlabel metal2 s 10782 0 10838 56 6 tap_o[195]
port 196 nsew default tristate
rlabel metal2 s 8666 0 8722 56 6 tap_o[196]
port 197 nsew default tristate
rlabel metal2 s 6550 0 6606 56 6 tap_o[197]
port 198 nsew default tristate
rlabel metal2 s 4434 0 4490 56 6 tap_o[198]
port 199 nsew default tristate
rlabel metal2 s 2318 0 2374 56 6 tap_o[199]
port 200 nsew default tristate
rlabel metal2 s 1030 8648 1086 8704 6 clk_i[0]
port 201 nsew default input
rlabel metal2 s 3146 8648 3202 8704 6 clk_i[1]
port 202 nsew default input
rlabel metal2 s 5262 8648 5318 8704 6 clk_i[2]
port 203 nsew default input
rlabel metal2 s 7378 8648 7434 8704 6 clk_i[3]
port 204 nsew default input
rlabel metal2 s 9494 8648 9550 8704 6 clk_i[4]
port 205 nsew default input
rlabel metal2 s 11610 8648 11666 8704 6 clk_i[5]
port 206 nsew default input
rlabel metal2 s 13726 8648 13782 8704 6 clk_i[6]
port 207 nsew default input
rlabel metal2 s 15842 8648 15898 8704 6 clk_i[7]
port 208 nsew default input
rlabel metal2 s 17958 8648 18014 8704 6 clk_i[8]
port 209 nsew default input
rlabel metal2 s 20074 8648 20130 8704 6 clk_i[9]
port 210 nsew default input
rlabel metal2 s 22190 8648 22246 8704 6 clk_i[10]
port 211 nsew default input
rlabel metal2 s 24306 8648 24362 8704 6 clk_i[11]
port 212 nsew default input
rlabel metal2 s 26422 8648 26478 8704 6 clk_i[12]
port 213 nsew default input
rlabel metal2 s 28538 8648 28594 8704 6 clk_i[13]
port 214 nsew default input
rlabel metal2 s 30654 8648 30710 8704 6 clk_i[14]
port 215 nsew default input
rlabel metal2 s 32770 8648 32826 8704 6 clk_i[15]
port 216 nsew default input
rlabel metal2 s 34886 8648 34942 8704 6 clk_i[16]
port 217 nsew default input
rlabel metal2 s 37002 8648 37058 8704 6 clk_i[17]
port 218 nsew default input
rlabel metal2 s 39118 8648 39174 8704 6 clk_i[18]
port 219 nsew default input
rlabel metal2 s 41234 8648 41290 8704 6 clk_i[19]
port 220 nsew default input
rlabel metal2 s 43350 8648 43406 8704 6 clk_i[20]
port 221 nsew default input
rlabel metal2 s 45466 8648 45522 8704 6 clk_i[21]
port 222 nsew default input
rlabel metal2 s 47582 8648 47638 8704 6 clk_i[22]
port 223 nsew default input
rlabel metal2 s 49698 8648 49754 8704 6 clk_i[23]
port 224 nsew default input
rlabel metal2 s 51814 8648 51870 8704 6 clk_i[24]
port 225 nsew default input
rlabel metal2 s 53930 8648 53986 8704 6 clk_i[25]
port 226 nsew default input
rlabel metal2 s 56046 8648 56102 8704 6 clk_i[26]
port 227 nsew default input
rlabel metal2 s 58162 8648 58218 8704 6 clk_i[27]
port 228 nsew default input
rlabel metal2 s 60278 8648 60334 8704 6 clk_i[28]
port 229 nsew default input
rlabel metal2 s 62394 8648 62450 8704 6 clk_i[29]
port 230 nsew default input
rlabel metal2 s 64510 8648 64566 8704 6 clk_i[30]
port 231 nsew default input
rlabel metal2 s 66626 8648 66682 8704 6 clk_i[31]
port 232 nsew default input
rlabel metal2 s 68742 8648 68798 8704 6 clk_i[32]
port 233 nsew default input
rlabel metal2 s 70858 8648 70914 8704 6 clk_i[33]
port 234 nsew default input
rlabel metal2 s 72974 8648 73030 8704 6 clk_i[34]
port 235 nsew default input
rlabel metal2 s 75090 8648 75146 8704 6 clk_i[35]
port 236 nsew default input
rlabel metal2 s 77206 8648 77262 8704 6 clk_i[36]
port 237 nsew default input
rlabel metal2 s 79322 8648 79378 8704 6 clk_i[37]
port 238 nsew default input
rlabel metal2 s 81438 8648 81494 8704 6 clk_i[38]
port 239 nsew default input
rlabel metal2 s 83554 8648 83610 8704 6 clk_i[39]
port 240 nsew default input
rlabel metal2 s 85670 8648 85726 8704 6 clk_i[40]
port 241 nsew default input
rlabel metal2 s 87786 8648 87842 8704 6 clk_i[41]
port 242 nsew default input
rlabel metal2 s 89902 8648 89958 8704 6 clk_i[42]
port 243 nsew default input
rlabel metal2 s 92018 8648 92074 8704 6 clk_i[43]
port 244 nsew default input
rlabel metal2 s 94134 8648 94190 8704 6 clk_i[44]
port 245 nsew default input
rlabel metal2 s 96250 8648 96306 8704 6 clk_i[45]
port 246 nsew default input
rlabel metal2 s 98366 8648 98422 8704 6 clk_i[46]
port 247 nsew default input
rlabel metal2 s 100482 8648 100538 8704 6 clk_i[47]
port 248 nsew default input
rlabel metal2 s 102598 8648 102654 8704 6 clk_i[48]
port 249 nsew default input
rlabel metal2 s 104714 8648 104770 8704 6 clk_i[49]
port 250 nsew default input
rlabel metal4 s 4004 1040 4324 7664 6 VPWR
port 251 nsew default input
rlabel metal4 s 19364 1040 19684 7664 6 VGND
port 252 nsew default input
<< properties >>
string FIXED_BBOX 0 0 108008 8704
<< end >>
