magic
tech sky130A
magscale 1 2
timestamp 1607274927
<< viali >>
rect 2751 26906 2785 26940
rect 2271 26832 2305 26866
rect 3999 26832 4033 26866
rect 2367 26758 2401 26792
rect 3327 26758 3361 26792
rect 2079 26684 2113 26718
rect 2751 26240 2785 26274
rect 2079 26018 2113 26052
rect 2367 25944 2401 25978
rect 3423 25944 3457 25978
rect 2271 25870 2305 25904
rect 3999 25870 4033 25904
rect 3999 25574 4033 25608
rect 3327 25426 3361 25460
rect 2751 24908 2785 24942
rect 2079 24686 2113 24720
rect 3423 24686 3457 24720
rect 5247 24686 5281 24720
rect 2367 24612 2401 24646
rect 4671 24612 4705 24646
rect 2271 24538 2305 24572
rect 3999 24538 4033 24572
rect 5247 24242 5281 24276
rect 3327 24020 3361 24054
rect 3999 24020 4033 24054
rect 4575 24020 4609 24054
rect 2751 23502 2785 23536
rect 2079 23354 2113 23388
rect 3423 23354 3457 23388
rect 5247 23354 5281 23388
rect 5919 23354 5953 23388
rect 7743 23354 7777 23388
rect 2367 23280 2401 23314
rect 4671 23280 4705 23314
rect 7167 23280 7201 23314
rect 2271 23206 2305 23240
rect 3999 23206 4033 23240
rect 6495 23206 6529 23240
rect 3327 22688 3361 22722
rect 3999 22688 4033 22722
rect 4575 22688 4609 22722
rect 5247 22688 5281 22722
rect 5823 22688 5857 22722
rect 6495 22688 6529 22722
rect 7071 22688 7105 22722
rect 7743 22688 7777 22722
rect 2751 22244 2785 22278
rect 6495 22170 6529 22204
rect 10239 22170 10273 22204
rect 5247 22096 5281 22130
rect 7743 22096 7777 22130
rect 8991 22096 9025 22130
rect 11487 22096 11521 22130
rect 2079 22022 2113 22056
rect 3423 22022 3457 22056
rect 4575 22022 4609 22056
rect 5919 22022 5953 22056
rect 7167 22022 7201 22056
rect 8415 22022 8449 22056
rect 9663 22022 9697 22056
rect 10911 22022 10945 22056
rect 12735 22022 12769 22056
rect 2367 21948 2401 21982
rect 12159 21948 12193 21982
rect 2271 21874 2305 21908
rect 3999 21874 4033 21908
rect 12735 21578 12769 21612
rect 3327 21356 3361 21390
rect 3999 21356 4033 21390
rect 4575 21356 4609 21390
rect 5247 21356 5281 21390
rect 5823 21356 5857 21390
rect 6495 21356 6529 21390
rect 7071 21356 7105 21390
rect 7743 21356 7777 21390
rect 8319 21356 8353 21390
rect 8991 21356 9025 21390
rect 9567 21356 9601 21390
rect 10239 21356 10273 21390
rect 10815 21356 10849 21390
rect 11487 21356 11521 21390
rect 12063 21356 12097 21390
rect 2751 20912 2785 20946
rect 2079 20690 2113 20724
rect 3423 20690 3457 20724
rect 5247 20690 5281 20724
rect 5919 20690 5953 20724
rect 7743 20690 7777 20724
rect 8991 20690 9025 20724
rect 9663 20690 9697 20724
rect 11487 20690 11521 20724
rect 12159 20690 12193 20724
rect 13983 20690 14017 20724
rect 14559 20690 14593 20724
rect 16479 20690 16513 20724
rect 17151 20690 17185 20724
rect 18975 20690 19009 20724
rect 19647 20690 19681 20724
rect 21471 20690 21505 20724
rect 2367 20616 2401 20650
rect 4671 20616 4705 20650
rect 7167 20616 7201 20650
rect 8415 20616 8449 20650
rect 10239 20616 10273 20650
rect 10911 20616 10945 20650
rect 12735 20616 12769 20650
rect 13407 20616 13441 20650
rect 15231 20616 15265 20650
rect 15903 20616 15937 20650
rect 17727 20616 17761 20650
rect 18399 20616 18433 20650
rect 20223 20616 20257 20650
rect 20895 20616 20929 20650
rect 22143 20616 22177 20650
rect 2271 20542 2305 20576
rect 3999 20542 4033 20576
rect 6495 20542 6529 20576
rect 22719 20542 22753 20576
rect 22719 20246 22753 20280
rect 3327 20098 3361 20132
rect 3999 20024 4033 20058
rect 4575 20024 4609 20058
rect 5247 20024 5281 20058
rect 5823 20024 5857 20058
rect 6495 20024 6529 20058
rect 7071 20024 7105 20058
rect 7743 20024 7777 20058
rect 8319 20024 8353 20058
rect 8991 20024 9025 20058
rect 9567 20024 9601 20058
rect 10239 20024 10273 20058
rect 10815 20024 10849 20058
rect 11487 20024 11521 20058
rect 12063 20024 12097 20058
rect 12735 20024 12769 20058
rect 13311 20024 13345 20058
rect 13983 20024 14017 20058
rect 14559 20024 14593 20058
rect 15231 20024 15265 20058
rect 15807 20024 15841 20058
rect 16479 20024 16513 20058
rect 17055 20024 17089 20058
rect 17727 20024 17761 20058
rect 18303 20024 18337 20058
rect 18975 20024 19009 20058
rect 19551 20024 19585 20058
rect 20223 20024 20257 20058
rect 20799 20024 20833 20058
rect 21471 20024 21505 20058
rect 22047 20024 22081 20058
rect 2751 19580 2785 19614
rect 2079 19358 2113 19392
rect 3423 19358 3457 19392
rect 5247 19358 5281 19392
rect 5919 19358 5953 19392
rect 7743 19358 7777 19392
rect 8991 19358 9025 19392
rect 9663 19358 9697 19392
rect 11487 19358 11521 19392
rect 12159 19358 12193 19392
rect 13983 19358 14017 19392
rect 14559 19358 14593 19392
rect 16479 19358 16513 19392
rect 17151 19358 17185 19392
rect 18975 19358 19009 19392
rect 19647 19358 19681 19392
rect 21471 19358 21505 19392
rect 2367 19284 2401 19318
rect 4671 19284 4705 19318
rect 7167 19284 7201 19318
rect 8415 19284 8449 19318
rect 10239 19284 10273 19318
rect 10911 19284 10945 19318
rect 12735 19284 12769 19318
rect 13407 19284 13441 19318
rect 15231 19284 15265 19318
rect 15903 19284 15937 19318
rect 17727 19284 17761 19318
rect 18399 19284 18433 19318
rect 20223 19284 20257 19318
rect 20895 19284 20929 19318
rect 22143 19284 22177 19318
rect 2271 19210 2305 19244
rect 3999 19210 4033 19244
rect 6495 19210 6529 19244
rect 22719 19210 22753 19244
rect 22719 18840 22753 18874
rect 3423 18692 3457 18726
rect 3999 18692 4033 18726
rect 4575 18692 4609 18726
rect 5247 18692 5281 18726
rect 5823 18692 5857 18726
rect 6495 18692 6529 18726
rect 7071 18692 7105 18726
rect 7743 18692 7777 18726
rect 8319 18692 8353 18726
rect 8991 18692 9025 18726
rect 9567 18692 9601 18726
rect 10239 18692 10273 18726
rect 10815 18692 10849 18726
rect 11487 18692 11521 18726
rect 12063 18692 12097 18726
rect 12735 18692 12769 18726
rect 13311 18692 13345 18726
rect 13983 18692 14017 18726
rect 14559 18692 14593 18726
rect 15231 18692 15265 18726
rect 15807 18692 15841 18726
rect 16479 18692 16513 18726
rect 17055 18692 17089 18726
rect 17727 18692 17761 18726
rect 18303 18692 18337 18726
rect 18975 18692 19009 18726
rect 19551 18692 19585 18726
rect 20223 18692 20257 18726
rect 20799 18692 20833 18726
rect 21471 18692 21505 18726
rect 22047 18692 22081 18726
rect 3999 18100 4033 18134
rect 3423 18026 3457 18060
rect 5247 18026 5281 18060
rect 5919 18026 5953 18060
rect 7743 18026 7777 18060
rect 8991 18026 9025 18060
rect 9663 18026 9697 18060
rect 11487 18026 11521 18060
rect 12159 18026 12193 18060
rect 13983 18026 14017 18060
rect 14559 18026 14593 18060
rect 16479 18026 16513 18060
rect 17151 18026 17185 18060
rect 18975 18026 19009 18060
rect 19647 18026 19681 18060
rect 21471 18026 21505 18060
rect 4671 17952 4705 17986
rect 7167 17952 7201 17986
rect 8415 17952 8449 17986
rect 10239 17952 10273 17986
rect 10911 17952 10945 17986
rect 12735 17952 12769 17986
rect 13407 17952 13441 17986
rect 15231 17952 15265 17986
rect 15903 17952 15937 17986
rect 17727 17952 17761 17986
rect 18399 17952 18433 17986
rect 20223 17952 20257 17986
rect 20895 17952 20929 17986
rect 22143 17952 22177 17986
rect 6495 17878 6529 17912
rect 22719 17878 22753 17912
rect 22719 17582 22753 17616
rect 3327 17434 3361 17468
rect 3999 17434 4033 17468
rect 4575 17434 4609 17468
rect 5247 17434 5281 17468
rect 5823 17434 5857 17468
rect 6495 17434 6529 17468
rect 7071 17434 7105 17468
rect 7743 17434 7777 17468
rect 8319 17434 8353 17468
rect 8991 17434 9025 17468
rect 9567 17434 9601 17468
rect 10239 17434 10273 17468
rect 10815 17434 10849 17468
rect 11487 17434 11521 17468
rect 12063 17434 12097 17468
rect 12735 17434 12769 17468
rect 13311 17434 13345 17468
rect 13983 17434 14017 17468
rect 14559 17434 14593 17468
rect 15231 17434 15265 17468
rect 15807 17434 15841 17468
rect 16479 17434 16513 17468
rect 17055 17434 17089 17468
rect 17727 17434 17761 17468
rect 18303 17434 18337 17468
rect 18975 17434 19009 17468
rect 19551 17434 19585 17468
rect 20223 17434 20257 17468
rect 20799 17434 20833 17468
rect 21471 17434 21505 17468
rect 22047 17434 22081 17468
rect 2751 16916 2785 16950
rect 6495 16768 6529 16802
rect 16479 16768 16513 16802
rect 21471 16768 21505 16802
rect 2079 16694 2113 16728
rect 3999 16694 4033 16728
rect 4671 16694 4705 16728
rect 7743 16694 7777 16728
rect 8415 16694 8449 16728
rect 10239 16694 10273 16728
rect 11487 16694 11521 16728
rect 12735 16694 12769 16728
rect 13407 16694 13441 16728
rect 15231 16694 15265 16728
rect 17727 16694 17761 16728
rect 18399 16694 18433 16728
rect 20223 16694 20257 16728
rect 22719 16694 22753 16728
rect 2367 16620 2401 16654
rect 2463 16620 2497 16654
rect 3423 16620 3457 16654
rect 5247 16620 5281 16654
rect 5919 16620 5953 16654
rect 7167 16620 7201 16654
rect 8991 16620 9025 16654
rect 9663 16620 9697 16654
rect 10911 16620 10945 16654
rect 12159 16620 12193 16654
rect 13983 16620 14017 16654
rect 14655 16620 14689 16654
rect 15903 16620 15937 16654
rect 17151 16620 17185 16654
rect 18975 16620 19009 16654
rect 19647 16620 19681 16654
rect 20895 16620 20929 16654
rect 22143 16620 22177 16654
rect 22719 16250 22753 16284
rect 3423 16028 3457 16062
rect 3999 16028 4033 16062
rect 4575 16028 4609 16062
rect 5247 16028 5281 16062
rect 5823 16028 5857 16062
rect 6495 16028 6529 16062
rect 7071 16028 7105 16062
rect 7743 16028 7777 16062
rect 8319 16028 8353 16062
rect 8991 16028 9025 16062
rect 9567 16028 9601 16062
rect 10239 16028 10273 16062
rect 10815 16028 10849 16062
rect 11487 16028 11521 16062
rect 12063 16028 12097 16062
rect 12735 16028 12769 16062
rect 13311 16028 13345 16062
rect 13983 16028 14017 16062
rect 14559 16028 14593 16062
rect 15231 16028 15265 16062
rect 15807 16028 15841 16062
rect 16479 16028 16513 16062
rect 17055 16028 17089 16062
rect 17727 16028 17761 16062
rect 18303 16028 18337 16062
rect 18975 16028 19009 16062
rect 19551 16028 19585 16062
rect 20223 16028 20257 16062
rect 20799 16028 20833 16062
rect 21471 16028 21505 16062
rect 22047 16028 22081 16062
rect 3999 15584 4033 15618
rect 3423 15362 3457 15396
rect 5247 15362 5281 15396
rect 5919 15362 5953 15396
rect 7743 15362 7777 15396
rect 8415 15362 8449 15396
rect 10239 15362 10273 15396
rect 12159 15362 12193 15396
rect 13983 15362 14017 15396
rect 14559 15362 14593 15396
rect 16479 15362 16513 15396
rect 17151 15362 17185 15396
rect 18975 15362 19009 15396
rect 19647 15362 19681 15396
rect 21471 15362 21505 15396
rect 4671 15288 4705 15322
rect 7167 15288 7201 15322
rect 8991 15288 9025 15322
rect 9567 15288 9601 15322
rect 10911 15288 10945 15322
rect 12735 15288 12769 15322
rect 13407 15288 13441 15322
rect 15231 15288 15265 15322
rect 15903 15288 15937 15322
rect 17727 15288 17761 15322
rect 18399 15288 18433 15322
rect 20223 15288 20257 15322
rect 20895 15288 20929 15322
rect 22143 15288 22177 15322
rect 6495 15214 6529 15248
rect 11487 15214 11521 15248
rect 22719 15214 22753 15248
rect 22719 14918 22753 14952
rect 3423 14696 3457 14730
rect 3999 14696 4033 14730
rect 4575 14696 4609 14730
rect 5247 14696 5281 14730
rect 5823 14696 5857 14730
rect 6495 14696 6529 14730
rect 7071 14696 7105 14730
rect 7743 14696 7777 14730
rect 8319 14696 8353 14730
rect 8991 14696 9025 14730
rect 9567 14696 9601 14730
rect 10239 14696 10273 14730
rect 10815 14696 10849 14730
rect 11487 14696 11521 14730
rect 12063 14696 12097 14730
rect 12735 14696 12769 14730
rect 13311 14696 13345 14730
rect 13983 14696 14017 14730
rect 14559 14696 14593 14730
rect 15231 14696 15265 14730
rect 15807 14696 15841 14730
rect 16479 14696 16513 14730
rect 17055 14696 17089 14730
rect 17727 14696 17761 14730
rect 18303 14696 18337 14730
rect 18975 14696 19009 14730
rect 19551 14696 19585 14730
rect 20223 14696 20257 14730
rect 20799 14696 20833 14730
rect 21471 14696 21505 14730
rect 22047 14696 22081 14730
rect 3999 14252 4033 14286
rect 3423 14030 3457 14064
rect 5247 14030 5281 14064
rect 5919 14030 5953 14064
rect 7743 14030 7777 14064
rect 8415 14030 8449 14064
rect 10239 14030 10273 14064
rect 12159 14030 12193 14064
rect 13983 14030 14017 14064
rect 14559 14030 14593 14064
rect 16479 14030 16513 14064
rect 17151 14030 17185 14064
rect 18975 14030 19009 14064
rect 19647 14030 19681 14064
rect 21471 14030 21505 14064
rect 4671 13956 4705 13990
rect 7167 13956 7201 13990
rect 8991 13956 9025 13990
rect 9567 13956 9601 13990
rect 10911 13956 10945 13990
rect 12735 13956 12769 13990
rect 13407 13956 13441 13990
rect 15231 13956 15265 13990
rect 15903 13956 15937 13990
rect 17727 13956 17761 13990
rect 18399 13956 18433 13990
rect 20223 13956 20257 13990
rect 20895 13956 20929 13990
rect 22143 13956 22177 13990
rect 6495 13882 6529 13916
rect 11487 13882 11521 13916
rect 22719 13882 22753 13916
rect 22719 13512 22753 13546
rect 3423 13364 3457 13398
rect 3999 13364 4033 13398
rect 4575 13364 4609 13398
rect 5247 13364 5281 13398
rect 5823 13364 5857 13398
rect 6495 13364 6529 13398
rect 7071 13364 7105 13398
rect 7743 13364 7777 13398
rect 8319 13364 8353 13398
rect 8991 13364 9025 13398
rect 9567 13364 9601 13398
rect 10239 13364 10273 13398
rect 10815 13364 10849 13398
rect 11487 13364 11521 13398
rect 12063 13364 12097 13398
rect 12735 13364 12769 13398
rect 13311 13364 13345 13398
rect 13983 13364 14017 13398
rect 14559 13364 14593 13398
rect 15231 13364 15265 13398
rect 15807 13364 15841 13398
rect 16479 13364 16513 13398
rect 17055 13364 17089 13398
rect 17727 13364 17761 13398
rect 18303 13364 18337 13398
rect 18975 13364 19009 13398
rect 19551 13364 19585 13398
rect 20223 13364 20257 13398
rect 20799 13364 20833 13398
rect 21471 13364 21505 13398
rect 22047 13364 22081 13398
rect 3999 12920 4033 12954
rect 3423 12698 3457 12732
rect 5247 12698 5281 12732
rect 5919 12698 5953 12732
rect 7743 12698 7777 12732
rect 8415 12698 8449 12732
rect 10239 12698 10273 12732
rect 12159 12698 12193 12732
rect 13983 12698 14017 12732
rect 14559 12698 14593 12732
rect 16479 12698 16513 12732
rect 17151 12698 17185 12732
rect 18975 12698 19009 12732
rect 19647 12698 19681 12732
rect 21471 12698 21505 12732
rect 4671 12624 4705 12658
rect 7167 12624 7201 12658
rect 8991 12624 9025 12658
rect 9567 12624 9601 12658
rect 10911 12624 10945 12658
rect 12735 12624 12769 12658
rect 13407 12624 13441 12658
rect 15231 12624 15265 12658
rect 15903 12624 15937 12658
rect 17727 12624 17761 12658
rect 18399 12624 18433 12658
rect 20223 12624 20257 12658
rect 20895 12624 20929 12658
rect 22143 12624 22177 12658
rect 6495 12550 6529 12584
rect 11487 12550 11521 12584
rect 22719 12550 22753 12584
rect 22719 12254 22753 12288
rect 3327 12106 3361 12140
rect 3999 12032 4033 12066
rect 4575 12032 4609 12066
rect 5247 12032 5281 12066
rect 5823 12032 5857 12066
rect 6495 12032 6529 12066
rect 7071 12032 7105 12066
rect 7743 12032 7777 12066
rect 8319 12032 8353 12066
rect 8991 12032 9025 12066
rect 9567 12032 9601 12066
rect 10239 12032 10273 12066
rect 10815 12032 10849 12066
rect 11487 12032 11521 12066
rect 12063 12032 12097 12066
rect 12735 12032 12769 12066
rect 13311 12032 13345 12066
rect 13983 12032 14017 12066
rect 14559 12032 14593 12066
rect 15231 12032 15265 12066
rect 15807 12032 15841 12066
rect 16479 12032 16513 12066
rect 17055 12032 17089 12066
rect 17727 12032 17761 12066
rect 18303 12032 18337 12066
rect 18975 12032 19009 12066
rect 19551 12032 19585 12066
rect 20223 12032 20257 12066
rect 20799 12032 20833 12066
rect 21471 12032 21505 12066
rect 22047 12032 22081 12066
rect 2751 11588 2785 11622
rect 21471 11440 21505 11474
rect 2079 11366 2113 11400
rect 3999 11366 4033 11400
rect 5247 11366 5281 11400
rect 6495 11366 6529 11400
rect 7743 11366 7777 11400
rect 8991 11366 9025 11400
rect 9663 11366 9697 11400
rect 11487 11366 11521 11400
rect 12159 11366 12193 11400
rect 13983 11366 14017 11400
rect 14559 11366 14593 11400
rect 16479 11366 16513 11400
rect 17727 11366 17761 11400
rect 18399 11366 18433 11400
rect 20223 11366 20257 11400
rect 22719 11366 22753 11400
rect 2367 11292 2401 11326
rect 2463 11292 2497 11326
rect 3423 11292 3457 11326
rect 4575 11292 4609 11326
rect 5919 11292 5953 11326
rect 7167 11292 7201 11326
rect 8415 11292 8449 11326
rect 10239 11292 10273 11326
rect 10911 11292 10945 11326
rect 12735 11292 12769 11326
rect 13407 11292 13441 11326
rect 15231 11292 15265 11326
rect 15903 11292 15937 11326
rect 17151 11292 17185 11326
rect 18975 11292 19009 11326
rect 19647 11292 19681 11326
rect 20895 11292 20929 11326
rect 22143 11292 22177 11326
rect 22719 10922 22753 10956
rect 3423 10700 3457 10734
rect 3999 10700 4033 10734
rect 4575 10700 4609 10734
rect 5247 10700 5281 10734
rect 5823 10700 5857 10734
rect 6495 10700 6529 10734
rect 7071 10700 7105 10734
rect 7743 10700 7777 10734
rect 8319 10700 8353 10734
rect 8991 10700 9025 10734
rect 9567 10700 9601 10734
rect 10239 10700 10273 10734
rect 10815 10700 10849 10734
rect 11487 10700 11521 10734
rect 12063 10700 12097 10734
rect 12735 10700 12769 10734
rect 13311 10700 13345 10734
rect 13983 10700 14017 10734
rect 14559 10700 14593 10734
rect 15231 10700 15265 10734
rect 15807 10700 15841 10734
rect 16479 10700 16513 10734
rect 17055 10700 17089 10734
rect 17727 10700 17761 10734
rect 18303 10700 18337 10734
rect 18975 10700 19009 10734
rect 19551 10700 19585 10734
rect 20223 10700 20257 10734
rect 20799 10700 20833 10734
rect 21471 10700 21505 10734
rect 22047 10700 22081 10734
rect 3999 10256 4033 10290
rect 4671 10034 4705 10068
rect 6495 10034 6529 10068
rect 8991 10034 9025 10068
rect 9663 10034 9697 10068
rect 11487 10034 11521 10068
rect 12159 10034 12193 10068
rect 13983 10034 14017 10068
rect 14559 10034 14593 10068
rect 16479 10034 16513 10068
rect 17151 10034 17185 10068
rect 18975 10034 19009 10068
rect 19647 10034 19681 10068
rect 21471 10034 21505 10068
rect 3423 9960 3457 9994
rect 5247 9960 5281 9994
rect 5919 9960 5953 9994
rect 7167 9960 7201 9994
rect 8415 9960 8449 9994
rect 10239 9960 10273 9994
rect 10911 9960 10945 9994
rect 12735 9960 12769 9994
rect 13407 9960 13441 9994
rect 15231 9960 15265 9994
rect 15903 9960 15937 9994
rect 17727 9960 17761 9994
rect 18399 9960 18433 9994
rect 20223 9960 20257 9994
rect 20895 9960 20929 9994
rect 22143 9960 22177 9994
rect 7743 9886 7777 9920
rect 22719 9886 22753 9920
rect 22719 9590 22753 9624
rect 3423 9368 3457 9402
rect 3999 9368 4033 9402
rect 4575 9368 4609 9402
rect 5247 9368 5281 9402
rect 5823 9368 5857 9402
rect 6495 9368 6529 9402
rect 7071 9368 7105 9402
rect 7743 9368 7777 9402
rect 8319 9368 8353 9402
rect 8991 9368 9025 9402
rect 9567 9368 9601 9402
rect 10239 9368 10273 9402
rect 10815 9368 10849 9402
rect 11487 9368 11521 9402
rect 12063 9368 12097 9402
rect 12735 9368 12769 9402
rect 13311 9368 13345 9402
rect 13983 9368 14017 9402
rect 14559 9368 14593 9402
rect 15231 9368 15265 9402
rect 15807 9368 15841 9402
rect 16479 9368 16513 9402
rect 17055 9368 17089 9402
rect 17727 9368 17761 9402
rect 18303 9368 18337 9402
rect 18975 9368 19009 9402
rect 19551 9368 19585 9402
rect 20223 9368 20257 9402
rect 20799 9368 20833 9402
rect 21471 9368 21505 9402
rect 22047 9368 22081 9402
rect 3999 8924 4033 8958
rect 3423 8702 3457 8736
rect 5247 8702 5281 8736
rect 5919 8702 5953 8736
rect 7743 8702 7777 8736
rect 8991 8702 9025 8736
rect 9663 8702 9697 8736
rect 11487 8702 11521 8736
rect 12159 8702 12193 8736
rect 13983 8702 14017 8736
rect 14559 8702 14593 8736
rect 16479 8702 16513 8736
rect 17151 8702 17185 8736
rect 18975 8702 19009 8736
rect 19647 8702 19681 8736
rect 21471 8702 21505 8736
rect 4671 8628 4705 8662
rect 7167 8628 7201 8662
rect 8415 8628 8449 8662
rect 10239 8628 10273 8662
rect 10911 8628 10945 8662
rect 12735 8628 12769 8662
rect 13407 8628 13441 8662
rect 15231 8628 15265 8662
rect 15903 8628 15937 8662
rect 17727 8628 17761 8662
rect 18399 8628 18433 8662
rect 20223 8628 20257 8662
rect 20895 8628 20929 8662
rect 22143 8628 22177 8662
rect 6495 8554 6529 8588
rect 22719 8554 22753 8588
rect 22719 8110 22753 8144
rect 3423 8036 3457 8070
rect 3999 8036 4033 8070
rect 4575 8036 4609 8070
rect 5247 8036 5281 8070
rect 5823 8036 5857 8070
rect 6495 8036 6529 8070
rect 7071 8036 7105 8070
rect 7743 8036 7777 8070
rect 8319 8036 8353 8070
rect 8991 8036 9025 8070
rect 9567 8036 9601 8070
rect 10239 8036 10273 8070
rect 10815 8036 10849 8070
rect 11487 8036 11521 8070
rect 12063 8036 12097 8070
rect 12735 8036 12769 8070
rect 13311 8036 13345 8070
rect 13983 8036 14017 8070
rect 14559 8036 14593 8070
rect 15231 8036 15265 8070
rect 15807 8036 15841 8070
rect 16479 8036 16513 8070
rect 17055 8036 17089 8070
rect 17727 8036 17761 8070
rect 18303 8036 18337 8070
rect 18975 8036 19009 8070
rect 19551 8036 19585 8070
rect 20223 8036 20257 8070
rect 20799 8036 20833 8070
rect 21471 8036 21505 8070
rect 22047 8036 22081 8070
rect 3999 7592 4033 7626
rect 3423 7370 3457 7404
rect 5247 7370 5281 7404
rect 5919 7370 5953 7404
rect 7743 7370 7777 7404
rect 8991 7370 9025 7404
rect 9663 7370 9697 7404
rect 11487 7370 11521 7404
rect 12159 7370 12193 7404
rect 13983 7370 14017 7404
rect 14559 7370 14593 7404
rect 16479 7370 16513 7404
rect 17151 7370 17185 7404
rect 18975 7370 19009 7404
rect 19647 7370 19681 7404
rect 21471 7370 21505 7404
rect 4671 7296 4705 7330
rect 7167 7296 7201 7330
rect 8415 7296 8449 7330
rect 10239 7296 10273 7330
rect 10911 7296 10945 7330
rect 12735 7296 12769 7330
rect 13407 7296 13441 7330
rect 15231 7296 15265 7330
rect 15903 7296 15937 7330
rect 17727 7296 17761 7330
rect 18399 7296 18433 7330
rect 20223 7296 20257 7330
rect 20895 7296 20929 7330
rect 22143 7296 22177 7330
rect 6495 7222 6529 7256
rect 22719 7222 22753 7256
rect 22719 6926 22753 6960
rect 3423 6704 3457 6738
rect 3999 6704 4033 6738
rect 4575 6704 4609 6738
rect 5247 6704 5281 6738
rect 5823 6704 5857 6738
rect 6495 6704 6529 6738
rect 7071 6704 7105 6738
rect 7743 6704 7777 6738
rect 8319 6704 8353 6738
rect 8991 6704 9025 6738
rect 9567 6704 9601 6738
rect 10239 6704 10273 6738
rect 10815 6704 10849 6738
rect 11487 6704 11521 6738
rect 12063 6704 12097 6738
rect 12735 6704 12769 6738
rect 13311 6704 13345 6738
rect 13983 6704 14017 6738
rect 14559 6704 14593 6738
rect 15231 6704 15265 6738
rect 15807 6704 15841 6738
rect 16479 6704 16513 6738
rect 17055 6704 17089 6738
rect 17727 6704 17761 6738
rect 18303 6704 18337 6738
rect 18975 6704 19009 6738
rect 19551 6704 19585 6738
rect 20223 6704 20257 6738
rect 20799 6704 20833 6738
rect 21471 6704 21505 6738
rect 22047 6704 22081 6738
rect 3999 6260 4033 6294
rect 21471 6112 21505 6146
rect 3423 6038 3457 6072
rect 5247 6038 5281 6072
rect 5919 6038 5953 6072
rect 7743 6038 7777 6072
rect 8991 6038 9025 6072
rect 9663 6038 9697 6072
rect 11487 6038 11521 6072
rect 12159 6038 12193 6072
rect 13983 6038 14017 6072
rect 14559 6038 14593 6072
rect 16479 6038 16513 6072
rect 18399 6038 18433 6072
rect 20223 6038 20257 6072
rect 4671 5964 4705 5998
rect 7167 5964 7201 5998
rect 8415 5964 8449 5998
rect 10239 5964 10273 5998
rect 10911 5964 10945 5998
rect 12735 5964 12769 5998
rect 13407 5964 13441 5998
rect 15231 5964 15265 5998
rect 15903 5964 15937 5998
rect 17151 5964 17185 5998
rect 18975 5964 19009 5998
rect 19647 5964 19681 5998
rect 20895 5964 20929 5998
rect 22143 5964 22177 5998
rect 6495 5890 6529 5924
rect 17727 5890 17761 5924
rect 22719 5890 22753 5924
rect 22719 5594 22753 5628
rect 3423 5372 3457 5406
rect 3999 5372 4033 5406
rect 4575 5372 4609 5406
rect 5247 5372 5281 5406
rect 5823 5372 5857 5406
rect 6495 5372 6529 5406
rect 7071 5372 7105 5406
rect 7743 5372 7777 5406
rect 8319 5372 8353 5406
rect 8991 5372 9025 5406
rect 9567 5372 9601 5406
rect 10239 5372 10273 5406
rect 10815 5372 10849 5406
rect 11487 5372 11521 5406
rect 12063 5372 12097 5406
rect 12735 5372 12769 5406
rect 13311 5372 13345 5406
rect 13983 5372 14017 5406
rect 14559 5372 14593 5406
rect 15231 5372 15265 5406
rect 15807 5372 15841 5406
rect 16479 5372 16513 5406
rect 17055 5372 17089 5406
rect 17727 5372 17761 5406
rect 18303 5372 18337 5406
rect 18975 5372 19009 5406
rect 19551 5372 19585 5406
rect 20223 5372 20257 5406
rect 20799 5372 20833 5406
rect 21471 5372 21505 5406
rect 22047 5372 22081 5406
rect 3999 4928 4033 4962
rect 4671 4706 4705 4740
rect 6495 4706 6529 4740
rect 8991 4706 9025 4740
rect 9663 4706 9697 4740
rect 11487 4706 11521 4740
rect 12159 4706 12193 4740
rect 13983 4706 14017 4740
rect 14559 4706 14593 4740
rect 16479 4706 16513 4740
rect 17151 4706 17185 4740
rect 18975 4706 19009 4740
rect 19647 4706 19681 4740
rect 21471 4706 21505 4740
rect 3423 4632 3457 4666
rect 5247 4632 5281 4666
rect 5919 4632 5953 4666
rect 7167 4632 7201 4666
rect 8415 4632 8449 4666
rect 10239 4632 10273 4666
rect 10911 4632 10945 4666
rect 12735 4632 12769 4666
rect 13407 4632 13441 4666
rect 15231 4632 15265 4666
rect 15903 4632 15937 4666
rect 17727 4632 17761 4666
rect 18399 4632 18433 4666
rect 20223 4632 20257 4666
rect 20895 4632 20929 4666
rect 22143 4632 22177 4666
rect 7743 4558 7777 4592
rect 22719 4558 22753 4592
rect 22719 4262 22753 4296
rect 3423 4040 3457 4074
rect 3999 4040 4033 4074
rect 4575 4040 4609 4074
rect 5247 4040 5281 4074
rect 5823 4040 5857 4074
rect 6495 4040 6529 4074
rect 7071 4040 7105 4074
rect 7743 4040 7777 4074
rect 8319 4040 8353 4074
rect 8991 4040 9025 4074
rect 9567 4040 9601 4074
rect 10239 4040 10273 4074
rect 10815 4040 10849 4074
rect 11487 4040 11521 4074
rect 12063 4040 12097 4074
rect 12735 4040 12769 4074
rect 13311 4040 13345 4074
rect 13983 4040 14017 4074
rect 14559 4040 14593 4074
rect 15231 4040 15265 4074
rect 15807 4040 15841 4074
rect 16479 4040 16513 4074
rect 17055 4040 17089 4074
rect 17727 4040 17761 4074
rect 18303 4040 18337 4074
rect 18975 4040 19009 4074
rect 19551 4040 19585 4074
rect 20223 4040 20257 4074
rect 20799 4040 20833 4074
rect 21471 4040 21505 4074
rect 22047 4040 22081 4074
rect 3999 3522 4033 3556
rect 3423 3374 3457 3408
rect 5247 3374 5281 3408
rect 5919 3374 5953 3408
rect 7743 3374 7777 3408
rect 8991 3374 9025 3408
rect 9663 3374 9697 3408
rect 11487 3374 11521 3408
rect 12159 3374 12193 3408
rect 13983 3374 14017 3408
rect 14559 3374 14593 3408
rect 16479 3374 16513 3408
rect 17151 3374 17185 3408
rect 18975 3374 19009 3408
rect 19647 3374 19681 3408
rect 21471 3374 21505 3408
rect 4671 3300 4705 3334
rect 7167 3300 7201 3334
rect 8415 3300 8449 3334
rect 10239 3300 10273 3334
rect 10911 3300 10945 3334
rect 12735 3300 12769 3334
rect 13407 3300 13441 3334
rect 15231 3300 15265 3334
rect 15903 3300 15937 3334
rect 17727 3300 17761 3334
rect 18399 3300 18433 3334
rect 20223 3300 20257 3334
rect 20895 3300 20929 3334
rect 22143 3300 22177 3334
rect 6495 3226 6529 3260
rect 22719 3226 22753 3260
rect 22719 2782 22753 2816
rect 3423 2708 3457 2742
rect 3999 2708 4033 2742
rect 4575 2708 4609 2742
rect 5247 2708 5281 2742
rect 5823 2708 5857 2742
rect 6495 2708 6529 2742
rect 7071 2708 7105 2742
rect 7743 2708 7777 2742
rect 8319 2708 8353 2742
rect 8991 2708 9025 2742
rect 9567 2708 9601 2742
rect 10239 2708 10273 2742
rect 10815 2708 10849 2742
rect 11487 2708 11521 2742
rect 12063 2708 12097 2742
rect 12735 2708 12769 2742
rect 13311 2708 13345 2742
rect 13983 2708 14017 2742
rect 14559 2708 14593 2742
rect 15231 2708 15265 2742
rect 15807 2708 15841 2742
rect 16479 2708 16513 2742
rect 17055 2708 17089 2742
rect 17727 2708 17761 2742
rect 18303 2708 18337 2742
rect 18975 2708 19009 2742
rect 19551 2708 19585 2742
rect 20223 2708 20257 2742
rect 20799 2708 20833 2742
rect 21471 2708 21505 2742
rect 22047 2708 22081 2742
rect 3999 2264 4033 2298
rect 3327 1968 3361 2002
rect 4671 1968 4705 2002
rect 5919 1968 5953 2002
rect 7167 1968 7201 2002
rect 8415 1968 8449 2002
rect 9663 1968 9697 2002
rect 10911 1968 10945 2002
rect 12063 1968 12097 2002
rect 12735 1968 12769 2002
rect 13407 1968 13441 2002
rect 14559 1968 14593 2002
rect 15231 1968 15265 2002
rect 15903 1968 15937 2002
rect 17151 1968 17185 2002
rect 18399 1968 18433 2002
rect 19647 1968 19681 2002
rect 20895 1968 20929 2002
rect 22143 1968 22177 2002
rect 6495 1894 6529 1928
rect 7743 1894 7777 1928
rect 10239 1894 10273 1928
rect 17727 1894 17761 1928
rect 20223 1894 20257 1928
rect 22719 1894 22753 1928
rect 5247 1820 5281 1854
rect 8991 1820 9025 1854
rect 11487 1820 11521 1854
rect 13983 1820 14017 1854
rect 16479 1820 16513 1854
rect 18975 1820 19009 1854
rect 21471 1820 21505 1854
rect 22719 1598 22753 1632
rect 3327 1376 3361 1410
rect 3999 1376 4033 1410
rect 4575 1376 4609 1410
rect 5247 1376 5281 1410
rect 5823 1376 5857 1410
rect 6495 1376 6529 1410
rect 7071 1376 7105 1410
rect 7743 1376 7777 1410
rect 8319 1376 8353 1410
rect 8991 1376 9025 1410
rect 9567 1376 9601 1410
rect 10239 1376 10273 1410
rect 10815 1376 10849 1410
rect 11487 1376 11521 1410
rect 12063 1376 12097 1410
rect 12735 1376 12769 1410
rect 13311 1376 13345 1410
rect 13983 1376 14017 1410
rect 14559 1376 14593 1410
rect 15231 1376 15265 1410
rect 15807 1376 15841 1410
rect 16479 1376 16513 1410
rect 17055 1376 17089 1410
rect 17727 1376 17761 1410
rect 18303 1376 18337 1410
rect 18975 1376 19009 1410
rect 19551 1376 19585 1410
rect 20223 1376 20257 1410
rect 20799 1376 20833 1410
rect 21471 1376 21505 1410
rect 22047 1376 22081 1410
<< metal1 >>
rect 1952 27060 23264 27082
rect 1952 27008 4494 27060
rect 4546 27008 4558 27060
rect 4610 27008 4622 27060
rect 4674 27008 4686 27060
rect 4738 27008 9822 27060
rect 9874 27008 9886 27060
rect 9938 27008 9950 27060
rect 10002 27008 10014 27060
rect 10066 27008 15150 27060
rect 15202 27008 15214 27060
rect 15266 27008 15278 27060
rect 15330 27008 15342 27060
rect 15394 27008 20478 27060
rect 20530 27008 20542 27060
rect 20594 27008 20606 27060
rect 20658 27008 20670 27060
rect 20722 27008 23264 27060
rect 1952 26986 23264 27008
rect 2736 26937 2742 26949
rect 2697 26909 2742 26937
rect 2736 26897 2742 26909
rect 2794 26897 2800 26949
rect 2259 26866 2317 26872
rect 2259 26832 2271 26866
rect 2305 26863 2317 26866
rect 3987 26866 4045 26872
rect 3987 26863 3999 26866
rect 2305 26835 3999 26863
rect 2305 26832 2317 26835
rect 2259 26826 2317 26832
rect 3987 26832 3999 26835
rect 4033 26832 4045 26866
rect 3987 26826 4045 26832
rect 2355 26792 2413 26798
rect 2355 26758 2367 26792
rect 2401 26789 2413 26792
rect 2736 26789 2742 26801
rect 2401 26761 2742 26789
rect 2401 26758 2413 26761
rect 2355 26752 2413 26758
rect 2736 26749 2742 26761
rect 2794 26789 2800 26801
rect 3315 26792 3373 26798
rect 3315 26789 3327 26792
rect 2794 26761 3327 26789
rect 2794 26749 2800 26761
rect 3315 26758 3327 26761
rect 3361 26758 3373 26792
rect 3315 26752 3373 26758
rect 2067 26718 2125 26724
rect 2067 26684 2079 26718
rect 2113 26715 2125 26718
rect 2113 26687 2398 26715
rect 2113 26684 2125 26687
rect 2067 26678 2125 26684
rect 2370 26653 2398 26687
rect 2352 26601 2358 26653
rect 2410 26601 2416 26653
rect 1952 26394 23264 26416
rect 1952 26342 7158 26394
rect 7210 26342 7222 26394
rect 7274 26342 7286 26394
rect 7338 26342 7350 26394
rect 7402 26342 12486 26394
rect 12538 26342 12550 26394
rect 12602 26342 12614 26394
rect 12666 26342 12678 26394
rect 12730 26342 17814 26394
rect 17866 26342 17878 26394
rect 17930 26342 17942 26394
rect 17994 26342 18006 26394
rect 18058 26342 23264 26394
rect 1952 26320 23264 26342
rect 2736 26271 2742 26283
rect 2697 26243 2742 26271
rect 2736 26231 2742 26243
rect 2794 26231 2800 26283
rect 2067 26052 2125 26058
rect 2067 26018 2079 26052
rect 2113 26049 2125 26052
rect 2448 26049 2454 26061
rect 2113 26021 2454 26049
rect 2113 26018 2125 26021
rect 2067 26012 2125 26018
rect 2448 26009 2454 26021
rect 2506 26009 2512 26061
rect 2352 25975 2358 25987
rect 2313 25947 2358 25975
rect 2352 25935 2358 25947
rect 2410 25935 2416 25987
rect 3411 25978 3469 25984
rect 3411 25944 3423 25978
rect 3457 25975 3469 25978
rect 3888 25975 3894 25987
rect 3457 25947 3894 25975
rect 3457 25944 3469 25947
rect 3411 25938 3469 25944
rect 3888 25935 3894 25947
rect 3946 25935 3952 25987
rect 2259 25904 2317 25910
rect 2259 25870 2271 25904
rect 2305 25901 2317 25904
rect 3987 25904 4045 25910
rect 3987 25901 3999 25904
rect 2305 25873 3999 25901
rect 2305 25870 2317 25873
rect 2259 25864 2317 25870
rect 3987 25870 3999 25873
rect 4033 25870 4045 25904
rect 3987 25864 4045 25870
rect 1952 25728 23264 25750
rect 1952 25676 4494 25728
rect 4546 25676 4558 25728
rect 4610 25676 4622 25728
rect 4674 25676 4686 25728
rect 4738 25676 9822 25728
rect 9874 25676 9886 25728
rect 9938 25676 9950 25728
rect 10002 25676 10014 25728
rect 10066 25676 15150 25728
rect 15202 25676 15214 25728
rect 15266 25676 15278 25728
rect 15330 25676 15342 25728
rect 15394 25676 20478 25728
rect 20530 25676 20542 25728
rect 20594 25676 20606 25728
rect 20658 25676 20670 25728
rect 20722 25676 23264 25728
rect 1952 25654 23264 25676
rect 3888 25565 3894 25617
rect 3946 25605 3952 25617
rect 3987 25608 4045 25614
rect 3987 25605 3999 25608
rect 3946 25577 3999 25605
rect 3946 25565 3952 25577
rect 3987 25574 3999 25577
rect 4033 25574 4045 25608
rect 3987 25568 4045 25574
rect 2352 25417 2358 25469
rect 2410 25457 2416 25469
rect 2736 25457 2742 25469
rect 2410 25429 2742 25457
rect 2410 25417 2416 25429
rect 2736 25417 2742 25429
rect 2794 25457 2800 25469
rect 3315 25460 3373 25466
rect 3315 25457 3327 25460
rect 2794 25429 3327 25457
rect 2794 25417 2800 25429
rect 3315 25426 3327 25429
rect 3361 25426 3373 25460
rect 3315 25420 3373 25426
rect 1952 25062 23264 25084
rect 1952 25010 7158 25062
rect 7210 25010 7222 25062
rect 7274 25010 7286 25062
rect 7338 25010 7350 25062
rect 7402 25010 12486 25062
rect 12538 25010 12550 25062
rect 12602 25010 12614 25062
rect 12666 25010 12678 25062
rect 12730 25010 17814 25062
rect 17866 25010 17878 25062
rect 17930 25010 17942 25062
rect 17994 25010 18006 25062
rect 18058 25010 23264 25062
rect 1952 24988 23264 25010
rect 2736 24939 2742 24951
rect 2697 24911 2742 24939
rect 2736 24899 2742 24911
rect 2794 24899 2800 24951
rect 2064 24717 2070 24729
rect 2025 24689 2070 24717
rect 2064 24677 2070 24689
rect 2122 24677 2128 24729
rect 3411 24720 3469 24726
rect 3411 24686 3423 24720
rect 3457 24717 3469 24720
rect 5235 24720 5293 24726
rect 5235 24717 5247 24720
rect 3457 24689 5247 24717
rect 3457 24686 3469 24689
rect 3411 24680 3469 24686
rect 5235 24686 5247 24689
rect 5281 24686 5293 24720
rect 5235 24680 5293 24686
rect 2355 24646 2413 24652
rect 2355 24612 2367 24646
rect 2401 24643 2413 24646
rect 2736 24643 2742 24655
rect 2401 24615 2742 24643
rect 2401 24612 2413 24615
rect 2355 24606 2413 24612
rect 2736 24603 2742 24615
rect 2794 24603 2800 24655
rect 4659 24646 4717 24652
rect 4659 24612 4671 24646
rect 4705 24643 4717 24646
rect 5136 24643 5142 24655
rect 4705 24615 5142 24643
rect 4705 24612 4717 24615
rect 4659 24606 4717 24612
rect 5136 24603 5142 24615
rect 5194 24603 5200 24655
rect 2259 24572 2317 24578
rect 2259 24538 2271 24572
rect 2305 24569 2317 24572
rect 3987 24572 4045 24578
rect 3987 24569 3999 24572
rect 2305 24541 3999 24569
rect 2305 24538 2317 24541
rect 2259 24532 2317 24538
rect 3987 24538 3999 24541
rect 4033 24538 4045 24572
rect 3987 24532 4045 24538
rect 1952 24396 23264 24418
rect 1952 24344 4494 24396
rect 4546 24344 4558 24396
rect 4610 24344 4622 24396
rect 4674 24344 4686 24396
rect 4738 24344 9822 24396
rect 9874 24344 9886 24396
rect 9938 24344 9950 24396
rect 10002 24344 10014 24396
rect 10066 24344 15150 24396
rect 15202 24344 15214 24396
rect 15266 24344 15278 24396
rect 15330 24344 15342 24396
rect 15394 24344 20478 24396
rect 20530 24344 20542 24396
rect 20594 24344 20606 24396
rect 20658 24344 20670 24396
rect 20722 24344 23264 24396
rect 1952 24322 23264 24344
rect 5136 24233 5142 24285
rect 5194 24273 5200 24285
rect 5235 24276 5293 24282
rect 5235 24273 5247 24276
rect 5194 24245 5247 24273
rect 5194 24233 5200 24245
rect 5235 24242 5247 24245
rect 5281 24242 5293 24276
rect 5235 24236 5293 24242
rect 2736 24011 2742 24063
rect 2794 24051 2800 24063
rect 3315 24054 3373 24060
rect 3315 24051 3327 24054
rect 2794 24023 3327 24051
rect 2794 24011 2800 24023
rect 3315 24020 3327 24023
rect 3361 24020 3373 24054
rect 3315 24014 3373 24020
rect 3987 24054 4045 24060
rect 3987 24020 3999 24054
rect 4033 24051 4045 24054
rect 4563 24054 4621 24060
rect 4563 24051 4575 24054
rect 4033 24023 4575 24051
rect 4033 24020 4045 24023
rect 3987 24014 4045 24020
rect 4563 24020 4575 24023
rect 4609 24020 4621 24054
rect 4563 24014 4621 24020
rect 1952 23730 23264 23752
rect 1952 23678 7158 23730
rect 7210 23678 7222 23730
rect 7274 23678 7286 23730
rect 7338 23678 7350 23730
rect 7402 23678 12486 23730
rect 12538 23678 12550 23730
rect 12602 23678 12614 23730
rect 12666 23678 12678 23730
rect 12730 23678 17814 23730
rect 17866 23678 17878 23730
rect 17930 23678 17942 23730
rect 17994 23678 18006 23730
rect 18058 23678 23264 23730
rect 1952 23656 23264 23678
rect 2736 23533 2742 23545
rect 2697 23505 2742 23533
rect 2736 23493 2742 23505
rect 2794 23493 2800 23545
rect 2064 23385 2070 23397
rect 2025 23357 2070 23385
rect 2064 23345 2070 23357
rect 2122 23345 2128 23397
rect 3411 23388 3469 23394
rect 3411 23354 3423 23388
rect 3457 23385 3469 23388
rect 5235 23388 5293 23394
rect 5235 23385 5247 23388
rect 3457 23357 5247 23385
rect 3457 23354 3469 23357
rect 3411 23348 3469 23354
rect 5235 23354 5247 23357
rect 5281 23354 5293 23388
rect 5235 23348 5293 23354
rect 5907 23388 5965 23394
rect 5907 23354 5919 23388
rect 5953 23385 5965 23388
rect 7731 23388 7789 23394
rect 7731 23385 7743 23388
rect 5953 23357 7743 23385
rect 5953 23354 5965 23357
rect 5907 23348 5965 23354
rect 7731 23354 7743 23357
rect 7777 23354 7789 23388
rect 7731 23348 7789 23354
rect 2355 23314 2413 23320
rect 2355 23280 2367 23314
rect 2401 23311 2413 23314
rect 2736 23311 2742 23323
rect 2401 23283 2742 23311
rect 2401 23280 2413 23283
rect 2355 23274 2413 23280
rect 2736 23271 2742 23283
rect 2794 23271 2800 23323
rect 4659 23314 4717 23320
rect 4659 23280 4671 23314
rect 4705 23280 4717 23314
rect 4659 23274 4717 23280
rect 7155 23314 7213 23320
rect 7155 23280 7167 23314
rect 7201 23311 7213 23314
rect 7201 23283 7774 23311
rect 7201 23280 7213 23283
rect 7155 23274 7213 23280
rect 2259 23240 2317 23246
rect 2259 23206 2271 23240
rect 2305 23237 2317 23240
rect 3987 23240 4045 23246
rect 3987 23237 3999 23240
rect 2305 23209 3999 23237
rect 2305 23206 2317 23209
rect 2259 23200 2317 23206
rect 3987 23206 3999 23209
rect 4033 23206 4045 23240
rect 4674 23237 4702 23274
rect 7746 23249 7774 23283
rect 6483 23240 6541 23246
rect 6483 23237 6495 23240
rect 4674 23209 6495 23237
rect 3987 23200 4045 23206
rect 6483 23206 6495 23209
rect 6529 23206 6541 23240
rect 6483 23200 6541 23206
rect 7728 23197 7734 23249
rect 7786 23197 7792 23249
rect 1952 23064 23264 23086
rect 1952 23012 4494 23064
rect 4546 23012 4558 23064
rect 4610 23012 4622 23064
rect 4674 23012 4686 23064
rect 4738 23012 9822 23064
rect 9874 23012 9886 23064
rect 9938 23012 9950 23064
rect 10002 23012 10014 23064
rect 10066 23012 15150 23064
rect 15202 23012 15214 23064
rect 15266 23012 15278 23064
rect 15330 23012 15342 23064
rect 15394 23012 20478 23064
rect 20530 23012 20542 23064
rect 20594 23012 20606 23064
rect 20658 23012 20670 23064
rect 20722 23012 23264 23064
rect 1952 22990 23264 23012
rect 2736 22679 2742 22731
rect 2794 22719 2800 22731
rect 3315 22722 3373 22728
rect 3315 22719 3327 22722
rect 2794 22691 3327 22719
rect 2794 22679 2800 22691
rect 3315 22688 3327 22691
rect 3361 22688 3373 22722
rect 3315 22682 3373 22688
rect 3987 22722 4045 22728
rect 3987 22688 3999 22722
rect 4033 22719 4045 22722
rect 4563 22722 4621 22728
rect 4563 22719 4575 22722
rect 4033 22691 4575 22719
rect 4033 22688 4045 22691
rect 3987 22682 4045 22688
rect 4563 22688 4575 22691
rect 4609 22688 4621 22722
rect 4563 22682 4621 22688
rect 5235 22722 5293 22728
rect 5235 22688 5247 22722
rect 5281 22719 5293 22722
rect 5811 22722 5869 22728
rect 5811 22719 5823 22722
rect 5281 22691 5823 22719
rect 5281 22688 5293 22691
rect 5235 22682 5293 22688
rect 5811 22688 5823 22691
rect 5857 22688 5869 22722
rect 5811 22682 5869 22688
rect 6483 22722 6541 22728
rect 6483 22688 6495 22722
rect 6529 22719 6541 22722
rect 7059 22722 7117 22728
rect 7059 22719 7071 22722
rect 6529 22691 7071 22719
rect 6529 22688 6541 22691
rect 6483 22682 6541 22688
rect 7059 22688 7071 22691
rect 7105 22688 7117 22722
rect 7059 22682 7117 22688
rect 7728 22679 7734 22731
rect 7786 22719 7792 22731
rect 7786 22691 7831 22719
rect 7786 22679 7792 22691
rect 1952 22398 23264 22420
rect 1952 22346 7158 22398
rect 7210 22346 7222 22398
rect 7274 22346 7286 22398
rect 7338 22346 7350 22398
rect 7402 22346 12486 22398
rect 12538 22346 12550 22398
rect 12602 22346 12614 22398
rect 12666 22346 12678 22398
rect 12730 22346 17814 22398
rect 17866 22346 17878 22398
rect 17930 22346 17942 22398
rect 17994 22346 18006 22398
rect 18058 22346 23264 22398
rect 1952 22324 23264 22346
rect 2736 22275 2742 22287
rect 2697 22247 2742 22275
rect 2736 22235 2742 22247
rect 2794 22235 2800 22287
rect 6483 22204 6541 22210
rect 6483 22201 6495 22204
rect 5538 22173 6495 22201
rect 5235 22130 5293 22136
rect 5235 22127 5247 22130
rect 3426 22099 5247 22127
rect 2064 22053 2070 22065
rect 2025 22025 2070 22053
rect 2064 22013 2070 22025
rect 2122 22013 2128 22065
rect 3426 22062 3454 22099
rect 5235 22096 5247 22099
rect 5281 22096 5293 22130
rect 5235 22090 5293 22096
rect 3411 22056 3469 22062
rect 3411 22022 3423 22056
rect 3457 22022 3469 22056
rect 3411 22016 3469 22022
rect 4563 22056 4621 22062
rect 4563 22022 4575 22056
rect 4609 22053 4621 22056
rect 5538 22053 5566 22173
rect 6483 22170 6495 22173
rect 6529 22170 6541 22204
rect 10227 22204 10285 22210
rect 10227 22201 10239 22204
rect 6483 22164 6541 22170
rect 9282 22173 10239 22201
rect 7731 22130 7789 22136
rect 7731 22127 7743 22130
rect 5922 22099 7743 22127
rect 5922 22062 5950 22099
rect 7731 22096 7743 22099
rect 7777 22096 7789 22130
rect 8979 22130 9037 22136
rect 8979 22127 8991 22130
rect 7731 22090 7789 22096
rect 8322 22099 8991 22127
rect 4609 22025 5566 22053
rect 5907 22056 5965 22062
rect 4609 22022 4621 22025
rect 4563 22016 4621 22022
rect 5907 22022 5919 22056
rect 5953 22022 5965 22056
rect 5907 22016 5965 22022
rect 7155 22056 7213 22062
rect 7155 22022 7167 22056
rect 7201 22053 7213 22056
rect 8322 22053 8350 22099
rect 8979 22096 8991 22099
rect 9025 22096 9037 22130
rect 8979 22090 9037 22096
rect 7201 22025 8350 22053
rect 8403 22056 8461 22062
rect 7201 22022 7213 22025
rect 7155 22016 7213 22022
rect 8403 22022 8415 22056
rect 8449 22053 8461 22056
rect 9282 22053 9310 22173
rect 10227 22170 10239 22173
rect 10273 22170 10285 22204
rect 10227 22164 10285 22170
rect 11475 22130 11533 22136
rect 11475 22127 11487 22130
rect 9666 22099 11487 22127
rect 9666 22062 9694 22099
rect 11475 22096 11487 22099
rect 11521 22096 11533 22130
rect 11475 22090 11533 22096
rect 8449 22025 9310 22053
rect 9651 22056 9709 22062
rect 8449 22022 8461 22025
rect 8403 22016 8461 22022
rect 9651 22022 9663 22056
rect 9697 22022 9709 22056
rect 9651 22016 9709 22022
rect 10899 22056 10957 22062
rect 10899 22022 10911 22056
rect 10945 22053 10957 22056
rect 12723 22056 12781 22062
rect 12723 22053 12735 22056
rect 10945 22025 12735 22053
rect 10945 22022 10957 22025
rect 10899 22016 10957 22022
rect 12723 22022 12735 22025
rect 12769 22022 12781 22056
rect 12723 22016 12781 22022
rect 2355 21982 2413 21988
rect 2355 21948 2367 21982
rect 2401 21979 2413 21982
rect 2736 21979 2742 21991
rect 2401 21951 2742 21979
rect 2401 21948 2413 21951
rect 2355 21942 2413 21948
rect 2736 21939 2742 21951
rect 2794 21939 2800 21991
rect 12147 21982 12205 21988
rect 12147 21948 12159 21982
rect 12193 21979 12205 21982
rect 12624 21979 12630 21991
rect 12193 21951 12630 21979
rect 12193 21948 12205 21951
rect 12147 21942 12205 21948
rect 12624 21939 12630 21951
rect 12682 21939 12688 21991
rect 2259 21908 2317 21914
rect 2259 21874 2271 21908
rect 2305 21905 2317 21908
rect 3987 21908 4045 21914
rect 3987 21905 3999 21908
rect 2305 21877 3999 21905
rect 2305 21874 2317 21877
rect 2259 21868 2317 21874
rect 3987 21874 3999 21877
rect 4033 21874 4045 21908
rect 3987 21868 4045 21874
rect 1952 21732 23264 21754
rect 1952 21680 4494 21732
rect 4546 21680 4558 21732
rect 4610 21680 4622 21732
rect 4674 21680 4686 21732
rect 4738 21680 9822 21732
rect 9874 21680 9886 21732
rect 9938 21680 9950 21732
rect 10002 21680 10014 21732
rect 10066 21680 15150 21732
rect 15202 21680 15214 21732
rect 15266 21680 15278 21732
rect 15330 21680 15342 21732
rect 15394 21680 20478 21732
rect 20530 21680 20542 21732
rect 20594 21680 20606 21732
rect 20658 21680 20670 21732
rect 20722 21680 23264 21732
rect 1952 21658 23264 21680
rect 12624 21569 12630 21621
rect 12682 21609 12688 21621
rect 12723 21612 12781 21618
rect 12723 21609 12735 21612
rect 12682 21581 12735 21609
rect 12682 21569 12688 21581
rect 12723 21578 12735 21581
rect 12769 21578 12781 21612
rect 12723 21572 12781 21578
rect 2736 21347 2742 21399
rect 2794 21387 2800 21399
rect 3315 21390 3373 21396
rect 3315 21387 3327 21390
rect 2794 21359 3327 21387
rect 2794 21347 2800 21359
rect 3315 21356 3327 21359
rect 3361 21356 3373 21390
rect 3315 21350 3373 21356
rect 3987 21390 4045 21396
rect 3987 21356 3999 21390
rect 4033 21387 4045 21390
rect 4563 21390 4621 21396
rect 4563 21387 4575 21390
rect 4033 21359 4575 21387
rect 4033 21356 4045 21359
rect 3987 21350 4045 21356
rect 4563 21356 4575 21359
rect 4609 21356 4621 21390
rect 4563 21350 4621 21356
rect 5235 21390 5293 21396
rect 5235 21356 5247 21390
rect 5281 21387 5293 21390
rect 5811 21390 5869 21396
rect 5811 21387 5823 21390
rect 5281 21359 5823 21387
rect 5281 21356 5293 21359
rect 5235 21350 5293 21356
rect 5811 21356 5823 21359
rect 5857 21356 5869 21390
rect 5811 21350 5869 21356
rect 6483 21390 6541 21396
rect 6483 21356 6495 21390
rect 6529 21387 6541 21390
rect 7059 21390 7117 21396
rect 7059 21387 7071 21390
rect 6529 21359 7071 21387
rect 6529 21356 6541 21359
rect 6483 21350 6541 21356
rect 7059 21356 7071 21359
rect 7105 21356 7117 21390
rect 7059 21350 7117 21356
rect 7731 21390 7789 21396
rect 7731 21356 7743 21390
rect 7777 21387 7789 21390
rect 8307 21390 8365 21396
rect 8307 21387 8319 21390
rect 7777 21359 8319 21387
rect 7777 21356 7789 21359
rect 7731 21350 7789 21356
rect 8307 21356 8319 21359
rect 8353 21356 8365 21390
rect 8307 21350 8365 21356
rect 8979 21390 9037 21396
rect 8979 21356 8991 21390
rect 9025 21387 9037 21390
rect 9555 21390 9613 21396
rect 9555 21387 9567 21390
rect 9025 21359 9567 21387
rect 9025 21356 9037 21359
rect 8979 21350 9037 21356
rect 9555 21356 9567 21359
rect 9601 21356 9613 21390
rect 9555 21350 9613 21356
rect 10227 21390 10285 21396
rect 10227 21356 10239 21390
rect 10273 21387 10285 21390
rect 10803 21390 10861 21396
rect 10803 21387 10815 21390
rect 10273 21359 10815 21387
rect 10273 21356 10285 21359
rect 10227 21350 10285 21356
rect 10803 21356 10815 21359
rect 10849 21356 10861 21390
rect 10803 21350 10861 21356
rect 11475 21390 11533 21396
rect 11475 21356 11487 21390
rect 11521 21387 11533 21390
rect 12051 21390 12109 21396
rect 12051 21387 12063 21390
rect 11521 21359 12063 21387
rect 11521 21356 11533 21359
rect 11475 21350 11533 21356
rect 12051 21356 12063 21359
rect 12097 21356 12109 21390
rect 12051 21350 12109 21356
rect 1952 21066 23264 21088
rect 1952 21014 7158 21066
rect 7210 21014 7222 21066
rect 7274 21014 7286 21066
rect 7338 21014 7350 21066
rect 7402 21014 12486 21066
rect 12538 21014 12550 21066
rect 12602 21014 12614 21066
rect 12666 21014 12678 21066
rect 12730 21014 17814 21066
rect 17866 21014 17878 21066
rect 17930 21014 17942 21066
rect 17994 21014 18006 21066
rect 18058 21014 23264 21066
rect 1952 20992 23264 21014
rect 2736 20943 2742 20955
rect 2697 20915 2742 20943
rect 2736 20903 2742 20915
rect 2794 20903 2800 20955
rect 2067 20724 2125 20730
rect 2067 20690 2079 20724
rect 2113 20721 2125 20724
rect 2448 20721 2454 20733
rect 2113 20693 2454 20721
rect 2113 20690 2125 20693
rect 2067 20684 2125 20690
rect 2448 20681 2454 20693
rect 2506 20681 2512 20733
rect 3411 20724 3469 20730
rect 3411 20690 3423 20724
rect 3457 20721 3469 20724
rect 5235 20724 5293 20730
rect 5235 20721 5247 20724
rect 3457 20693 5247 20721
rect 3457 20690 3469 20693
rect 3411 20684 3469 20690
rect 5235 20690 5247 20693
rect 5281 20690 5293 20724
rect 5235 20684 5293 20690
rect 5907 20724 5965 20730
rect 5907 20690 5919 20724
rect 5953 20721 5965 20724
rect 7731 20724 7789 20730
rect 7731 20721 7743 20724
rect 5953 20693 7743 20721
rect 5953 20690 5965 20693
rect 5907 20684 5965 20690
rect 7731 20690 7743 20693
rect 7777 20690 7789 20724
rect 8979 20724 9037 20730
rect 8979 20721 8991 20724
rect 7731 20684 7789 20690
rect 8322 20693 8991 20721
rect 2352 20647 2358 20659
rect 2313 20619 2358 20647
rect 2352 20607 2358 20619
rect 2410 20607 2416 20659
rect 4659 20650 4717 20656
rect 4659 20616 4671 20650
rect 4705 20616 4717 20650
rect 4659 20610 4717 20616
rect 7155 20650 7213 20656
rect 7155 20616 7167 20650
rect 7201 20647 7213 20650
rect 8322 20647 8350 20693
rect 8979 20690 8991 20693
rect 9025 20690 9037 20724
rect 8979 20684 9037 20690
rect 9651 20724 9709 20730
rect 9651 20690 9663 20724
rect 9697 20721 9709 20724
rect 11475 20724 11533 20730
rect 11475 20721 11487 20724
rect 9697 20693 11487 20721
rect 9697 20690 9709 20693
rect 9651 20684 9709 20690
rect 11475 20690 11487 20693
rect 11521 20690 11533 20724
rect 11475 20684 11533 20690
rect 12147 20724 12205 20730
rect 12147 20690 12159 20724
rect 12193 20721 12205 20724
rect 13971 20724 14029 20730
rect 13971 20721 13983 20724
rect 12193 20693 13983 20721
rect 12193 20690 12205 20693
rect 12147 20684 12205 20690
rect 13971 20690 13983 20693
rect 14017 20690 14029 20724
rect 13971 20684 14029 20690
rect 14547 20724 14605 20730
rect 14547 20690 14559 20724
rect 14593 20721 14605 20724
rect 16467 20724 16525 20730
rect 16467 20721 16479 20724
rect 14593 20693 16479 20721
rect 14593 20690 14605 20693
rect 14547 20684 14605 20690
rect 16467 20690 16479 20693
rect 16513 20690 16525 20724
rect 16467 20684 16525 20690
rect 17139 20724 17197 20730
rect 17139 20690 17151 20724
rect 17185 20721 17197 20724
rect 18963 20724 19021 20730
rect 18963 20721 18975 20724
rect 17185 20693 18975 20721
rect 17185 20690 17197 20693
rect 17139 20684 17197 20690
rect 18963 20690 18975 20693
rect 19009 20690 19021 20724
rect 18963 20684 19021 20690
rect 19635 20724 19693 20730
rect 19635 20690 19647 20724
rect 19681 20721 19693 20724
rect 21459 20724 21517 20730
rect 21459 20721 21471 20724
rect 19681 20693 21471 20721
rect 19681 20690 19693 20693
rect 19635 20684 19693 20690
rect 21459 20690 21471 20693
rect 21505 20690 21517 20724
rect 21459 20684 21517 20690
rect 7201 20619 8350 20647
rect 8403 20650 8461 20656
rect 7201 20616 7213 20619
rect 7155 20610 7213 20616
rect 8403 20616 8415 20650
rect 8449 20647 8461 20650
rect 10227 20650 10285 20656
rect 10227 20647 10239 20650
rect 8449 20619 10239 20647
rect 8449 20616 8461 20619
rect 8403 20610 8461 20616
rect 10227 20616 10239 20619
rect 10273 20616 10285 20650
rect 10227 20610 10285 20616
rect 10899 20650 10957 20656
rect 10899 20616 10911 20650
rect 10945 20647 10957 20650
rect 12723 20650 12781 20656
rect 12723 20647 12735 20650
rect 10945 20619 12735 20647
rect 10945 20616 10957 20619
rect 10899 20610 10957 20616
rect 12723 20616 12735 20619
rect 12769 20616 12781 20650
rect 12723 20610 12781 20616
rect 13395 20650 13453 20656
rect 13395 20616 13407 20650
rect 13441 20647 13453 20650
rect 15219 20650 15277 20656
rect 15219 20647 15231 20650
rect 13441 20619 15231 20647
rect 13441 20616 13453 20619
rect 13395 20610 13453 20616
rect 15219 20616 15231 20619
rect 15265 20616 15277 20650
rect 15219 20610 15277 20616
rect 15891 20650 15949 20656
rect 15891 20616 15903 20650
rect 15937 20647 15949 20650
rect 17715 20650 17773 20656
rect 17715 20647 17727 20650
rect 15937 20619 17727 20647
rect 15937 20616 15949 20619
rect 15891 20610 15949 20616
rect 17715 20616 17727 20619
rect 17761 20616 17773 20650
rect 17715 20610 17773 20616
rect 18387 20650 18445 20656
rect 18387 20616 18399 20650
rect 18433 20647 18445 20650
rect 20211 20650 20269 20656
rect 20211 20647 20223 20650
rect 18433 20619 20223 20647
rect 18433 20616 18445 20619
rect 18387 20610 18445 20616
rect 20211 20616 20223 20619
rect 20257 20616 20269 20650
rect 20211 20610 20269 20616
rect 20883 20650 20941 20656
rect 20883 20616 20895 20650
rect 20929 20616 20941 20650
rect 20883 20610 20941 20616
rect 22131 20650 22189 20656
rect 22131 20616 22143 20650
rect 22177 20647 22189 20650
rect 22608 20647 22614 20659
rect 22177 20619 22614 20647
rect 22177 20616 22189 20619
rect 22131 20610 22189 20616
rect 2259 20576 2317 20582
rect 2259 20542 2271 20576
rect 2305 20573 2317 20576
rect 3987 20576 4045 20582
rect 3987 20573 3999 20576
rect 2305 20545 3999 20573
rect 2305 20542 2317 20545
rect 2259 20536 2317 20542
rect 3987 20542 3999 20545
rect 4033 20542 4045 20576
rect 4674 20573 4702 20610
rect 6483 20576 6541 20582
rect 6483 20573 6495 20576
rect 4674 20545 6495 20573
rect 3987 20536 4045 20542
rect 6483 20542 6495 20545
rect 6529 20542 6541 20576
rect 20898 20573 20926 20610
rect 22608 20607 22614 20619
rect 22666 20607 22672 20659
rect 22707 20576 22765 20582
rect 22707 20573 22719 20576
rect 20898 20545 22719 20573
rect 6483 20536 6541 20542
rect 22707 20542 22719 20545
rect 22753 20542 22765 20576
rect 22707 20536 22765 20542
rect 1952 20400 23264 20422
rect 1952 20348 4494 20400
rect 4546 20348 4558 20400
rect 4610 20348 4622 20400
rect 4674 20348 4686 20400
rect 4738 20348 9822 20400
rect 9874 20348 9886 20400
rect 9938 20348 9950 20400
rect 10002 20348 10014 20400
rect 10066 20348 15150 20400
rect 15202 20348 15214 20400
rect 15266 20348 15278 20400
rect 15330 20348 15342 20400
rect 15394 20348 20478 20400
rect 20530 20348 20542 20400
rect 20594 20348 20606 20400
rect 20658 20348 20670 20400
rect 20722 20348 23264 20400
rect 1952 20326 23264 20348
rect 22608 20237 22614 20289
rect 22666 20277 22672 20289
rect 22707 20280 22765 20286
rect 22707 20277 22719 20280
rect 22666 20249 22719 20277
rect 22666 20237 22672 20249
rect 22707 20246 22719 20249
rect 22753 20246 22765 20280
rect 22707 20240 22765 20246
rect 2352 20089 2358 20141
rect 2410 20129 2416 20141
rect 2736 20129 2742 20141
rect 2410 20101 2742 20129
rect 2410 20089 2416 20101
rect 2736 20089 2742 20101
rect 2794 20129 2800 20141
rect 3315 20132 3373 20138
rect 3315 20129 3327 20132
rect 2794 20101 3327 20129
rect 2794 20089 2800 20101
rect 3315 20098 3327 20101
rect 3361 20098 3373 20132
rect 3315 20092 3373 20098
rect 3987 20058 4045 20064
rect 3987 20024 3999 20058
rect 4033 20055 4045 20058
rect 4563 20058 4621 20064
rect 4563 20055 4575 20058
rect 4033 20027 4575 20055
rect 4033 20024 4045 20027
rect 3987 20018 4045 20024
rect 4563 20024 4575 20027
rect 4609 20024 4621 20058
rect 4563 20018 4621 20024
rect 5235 20058 5293 20064
rect 5235 20024 5247 20058
rect 5281 20055 5293 20058
rect 5811 20058 5869 20064
rect 5811 20055 5823 20058
rect 5281 20027 5823 20055
rect 5281 20024 5293 20027
rect 5235 20018 5293 20024
rect 5811 20024 5823 20027
rect 5857 20024 5869 20058
rect 5811 20018 5869 20024
rect 6483 20058 6541 20064
rect 6483 20024 6495 20058
rect 6529 20055 6541 20058
rect 7059 20058 7117 20064
rect 7059 20055 7071 20058
rect 6529 20027 7071 20055
rect 6529 20024 6541 20027
rect 6483 20018 6541 20024
rect 7059 20024 7071 20027
rect 7105 20024 7117 20058
rect 7059 20018 7117 20024
rect 7731 20058 7789 20064
rect 7731 20024 7743 20058
rect 7777 20055 7789 20058
rect 8307 20058 8365 20064
rect 8307 20055 8319 20058
rect 7777 20027 8319 20055
rect 7777 20024 7789 20027
rect 7731 20018 7789 20024
rect 8307 20024 8319 20027
rect 8353 20024 8365 20058
rect 8307 20018 8365 20024
rect 8979 20058 9037 20064
rect 8979 20024 8991 20058
rect 9025 20055 9037 20058
rect 9555 20058 9613 20064
rect 9555 20055 9567 20058
rect 9025 20027 9567 20055
rect 9025 20024 9037 20027
rect 8979 20018 9037 20024
rect 9555 20024 9567 20027
rect 9601 20024 9613 20058
rect 9555 20018 9613 20024
rect 10227 20058 10285 20064
rect 10227 20024 10239 20058
rect 10273 20055 10285 20058
rect 10803 20058 10861 20064
rect 10803 20055 10815 20058
rect 10273 20027 10815 20055
rect 10273 20024 10285 20027
rect 10227 20018 10285 20024
rect 10803 20024 10815 20027
rect 10849 20024 10861 20058
rect 10803 20018 10861 20024
rect 11475 20058 11533 20064
rect 11475 20024 11487 20058
rect 11521 20055 11533 20058
rect 12051 20058 12109 20064
rect 12051 20055 12063 20058
rect 11521 20027 12063 20055
rect 11521 20024 11533 20027
rect 11475 20018 11533 20024
rect 12051 20024 12063 20027
rect 12097 20024 12109 20058
rect 12051 20018 12109 20024
rect 12723 20058 12781 20064
rect 12723 20024 12735 20058
rect 12769 20055 12781 20058
rect 13299 20058 13357 20064
rect 13299 20055 13311 20058
rect 12769 20027 13311 20055
rect 12769 20024 12781 20027
rect 12723 20018 12781 20024
rect 13299 20024 13311 20027
rect 13345 20024 13357 20058
rect 13299 20018 13357 20024
rect 13971 20058 14029 20064
rect 13971 20024 13983 20058
rect 14017 20055 14029 20058
rect 14547 20058 14605 20064
rect 14547 20055 14559 20058
rect 14017 20027 14559 20055
rect 14017 20024 14029 20027
rect 13971 20018 14029 20024
rect 14547 20024 14559 20027
rect 14593 20024 14605 20058
rect 14547 20018 14605 20024
rect 15219 20058 15277 20064
rect 15219 20024 15231 20058
rect 15265 20055 15277 20058
rect 15795 20058 15853 20064
rect 15795 20055 15807 20058
rect 15265 20027 15807 20055
rect 15265 20024 15277 20027
rect 15219 20018 15277 20024
rect 15795 20024 15807 20027
rect 15841 20024 15853 20058
rect 15795 20018 15853 20024
rect 16467 20058 16525 20064
rect 16467 20024 16479 20058
rect 16513 20055 16525 20058
rect 17043 20058 17101 20064
rect 17043 20055 17055 20058
rect 16513 20027 17055 20055
rect 16513 20024 16525 20027
rect 16467 20018 16525 20024
rect 17043 20024 17055 20027
rect 17089 20024 17101 20058
rect 17043 20018 17101 20024
rect 17715 20058 17773 20064
rect 17715 20024 17727 20058
rect 17761 20055 17773 20058
rect 18291 20058 18349 20064
rect 18291 20055 18303 20058
rect 17761 20027 18303 20055
rect 17761 20024 17773 20027
rect 17715 20018 17773 20024
rect 18291 20024 18303 20027
rect 18337 20024 18349 20058
rect 18291 20018 18349 20024
rect 18963 20058 19021 20064
rect 18963 20024 18975 20058
rect 19009 20055 19021 20058
rect 19539 20058 19597 20064
rect 19539 20055 19551 20058
rect 19009 20027 19551 20055
rect 19009 20024 19021 20027
rect 18963 20018 19021 20024
rect 19539 20024 19551 20027
rect 19585 20024 19597 20058
rect 19539 20018 19597 20024
rect 20211 20058 20269 20064
rect 20211 20024 20223 20058
rect 20257 20055 20269 20058
rect 20787 20058 20845 20064
rect 20787 20055 20799 20058
rect 20257 20027 20799 20055
rect 20257 20024 20269 20027
rect 20211 20018 20269 20024
rect 20787 20024 20799 20027
rect 20833 20024 20845 20058
rect 20787 20018 20845 20024
rect 21459 20058 21517 20064
rect 21459 20024 21471 20058
rect 21505 20055 21517 20058
rect 22035 20058 22093 20064
rect 22035 20055 22047 20058
rect 21505 20027 22047 20055
rect 21505 20024 21517 20027
rect 21459 20018 21517 20024
rect 22035 20024 22047 20027
rect 22081 20024 22093 20058
rect 22035 20018 22093 20024
rect 1952 19734 23264 19756
rect 1952 19682 7158 19734
rect 7210 19682 7222 19734
rect 7274 19682 7286 19734
rect 7338 19682 7350 19734
rect 7402 19682 12486 19734
rect 12538 19682 12550 19734
rect 12602 19682 12614 19734
rect 12666 19682 12678 19734
rect 12730 19682 17814 19734
rect 17866 19682 17878 19734
rect 17930 19682 17942 19734
rect 17994 19682 18006 19734
rect 18058 19682 23264 19734
rect 1952 19660 23264 19682
rect 2736 19611 2742 19623
rect 2697 19583 2742 19611
rect 2736 19571 2742 19583
rect 2794 19571 2800 19623
rect 2064 19389 2070 19401
rect 2025 19361 2070 19389
rect 2064 19349 2070 19361
rect 2122 19349 2128 19401
rect 3411 19392 3469 19398
rect 3411 19358 3423 19392
rect 3457 19389 3469 19392
rect 5235 19392 5293 19398
rect 5235 19389 5247 19392
rect 3457 19361 5247 19389
rect 3457 19358 3469 19361
rect 3411 19352 3469 19358
rect 5235 19358 5247 19361
rect 5281 19358 5293 19392
rect 5235 19352 5293 19358
rect 5907 19392 5965 19398
rect 5907 19358 5919 19392
rect 5953 19389 5965 19392
rect 7731 19392 7789 19398
rect 7731 19389 7743 19392
rect 5953 19361 7743 19389
rect 5953 19358 5965 19361
rect 5907 19352 5965 19358
rect 7731 19358 7743 19361
rect 7777 19358 7789 19392
rect 8979 19392 9037 19398
rect 8979 19389 8991 19392
rect 7731 19352 7789 19358
rect 8322 19361 8991 19389
rect 2352 19315 2358 19327
rect 2313 19287 2358 19315
rect 2352 19275 2358 19287
rect 2410 19275 2416 19327
rect 4659 19318 4717 19324
rect 4659 19284 4671 19318
rect 4705 19284 4717 19318
rect 4659 19278 4717 19284
rect 7155 19318 7213 19324
rect 7155 19284 7167 19318
rect 7201 19315 7213 19318
rect 8322 19315 8350 19361
rect 8979 19358 8991 19361
rect 9025 19358 9037 19392
rect 8979 19352 9037 19358
rect 9651 19392 9709 19398
rect 9651 19358 9663 19392
rect 9697 19389 9709 19392
rect 11475 19392 11533 19398
rect 11475 19389 11487 19392
rect 9697 19361 11487 19389
rect 9697 19358 9709 19361
rect 9651 19352 9709 19358
rect 11475 19358 11487 19361
rect 11521 19358 11533 19392
rect 11475 19352 11533 19358
rect 12147 19392 12205 19398
rect 12147 19358 12159 19392
rect 12193 19389 12205 19392
rect 13971 19392 14029 19398
rect 13971 19389 13983 19392
rect 12193 19361 13983 19389
rect 12193 19358 12205 19361
rect 12147 19352 12205 19358
rect 13971 19358 13983 19361
rect 14017 19358 14029 19392
rect 13971 19352 14029 19358
rect 14547 19392 14605 19398
rect 14547 19358 14559 19392
rect 14593 19389 14605 19392
rect 16467 19392 16525 19398
rect 16467 19389 16479 19392
rect 14593 19361 16479 19389
rect 14593 19358 14605 19361
rect 14547 19352 14605 19358
rect 16467 19358 16479 19361
rect 16513 19358 16525 19392
rect 16467 19352 16525 19358
rect 17139 19392 17197 19398
rect 17139 19358 17151 19392
rect 17185 19389 17197 19392
rect 18963 19392 19021 19398
rect 18963 19389 18975 19392
rect 17185 19361 18975 19389
rect 17185 19358 17197 19361
rect 17139 19352 17197 19358
rect 18963 19358 18975 19361
rect 19009 19358 19021 19392
rect 18963 19352 19021 19358
rect 19635 19392 19693 19398
rect 19635 19358 19647 19392
rect 19681 19389 19693 19392
rect 21459 19392 21517 19398
rect 21459 19389 21471 19392
rect 19681 19361 21471 19389
rect 19681 19358 19693 19361
rect 19635 19352 19693 19358
rect 21459 19358 21471 19361
rect 21505 19358 21517 19392
rect 21459 19352 21517 19358
rect 7201 19287 8350 19315
rect 8403 19318 8461 19324
rect 7201 19284 7213 19287
rect 7155 19278 7213 19284
rect 8403 19284 8415 19318
rect 8449 19315 8461 19318
rect 10227 19318 10285 19324
rect 10227 19315 10239 19318
rect 8449 19287 10239 19315
rect 8449 19284 8461 19287
rect 8403 19278 8461 19284
rect 10227 19284 10239 19287
rect 10273 19284 10285 19318
rect 10227 19278 10285 19284
rect 10899 19318 10957 19324
rect 10899 19284 10911 19318
rect 10945 19315 10957 19318
rect 12723 19318 12781 19324
rect 12723 19315 12735 19318
rect 10945 19287 12735 19315
rect 10945 19284 10957 19287
rect 10899 19278 10957 19284
rect 12723 19284 12735 19287
rect 12769 19284 12781 19318
rect 12723 19278 12781 19284
rect 13395 19318 13453 19324
rect 13395 19284 13407 19318
rect 13441 19315 13453 19318
rect 15219 19318 15277 19324
rect 15219 19315 15231 19318
rect 13441 19287 15231 19315
rect 13441 19284 13453 19287
rect 13395 19278 13453 19284
rect 15219 19284 15231 19287
rect 15265 19284 15277 19318
rect 15219 19278 15277 19284
rect 15891 19318 15949 19324
rect 15891 19284 15903 19318
rect 15937 19315 15949 19318
rect 17715 19318 17773 19324
rect 17715 19315 17727 19318
rect 15937 19287 17727 19315
rect 15937 19284 15949 19287
rect 15891 19278 15949 19284
rect 17715 19284 17727 19287
rect 17761 19284 17773 19318
rect 17715 19278 17773 19284
rect 18387 19318 18445 19324
rect 18387 19284 18399 19318
rect 18433 19315 18445 19318
rect 20211 19318 20269 19324
rect 20211 19315 20223 19318
rect 18433 19287 20223 19315
rect 18433 19284 18445 19287
rect 18387 19278 18445 19284
rect 20211 19284 20223 19287
rect 20257 19284 20269 19318
rect 20211 19278 20269 19284
rect 20883 19318 20941 19324
rect 20883 19284 20895 19318
rect 20929 19284 20941 19318
rect 20883 19278 20941 19284
rect 22131 19318 22189 19324
rect 22131 19284 22143 19318
rect 22177 19315 22189 19318
rect 22608 19315 22614 19327
rect 22177 19287 22614 19315
rect 22177 19284 22189 19287
rect 22131 19278 22189 19284
rect 2259 19244 2317 19250
rect 2259 19210 2271 19244
rect 2305 19241 2317 19244
rect 3987 19244 4045 19250
rect 3987 19241 3999 19244
rect 2305 19213 3999 19241
rect 2305 19210 2317 19213
rect 2259 19204 2317 19210
rect 3987 19210 3999 19213
rect 4033 19210 4045 19244
rect 4674 19241 4702 19278
rect 6483 19244 6541 19250
rect 6483 19241 6495 19244
rect 4674 19213 6495 19241
rect 3987 19204 4045 19210
rect 6483 19210 6495 19213
rect 6529 19210 6541 19244
rect 20898 19241 20926 19278
rect 22608 19275 22614 19287
rect 22666 19275 22672 19327
rect 22707 19244 22765 19250
rect 22707 19241 22719 19244
rect 20898 19213 22719 19241
rect 6483 19204 6541 19210
rect 22707 19210 22719 19213
rect 22753 19210 22765 19244
rect 22707 19204 22765 19210
rect 1952 19068 23264 19090
rect 1952 19016 4494 19068
rect 4546 19016 4558 19068
rect 4610 19016 4622 19068
rect 4674 19016 4686 19068
rect 4738 19016 9822 19068
rect 9874 19016 9886 19068
rect 9938 19016 9950 19068
rect 10002 19016 10014 19068
rect 10066 19016 15150 19068
rect 15202 19016 15214 19068
rect 15266 19016 15278 19068
rect 15330 19016 15342 19068
rect 15394 19016 20478 19068
rect 20530 19016 20542 19068
rect 20594 19016 20606 19068
rect 20658 19016 20670 19068
rect 20722 19016 23264 19068
rect 1952 18994 23264 19016
rect 22608 18831 22614 18883
rect 22666 18871 22672 18883
rect 22707 18874 22765 18880
rect 22707 18871 22719 18874
rect 22666 18843 22719 18871
rect 22666 18831 22672 18843
rect 22707 18840 22719 18843
rect 22753 18840 22765 18874
rect 22707 18834 22765 18840
rect 3411 18726 3469 18732
rect 3411 18692 3423 18726
rect 3457 18723 3469 18726
rect 3888 18723 3894 18735
rect 3457 18695 3894 18723
rect 3457 18692 3469 18695
rect 3411 18686 3469 18692
rect 3888 18683 3894 18695
rect 3946 18683 3952 18735
rect 3987 18726 4045 18732
rect 3987 18692 3999 18726
rect 4033 18723 4045 18726
rect 4563 18726 4621 18732
rect 4563 18723 4575 18726
rect 4033 18695 4575 18723
rect 4033 18692 4045 18695
rect 3987 18686 4045 18692
rect 4563 18692 4575 18695
rect 4609 18692 4621 18726
rect 4563 18686 4621 18692
rect 5235 18726 5293 18732
rect 5235 18692 5247 18726
rect 5281 18723 5293 18726
rect 5811 18726 5869 18732
rect 5811 18723 5823 18726
rect 5281 18695 5823 18723
rect 5281 18692 5293 18695
rect 5235 18686 5293 18692
rect 5811 18692 5823 18695
rect 5857 18692 5869 18726
rect 5811 18686 5869 18692
rect 6483 18726 6541 18732
rect 6483 18692 6495 18726
rect 6529 18723 6541 18726
rect 7059 18726 7117 18732
rect 7059 18723 7071 18726
rect 6529 18695 7071 18723
rect 6529 18692 6541 18695
rect 6483 18686 6541 18692
rect 7059 18692 7071 18695
rect 7105 18692 7117 18726
rect 7059 18686 7117 18692
rect 7731 18726 7789 18732
rect 7731 18692 7743 18726
rect 7777 18723 7789 18726
rect 8307 18726 8365 18732
rect 8307 18723 8319 18726
rect 7777 18695 8319 18723
rect 7777 18692 7789 18695
rect 7731 18686 7789 18692
rect 8307 18692 8319 18695
rect 8353 18692 8365 18726
rect 8307 18686 8365 18692
rect 8979 18726 9037 18732
rect 8979 18692 8991 18726
rect 9025 18723 9037 18726
rect 9555 18726 9613 18732
rect 9555 18723 9567 18726
rect 9025 18695 9567 18723
rect 9025 18692 9037 18695
rect 8979 18686 9037 18692
rect 9555 18692 9567 18695
rect 9601 18692 9613 18726
rect 9555 18686 9613 18692
rect 10227 18726 10285 18732
rect 10227 18692 10239 18726
rect 10273 18723 10285 18726
rect 10803 18726 10861 18732
rect 10803 18723 10815 18726
rect 10273 18695 10815 18723
rect 10273 18692 10285 18695
rect 10227 18686 10285 18692
rect 10803 18692 10815 18695
rect 10849 18692 10861 18726
rect 10803 18686 10861 18692
rect 11475 18726 11533 18732
rect 11475 18692 11487 18726
rect 11521 18723 11533 18726
rect 12051 18726 12109 18732
rect 12051 18723 12063 18726
rect 11521 18695 12063 18723
rect 11521 18692 11533 18695
rect 11475 18686 11533 18692
rect 12051 18692 12063 18695
rect 12097 18692 12109 18726
rect 12051 18686 12109 18692
rect 12723 18726 12781 18732
rect 12723 18692 12735 18726
rect 12769 18723 12781 18726
rect 13299 18726 13357 18732
rect 13299 18723 13311 18726
rect 12769 18695 13311 18723
rect 12769 18692 12781 18695
rect 12723 18686 12781 18692
rect 13299 18692 13311 18695
rect 13345 18692 13357 18726
rect 13299 18686 13357 18692
rect 13971 18726 14029 18732
rect 13971 18692 13983 18726
rect 14017 18723 14029 18726
rect 14547 18726 14605 18732
rect 14547 18723 14559 18726
rect 14017 18695 14559 18723
rect 14017 18692 14029 18695
rect 13971 18686 14029 18692
rect 14547 18692 14559 18695
rect 14593 18692 14605 18726
rect 14547 18686 14605 18692
rect 15219 18726 15277 18732
rect 15219 18692 15231 18726
rect 15265 18723 15277 18726
rect 15795 18726 15853 18732
rect 15795 18723 15807 18726
rect 15265 18695 15807 18723
rect 15265 18692 15277 18695
rect 15219 18686 15277 18692
rect 15795 18692 15807 18695
rect 15841 18692 15853 18726
rect 15795 18686 15853 18692
rect 16467 18726 16525 18732
rect 16467 18692 16479 18726
rect 16513 18723 16525 18726
rect 17043 18726 17101 18732
rect 17043 18723 17055 18726
rect 16513 18695 17055 18723
rect 16513 18692 16525 18695
rect 16467 18686 16525 18692
rect 17043 18692 17055 18695
rect 17089 18692 17101 18726
rect 17043 18686 17101 18692
rect 17715 18726 17773 18732
rect 17715 18692 17727 18726
rect 17761 18723 17773 18726
rect 18291 18726 18349 18732
rect 18291 18723 18303 18726
rect 17761 18695 18303 18723
rect 17761 18692 17773 18695
rect 17715 18686 17773 18692
rect 18291 18692 18303 18695
rect 18337 18692 18349 18726
rect 18291 18686 18349 18692
rect 18963 18726 19021 18732
rect 18963 18692 18975 18726
rect 19009 18723 19021 18726
rect 19539 18726 19597 18732
rect 19539 18723 19551 18726
rect 19009 18695 19551 18723
rect 19009 18692 19021 18695
rect 18963 18686 19021 18692
rect 19539 18692 19551 18695
rect 19585 18692 19597 18726
rect 19539 18686 19597 18692
rect 20211 18726 20269 18732
rect 20211 18692 20223 18726
rect 20257 18723 20269 18726
rect 20787 18726 20845 18732
rect 20787 18723 20799 18726
rect 20257 18695 20799 18723
rect 20257 18692 20269 18695
rect 20211 18686 20269 18692
rect 20787 18692 20799 18695
rect 20833 18692 20845 18726
rect 20787 18686 20845 18692
rect 21459 18726 21517 18732
rect 21459 18692 21471 18726
rect 21505 18723 21517 18726
rect 22035 18726 22093 18732
rect 22035 18723 22047 18726
rect 21505 18695 22047 18723
rect 21505 18692 21517 18695
rect 21459 18686 21517 18692
rect 22035 18692 22047 18695
rect 22081 18692 22093 18726
rect 22035 18686 22093 18692
rect 1952 18402 23264 18424
rect 1952 18350 7158 18402
rect 7210 18350 7222 18402
rect 7274 18350 7286 18402
rect 7338 18350 7350 18402
rect 7402 18350 12486 18402
rect 12538 18350 12550 18402
rect 12602 18350 12614 18402
rect 12666 18350 12678 18402
rect 12730 18350 17814 18402
rect 17866 18350 17878 18402
rect 17930 18350 17942 18402
rect 17994 18350 18006 18402
rect 18058 18350 23264 18402
rect 1952 18328 23264 18350
rect 3888 18091 3894 18143
rect 3946 18131 3952 18143
rect 3987 18134 4045 18140
rect 3987 18131 3999 18134
rect 3946 18103 3999 18131
rect 3946 18091 3952 18103
rect 3987 18100 3999 18103
rect 4033 18100 4045 18134
rect 3987 18094 4045 18100
rect 3411 18060 3469 18066
rect 3411 18026 3423 18060
rect 3457 18057 3469 18060
rect 5235 18060 5293 18066
rect 5235 18057 5247 18060
rect 3457 18029 5247 18057
rect 3457 18026 3469 18029
rect 3411 18020 3469 18026
rect 5235 18026 5247 18029
rect 5281 18026 5293 18060
rect 5235 18020 5293 18026
rect 5907 18060 5965 18066
rect 5907 18026 5919 18060
rect 5953 18057 5965 18060
rect 7731 18060 7789 18066
rect 7731 18057 7743 18060
rect 5953 18029 7743 18057
rect 5953 18026 5965 18029
rect 5907 18020 5965 18026
rect 7731 18026 7743 18029
rect 7777 18026 7789 18060
rect 8979 18060 9037 18066
rect 8979 18057 8991 18060
rect 7731 18020 7789 18026
rect 8322 18029 8991 18057
rect 4659 17986 4717 17992
rect 4659 17952 4671 17986
rect 4705 17952 4717 17986
rect 4659 17946 4717 17952
rect 7155 17986 7213 17992
rect 7155 17952 7167 17986
rect 7201 17983 7213 17986
rect 8322 17983 8350 18029
rect 8979 18026 8991 18029
rect 9025 18026 9037 18060
rect 8979 18020 9037 18026
rect 9651 18060 9709 18066
rect 9651 18026 9663 18060
rect 9697 18057 9709 18060
rect 11475 18060 11533 18066
rect 11475 18057 11487 18060
rect 9697 18029 11487 18057
rect 9697 18026 9709 18029
rect 9651 18020 9709 18026
rect 11475 18026 11487 18029
rect 11521 18026 11533 18060
rect 11475 18020 11533 18026
rect 12147 18060 12205 18066
rect 12147 18026 12159 18060
rect 12193 18057 12205 18060
rect 13971 18060 14029 18066
rect 13971 18057 13983 18060
rect 12193 18029 13983 18057
rect 12193 18026 12205 18029
rect 12147 18020 12205 18026
rect 13971 18026 13983 18029
rect 14017 18026 14029 18060
rect 13971 18020 14029 18026
rect 14547 18060 14605 18066
rect 14547 18026 14559 18060
rect 14593 18057 14605 18060
rect 16467 18060 16525 18066
rect 16467 18057 16479 18060
rect 14593 18029 16479 18057
rect 14593 18026 14605 18029
rect 14547 18020 14605 18026
rect 16467 18026 16479 18029
rect 16513 18026 16525 18060
rect 16467 18020 16525 18026
rect 17139 18060 17197 18066
rect 17139 18026 17151 18060
rect 17185 18057 17197 18060
rect 18963 18060 19021 18066
rect 18963 18057 18975 18060
rect 17185 18029 18975 18057
rect 17185 18026 17197 18029
rect 17139 18020 17197 18026
rect 18963 18026 18975 18029
rect 19009 18026 19021 18060
rect 18963 18020 19021 18026
rect 19635 18060 19693 18066
rect 19635 18026 19647 18060
rect 19681 18057 19693 18060
rect 21459 18060 21517 18066
rect 21459 18057 21471 18060
rect 19681 18029 21471 18057
rect 19681 18026 19693 18029
rect 19635 18020 19693 18026
rect 21459 18026 21471 18029
rect 21505 18026 21517 18060
rect 21459 18020 21517 18026
rect 7201 17955 8350 17983
rect 8403 17986 8461 17992
rect 7201 17952 7213 17955
rect 7155 17946 7213 17952
rect 8403 17952 8415 17986
rect 8449 17983 8461 17986
rect 10227 17986 10285 17992
rect 10227 17983 10239 17986
rect 8449 17955 10239 17983
rect 8449 17952 8461 17955
rect 8403 17946 8461 17952
rect 10227 17952 10239 17955
rect 10273 17952 10285 17986
rect 10227 17946 10285 17952
rect 10899 17986 10957 17992
rect 10899 17952 10911 17986
rect 10945 17983 10957 17986
rect 12723 17986 12781 17992
rect 12723 17983 12735 17986
rect 10945 17955 12735 17983
rect 10945 17952 10957 17955
rect 10899 17946 10957 17952
rect 12723 17952 12735 17955
rect 12769 17952 12781 17986
rect 12723 17946 12781 17952
rect 13395 17986 13453 17992
rect 13395 17952 13407 17986
rect 13441 17983 13453 17986
rect 15219 17986 15277 17992
rect 15219 17983 15231 17986
rect 13441 17955 15231 17983
rect 13441 17952 13453 17955
rect 13395 17946 13453 17952
rect 15219 17952 15231 17955
rect 15265 17952 15277 17986
rect 15219 17946 15277 17952
rect 15891 17986 15949 17992
rect 15891 17952 15903 17986
rect 15937 17983 15949 17986
rect 17715 17986 17773 17992
rect 17715 17983 17727 17986
rect 15937 17955 17727 17983
rect 15937 17952 15949 17955
rect 15891 17946 15949 17952
rect 17715 17952 17727 17955
rect 17761 17952 17773 17986
rect 17715 17946 17773 17952
rect 18387 17986 18445 17992
rect 18387 17952 18399 17986
rect 18433 17983 18445 17986
rect 20211 17986 20269 17992
rect 20211 17983 20223 17986
rect 18433 17955 20223 17983
rect 18433 17952 18445 17955
rect 18387 17946 18445 17952
rect 20211 17952 20223 17955
rect 20257 17952 20269 17986
rect 20211 17946 20269 17952
rect 20883 17986 20941 17992
rect 20883 17952 20895 17986
rect 20929 17952 20941 17986
rect 22128 17983 22134 17995
rect 22089 17955 22134 17983
rect 20883 17946 20941 17952
rect 4674 17909 4702 17946
rect 6483 17912 6541 17918
rect 6483 17909 6495 17912
rect 4674 17881 6495 17909
rect 6483 17878 6495 17881
rect 6529 17878 6541 17912
rect 20898 17909 20926 17946
rect 22128 17943 22134 17955
rect 22186 17943 22192 17995
rect 22707 17912 22765 17918
rect 22707 17909 22719 17912
rect 20898 17881 22719 17909
rect 6483 17872 6541 17878
rect 22707 17878 22719 17881
rect 22753 17878 22765 17912
rect 22707 17872 22765 17878
rect 1952 17736 23264 17758
rect 1952 17684 4494 17736
rect 4546 17684 4558 17736
rect 4610 17684 4622 17736
rect 4674 17684 4686 17736
rect 4738 17684 9822 17736
rect 9874 17684 9886 17736
rect 9938 17684 9950 17736
rect 10002 17684 10014 17736
rect 10066 17684 15150 17736
rect 15202 17684 15214 17736
rect 15266 17684 15278 17736
rect 15330 17684 15342 17736
rect 15394 17684 20478 17736
rect 20530 17684 20542 17736
rect 20594 17684 20606 17736
rect 20658 17684 20670 17736
rect 20722 17684 23264 17736
rect 1952 17662 23264 17684
rect 22128 17573 22134 17625
rect 22186 17613 22192 17625
rect 22707 17616 22765 17622
rect 22707 17613 22719 17616
rect 22186 17585 22719 17613
rect 22186 17573 22192 17585
rect 22707 17582 22719 17585
rect 22753 17582 22765 17616
rect 22707 17576 22765 17582
rect 2352 17425 2358 17477
rect 2410 17465 2416 17477
rect 3315 17468 3373 17474
rect 3315 17465 3327 17468
rect 2410 17437 3327 17465
rect 2410 17425 2416 17437
rect 3315 17434 3327 17437
rect 3361 17434 3373 17468
rect 3315 17428 3373 17434
rect 3987 17468 4045 17474
rect 3987 17434 3999 17468
rect 4033 17465 4045 17468
rect 4563 17468 4621 17474
rect 4563 17465 4575 17468
rect 4033 17437 4575 17465
rect 4033 17434 4045 17437
rect 3987 17428 4045 17434
rect 4563 17434 4575 17437
rect 4609 17434 4621 17468
rect 4563 17428 4621 17434
rect 5235 17468 5293 17474
rect 5235 17434 5247 17468
rect 5281 17465 5293 17468
rect 5811 17468 5869 17474
rect 5811 17465 5823 17468
rect 5281 17437 5823 17465
rect 5281 17434 5293 17437
rect 5235 17428 5293 17434
rect 5811 17434 5823 17437
rect 5857 17434 5869 17468
rect 5811 17428 5869 17434
rect 6483 17468 6541 17474
rect 6483 17434 6495 17468
rect 6529 17465 6541 17468
rect 7059 17468 7117 17474
rect 7059 17465 7071 17468
rect 6529 17437 7071 17465
rect 6529 17434 6541 17437
rect 6483 17428 6541 17434
rect 7059 17434 7071 17437
rect 7105 17434 7117 17468
rect 7059 17428 7117 17434
rect 7731 17468 7789 17474
rect 7731 17434 7743 17468
rect 7777 17465 7789 17468
rect 8307 17468 8365 17474
rect 8307 17465 8319 17468
rect 7777 17437 8319 17465
rect 7777 17434 7789 17437
rect 7731 17428 7789 17434
rect 8307 17434 8319 17437
rect 8353 17434 8365 17468
rect 8307 17428 8365 17434
rect 8979 17468 9037 17474
rect 8979 17434 8991 17468
rect 9025 17465 9037 17468
rect 9555 17468 9613 17474
rect 9555 17465 9567 17468
rect 9025 17437 9567 17465
rect 9025 17434 9037 17437
rect 8979 17428 9037 17434
rect 9555 17434 9567 17437
rect 9601 17434 9613 17468
rect 9555 17428 9613 17434
rect 10227 17468 10285 17474
rect 10227 17434 10239 17468
rect 10273 17465 10285 17468
rect 10803 17468 10861 17474
rect 10803 17465 10815 17468
rect 10273 17437 10815 17465
rect 10273 17434 10285 17437
rect 10227 17428 10285 17434
rect 10803 17434 10815 17437
rect 10849 17434 10861 17468
rect 10803 17428 10861 17434
rect 11475 17468 11533 17474
rect 11475 17434 11487 17468
rect 11521 17465 11533 17468
rect 12051 17468 12109 17474
rect 12051 17465 12063 17468
rect 11521 17437 12063 17465
rect 11521 17434 11533 17437
rect 11475 17428 11533 17434
rect 12051 17434 12063 17437
rect 12097 17434 12109 17468
rect 12051 17428 12109 17434
rect 12723 17468 12781 17474
rect 12723 17434 12735 17468
rect 12769 17465 12781 17468
rect 13299 17468 13357 17474
rect 13299 17465 13311 17468
rect 12769 17437 13311 17465
rect 12769 17434 12781 17437
rect 12723 17428 12781 17434
rect 13299 17434 13311 17437
rect 13345 17434 13357 17468
rect 13299 17428 13357 17434
rect 13971 17468 14029 17474
rect 13971 17434 13983 17468
rect 14017 17465 14029 17468
rect 14547 17468 14605 17474
rect 14547 17465 14559 17468
rect 14017 17437 14559 17465
rect 14017 17434 14029 17437
rect 13971 17428 14029 17434
rect 14547 17434 14559 17437
rect 14593 17434 14605 17468
rect 14547 17428 14605 17434
rect 15219 17468 15277 17474
rect 15219 17434 15231 17468
rect 15265 17465 15277 17468
rect 15795 17468 15853 17474
rect 15795 17465 15807 17468
rect 15265 17437 15807 17465
rect 15265 17434 15277 17437
rect 15219 17428 15277 17434
rect 15795 17434 15807 17437
rect 15841 17434 15853 17468
rect 15795 17428 15853 17434
rect 16467 17468 16525 17474
rect 16467 17434 16479 17468
rect 16513 17465 16525 17468
rect 17043 17468 17101 17474
rect 17043 17465 17055 17468
rect 16513 17437 17055 17465
rect 16513 17434 16525 17437
rect 16467 17428 16525 17434
rect 17043 17434 17055 17437
rect 17089 17434 17101 17468
rect 17043 17428 17101 17434
rect 17715 17468 17773 17474
rect 17715 17434 17727 17468
rect 17761 17465 17773 17468
rect 18291 17468 18349 17474
rect 18291 17465 18303 17468
rect 17761 17437 18303 17465
rect 17761 17434 17773 17437
rect 17715 17428 17773 17434
rect 18291 17434 18303 17437
rect 18337 17434 18349 17468
rect 18291 17428 18349 17434
rect 18963 17468 19021 17474
rect 18963 17434 18975 17468
rect 19009 17465 19021 17468
rect 19539 17468 19597 17474
rect 19539 17465 19551 17468
rect 19009 17437 19551 17465
rect 19009 17434 19021 17437
rect 18963 17428 19021 17434
rect 19539 17434 19551 17437
rect 19585 17434 19597 17468
rect 19539 17428 19597 17434
rect 20211 17468 20269 17474
rect 20211 17434 20223 17468
rect 20257 17465 20269 17468
rect 20787 17468 20845 17474
rect 20787 17465 20799 17468
rect 20257 17437 20799 17465
rect 20257 17434 20269 17437
rect 20211 17428 20269 17434
rect 20787 17434 20799 17437
rect 20833 17434 20845 17468
rect 20787 17428 20845 17434
rect 21459 17468 21517 17474
rect 21459 17434 21471 17468
rect 21505 17465 21517 17468
rect 22035 17468 22093 17474
rect 22035 17465 22047 17468
rect 21505 17437 22047 17465
rect 21505 17434 21517 17437
rect 21459 17428 21517 17434
rect 22035 17434 22047 17437
rect 22081 17434 22093 17468
rect 22035 17428 22093 17434
rect 1952 17070 23264 17092
rect 1952 17018 7158 17070
rect 7210 17018 7222 17070
rect 7274 17018 7286 17070
rect 7338 17018 7350 17070
rect 7402 17018 12486 17070
rect 12538 17018 12550 17070
rect 12602 17018 12614 17070
rect 12666 17018 12678 17070
rect 12730 17018 17814 17070
rect 17866 17018 17878 17070
rect 17930 17018 17942 17070
rect 17994 17018 18006 17070
rect 18058 17018 23264 17070
rect 1952 16996 23264 17018
rect 2352 16907 2358 16959
rect 2410 16947 2416 16959
rect 2739 16950 2797 16956
rect 2739 16947 2751 16950
rect 2410 16919 2751 16947
rect 2410 16907 2416 16919
rect 2739 16916 2751 16919
rect 2785 16916 2797 16950
rect 2739 16910 2797 16916
rect 6483 16802 6541 16808
rect 6483 16799 6495 16802
rect 4674 16771 6495 16799
rect 2064 16725 2070 16737
rect 2025 16697 2070 16725
rect 2064 16685 2070 16697
rect 2122 16685 2128 16737
rect 4674 16734 4702 16771
rect 6483 16768 6495 16771
rect 6529 16768 6541 16802
rect 16467 16802 16525 16808
rect 16467 16799 16479 16802
rect 6483 16762 6541 16768
rect 15426 16771 16479 16799
rect 3987 16728 4045 16734
rect 3987 16725 3999 16728
rect 2466 16697 3999 16725
rect 2352 16651 2358 16663
rect 2313 16623 2358 16651
rect 2352 16611 2358 16623
rect 2410 16611 2416 16663
rect 2466 16660 2494 16697
rect 3987 16694 3999 16697
rect 4033 16694 4045 16728
rect 3987 16688 4045 16694
rect 4659 16728 4717 16734
rect 4659 16694 4671 16728
rect 4705 16694 4717 16728
rect 7731 16728 7789 16734
rect 7731 16725 7743 16728
rect 4659 16688 4717 16694
rect 6786 16697 7743 16725
rect 2451 16654 2509 16660
rect 2451 16620 2463 16654
rect 2497 16620 2509 16654
rect 2451 16614 2509 16620
rect 3411 16654 3469 16660
rect 3411 16620 3423 16654
rect 3457 16651 3469 16654
rect 5235 16654 5293 16660
rect 5235 16651 5247 16654
rect 3457 16623 5247 16651
rect 3457 16620 3469 16623
rect 3411 16614 3469 16620
rect 5235 16620 5247 16623
rect 5281 16620 5293 16654
rect 5235 16614 5293 16620
rect 5907 16654 5965 16660
rect 5907 16620 5919 16654
rect 5953 16651 5965 16654
rect 6786 16651 6814 16697
rect 7731 16694 7743 16697
rect 7777 16694 7789 16728
rect 7731 16688 7789 16694
rect 8403 16728 8461 16734
rect 8403 16694 8415 16728
rect 8449 16725 8461 16728
rect 10227 16728 10285 16734
rect 10227 16725 10239 16728
rect 8449 16697 10239 16725
rect 8449 16694 8461 16697
rect 8403 16688 8461 16694
rect 10227 16694 10239 16697
rect 10273 16694 10285 16728
rect 11475 16728 11533 16734
rect 11475 16725 11487 16728
rect 10227 16688 10285 16694
rect 10722 16697 11487 16725
rect 5953 16623 6814 16651
rect 7155 16654 7213 16660
rect 5953 16620 5965 16623
rect 5907 16614 5965 16620
rect 7155 16620 7167 16654
rect 7201 16651 7213 16654
rect 8979 16654 9037 16660
rect 8979 16651 8991 16654
rect 7201 16623 8991 16651
rect 7201 16620 7213 16623
rect 7155 16614 7213 16620
rect 8979 16620 8991 16623
rect 9025 16620 9037 16654
rect 8979 16614 9037 16620
rect 9651 16654 9709 16660
rect 9651 16620 9663 16654
rect 9697 16651 9709 16654
rect 10722 16651 10750 16697
rect 11475 16694 11487 16697
rect 11521 16694 11533 16728
rect 12723 16728 12781 16734
rect 12723 16725 12735 16728
rect 11475 16688 11533 16694
rect 11778 16697 12735 16725
rect 9697 16623 10750 16651
rect 10899 16654 10957 16660
rect 9697 16620 9709 16623
rect 9651 16614 9709 16620
rect 10899 16620 10911 16654
rect 10945 16651 10957 16654
rect 11778 16651 11806 16697
rect 12723 16694 12735 16697
rect 12769 16694 12781 16728
rect 12723 16688 12781 16694
rect 13395 16728 13453 16734
rect 13395 16694 13407 16728
rect 13441 16725 13453 16728
rect 15219 16728 15277 16734
rect 15219 16725 15231 16728
rect 13441 16697 15231 16725
rect 13441 16694 13453 16697
rect 13395 16688 13453 16694
rect 15219 16694 15231 16697
rect 15265 16694 15277 16728
rect 15219 16688 15277 16694
rect 10945 16623 11806 16651
rect 12147 16654 12205 16660
rect 10945 16620 10957 16623
rect 10899 16614 10957 16620
rect 12147 16620 12159 16654
rect 12193 16651 12205 16654
rect 13971 16654 14029 16660
rect 13971 16651 13983 16654
rect 12193 16623 13983 16651
rect 12193 16620 12205 16623
rect 12147 16614 12205 16620
rect 13971 16620 13983 16623
rect 14017 16620 14029 16654
rect 13971 16614 14029 16620
rect 14643 16654 14701 16660
rect 14643 16620 14655 16654
rect 14689 16651 14701 16654
rect 15426 16651 15454 16771
rect 16467 16768 16479 16771
rect 16513 16768 16525 16802
rect 21459 16802 21517 16808
rect 21459 16799 21471 16802
rect 16467 16762 16525 16768
rect 20802 16771 21471 16799
rect 17715 16728 17773 16734
rect 17715 16725 17727 16728
rect 16770 16697 17727 16725
rect 14689 16623 15454 16651
rect 15891 16654 15949 16660
rect 14689 16620 14701 16623
rect 14643 16614 14701 16620
rect 15891 16620 15903 16654
rect 15937 16651 15949 16654
rect 16770 16651 16798 16697
rect 17715 16694 17727 16697
rect 17761 16694 17773 16728
rect 17715 16688 17773 16694
rect 18387 16728 18445 16734
rect 18387 16694 18399 16728
rect 18433 16725 18445 16728
rect 20211 16728 20269 16734
rect 20211 16725 20223 16728
rect 18433 16697 20223 16725
rect 18433 16694 18445 16697
rect 18387 16688 18445 16694
rect 20211 16694 20223 16697
rect 20257 16694 20269 16728
rect 20211 16688 20269 16694
rect 15937 16623 16798 16651
rect 17139 16654 17197 16660
rect 15937 16620 15949 16623
rect 15891 16614 15949 16620
rect 17139 16620 17151 16654
rect 17185 16651 17197 16654
rect 18963 16654 19021 16660
rect 18963 16651 18975 16654
rect 17185 16623 18975 16651
rect 17185 16620 17197 16623
rect 17139 16614 17197 16620
rect 18963 16620 18975 16623
rect 19009 16620 19021 16654
rect 18963 16614 19021 16620
rect 19635 16654 19693 16660
rect 19635 16620 19647 16654
rect 19681 16651 19693 16654
rect 20802 16651 20830 16771
rect 21459 16768 21471 16771
rect 21505 16768 21517 16802
rect 21459 16762 21517 16768
rect 22707 16728 22765 16734
rect 22707 16725 22719 16728
rect 21762 16697 22719 16725
rect 19681 16623 20830 16651
rect 20883 16654 20941 16660
rect 19681 16620 19693 16623
rect 19635 16614 19693 16620
rect 20883 16620 20895 16654
rect 20929 16651 20941 16654
rect 21762 16651 21790 16697
rect 22707 16694 22719 16697
rect 22753 16694 22765 16728
rect 22707 16688 22765 16694
rect 20929 16623 21790 16651
rect 22131 16654 22189 16660
rect 20929 16620 20941 16623
rect 20883 16614 20941 16620
rect 22131 16620 22143 16654
rect 22177 16651 22189 16654
rect 22608 16651 22614 16663
rect 22177 16623 22614 16651
rect 22177 16620 22189 16623
rect 22131 16614 22189 16620
rect 22608 16611 22614 16623
rect 22666 16611 22672 16663
rect 1952 16404 23264 16426
rect 1952 16352 4494 16404
rect 4546 16352 4558 16404
rect 4610 16352 4622 16404
rect 4674 16352 4686 16404
rect 4738 16352 9822 16404
rect 9874 16352 9886 16404
rect 9938 16352 9950 16404
rect 10002 16352 10014 16404
rect 10066 16352 15150 16404
rect 15202 16352 15214 16404
rect 15266 16352 15278 16404
rect 15330 16352 15342 16404
rect 15394 16352 20478 16404
rect 20530 16352 20542 16404
rect 20594 16352 20606 16404
rect 20658 16352 20670 16404
rect 20722 16352 23264 16404
rect 1952 16330 23264 16352
rect 22608 16241 22614 16293
rect 22666 16281 22672 16293
rect 22707 16284 22765 16290
rect 22707 16281 22719 16284
rect 22666 16253 22719 16281
rect 22666 16241 22672 16253
rect 22707 16250 22719 16253
rect 22753 16250 22765 16284
rect 22707 16244 22765 16250
rect 3411 16062 3469 16068
rect 3411 16028 3423 16062
rect 3457 16059 3469 16062
rect 3888 16059 3894 16071
rect 3457 16031 3894 16059
rect 3457 16028 3469 16031
rect 3411 16022 3469 16028
rect 3888 16019 3894 16031
rect 3946 16019 3952 16071
rect 3987 16062 4045 16068
rect 3987 16028 3999 16062
rect 4033 16059 4045 16062
rect 4563 16062 4621 16068
rect 4563 16059 4575 16062
rect 4033 16031 4575 16059
rect 4033 16028 4045 16031
rect 3987 16022 4045 16028
rect 4563 16028 4575 16031
rect 4609 16028 4621 16062
rect 4563 16022 4621 16028
rect 5235 16062 5293 16068
rect 5235 16028 5247 16062
rect 5281 16059 5293 16062
rect 5811 16062 5869 16068
rect 5811 16059 5823 16062
rect 5281 16031 5823 16059
rect 5281 16028 5293 16031
rect 5235 16022 5293 16028
rect 5811 16028 5823 16031
rect 5857 16028 5869 16062
rect 5811 16022 5869 16028
rect 6483 16062 6541 16068
rect 6483 16028 6495 16062
rect 6529 16059 6541 16062
rect 7059 16062 7117 16068
rect 7059 16059 7071 16062
rect 6529 16031 7071 16059
rect 6529 16028 6541 16031
rect 6483 16022 6541 16028
rect 7059 16028 7071 16031
rect 7105 16028 7117 16062
rect 7059 16022 7117 16028
rect 7731 16062 7789 16068
rect 7731 16028 7743 16062
rect 7777 16059 7789 16062
rect 8307 16062 8365 16068
rect 8307 16059 8319 16062
rect 7777 16031 8319 16059
rect 7777 16028 7789 16031
rect 7731 16022 7789 16028
rect 8307 16028 8319 16031
rect 8353 16028 8365 16062
rect 8307 16022 8365 16028
rect 8979 16062 9037 16068
rect 8979 16028 8991 16062
rect 9025 16059 9037 16062
rect 9555 16062 9613 16068
rect 9555 16059 9567 16062
rect 9025 16031 9567 16059
rect 9025 16028 9037 16031
rect 8979 16022 9037 16028
rect 9555 16028 9567 16031
rect 9601 16028 9613 16062
rect 9555 16022 9613 16028
rect 10227 16062 10285 16068
rect 10227 16028 10239 16062
rect 10273 16059 10285 16062
rect 10803 16062 10861 16068
rect 10803 16059 10815 16062
rect 10273 16031 10815 16059
rect 10273 16028 10285 16031
rect 10227 16022 10285 16028
rect 10803 16028 10815 16031
rect 10849 16028 10861 16062
rect 10803 16022 10861 16028
rect 11475 16062 11533 16068
rect 11475 16028 11487 16062
rect 11521 16059 11533 16062
rect 12051 16062 12109 16068
rect 12051 16059 12063 16062
rect 11521 16031 12063 16059
rect 11521 16028 11533 16031
rect 11475 16022 11533 16028
rect 12051 16028 12063 16031
rect 12097 16028 12109 16062
rect 12051 16022 12109 16028
rect 12723 16062 12781 16068
rect 12723 16028 12735 16062
rect 12769 16059 12781 16062
rect 13299 16062 13357 16068
rect 13299 16059 13311 16062
rect 12769 16031 13311 16059
rect 12769 16028 12781 16031
rect 12723 16022 12781 16028
rect 13299 16028 13311 16031
rect 13345 16028 13357 16062
rect 13299 16022 13357 16028
rect 13971 16062 14029 16068
rect 13971 16028 13983 16062
rect 14017 16059 14029 16062
rect 14547 16062 14605 16068
rect 14547 16059 14559 16062
rect 14017 16031 14559 16059
rect 14017 16028 14029 16031
rect 13971 16022 14029 16028
rect 14547 16028 14559 16031
rect 14593 16028 14605 16062
rect 14547 16022 14605 16028
rect 15219 16062 15277 16068
rect 15219 16028 15231 16062
rect 15265 16059 15277 16062
rect 15795 16062 15853 16068
rect 15795 16059 15807 16062
rect 15265 16031 15807 16059
rect 15265 16028 15277 16031
rect 15219 16022 15277 16028
rect 15795 16028 15807 16031
rect 15841 16028 15853 16062
rect 15795 16022 15853 16028
rect 16467 16062 16525 16068
rect 16467 16028 16479 16062
rect 16513 16059 16525 16062
rect 17043 16062 17101 16068
rect 17043 16059 17055 16062
rect 16513 16031 17055 16059
rect 16513 16028 16525 16031
rect 16467 16022 16525 16028
rect 17043 16028 17055 16031
rect 17089 16028 17101 16062
rect 17043 16022 17101 16028
rect 17715 16062 17773 16068
rect 17715 16028 17727 16062
rect 17761 16059 17773 16062
rect 18291 16062 18349 16068
rect 18291 16059 18303 16062
rect 17761 16031 18303 16059
rect 17761 16028 17773 16031
rect 17715 16022 17773 16028
rect 18291 16028 18303 16031
rect 18337 16028 18349 16062
rect 18291 16022 18349 16028
rect 18963 16062 19021 16068
rect 18963 16028 18975 16062
rect 19009 16059 19021 16062
rect 19539 16062 19597 16068
rect 19539 16059 19551 16062
rect 19009 16031 19551 16059
rect 19009 16028 19021 16031
rect 18963 16022 19021 16028
rect 19539 16028 19551 16031
rect 19585 16028 19597 16062
rect 19539 16022 19597 16028
rect 20211 16062 20269 16068
rect 20211 16028 20223 16062
rect 20257 16059 20269 16062
rect 20787 16062 20845 16068
rect 20787 16059 20799 16062
rect 20257 16031 20799 16059
rect 20257 16028 20269 16031
rect 20211 16022 20269 16028
rect 20787 16028 20799 16031
rect 20833 16028 20845 16062
rect 20787 16022 20845 16028
rect 21459 16062 21517 16068
rect 21459 16028 21471 16062
rect 21505 16059 21517 16062
rect 22035 16062 22093 16068
rect 22035 16059 22047 16062
rect 21505 16031 22047 16059
rect 21505 16028 21517 16031
rect 21459 16022 21517 16028
rect 22035 16028 22047 16031
rect 22081 16028 22093 16062
rect 22035 16022 22093 16028
rect 1952 15738 23264 15760
rect 1952 15686 7158 15738
rect 7210 15686 7222 15738
rect 7274 15686 7286 15738
rect 7338 15686 7350 15738
rect 7402 15686 12486 15738
rect 12538 15686 12550 15738
rect 12602 15686 12614 15738
rect 12666 15686 12678 15738
rect 12730 15686 17814 15738
rect 17866 15686 17878 15738
rect 17930 15686 17942 15738
rect 17994 15686 18006 15738
rect 18058 15686 23264 15738
rect 1952 15664 23264 15686
rect 3888 15575 3894 15627
rect 3946 15615 3952 15627
rect 3987 15618 4045 15624
rect 3987 15615 3999 15618
rect 3946 15587 3999 15615
rect 3946 15575 3952 15587
rect 3987 15584 3999 15587
rect 4033 15584 4045 15618
rect 3987 15578 4045 15584
rect 3411 15396 3469 15402
rect 3411 15362 3423 15396
rect 3457 15393 3469 15396
rect 5235 15396 5293 15402
rect 5235 15393 5247 15396
rect 3457 15365 5247 15393
rect 3457 15362 3469 15365
rect 3411 15356 3469 15362
rect 5235 15362 5247 15365
rect 5281 15362 5293 15396
rect 5235 15356 5293 15362
rect 5907 15396 5965 15402
rect 5907 15362 5919 15396
rect 5953 15393 5965 15396
rect 7731 15396 7789 15402
rect 7731 15393 7743 15396
rect 5953 15365 7743 15393
rect 5953 15362 5965 15365
rect 5907 15356 5965 15362
rect 7731 15362 7743 15365
rect 7777 15362 7789 15396
rect 7731 15356 7789 15362
rect 8403 15396 8461 15402
rect 8403 15362 8415 15396
rect 8449 15393 8461 15396
rect 10227 15396 10285 15402
rect 10227 15393 10239 15396
rect 8449 15365 10239 15393
rect 8449 15362 8461 15365
rect 8403 15356 8461 15362
rect 10227 15362 10239 15365
rect 10273 15362 10285 15396
rect 10227 15356 10285 15362
rect 12147 15396 12205 15402
rect 12147 15362 12159 15396
rect 12193 15393 12205 15396
rect 13971 15396 14029 15402
rect 13971 15393 13983 15396
rect 12193 15365 13983 15393
rect 12193 15362 12205 15365
rect 12147 15356 12205 15362
rect 13971 15362 13983 15365
rect 14017 15362 14029 15396
rect 13971 15356 14029 15362
rect 14547 15396 14605 15402
rect 14547 15362 14559 15396
rect 14593 15393 14605 15396
rect 16467 15396 16525 15402
rect 16467 15393 16479 15396
rect 14593 15365 16479 15393
rect 14593 15362 14605 15365
rect 14547 15356 14605 15362
rect 16467 15362 16479 15365
rect 16513 15362 16525 15396
rect 16467 15356 16525 15362
rect 17139 15396 17197 15402
rect 17139 15362 17151 15396
rect 17185 15393 17197 15396
rect 18963 15396 19021 15402
rect 18963 15393 18975 15396
rect 17185 15365 18975 15393
rect 17185 15362 17197 15365
rect 17139 15356 17197 15362
rect 18963 15362 18975 15365
rect 19009 15362 19021 15396
rect 18963 15356 19021 15362
rect 19635 15396 19693 15402
rect 19635 15362 19647 15396
rect 19681 15393 19693 15396
rect 21459 15396 21517 15402
rect 21459 15393 21471 15396
rect 19681 15365 21471 15393
rect 19681 15362 19693 15365
rect 19635 15356 19693 15362
rect 21459 15362 21471 15365
rect 21505 15362 21517 15396
rect 21459 15356 21517 15362
rect 4659 15322 4717 15328
rect 4659 15288 4671 15322
rect 4705 15288 4717 15322
rect 4659 15282 4717 15288
rect 7155 15322 7213 15328
rect 7155 15288 7167 15322
rect 7201 15319 7213 15322
rect 8979 15322 9037 15328
rect 8979 15319 8991 15322
rect 7201 15291 8991 15319
rect 7201 15288 7213 15291
rect 7155 15282 7213 15288
rect 8979 15288 8991 15291
rect 9025 15288 9037 15322
rect 8979 15282 9037 15288
rect 9555 15322 9613 15328
rect 9555 15288 9567 15322
rect 9601 15288 9613 15322
rect 9555 15282 9613 15288
rect 10899 15322 10957 15328
rect 10899 15288 10911 15322
rect 10945 15319 10957 15322
rect 12723 15322 12781 15328
rect 12723 15319 12735 15322
rect 10945 15291 12735 15319
rect 10945 15288 10957 15291
rect 10899 15282 10957 15288
rect 12723 15288 12735 15291
rect 12769 15288 12781 15322
rect 12723 15282 12781 15288
rect 13395 15322 13453 15328
rect 13395 15288 13407 15322
rect 13441 15319 13453 15322
rect 15219 15322 15277 15328
rect 15219 15319 15231 15322
rect 13441 15291 15231 15319
rect 13441 15288 13453 15291
rect 13395 15282 13453 15288
rect 15219 15288 15231 15291
rect 15265 15288 15277 15322
rect 15219 15282 15277 15288
rect 15891 15322 15949 15328
rect 15891 15288 15903 15322
rect 15937 15319 15949 15322
rect 17715 15322 17773 15328
rect 17715 15319 17727 15322
rect 15937 15291 17727 15319
rect 15937 15288 15949 15291
rect 15891 15282 15949 15288
rect 17715 15288 17727 15291
rect 17761 15288 17773 15322
rect 17715 15282 17773 15288
rect 18387 15322 18445 15328
rect 18387 15288 18399 15322
rect 18433 15319 18445 15322
rect 20211 15322 20269 15328
rect 20211 15319 20223 15322
rect 18433 15291 20223 15319
rect 18433 15288 18445 15291
rect 18387 15282 18445 15288
rect 20211 15288 20223 15291
rect 20257 15288 20269 15322
rect 20211 15282 20269 15288
rect 20883 15322 20941 15328
rect 20883 15288 20895 15322
rect 20929 15288 20941 15322
rect 20883 15282 20941 15288
rect 22131 15322 22189 15328
rect 22131 15288 22143 15322
rect 22177 15319 22189 15322
rect 22608 15319 22614 15331
rect 22177 15291 22614 15319
rect 22177 15288 22189 15291
rect 22131 15282 22189 15288
rect 4674 15245 4702 15282
rect 6483 15248 6541 15254
rect 6483 15245 6495 15248
rect 4674 15217 6495 15245
rect 6483 15214 6495 15217
rect 6529 15214 6541 15248
rect 9570 15245 9598 15282
rect 11475 15248 11533 15254
rect 11475 15245 11487 15248
rect 9570 15217 11487 15245
rect 6483 15208 6541 15214
rect 11475 15214 11487 15217
rect 11521 15214 11533 15248
rect 20898 15245 20926 15282
rect 22608 15279 22614 15291
rect 22666 15279 22672 15331
rect 22707 15248 22765 15254
rect 22707 15245 22719 15248
rect 20898 15217 22719 15245
rect 11475 15208 11533 15214
rect 22707 15214 22719 15217
rect 22753 15214 22765 15248
rect 22707 15208 22765 15214
rect 1952 15072 23264 15094
rect 1952 15020 4494 15072
rect 4546 15020 4558 15072
rect 4610 15020 4622 15072
rect 4674 15020 4686 15072
rect 4738 15020 9822 15072
rect 9874 15020 9886 15072
rect 9938 15020 9950 15072
rect 10002 15020 10014 15072
rect 10066 15020 15150 15072
rect 15202 15020 15214 15072
rect 15266 15020 15278 15072
rect 15330 15020 15342 15072
rect 15394 15020 20478 15072
rect 20530 15020 20542 15072
rect 20594 15020 20606 15072
rect 20658 15020 20670 15072
rect 20722 15020 23264 15072
rect 1952 14998 23264 15020
rect 22608 14909 22614 14961
rect 22666 14949 22672 14961
rect 22707 14952 22765 14958
rect 22707 14949 22719 14952
rect 22666 14921 22719 14949
rect 22666 14909 22672 14921
rect 22707 14918 22719 14921
rect 22753 14918 22765 14952
rect 22707 14912 22765 14918
rect 3411 14730 3469 14736
rect 3411 14696 3423 14730
rect 3457 14727 3469 14730
rect 3888 14727 3894 14739
rect 3457 14699 3894 14727
rect 3457 14696 3469 14699
rect 3411 14690 3469 14696
rect 3888 14687 3894 14699
rect 3946 14687 3952 14739
rect 3987 14730 4045 14736
rect 3987 14696 3999 14730
rect 4033 14727 4045 14730
rect 4563 14730 4621 14736
rect 4563 14727 4575 14730
rect 4033 14699 4575 14727
rect 4033 14696 4045 14699
rect 3987 14690 4045 14696
rect 4563 14696 4575 14699
rect 4609 14696 4621 14730
rect 4563 14690 4621 14696
rect 5235 14730 5293 14736
rect 5235 14696 5247 14730
rect 5281 14727 5293 14730
rect 5811 14730 5869 14736
rect 5811 14727 5823 14730
rect 5281 14699 5823 14727
rect 5281 14696 5293 14699
rect 5235 14690 5293 14696
rect 5811 14696 5823 14699
rect 5857 14696 5869 14730
rect 5811 14690 5869 14696
rect 6483 14730 6541 14736
rect 6483 14696 6495 14730
rect 6529 14727 6541 14730
rect 7059 14730 7117 14736
rect 7059 14727 7071 14730
rect 6529 14699 7071 14727
rect 6529 14696 6541 14699
rect 6483 14690 6541 14696
rect 7059 14696 7071 14699
rect 7105 14696 7117 14730
rect 7059 14690 7117 14696
rect 7731 14730 7789 14736
rect 7731 14696 7743 14730
rect 7777 14727 7789 14730
rect 8307 14730 8365 14736
rect 8307 14727 8319 14730
rect 7777 14699 8319 14727
rect 7777 14696 7789 14699
rect 7731 14690 7789 14696
rect 8307 14696 8319 14699
rect 8353 14696 8365 14730
rect 8307 14690 8365 14696
rect 8979 14730 9037 14736
rect 8979 14696 8991 14730
rect 9025 14727 9037 14730
rect 9555 14730 9613 14736
rect 9555 14727 9567 14730
rect 9025 14699 9567 14727
rect 9025 14696 9037 14699
rect 8979 14690 9037 14696
rect 9555 14696 9567 14699
rect 9601 14696 9613 14730
rect 9555 14690 9613 14696
rect 10227 14730 10285 14736
rect 10227 14696 10239 14730
rect 10273 14727 10285 14730
rect 10803 14730 10861 14736
rect 10803 14727 10815 14730
rect 10273 14699 10815 14727
rect 10273 14696 10285 14699
rect 10227 14690 10285 14696
rect 10803 14696 10815 14699
rect 10849 14696 10861 14730
rect 10803 14690 10861 14696
rect 11475 14730 11533 14736
rect 11475 14696 11487 14730
rect 11521 14727 11533 14730
rect 12051 14730 12109 14736
rect 12051 14727 12063 14730
rect 11521 14699 12063 14727
rect 11521 14696 11533 14699
rect 11475 14690 11533 14696
rect 12051 14696 12063 14699
rect 12097 14696 12109 14730
rect 12051 14690 12109 14696
rect 12723 14730 12781 14736
rect 12723 14696 12735 14730
rect 12769 14727 12781 14730
rect 13299 14730 13357 14736
rect 13299 14727 13311 14730
rect 12769 14699 13311 14727
rect 12769 14696 12781 14699
rect 12723 14690 12781 14696
rect 13299 14696 13311 14699
rect 13345 14696 13357 14730
rect 13299 14690 13357 14696
rect 13971 14730 14029 14736
rect 13971 14696 13983 14730
rect 14017 14727 14029 14730
rect 14547 14730 14605 14736
rect 14547 14727 14559 14730
rect 14017 14699 14559 14727
rect 14017 14696 14029 14699
rect 13971 14690 14029 14696
rect 14547 14696 14559 14699
rect 14593 14696 14605 14730
rect 14547 14690 14605 14696
rect 15219 14730 15277 14736
rect 15219 14696 15231 14730
rect 15265 14727 15277 14730
rect 15795 14730 15853 14736
rect 15795 14727 15807 14730
rect 15265 14699 15807 14727
rect 15265 14696 15277 14699
rect 15219 14690 15277 14696
rect 15795 14696 15807 14699
rect 15841 14696 15853 14730
rect 15795 14690 15853 14696
rect 16467 14730 16525 14736
rect 16467 14696 16479 14730
rect 16513 14727 16525 14730
rect 17043 14730 17101 14736
rect 17043 14727 17055 14730
rect 16513 14699 17055 14727
rect 16513 14696 16525 14699
rect 16467 14690 16525 14696
rect 17043 14696 17055 14699
rect 17089 14696 17101 14730
rect 17043 14690 17101 14696
rect 17715 14730 17773 14736
rect 17715 14696 17727 14730
rect 17761 14727 17773 14730
rect 18291 14730 18349 14736
rect 18291 14727 18303 14730
rect 17761 14699 18303 14727
rect 17761 14696 17773 14699
rect 17715 14690 17773 14696
rect 18291 14696 18303 14699
rect 18337 14696 18349 14730
rect 18291 14690 18349 14696
rect 18963 14730 19021 14736
rect 18963 14696 18975 14730
rect 19009 14727 19021 14730
rect 19539 14730 19597 14736
rect 19539 14727 19551 14730
rect 19009 14699 19551 14727
rect 19009 14696 19021 14699
rect 18963 14690 19021 14696
rect 19539 14696 19551 14699
rect 19585 14696 19597 14730
rect 19539 14690 19597 14696
rect 20211 14730 20269 14736
rect 20211 14696 20223 14730
rect 20257 14727 20269 14730
rect 20787 14730 20845 14736
rect 20787 14727 20799 14730
rect 20257 14699 20799 14727
rect 20257 14696 20269 14699
rect 20211 14690 20269 14696
rect 20787 14696 20799 14699
rect 20833 14696 20845 14730
rect 20787 14690 20845 14696
rect 21459 14730 21517 14736
rect 21459 14696 21471 14730
rect 21505 14727 21517 14730
rect 22035 14730 22093 14736
rect 22035 14727 22047 14730
rect 21505 14699 22047 14727
rect 21505 14696 21517 14699
rect 21459 14690 21517 14696
rect 22035 14696 22047 14699
rect 22081 14696 22093 14730
rect 22035 14690 22093 14696
rect 1952 14406 23264 14428
rect 1952 14354 7158 14406
rect 7210 14354 7222 14406
rect 7274 14354 7286 14406
rect 7338 14354 7350 14406
rect 7402 14354 12486 14406
rect 12538 14354 12550 14406
rect 12602 14354 12614 14406
rect 12666 14354 12678 14406
rect 12730 14354 17814 14406
rect 17866 14354 17878 14406
rect 17930 14354 17942 14406
rect 17994 14354 18006 14406
rect 18058 14354 23264 14406
rect 1952 14332 23264 14354
rect 3888 14243 3894 14295
rect 3946 14283 3952 14295
rect 3987 14286 4045 14292
rect 3987 14283 3999 14286
rect 3946 14255 3999 14283
rect 3946 14243 3952 14255
rect 3987 14252 3999 14255
rect 4033 14252 4045 14286
rect 3987 14246 4045 14252
rect 3411 14064 3469 14070
rect 3411 14030 3423 14064
rect 3457 14061 3469 14064
rect 5235 14064 5293 14070
rect 5235 14061 5247 14064
rect 3457 14033 5247 14061
rect 3457 14030 3469 14033
rect 3411 14024 3469 14030
rect 5235 14030 5247 14033
rect 5281 14030 5293 14064
rect 5235 14024 5293 14030
rect 5907 14064 5965 14070
rect 5907 14030 5919 14064
rect 5953 14061 5965 14064
rect 7731 14064 7789 14070
rect 7731 14061 7743 14064
rect 5953 14033 7743 14061
rect 5953 14030 5965 14033
rect 5907 14024 5965 14030
rect 7731 14030 7743 14033
rect 7777 14030 7789 14064
rect 7731 14024 7789 14030
rect 8403 14064 8461 14070
rect 8403 14030 8415 14064
rect 8449 14061 8461 14064
rect 10227 14064 10285 14070
rect 10227 14061 10239 14064
rect 8449 14033 10239 14061
rect 8449 14030 8461 14033
rect 8403 14024 8461 14030
rect 10227 14030 10239 14033
rect 10273 14030 10285 14064
rect 10227 14024 10285 14030
rect 12147 14064 12205 14070
rect 12147 14030 12159 14064
rect 12193 14061 12205 14064
rect 13971 14064 14029 14070
rect 13971 14061 13983 14064
rect 12193 14033 13983 14061
rect 12193 14030 12205 14033
rect 12147 14024 12205 14030
rect 13971 14030 13983 14033
rect 14017 14030 14029 14064
rect 13971 14024 14029 14030
rect 14547 14064 14605 14070
rect 14547 14030 14559 14064
rect 14593 14061 14605 14064
rect 16467 14064 16525 14070
rect 16467 14061 16479 14064
rect 14593 14033 16479 14061
rect 14593 14030 14605 14033
rect 14547 14024 14605 14030
rect 16467 14030 16479 14033
rect 16513 14030 16525 14064
rect 16467 14024 16525 14030
rect 17139 14064 17197 14070
rect 17139 14030 17151 14064
rect 17185 14061 17197 14064
rect 18963 14064 19021 14070
rect 18963 14061 18975 14064
rect 17185 14033 18975 14061
rect 17185 14030 17197 14033
rect 17139 14024 17197 14030
rect 18963 14030 18975 14033
rect 19009 14030 19021 14064
rect 18963 14024 19021 14030
rect 19635 14064 19693 14070
rect 19635 14030 19647 14064
rect 19681 14061 19693 14064
rect 21459 14064 21517 14070
rect 21459 14061 21471 14064
rect 19681 14033 21471 14061
rect 19681 14030 19693 14033
rect 19635 14024 19693 14030
rect 21459 14030 21471 14033
rect 21505 14030 21517 14064
rect 21459 14024 21517 14030
rect 4659 13990 4717 13996
rect 4659 13956 4671 13990
rect 4705 13956 4717 13990
rect 4659 13950 4717 13956
rect 7155 13990 7213 13996
rect 7155 13956 7167 13990
rect 7201 13987 7213 13990
rect 8979 13990 9037 13996
rect 8979 13987 8991 13990
rect 7201 13959 8991 13987
rect 7201 13956 7213 13959
rect 7155 13950 7213 13956
rect 8979 13956 8991 13959
rect 9025 13956 9037 13990
rect 8979 13950 9037 13956
rect 9555 13990 9613 13996
rect 9555 13956 9567 13990
rect 9601 13956 9613 13990
rect 9555 13950 9613 13956
rect 10899 13990 10957 13996
rect 10899 13956 10911 13990
rect 10945 13987 10957 13990
rect 12723 13990 12781 13996
rect 12723 13987 12735 13990
rect 10945 13959 12735 13987
rect 10945 13956 10957 13959
rect 10899 13950 10957 13956
rect 12723 13956 12735 13959
rect 12769 13956 12781 13990
rect 12723 13950 12781 13956
rect 13395 13990 13453 13996
rect 13395 13956 13407 13990
rect 13441 13987 13453 13990
rect 15219 13990 15277 13996
rect 15219 13987 15231 13990
rect 13441 13959 15231 13987
rect 13441 13956 13453 13959
rect 13395 13950 13453 13956
rect 15219 13956 15231 13959
rect 15265 13956 15277 13990
rect 15219 13950 15277 13956
rect 15891 13990 15949 13996
rect 15891 13956 15903 13990
rect 15937 13987 15949 13990
rect 17715 13990 17773 13996
rect 17715 13987 17727 13990
rect 15937 13959 17727 13987
rect 15937 13956 15949 13959
rect 15891 13950 15949 13956
rect 17715 13956 17727 13959
rect 17761 13956 17773 13990
rect 17715 13950 17773 13956
rect 18387 13990 18445 13996
rect 18387 13956 18399 13990
rect 18433 13987 18445 13990
rect 20211 13990 20269 13996
rect 20211 13987 20223 13990
rect 18433 13959 20223 13987
rect 18433 13956 18445 13959
rect 18387 13950 18445 13956
rect 20211 13956 20223 13959
rect 20257 13956 20269 13990
rect 20211 13950 20269 13956
rect 20883 13990 20941 13996
rect 20883 13956 20895 13990
rect 20929 13956 20941 13990
rect 20883 13950 20941 13956
rect 22131 13990 22189 13996
rect 22131 13956 22143 13990
rect 22177 13987 22189 13990
rect 22608 13987 22614 13999
rect 22177 13959 22614 13987
rect 22177 13956 22189 13959
rect 22131 13950 22189 13956
rect 4674 13913 4702 13950
rect 6483 13916 6541 13922
rect 6483 13913 6495 13916
rect 4674 13885 6495 13913
rect 6483 13882 6495 13885
rect 6529 13882 6541 13916
rect 9570 13913 9598 13950
rect 11475 13916 11533 13922
rect 11475 13913 11487 13916
rect 9570 13885 11487 13913
rect 6483 13876 6541 13882
rect 11475 13882 11487 13885
rect 11521 13882 11533 13916
rect 20898 13913 20926 13950
rect 22608 13947 22614 13959
rect 22666 13947 22672 13999
rect 22707 13916 22765 13922
rect 22707 13913 22719 13916
rect 20898 13885 22719 13913
rect 11475 13876 11533 13882
rect 22707 13882 22719 13885
rect 22753 13882 22765 13916
rect 22707 13876 22765 13882
rect 1952 13740 23264 13762
rect 1952 13688 4494 13740
rect 4546 13688 4558 13740
rect 4610 13688 4622 13740
rect 4674 13688 4686 13740
rect 4738 13688 9822 13740
rect 9874 13688 9886 13740
rect 9938 13688 9950 13740
rect 10002 13688 10014 13740
rect 10066 13688 15150 13740
rect 15202 13688 15214 13740
rect 15266 13688 15278 13740
rect 15330 13688 15342 13740
rect 15394 13688 20478 13740
rect 20530 13688 20542 13740
rect 20594 13688 20606 13740
rect 20658 13688 20670 13740
rect 20722 13688 23264 13740
rect 1952 13666 23264 13688
rect 22608 13503 22614 13555
rect 22666 13543 22672 13555
rect 22707 13546 22765 13552
rect 22707 13543 22719 13546
rect 22666 13515 22719 13543
rect 22666 13503 22672 13515
rect 22707 13512 22719 13515
rect 22753 13512 22765 13546
rect 22707 13506 22765 13512
rect 3411 13398 3469 13404
rect 3411 13364 3423 13398
rect 3457 13395 3469 13398
rect 3888 13395 3894 13407
rect 3457 13367 3894 13395
rect 3457 13364 3469 13367
rect 3411 13358 3469 13364
rect 3888 13355 3894 13367
rect 3946 13355 3952 13407
rect 3987 13398 4045 13404
rect 3987 13364 3999 13398
rect 4033 13395 4045 13398
rect 4563 13398 4621 13404
rect 4563 13395 4575 13398
rect 4033 13367 4575 13395
rect 4033 13364 4045 13367
rect 3987 13358 4045 13364
rect 4563 13364 4575 13367
rect 4609 13364 4621 13398
rect 4563 13358 4621 13364
rect 5235 13398 5293 13404
rect 5235 13364 5247 13398
rect 5281 13395 5293 13398
rect 5811 13398 5869 13404
rect 5811 13395 5823 13398
rect 5281 13367 5823 13395
rect 5281 13364 5293 13367
rect 5235 13358 5293 13364
rect 5811 13364 5823 13367
rect 5857 13364 5869 13398
rect 5811 13358 5869 13364
rect 6483 13398 6541 13404
rect 6483 13364 6495 13398
rect 6529 13395 6541 13398
rect 7059 13398 7117 13404
rect 7059 13395 7071 13398
rect 6529 13367 7071 13395
rect 6529 13364 6541 13367
rect 6483 13358 6541 13364
rect 7059 13364 7071 13367
rect 7105 13364 7117 13398
rect 7059 13358 7117 13364
rect 7731 13398 7789 13404
rect 7731 13364 7743 13398
rect 7777 13395 7789 13398
rect 8307 13398 8365 13404
rect 8307 13395 8319 13398
rect 7777 13367 8319 13395
rect 7777 13364 7789 13367
rect 7731 13358 7789 13364
rect 8307 13364 8319 13367
rect 8353 13364 8365 13398
rect 8307 13358 8365 13364
rect 8979 13398 9037 13404
rect 8979 13364 8991 13398
rect 9025 13395 9037 13398
rect 9555 13398 9613 13404
rect 9555 13395 9567 13398
rect 9025 13367 9567 13395
rect 9025 13364 9037 13367
rect 8979 13358 9037 13364
rect 9555 13364 9567 13367
rect 9601 13364 9613 13398
rect 9555 13358 9613 13364
rect 10227 13398 10285 13404
rect 10227 13364 10239 13398
rect 10273 13395 10285 13398
rect 10803 13398 10861 13404
rect 10803 13395 10815 13398
rect 10273 13367 10815 13395
rect 10273 13364 10285 13367
rect 10227 13358 10285 13364
rect 10803 13364 10815 13367
rect 10849 13364 10861 13398
rect 10803 13358 10861 13364
rect 11475 13398 11533 13404
rect 11475 13364 11487 13398
rect 11521 13395 11533 13398
rect 12051 13398 12109 13404
rect 12051 13395 12063 13398
rect 11521 13367 12063 13395
rect 11521 13364 11533 13367
rect 11475 13358 11533 13364
rect 12051 13364 12063 13367
rect 12097 13364 12109 13398
rect 12051 13358 12109 13364
rect 12723 13398 12781 13404
rect 12723 13364 12735 13398
rect 12769 13395 12781 13398
rect 13299 13398 13357 13404
rect 13299 13395 13311 13398
rect 12769 13367 13311 13395
rect 12769 13364 12781 13367
rect 12723 13358 12781 13364
rect 13299 13364 13311 13367
rect 13345 13364 13357 13398
rect 13299 13358 13357 13364
rect 13971 13398 14029 13404
rect 13971 13364 13983 13398
rect 14017 13395 14029 13398
rect 14547 13398 14605 13404
rect 14547 13395 14559 13398
rect 14017 13367 14559 13395
rect 14017 13364 14029 13367
rect 13971 13358 14029 13364
rect 14547 13364 14559 13367
rect 14593 13364 14605 13398
rect 14547 13358 14605 13364
rect 15219 13398 15277 13404
rect 15219 13364 15231 13398
rect 15265 13395 15277 13398
rect 15795 13398 15853 13404
rect 15795 13395 15807 13398
rect 15265 13367 15807 13395
rect 15265 13364 15277 13367
rect 15219 13358 15277 13364
rect 15795 13364 15807 13367
rect 15841 13364 15853 13398
rect 15795 13358 15853 13364
rect 16467 13398 16525 13404
rect 16467 13364 16479 13398
rect 16513 13395 16525 13398
rect 17043 13398 17101 13404
rect 17043 13395 17055 13398
rect 16513 13367 17055 13395
rect 16513 13364 16525 13367
rect 16467 13358 16525 13364
rect 17043 13364 17055 13367
rect 17089 13364 17101 13398
rect 17043 13358 17101 13364
rect 17715 13398 17773 13404
rect 17715 13364 17727 13398
rect 17761 13395 17773 13398
rect 18291 13398 18349 13404
rect 18291 13395 18303 13398
rect 17761 13367 18303 13395
rect 17761 13364 17773 13367
rect 17715 13358 17773 13364
rect 18291 13364 18303 13367
rect 18337 13364 18349 13398
rect 18291 13358 18349 13364
rect 18963 13398 19021 13404
rect 18963 13364 18975 13398
rect 19009 13395 19021 13398
rect 19539 13398 19597 13404
rect 19539 13395 19551 13398
rect 19009 13367 19551 13395
rect 19009 13364 19021 13367
rect 18963 13358 19021 13364
rect 19539 13364 19551 13367
rect 19585 13364 19597 13398
rect 19539 13358 19597 13364
rect 20211 13398 20269 13404
rect 20211 13364 20223 13398
rect 20257 13395 20269 13398
rect 20787 13398 20845 13404
rect 20787 13395 20799 13398
rect 20257 13367 20799 13395
rect 20257 13364 20269 13367
rect 20211 13358 20269 13364
rect 20787 13364 20799 13367
rect 20833 13364 20845 13398
rect 20787 13358 20845 13364
rect 21459 13398 21517 13404
rect 21459 13364 21471 13398
rect 21505 13395 21517 13398
rect 22035 13398 22093 13404
rect 22035 13395 22047 13398
rect 21505 13367 22047 13395
rect 21505 13364 21517 13367
rect 21459 13358 21517 13364
rect 22035 13364 22047 13367
rect 22081 13364 22093 13398
rect 22035 13358 22093 13364
rect 1952 13074 23264 13096
rect 1952 13022 7158 13074
rect 7210 13022 7222 13074
rect 7274 13022 7286 13074
rect 7338 13022 7350 13074
rect 7402 13022 12486 13074
rect 12538 13022 12550 13074
rect 12602 13022 12614 13074
rect 12666 13022 12678 13074
rect 12730 13022 17814 13074
rect 17866 13022 17878 13074
rect 17930 13022 17942 13074
rect 17994 13022 18006 13074
rect 18058 13022 23264 13074
rect 1952 13000 23264 13022
rect 3888 12911 3894 12963
rect 3946 12951 3952 12963
rect 3987 12954 4045 12960
rect 3987 12951 3999 12954
rect 3946 12923 3999 12951
rect 3946 12911 3952 12923
rect 3987 12920 3999 12923
rect 4033 12920 4045 12954
rect 3987 12914 4045 12920
rect 3411 12732 3469 12738
rect 3411 12698 3423 12732
rect 3457 12729 3469 12732
rect 5235 12732 5293 12738
rect 5235 12729 5247 12732
rect 3457 12701 5247 12729
rect 3457 12698 3469 12701
rect 3411 12692 3469 12698
rect 5235 12698 5247 12701
rect 5281 12698 5293 12732
rect 5235 12692 5293 12698
rect 5907 12732 5965 12738
rect 5907 12698 5919 12732
rect 5953 12729 5965 12732
rect 7731 12732 7789 12738
rect 7731 12729 7743 12732
rect 5953 12701 7743 12729
rect 5953 12698 5965 12701
rect 5907 12692 5965 12698
rect 7731 12698 7743 12701
rect 7777 12698 7789 12732
rect 7731 12692 7789 12698
rect 8403 12732 8461 12738
rect 8403 12698 8415 12732
rect 8449 12729 8461 12732
rect 10227 12732 10285 12738
rect 10227 12729 10239 12732
rect 8449 12701 10239 12729
rect 8449 12698 8461 12701
rect 8403 12692 8461 12698
rect 10227 12698 10239 12701
rect 10273 12698 10285 12732
rect 10227 12692 10285 12698
rect 12147 12732 12205 12738
rect 12147 12698 12159 12732
rect 12193 12729 12205 12732
rect 13971 12732 14029 12738
rect 13971 12729 13983 12732
rect 12193 12701 13983 12729
rect 12193 12698 12205 12701
rect 12147 12692 12205 12698
rect 13971 12698 13983 12701
rect 14017 12698 14029 12732
rect 13971 12692 14029 12698
rect 14547 12732 14605 12738
rect 14547 12698 14559 12732
rect 14593 12729 14605 12732
rect 16467 12732 16525 12738
rect 16467 12729 16479 12732
rect 14593 12701 16479 12729
rect 14593 12698 14605 12701
rect 14547 12692 14605 12698
rect 16467 12698 16479 12701
rect 16513 12698 16525 12732
rect 16467 12692 16525 12698
rect 17139 12732 17197 12738
rect 17139 12698 17151 12732
rect 17185 12729 17197 12732
rect 18963 12732 19021 12738
rect 18963 12729 18975 12732
rect 17185 12701 18975 12729
rect 17185 12698 17197 12701
rect 17139 12692 17197 12698
rect 18963 12698 18975 12701
rect 19009 12698 19021 12732
rect 18963 12692 19021 12698
rect 19635 12732 19693 12738
rect 19635 12698 19647 12732
rect 19681 12729 19693 12732
rect 21459 12732 21517 12738
rect 21459 12729 21471 12732
rect 19681 12701 21471 12729
rect 19681 12698 19693 12701
rect 19635 12692 19693 12698
rect 21459 12698 21471 12701
rect 21505 12698 21517 12732
rect 21459 12692 21517 12698
rect 4659 12658 4717 12664
rect 4659 12624 4671 12658
rect 4705 12624 4717 12658
rect 4659 12618 4717 12624
rect 7155 12658 7213 12664
rect 7155 12624 7167 12658
rect 7201 12655 7213 12658
rect 8979 12658 9037 12664
rect 8979 12655 8991 12658
rect 7201 12627 8991 12655
rect 7201 12624 7213 12627
rect 7155 12618 7213 12624
rect 8979 12624 8991 12627
rect 9025 12624 9037 12658
rect 8979 12618 9037 12624
rect 9555 12658 9613 12664
rect 9555 12624 9567 12658
rect 9601 12624 9613 12658
rect 9555 12618 9613 12624
rect 10899 12658 10957 12664
rect 10899 12624 10911 12658
rect 10945 12655 10957 12658
rect 12723 12658 12781 12664
rect 12723 12655 12735 12658
rect 10945 12627 12735 12655
rect 10945 12624 10957 12627
rect 10899 12618 10957 12624
rect 12723 12624 12735 12627
rect 12769 12624 12781 12658
rect 12723 12618 12781 12624
rect 13395 12658 13453 12664
rect 13395 12624 13407 12658
rect 13441 12655 13453 12658
rect 15219 12658 15277 12664
rect 15219 12655 15231 12658
rect 13441 12627 15231 12655
rect 13441 12624 13453 12627
rect 13395 12618 13453 12624
rect 15219 12624 15231 12627
rect 15265 12624 15277 12658
rect 15219 12618 15277 12624
rect 15891 12658 15949 12664
rect 15891 12624 15903 12658
rect 15937 12655 15949 12658
rect 17715 12658 17773 12664
rect 17715 12655 17727 12658
rect 15937 12627 17727 12655
rect 15937 12624 15949 12627
rect 15891 12618 15949 12624
rect 17715 12624 17727 12627
rect 17761 12624 17773 12658
rect 17715 12618 17773 12624
rect 18387 12658 18445 12664
rect 18387 12624 18399 12658
rect 18433 12655 18445 12658
rect 20211 12658 20269 12664
rect 20211 12655 20223 12658
rect 18433 12627 20223 12655
rect 18433 12624 18445 12627
rect 18387 12618 18445 12624
rect 20211 12624 20223 12627
rect 20257 12624 20269 12658
rect 20211 12618 20269 12624
rect 20883 12658 20941 12664
rect 20883 12624 20895 12658
rect 20929 12624 20941 12658
rect 22128 12655 22134 12667
rect 22089 12627 22134 12655
rect 20883 12618 20941 12624
rect 4674 12581 4702 12618
rect 6483 12584 6541 12590
rect 6483 12581 6495 12584
rect 4674 12553 6495 12581
rect 6483 12550 6495 12553
rect 6529 12550 6541 12584
rect 9570 12581 9598 12618
rect 11475 12584 11533 12590
rect 11475 12581 11487 12584
rect 9570 12553 11487 12581
rect 6483 12544 6541 12550
rect 11475 12550 11487 12553
rect 11521 12550 11533 12584
rect 20898 12581 20926 12618
rect 22128 12615 22134 12627
rect 22186 12615 22192 12667
rect 22707 12584 22765 12590
rect 22707 12581 22719 12584
rect 20898 12553 22719 12581
rect 11475 12544 11533 12550
rect 22707 12550 22719 12553
rect 22753 12550 22765 12584
rect 22707 12544 22765 12550
rect 1952 12408 23264 12430
rect 1952 12356 4494 12408
rect 4546 12356 4558 12408
rect 4610 12356 4622 12408
rect 4674 12356 4686 12408
rect 4738 12356 9822 12408
rect 9874 12356 9886 12408
rect 9938 12356 9950 12408
rect 10002 12356 10014 12408
rect 10066 12356 15150 12408
rect 15202 12356 15214 12408
rect 15266 12356 15278 12408
rect 15330 12356 15342 12408
rect 15394 12356 20478 12408
rect 20530 12356 20542 12408
rect 20594 12356 20606 12408
rect 20658 12356 20670 12408
rect 20722 12356 23264 12408
rect 1952 12334 23264 12356
rect 22128 12245 22134 12297
rect 22186 12285 22192 12297
rect 22707 12288 22765 12294
rect 22707 12285 22719 12288
rect 22186 12257 22719 12285
rect 22186 12245 22192 12257
rect 22707 12254 22719 12257
rect 22753 12254 22765 12288
rect 22707 12248 22765 12254
rect 2352 12097 2358 12149
rect 2410 12137 2416 12149
rect 3315 12140 3373 12146
rect 3315 12137 3327 12140
rect 2410 12109 3327 12137
rect 2410 12097 2416 12109
rect 3315 12106 3327 12109
rect 3361 12106 3373 12140
rect 3315 12100 3373 12106
rect 3987 12066 4045 12072
rect 3987 12032 3999 12066
rect 4033 12063 4045 12066
rect 4563 12066 4621 12072
rect 4563 12063 4575 12066
rect 4033 12035 4575 12063
rect 4033 12032 4045 12035
rect 3987 12026 4045 12032
rect 4563 12032 4575 12035
rect 4609 12032 4621 12066
rect 4563 12026 4621 12032
rect 5235 12066 5293 12072
rect 5235 12032 5247 12066
rect 5281 12063 5293 12066
rect 5811 12066 5869 12072
rect 5811 12063 5823 12066
rect 5281 12035 5823 12063
rect 5281 12032 5293 12035
rect 5235 12026 5293 12032
rect 5811 12032 5823 12035
rect 5857 12032 5869 12066
rect 5811 12026 5869 12032
rect 6483 12066 6541 12072
rect 6483 12032 6495 12066
rect 6529 12063 6541 12066
rect 7059 12066 7117 12072
rect 7059 12063 7071 12066
rect 6529 12035 7071 12063
rect 6529 12032 6541 12035
rect 6483 12026 6541 12032
rect 7059 12032 7071 12035
rect 7105 12032 7117 12066
rect 7059 12026 7117 12032
rect 7731 12066 7789 12072
rect 7731 12032 7743 12066
rect 7777 12063 7789 12066
rect 8307 12066 8365 12072
rect 8307 12063 8319 12066
rect 7777 12035 8319 12063
rect 7777 12032 7789 12035
rect 7731 12026 7789 12032
rect 8307 12032 8319 12035
rect 8353 12032 8365 12066
rect 8307 12026 8365 12032
rect 8979 12066 9037 12072
rect 8979 12032 8991 12066
rect 9025 12063 9037 12066
rect 9555 12066 9613 12072
rect 9555 12063 9567 12066
rect 9025 12035 9567 12063
rect 9025 12032 9037 12035
rect 8979 12026 9037 12032
rect 9555 12032 9567 12035
rect 9601 12032 9613 12066
rect 9555 12026 9613 12032
rect 10227 12066 10285 12072
rect 10227 12032 10239 12066
rect 10273 12063 10285 12066
rect 10803 12066 10861 12072
rect 10803 12063 10815 12066
rect 10273 12035 10815 12063
rect 10273 12032 10285 12035
rect 10227 12026 10285 12032
rect 10803 12032 10815 12035
rect 10849 12032 10861 12066
rect 10803 12026 10861 12032
rect 11475 12066 11533 12072
rect 11475 12032 11487 12066
rect 11521 12063 11533 12066
rect 12051 12066 12109 12072
rect 12051 12063 12063 12066
rect 11521 12035 12063 12063
rect 11521 12032 11533 12035
rect 11475 12026 11533 12032
rect 12051 12032 12063 12035
rect 12097 12032 12109 12066
rect 12051 12026 12109 12032
rect 12723 12066 12781 12072
rect 12723 12032 12735 12066
rect 12769 12063 12781 12066
rect 13299 12066 13357 12072
rect 13299 12063 13311 12066
rect 12769 12035 13311 12063
rect 12769 12032 12781 12035
rect 12723 12026 12781 12032
rect 13299 12032 13311 12035
rect 13345 12032 13357 12066
rect 13299 12026 13357 12032
rect 13971 12066 14029 12072
rect 13971 12032 13983 12066
rect 14017 12063 14029 12066
rect 14547 12066 14605 12072
rect 14547 12063 14559 12066
rect 14017 12035 14559 12063
rect 14017 12032 14029 12035
rect 13971 12026 14029 12032
rect 14547 12032 14559 12035
rect 14593 12032 14605 12066
rect 14547 12026 14605 12032
rect 15219 12066 15277 12072
rect 15219 12032 15231 12066
rect 15265 12063 15277 12066
rect 15795 12066 15853 12072
rect 15795 12063 15807 12066
rect 15265 12035 15807 12063
rect 15265 12032 15277 12035
rect 15219 12026 15277 12032
rect 15795 12032 15807 12035
rect 15841 12032 15853 12066
rect 15795 12026 15853 12032
rect 16467 12066 16525 12072
rect 16467 12032 16479 12066
rect 16513 12063 16525 12066
rect 17043 12066 17101 12072
rect 17043 12063 17055 12066
rect 16513 12035 17055 12063
rect 16513 12032 16525 12035
rect 16467 12026 16525 12032
rect 17043 12032 17055 12035
rect 17089 12032 17101 12066
rect 17043 12026 17101 12032
rect 17715 12066 17773 12072
rect 17715 12032 17727 12066
rect 17761 12063 17773 12066
rect 18291 12066 18349 12072
rect 18291 12063 18303 12066
rect 17761 12035 18303 12063
rect 17761 12032 17773 12035
rect 17715 12026 17773 12032
rect 18291 12032 18303 12035
rect 18337 12032 18349 12066
rect 18291 12026 18349 12032
rect 18963 12066 19021 12072
rect 18963 12032 18975 12066
rect 19009 12063 19021 12066
rect 19539 12066 19597 12072
rect 19539 12063 19551 12066
rect 19009 12035 19551 12063
rect 19009 12032 19021 12035
rect 18963 12026 19021 12032
rect 19539 12032 19551 12035
rect 19585 12032 19597 12066
rect 19539 12026 19597 12032
rect 20211 12066 20269 12072
rect 20211 12032 20223 12066
rect 20257 12063 20269 12066
rect 20787 12066 20845 12072
rect 20787 12063 20799 12066
rect 20257 12035 20799 12063
rect 20257 12032 20269 12035
rect 20211 12026 20269 12032
rect 20787 12032 20799 12035
rect 20833 12032 20845 12066
rect 20787 12026 20845 12032
rect 21459 12066 21517 12072
rect 21459 12032 21471 12066
rect 21505 12063 21517 12066
rect 22035 12066 22093 12072
rect 22035 12063 22047 12066
rect 21505 12035 22047 12063
rect 21505 12032 21517 12035
rect 21459 12026 21517 12032
rect 22035 12032 22047 12035
rect 22081 12032 22093 12066
rect 22035 12026 22093 12032
rect 1952 11742 23264 11764
rect 1952 11690 7158 11742
rect 7210 11690 7222 11742
rect 7274 11690 7286 11742
rect 7338 11690 7350 11742
rect 7402 11690 12486 11742
rect 12538 11690 12550 11742
rect 12602 11690 12614 11742
rect 12666 11690 12678 11742
rect 12730 11690 17814 11742
rect 17866 11690 17878 11742
rect 17930 11690 17942 11742
rect 17994 11690 18006 11742
rect 18058 11690 23264 11742
rect 1952 11668 23264 11690
rect 2352 11579 2358 11631
rect 2410 11619 2416 11631
rect 2739 11622 2797 11628
rect 2739 11619 2751 11622
rect 2410 11591 2751 11619
rect 2410 11579 2416 11591
rect 2739 11588 2751 11591
rect 2785 11588 2797 11622
rect 2739 11582 2797 11588
rect 21459 11474 21517 11480
rect 21459 11471 21471 11474
rect 20802 11443 21471 11471
rect 2064 11397 2070 11409
rect 2025 11369 2070 11397
rect 2064 11357 2070 11369
rect 2122 11357 2128 11409
rect 3987 11400 4045 11406
rect 3987 11397 3999 11400
rect 2466 11369 3999 11397
rect 2352 11323 2358 11335
rect 2313 11295 2358 11323
rect 2352 11283 2358 11295
rect 2410 11283 2416 11335
rect 2466 11332 2494 11369
rect 3987 11366 3999 11369
rect 4033 11366 4045 11400
rect 5235 11400 5293 11406
rect 5235 11397 5247 11400
rect 3987 11360 4045 11366
rect 4098 11369 5247 11397
rect 2451 11326 2509 11332
rect 2451 11292 2463 11326
rect 2497 11292 2509 11326
rect 2451 11286 2509 11292
rect 3411 11326 3469 11332
rect 3411 11292 3423 11326
rect 3457 11323 3469 11326
rect 4098 11323 4126 11369
rect 5235 11366 5247 11369
rect 5281 11366 5293 11400
rect 6483 11400 6541 11406
rect 6483 11397 6495 11400
rect 5235 11360 5293 11366
rect 5538 11369 6495 11397
rect 3457 11295 4126 11323
rect 4563 11326 4621 11332
rect 3457 11292 3469 11295
rect 3411 11286 3469 11292
rect 4563 11292 4575 11326
rect 4609 11323 4621 11326
rect 5538 11323 5566 11369
rect 6483 11366 6495 11369
rect 6529 11366 6541 11400
rect 7731 11400 7789 11406
rect 7731 11397 7743 11400
rect 6483 11360 6541 11366
rect 6594 11369 7743 11397
rect 4609 11295 5566 11323
rect 5907 11326 5965 11332
rect 4609 11292 4621 11295
rect 4563 11286 4621 11292
rect 5907 11292 5919 11326
rect 5953 11323 5965 11326
rect 6594 11323 6622 11369
rect 7731 11366 7743 11369
rect 7777 11366 7789 11400
rect 8979 11400 9037 11406
rect 8979 11397 8991 11400
rect 7731 11360 7789 11366
rect 8226 11369 8991 11397
rect 5953 11295 6622 11323
rect 7155 11326 7213 11332
rect 5953 11292 5965 11295
rect 5907 11286 5965 11292
rect 7155 11292 7167 11326
rect 7201 11323 7213 11326
rect 8226 11323 8254 11369
rect 8979 11366 8991 11369
rect 9025 11366 9037 11400
rect 8979 11360 9037 11366
rect 9651 11400 9709 11406
rect 9651 11366 9663 11400
rect 9697 11397 9709 11400
rect 11475 11400 11533 11406
rect 11475 11397 11487 11400
rect 9697 11369 11487 11397
rect 9697 11366 9709 11369
rect 9651 11360 9709 11366
rect 11475 11366 11487 11369
rect 11521 11366 11533 11400
rect 11475 11360 11533 11366
rect 12147 11400 12205 11406
rect 12147 11366 12159 11400
rect 12193 11397 12205 11400
rect 13971 11400 14029 11406
rect 13971 11397 13983 11400
rect 12193 11369 13983 11397
rect 12193 11366 12205 11369
rect 12147 11360 12205 11366
rect 13971 11366 13983 11369
rect 14017 11366 14029 11400
rect 13971 11360 14029 11366
rect 14547 11400 14605 11406
rect 14547 11366 14559 11400
rect 14593 11397 14605 11400
rect 16467 11400 16525 11406
rect 16467 11397 16479 11400
rect 14593 11369 16479 11397
rect 14593 11366 14605 11369
rect 14547 11360 14605 11366
rect 16467 11366 16479 11369
rect 16513 11366 16525 11400
rect 17715 11400 17773 11406
rect 17715 11397 17727 11400
rect 16467 11360 16525 11366
rect 16770 11369 17727 11397
rect 7201 11295 8254 11323
rect 8403 11326 8461 11332
rect 7201 11292 7213 11295
rect 7155 11286 7213 11292
rect 8403 11292 8415 11326
rect 8449 11323 8461 11326
rect 10227 11326 10285 11332
rect 10227 11323 10239 11326
rect 8449 11295 10239 11323
rect 8449 11292 8461 11295
rect 8403 11286 8461 11292
rect 10227 11292 10239 11295
rect 10273 11292 10285 11326
rect 10227 11286 10285 11292
rect 10899 11326 10957 11332
rect 10899 11292 10911 11326
rect 10945 11323 10957 11326
rect 12723 11326 12781 11332
rect 12723 11323 12735 11326
rect 10945 11295 12735 11323
rect 10945 11292 10957 11295
rect 10899 11286 10957 11292
rect 12723 11292 12735 11295
rect 12769 11292 12781 11326
rect 12723 11286 12781 11292
rect 13395 11326 13453 11332
rect 13395 11292 13407 11326
rect 13441 11323 13453 11326
rect 15219 11326 15277 11332
rect 15219 11323 15231 11326
rect 13441 11295 15231 11323
rect 13441 11292 13453 11295
rect 13395 11286 13453 11292
rect 15219 11292 15231 11295
rect 15265 11292 15277 11326
rect 15219 11286 15277 11292
rect 15891 11326 15949 11332
rect 15891 11292 15903 11326
rect 15937 11323 15949 11326
rect 16770 11323 16798 11369
rect 17715 11366 17727 11369
rect 17761 11366 17773 11400
rect 17715 11360 17773 11366
rect 18387 11400 18445 11406
rect 18387 11366 18399 11400
rect 18433 11397 18445 11400
rect 20211 11400 20269 11406
rect 20211 11397 20223 11400
rect 18433 11369 20223 11397
rect 18433 11366 18445 11369
rect 18387 11360 18445 11366
rect 20211 11366 20223 11369
rect 20257 11366 20269 11400
rect 20211 11360 20269 11366
rect 15937 11295 16798 11323
rect 17139 11326 17197 11332
rect 15937 11292 15949 11295
rect 15891 11286 15949 11292
rect 17139 11292 17151 11326
rect 17185 11323 17197 11326
rect 18963 11326 19021 11332
rect 18963 11323 18975 11326
rect 17185 11295 18975 11323
rect 17185 11292 17197 11295
rect 17139 11286 17197 11292
rect 18963 11292 18975 11295
rect 19009 11292 19021 11326
rect 18963 11286 19021 11292
rect 19635 11326 19693 11332
rect 19635 11292 19647 11326
rect 19681 11323 19693 11326
rect 20802 11323 20830 11443
rect 21459 11440 21471 11443
rect 21505 11440 21517 11474
rect 21459 11434 21517 11440
rect 22707 11400 22765 11406
rect 22707 11397 22719 11400
rect 21762 11369 22719 11397
rect 19681 11295 20830 11323
rect 20883 11326 20941 11332
rect 19681 11292 19693 11295
rect 19635 11286 19693 11292
rect 20883 11292 20895 11326
rect 20929 11323 20941 11326
rect 21762 11323 21790 11369
rect 22707 11366 22719 11369
rect 22753 11366 22765 11400
rect 22707 11360 22765 11366
rect 20929 11295 21790 11323
rect 22131 11326 22189 11332
rect 20929 11292 20941 11295
rect 20883 11286 20941 11292
rect 22131 11292 22143 11326
rect 22177 11323 22189 11326
rect 22608 11323 22614 11335
rect 22177 11295 22614 11323
rect 22177 11292 22189 11295
rect 22131 11286 22189 11292
rect 22608 11283 22614 11295
rect 22666 11283 22672 11335
rect 1952 11076 23264 11098
rect 1952 11024 4494 11076
rect 4546 11024 4558 11076
rect 4610 11024 4622 11076
rect 4674 11024 4686 11076
rect 4738 11024 9822 11076
rect 9874 11024 9886 11076
rect 9938 11024 9950 11076
rect 10002 11024 10014 11076
rect 10066 11024 15150 11076
rect 15202 11024 15214 11076
rect 15266 11024 15278 11076
rect 15330 11024 15342 11076
rect 15394 11024 20478 11076
rect 20530 11024 20542 11076
rect 20594 11024 20606 11076
rect 20658 11024 20670 11076
rect 20722 11024 23264 11076
rect 1952 11002 23264 11024
rect 22608 10913 22614 10965
rect 22666 10953 22672 10965
rect 22707 10956 22765 10962
rect 22707 10953 22719 10956
rect 22666 10925 22719 10953
rect 22666 10913 22672 10925
rect 22707 10922 22719 10925
rect 22753 10922 22765 10956
rect 22707 10916 22765 10922
rect 3411 10734 3469 10740
rect 3411 10700 3423 10734
rect 3457 10731 3469 10734
rect 3888 10731 3894 10743
rect 3457 10703 3894 10731
rect 3457 10700 3469 10703
rect 3411 10694 3469 10700
rect 3888 10691 3894 10703
rect 3946 10691 3952 10743
rect 3987 10734 4045 10740
rect 3987 10700 3999 10734
rect 4033 10731 4045 10734
rect 4563 10734 4621 10740
rect 4563 10731 4575 10734
rect 4033 10703 4575 10731
rect 4033 10700 4045 10703
rect 3987 10694 4045 10700
rect 4563 10700 4575 10703
rect 4609 10700 4621 10734
rect 4563 10694 4621 10700
rect 5235 10734 5293 10740
rect 5235 10700 5247 10734
rect 5281 10731 5293 10734
rect 5811 10734 5869 10740
rect 5811 10731 5823 10734
rect 5281 10703 5823 10731
rect 5281 10700 5293 10703
rect 5235 10694 5293 10700
rect 5811 10700 5823 10703
rect 5857 10700 5869 10734
rect 5811 10694 5869 10700
rect 6483 10734 6541 10740
rect 6483 10700 6495 10734
rect 6529 10731 6541 10734
rect 7059 10734 7117 10740
rect 7059 10731 7071 10734
rect 6529 10703 7071 10731
rect 6529 10700 6541 10703
rect 6483 10694 6541 10700
rect 7059 10700 7071 10703
rect 7105 10700 7117 10734
rect 7059 10694 7117 10700
rect 7731 10734 7789 10740
rect 7731 10700 7743 10734
rect 7777 10731 7789 10734
rect 8307 10734 8365 10740
rect 8307 10731 8319 10734
rect 7777 10703 8319 10731
rect 7777 10700 7789 10703
rect 7731 10694 7789 10700
rect 8307 10700 8319 10703
rect 8353 10700 8365 10734
rect 8307 10694 8365 10700
rect 8979 10734 9037 10740
rect 8979 10700 8991 10734
rect 9025 10731 9037 10734
rect 9555 10734 9613 10740
rect 9555 10731 9567 10734
rect 9025 10703 9567 10731
rect 9025 10700 9037 10703
rect 8979 10694 9037 10700
rect 9555 10700 9567 10703
rect 9601 10700 9613 10734
rect 9555 10694 9613 10700
rect 10227 10734 10285 10740
rect 10227 10700 10239 10734
rect 10273 10731 10285 10734
rect 10803 10734 10861 10740
rect 10803 10731 10815 10734
rect 10273 10703 10815 10731
rect 10273 10700 10285 10703
rect 10227 10694 10285 10700
rect 10803 10700 10815 10703
rect 10849 10700 10861 10734
rect 10803 10694 10861 10700
rect 11475 10734 11533 10740
rect 11475 10700 11487 10734
rect 11521 10731 11533 10734
rect 12051 10734 12109 10740
rect 12051 10731 12063 10734
rect 11521 10703 12063 10731
rect 11521 10700 11533 10703
rect 11475 10694 11533 10700
rect 12051 10700 12063 10703
rect 12097 10700 12109 10734
rect 12051 10694 12109 10700
rect 12723 10734 12781 10740
rect 12723 10700 12735 10734
rect 12769 10731 12781 10734
rect 13299 10734 13357 10740
rect 13299 10731 13311 10734
rect 12769 10703 13311 10731
rect 12769 10700 12781 10703
rect 12723 10694 12781 10700
rect 13299 10700 13311 10703
rect 13345 10700 13357 10734
rect 13299 10694 13357 10700
rect 13971 10734 14029 10740
rect 13971 10700 13983 10734
rect 14017 10731 14029 10734
rect 14547 10734 14605 10740
rect 14547 10731 14559 10734
rect 14017 10703 14559 10731
rect 14017 10700 14029 10703
rect 13971 10694 14029 10700
rect 14547 10700 14559 10703
rect 14593 10700 14605 10734
rect 14547 10694 14605 10700
rect 15219 10734 15277 10740
rect 15219 10700 15231 10734
rect 15265 10731 15277 10734
rect 15795 10734 15853 10740
rect 15795 10731 15807 10734
rect 15265 10703 15807 10731
rect 15265 10700 15277 10703
rect 15219 10694 15277 10700
rect 15795 10700 15807 10703
rect 15841 10700 15853 10734
rect 15795 10694 15853 10700
rect 16467 10734 16525 10740
rect 16467 10700 16479 10734
rect 16513 10731 16525 10734
rect 17043 10734 17101 10740
rect 17043 10731 17055 10734
rect 16513 10703 17055 10731
rect 16513 10700 16525 10703
rect 16467 10694 16525 10700
rect 17043 10700 17055 10703
rect 17089 10700 17101 10734
rect 17043 10694 17101 10700
rect 17715 10734 17773 10740
rect 17715 10700 17727 10734
rect 17761 10731 17773 10734
rect 18291 10734 18349 10740
rect 18291 10731 18303 10734
rect 17761 10703 18303 10731
rect 17761 10700 17773 10703
rect 17715 10694 17773 10700
rect 18291 10700 18303 10703
rect 18337 10700 18349 10734
rect 18291 10694 18349 10700
rect 18963 10734 19021 10740
rect 18963 10700 18975 10734
rect 19009 10731 19021 10734
rect 19539 10734 19597 10740
rect 19539 10731 19551 10734
rect 19009 10703 19551 10731
rect 19009 10700 19021 10703
rect 18963 10694 19021 10700
rect 19539 10700 19551 10703
rect 19585 10700 19597 10734
rect 19539 10694 19597 10700
rect 20211 10734 20269 10740
rect 20211 10700 20223 10734
rect 20257 10731 20269 10734
rect 20787 10734 20845 10740
rect 20787 10731 20799 10734
rect 20257 10703 20799 10731
rect 20257 10700 20269 10703
rect 20211 10694 20269 10700
rect 20787 10700 20799 10703
rect 20833 10700 20845 10734
rect 20787 10694 20845 10700
rect 21459 10734 21517 10740
rect 21459 10700 21471 10734
rect 21505 10731 21517 10734
rect 22035 10734 22093 10740
rect 22035 10731 22047 10734
rect 21505 10703 22047 10731
rect 21505 10700 21517 10703
rect 21459 10694 21517 10700
rect 22035 10700 22047 10703
rect 22081 10700 22093 10734
rect 22035 10694 22093 10700
rect 1952 10410 23264 10432
rect 1952 10358 7158 10410
rect 7210 10358 7222 10410
rect 7274 10358 7286 10410
rect 7338 10358 7350 10410
rect 7402 10358 12486 10410
rect 12538 10358 12550 10410
rect 12602 10358 12614 10410
rect 12666 10358 12678 10410
rect 12730 10358 17814 10410
rect 17866 10358 17878 10410
rect 17930 10358 17942 10410
rect 17994 10358 18006 10410
rect 18058 10358 23264 10410
rect 1952 10336 23264 10358
rect 3888 10247 3894 10299
rect 3946 10287 3952 10299
rect 3987 10290 4045 10296
rect 3987 10287 3999 10290
rect 3946 10259 3999 10287
rect 3946 10247 3952 10259
rect 3987 10256 3999 10259
rect 4033 10256 4045 10290
rect 3987 10250 4045 10256
rect 4659 10068 4717 10074
rect 4659 10034 4671 10068
rect 4705 10065 4717 10068
rect 6483 10068 6541 10074
rect 6483 10065 6495 10068
rect 4705 10037 6495 10065
rect 4705 10034 4717 10037
rect 4659 10028 4717 10034
rect 6483 10034 6495 10037
rect 6529 10034 6541 10068
rect 8979 10068 9037 10074
rect 8979 10065 8991 10068
rect 6483 10028 6541 10034
rect 8322 10037 8991 10065
rect 3411 9994 3469 10000
rect 3411 9960 3423 9994
rect 3457 9991 3469 9994
rect 5235 9994 5293 10000
rect 5235 9991 5247 9994
rect 3457 9963 5247 9991
rect 3457 9960 3469 9963
rect 3411 9954 3469 9960
rect 5235 9960 5247 9963
rect 5281 9960 5293 9994
rect 5235 9954 5293 9960
rect 5907 9994 5965 10000
rect 5907 9960 5919 9994
rect 5953 9960 5965 9994
rect 5907 9954 5965 9960
rect 7155 9994 7213 10000
rect 7155 9960 7167 9994
rect 7201 9991 7213 9994
rect 8322 9991 8350 10037
rect 8979 10034 8991 10037
rect 9025 10034 9037 10068
rect 8979 10028 9037 10034
rect 9651 10068 9709 10074
rect 9651 10034 9663 10068
rect 9697 10065 9709 10068
rect 11475 10068 11533 10074
rect 11475 10065 11487 10068
rect 9697 10037 11487 10065
rect 9697 10034 9709 10037
rect 9651 10028 9709 10034
rect 11475 10034 11487 10037
rect 11521 10034 11533 10068
rect 11475 10028 11533 10034
rect 12147 10068 12205 10074
rect 12147 10034 12159 10068
rect 12193 10065 12205 10068
rect 13971 10068 14029 10074
rect 13971 10065 13983 10068
rect 12193 10037 13983 10065
rect 12193 10034 12205 10037
rect 12147 10028 12205 10034
rect 13971 10034 13983 10037
rect 14017 10034 14029 10068
rect 13971 10028 14029 10034
rect 14547 10068 14605 10074
rect 14547 10034 14559 10068
rect 14593 10065 14605 10068
rect 16467 10068 16525 10074
rect 16467 10065 16479 10068
rect 14593 10037 16479 10065
rect 14593 10034 14605 10037
rect 14547 10028 14605 10034
rect 16467 10034 16479 10037
rect 16513 10034 16525 10068
rect 16467 10028 16525 10034
rect 17139 10068 17197 10074
rect 17139 10034 17151 10068
rect 17185 10065 17197 10068
rect 18963 10068 19021 10074
rect 18963 10065 18975 10068
rect 17185 10037 18975 10065
rect 17185 10034 17197 10037
rect 17139 10028 17197 10034
rect 18963 10034 18975 10037
rect 19009 10034 19021 10068
rect 18963 10028 19021 10034
rect 19635 10068 19693 10074
rect 19635 10034 19647 10068
rect 19681 10065 19693 10068
rect 21459 10068 21517 10074
rect 21459 10065 21471 10068
rect 19681 10037 21471 10065
rect 19681 10034 19693 10037
rect 19635 10028 19693 10034
rect 21459 10034 21471 10037
rect 21505 10034 21517 10068
rect 21459 10028 21517 10034
rect 7201 9963 8350 9991
rect 8403 9994 8461 10000
rect 7201 9960 7213 9963
rect 7155 9954 7213 9960
rect 8403 9960 8415 9994
rect 8449 9991 8461 9994
rect 10227 9994 10285 10000
rect 10227 9991 10239 9994
rect 8449 9963 10239 9991
rect 8449 9960 8461 9963
rect 8403 9954 8461 9960
rect 10227 9960 10239 9963
rect 10273 9960 10285 9994
rect 10227 9954 10285 9960
rect 10899 9994 10957 10000
rect 10899 9960 10911 9994
rect 10945 9991 10957 9994
rect 12723 9994 12781 10000
rect 12723 9991 12735 9994
rect 10945 9963 12735 9991
rect 10945 9960 10957 9963
rect 10899 9954 10957 9960
rect 12723 9960 12735 9963
rect 12769 9960 12781 9994
rect 12723 9954 12781 9960
rect 13395 9994 13453 10000
rect 13395 9960 13407 9994
rect 13441 9991 13453 9994
rect 15219 9994 15277 10000
rect 15219 9991 15231 9994
rect 13441 9963 15231 9991
rect 13441 9960 13453 9963
rect 13395 9954 13453 9960
rect 15219 9960 15231 9963
rect 15265 9960 15277 9994
rect 15219 9954 15277 9960
rect 15891 9994 15949 10000
rect 15891 9960 15903 9994
rect 15937 9991 15949 9994
rect 17715 9994 17773 10000
rect 17715 9991 17727 9994
rect 15937 9963 17727 9991
rect 15937 9960 15949 9963
rect 15891 9954 15949 9960
rect 17715 9960 17727 9963
rect 17761 9960 17773 9994
rect 17715 9954 17773 9960
rect 18387 9994 18445 10000
rect 18387 9960 18399 9994
rect 18433 9991 18445 9994
rect 20211 9994 20269 10000
rect 20211 9991 20223 9994
rect 18433 9963 20223 9991
rect 18433 9960 18445 9963
rect 18387 9954 18445 9960
rect 20211 9960 20223 9963
rect 20257 9960 20269 9994
rect 20211 9954 20269 9960
rect 20883 9994 20941 10000
rect 20883 9960 20895 9994
rect 20929 9960 20941 9994
rect 20883 9954 20941 9960
rect 22131 9994 22189 10000
rect 22131 9960 22143 9994
rect 22177 9991 22189 9994
rect 22608 9991 22614 10003
rect 22177 9963 22614 9991
rect 22177 9960 22189 9963
rect 22131 9954 22189 9960
rect 5922 9917 5950 9954
rect 7731 9920 7789 9926
rect 7731 9917 7743 9920
rect 5922 9889 7743 9917
rect 7731 9886 7743 9889
rect 7777 9886 7789 9920
rect 20898 9917 20926 9954
rect 22608 9951 22614 9963
rect 22666 9951 22672 10003
rect 22707 9920 22765 9926
rect 22707 9917 22719 9920
rect 20898 9889 22719 9917
rect 7731 9880 7789 9886
rect 22707 9886 22719 9889
rect 22753 9886 22765 9920
rect 22707 9880 22765 9886
rect 1952 9744 23264 9766
rect 1952 9692 4494 9744
rect 4546 9692 4558 9744
rect 4610 9692 4622 9744
rect 4674 9692 4686 9744
rect 4738 9692 9822 9744
rect 9874 9692 9886 9744
rect 9938 9692 9950 9744
rect 10002 9692 10014 9744
rect 10066 9692 15150 9744
rect 15202 9692 15214 9744
rect 15266 9692 15278 9744
rect 15330 9692 15342 9744
rect 15394 9692 20478 9744
rect 20530 9692 20542 9744
rect 20594 9692 20606 9744
rect 20658 9692 20670 9744
rect 20722 9692 23264 9744
rect 1952 9670 23264 9692
rect 22608 9581 22614 9633
rect 22666 9621 22672 9633
rect 22707 9624 22765 9630
rect 22707 9621 22719 9624
rect 22666 9593 22719 9621
rect 22666 9581 22672 9593
rect 22707 9590 22719 9593
rect 22753 9590 22765 9624
rect 22707 9584 22765 9590
rect 3411 9402 3469 9408
rect 3411 9368 3423 9402
rect 3457 9399 3469 9402
rect 3888 9399 3894 9411
rect 3457 9371 3894 9399
rect 3457 9368 3469 9371
rect 3411 9362 3469 9368
rect 3888 9359 3894 9371
rect 3946 9359 3952 9411
rect 3987 9402 4045 9408
rect 3987 9368 3999 9402
rect 4033 9399 4045 9402
rect 4563 9402 4621 9408
rect 4563 9399 4575 9402
rect 4033 9371 4575 9399
rect 4033 9368 4045 9371
rect 3987 9362 4045 9368
rect 4563 9368 4575 9371
rect 4609 9368 4621 9402
rect 4563 9362 4621 9368
rect 5235 9402 5293 9408
rect 5235 9368 5247 9402
rect 5281 9399 5293 9402
rect 5811 9402 5869 9408
rect 5811 9399 5823 9402
rect 5281 9371 5823 9399
rect 5281 9368 5293 9371
rect 5235 9362 5293 9368
rect 5811 9368 5823 9371
rect 5857 9368 5869 9402
rect 5811 9362 5869 9368
rect 6483 9402 6541 9408
rect 6483 9368 6495 9402
rect 6529 9399 6541 9402
rect 7059 9402 7117 9408
rect 7059 9399 7071 9402
rect 6529 9371 7071 9399
rect 6529 9368 6541 9371
rect 6483 9362 6541 9368
rect 7059 9368 7071 9371
rect 7105 9368 7117 9402
rect 7059 9362 7117 9368
rect 7731 9402 7789 9408
rect 7731 9368 7743 9402
rect 7777 9399 7789 9402
rect 8307 9402 8365 9408
rect 8307 9399 8319 9402
rect 7777 9371 8319 9399
rect 7777 9368 7789 9371
rect 7731 9362 7789 9368
rect 8307 9368 8319 9371
rect 8353 9368 8365 9402
rect 8307 9362 8365 9368
rect 8979 9402 9037 9408
rect 8979 9368 8991 9402
rect 9025 9399 9037 9402
rect 9555 9402 9613 9408
rect 9555 9399 9567 9402
rect 9025 9371 9567 9399
rect 9025 9368 9037 9371
rect 8979 9362 9037 9368
rect 9555 9368 9567 9371
rect 9601 9368 9613 9402
rect 9555 9362 9613 9368
rect 10227 9402 10285 9408
rect 10227 9368 10239 9402
rect 10273 9399 10285 9402
rect 10803 9402 10861 9408
rect 10803 9399 10815 9402
rect 10273 9371 10815 9399
rect 10273 9368 10285 9371
rect 10227 9362 10285 9368
rect 10803 9368 10815 9371
rect 10849 9368 10861 9402
rect 10803 9362 10861 9368
rect 11475 9402 11533 9408
rect 11475 9368 11487 9402
rect 11521 9399 11533 9402
rect 12051 9402 12109 9408
rect 12051 9399 12063 9402
rect 11521 9371 12063 9399
rect 11521 9368 11533 9371
rect 11475 9362 11533 9368
rect 12051 9368 12063 9371
rect 12097 9368 12109 9402
rect 12051 9362 12109 9368
rect 12723 9402 12781 9408
rect 12723 9368 12735 9402
rect 12769 9399 12781 9402
rect 13299 9402 13357 9408
rect 13299 9399 13311 9402
rect 12769 9371 13311 9399
rect 12769 9368 12781 9371
rect 12723 9362 12781 9368
rect 13299 9368 13311 9371
rect 13345 9368 13357 9402
rect 13299 9362 13357 9368
rect 13971 9402 14029 9408
rect 13971 9368 13983 9402
rect 14017 9399 14029 9402
rect 14547 9402 14605 9408
rect 14547 9399 14559 9402
rect 14017 9371 14559 9399
rect 14017 9368 14029 9371
rect 13971 9362 14029 9368
rect 14547 9368 14559 9371
rect 14593 9368 14605 9402
rect 14547 9362 14605 9368
rect 15219 9402 15277 9408
rect 15219 9368 15231 9402
rect 15265 9399 15277 9402
rect 15795 9402 15853 9408
rect 15795 9399 15807 9402
rect 15265 9371 15807 9399
rect 15265 9368 15277 9371
rect 15219 9362 15277 9368
rect 15795 9368 15807 9371
rect 15841 9368 15853 9402
rect 15795 9362 15853 9368
rect 16467 9402 16525 9408
rect 16467 9368 16479 9402
rect 16513 9399 16525 9402
rect 17043 9402 17101 9408
rect 17043 9399 17055 9402
rect 16513 9371 17055 9399
rect 16513 9368 16525 9371
rect 16467 9362 16525 9368
rect 17043 9368 17055 9371
rect 17089 9368 17101 9402
rect 17043 9362 17101 9368
rect 17715 9402 17773 9408
rect 17715 9368 17727 9402
rect 17761 9399 17773 9402
rect 18291 9402 18349 9408
rect 18291 9399 18303 9402
rect 17761 9371 18303 9399
rect 17761 9368 17773 9371
rect 17715 9362 17773 9368
rect 18291 9368 18303 9371
rect 18337 9368 18349 9402
rect 18291 9362 18349 9368
rect 18963 9402 19021 9408
rect 18963 9368 18975 9402
rect 19009 9399 19021 9402
rect 19539 9402 19597 9408
rect 19539 9399 19551 9402
rect 19009 9371 19551 9399
rect 19009 9368 19021 9371
rect 18963 9362 19021 9368
rect 19539 9368 19551 9371
rect 19585 9368 19597 9402
rect 19539 9362 19597 9368
rect 20211 9402 20269 9408
rect 20211 9368 20223 9402
rect 20257 9399 20269 9402
rect 20787 9402 20845 9408
rect 20787 9399 20799 9402
rect 20257 9371 20799 9399
rect 20257 9368 20269 9371
rect 20211 9362 20269 9368
rect 20787 9368 20799 9371
rect 20833 9368 20845 9402
rect 20787 9362 20845 9368
rect 21459 9402 21517 9408
rect 21459 9368 21471 9402
rect 21505 9399 21517 9402
rect 22035 9402 22093 9408
rect 22035 9399 22047 9402
rect 21505 9371 22047 9399
rect 21505 9368 21517 9371
rect 21459 9362 21517 9368
rect 22035 9368 22047 9371
rect 22081 9368 22093 9402
rect 22035 9362 22093 9368
rect 1952 9078 23264 9100
rect 1952 9026 7158 9078
rect 7210 9026 7222 9078
rect 7274 9026 7286 9078
rect 7338 9026 7350 9078
rect 7402 9026 12486 9078
rect 12538 9026 12550 9078
rect 12602 9026 12614 9078
rect 12666 9026 12678 9078
rect 12730 9026 17814 9078
rect 17866 9026 17878 9078
rect 17930 9026 17942 9078
rect 17994 9026 18006 9078
rect 18058 9026 23264 9078
rect 1952 9004 23264 9026
rect 3888 8915 3894 8967
rect 3946 8955 3952 8967
rect 3987 8958 4045 8964
rect 3987 8955 3999 8958
rect 3946 8927 3999 8955
rect 3946 8915 3952 8927
rect 3987 8924 3999 8927
rect 4033 8924 4045 8958
rect 3987 8918 4045 8924
rect 3411 8736 3469 8742
rect 3411 8702 3423 8736
rect 3457 8733 3469 8736
rect 5235 8736 5293 8742
rect 5235 8733 5247 8736
rect 3457 8705 5247 8733
rect 3457 8702 3469 8705
rect 3411 8696 3469 8702
rect 5235 8702 5247 8705
rect 5281 8702 5293 8736
rect 5235 8696 5293 8702
rect 5907 8736 5965 8742
rect 5907 8702 5919 8736
rect 5953 8733 5965 8736
rect 7731 8736 7789 8742
rect 7731 8733 7743 8736
rect 5953 8705 7743 8733
rect 5953 8702 5965 8705
rect 5907 8696 5965 8702
rect 7731 8702 7743 8705
rect 7777 8702 7789 8736
rect 8979 8736 9037 8742
rect 8979 8733 8991 8736
rect 7731 8696 7789 8702
rect 8322 8705 8991 8733
rect 4659 8662 4717 8668
rect 4659 8628 4671 8662
rect 4705 8628 4717 8662
rect 4659 8622 4717 8628
rect 7155 8662 7213 8668
rect 7155 8628 7167 8662
rect 7201 8659 7213 8662
rect 8322 8659 8350 8705
rect 8979 8702 8991 8705
rect 9025 8702 9037 8736
rect 8979 8696 9037 8702
rect 9651 8736 9709 8742
rect 9651 8702 9663 8736
rect 9697 8733 9709 8736
rect 11475 8736 11533 8742
rect 11475 8733 11487 8736
rect 9697 8705 11487 8733
rect 9697 8702 9709 8705
rect 9651 8696 9709 8702
rect 11475 8702 11487 8705
rect 11521 8702 11533 8736
rect 11475 8696 11533 8702
rect 12147 8736 12205 8742
rect 12147 8702 12159 8736
rect 12193 8733 12205 8736
rect 13971 8736 14029 8742
rect 13971 8733 13983 8736
rect 12193 8705 13983 8733
rect 12193 8702 12205 8705
rect 12147 8696 12205 8702
rect 13971 8702 13983 8705
rect 14017 8702 14029 8736
rect 13971 8696 14029 8702
rect 14547 8736 14605 8742
rect 14547 8702 14559 8736
rect 14593 8733 14605 8736
rect 16467 8736 16525 8742
rect 16467 8733 16479 8736
rect 14593 8705 16479 8733
rect 14593 8702 14605 8705
rect 14547 8696 14605 8702
rect 16467 8702 16479 8705
rect 16513 8702 16525 8736
rect 16467 8696 16525 8702
rect 17139 8736 17197 8742
rect 17139 8702 17151 8736
rect 17185 8733 17197 8736
rect 18963 8736 19021 8742
rect 18963 8733 18975 8736
rect 17185 8705 18975 8733
rect 17185 8702 17197 8705
rect 17139 8696 17197 8702
rect 18963 8702 18975 8705
rect 19009 8702 19021 8736
rect 18963 8696 19021 8702
rect 19635 8736 19693 8742
rect 19635 8702 19647 8736
rect 19681 8733 19693 8736
rect 21459 8736 21517 8742
rect 21459 8733 21471 8736
rect 19681 8705 21471 8733
rect 19681 8702 19693 8705
rect 19635 8696 19693 8702
rect 21459 8702 21471 8705
rect 21505 8702 21517 8736
rect 21459 8696 21517 8702
rect 7201 8631 8350 8659
rect 8403 8662 8461 8668
rect 7201 8628 7213 8631
rect 7155 8622 7213 8628
rect 8403 8628 8415 8662
rect 8449 8659 8461 8662
rect 10227 8662 10285 8668
rect 10227 8659 10239 8662
rect 8449 8631 10239 8659
rect 8449 8628 8461 8631
rect 8403 8622 8461 8628
rect 10227 8628 10239 8631
rect 10273 8628 10285 8662
rect 10227 8622 10285 8628
rect 10899 8662 10957 8668
rect 10899 8628 10911 8662
rect 10945 8659 10957 8662
rect 12723 8662 12781 8668
rect 12723 8659 12735 8662
rect 10945 8631 12735 8659
rect 10945 8628 10957 8631
rect 10899 8622 10957 8628
rect 12723 8628 12735 8631
rect 12769 8628 12781 8662
rect 12723 8622 12781 8628
rect 13395 8662 13453 8668
rect 13395 8628 13407 8662
rect 13441 8659 13453 8662
rect 15219 8662 15277 8668
rect 15219 8659 15231 8662
rect 13441 8631 15231 8659
rect 13441 8628 13453 8631
rect 13395 8622 13453 8628
rect 15219 8628 15231 8631
rect 15265 8628 15277 8662
rect 15219 8622 15277 8628
rect 15891 8662 15949 8668
rect 15891 8628 15903 8662
rect 15937 8659 15949 8662
rect 17715 8662 17773 8668
rect 17715 8659 17727 8662
rect 15937 8631 17727 8659
rect 15937 8628 15949 8631
rect 15891 8622 15949 8628
rect 17715 8628 17727 8631
rect 17761 8628 17773 8662
rect 17715 8622 17773 8628
rect 18387 8662 18445 8668
rect 18387 8628 18399 8662
rect 18433 8659 18445 8662
rect 20211 8662 20269 8668
rect 20211 8659 20223 8662
rect 18433 8631 20223 8659
rect 18433 8628 18445 8631
rect 18387 8622 18445 8628
rect 20211 8628 20223 8631
rect 20257 8628 20269 8662
rect 20211 8622 20269 8628
rect 20883 8662 20941 8668
rect 20883 8628 20895 8662
rect 20929 8628 20941 8662
rect 20883 8622 20941 8628
rect 22131 8662 22189 8668
rect 22131 8628 22143 8662
rect 22177 8659 22189 8662
rect 22608 8659 22614 8671
rect 22177 8631 22614 8659
rect 22177 8628 22189 8631
rect 22131 8622 22189 8628
rect 4674 8585 4702 8622
rect 6483 8588 6541 8594
rect 6483 8585 6495 8588
rect 4674 8557 6495 8585
rect 6483 8554 6495 8557
rect 6529 8554 6541 8588
rect 20898 8585 20926 8622
rect 22608 8619 22614 8631
rect 22666 8619 22672 8671
rect 22707 8588 22765 8594
rect 22707 8585 22719 8588
rect 20898 8557 22719 8585
rect 6483 8548 6541 8554
rect 22707 8554 22719 8557
rect 22753 8554 22765 8588
rect 22707 8548 22765 8554
rect 1952 8412 23264 8434
rect 1952 8360 4494 8412
rect 4546 8360 4558 8412
rect 4610 8360 4622 8412
rect 4674 8360 4686 8412
rect 4738 8360 9822 8412
rect 9874 8360 9886 8412
rect 9938 8360 9950 8412
rect 10002 8360 10014 8412
rect 10066 8360 15150 8412
rect 15202 8360 15214 8412
rect 15266 8360 15278 8412
rect 15330 8360 15342 8412
rect 15394 8360 20478 8412
rect 20530 8360 20542 8412
rect 20594 8360 20606 8412
rect 20658 8360 20670 8412
rect 20722 8360 23264 8412
rect 1952 8338 23264 8360
rect 22608 8101 22614 8153
rect 22666 8141 22672 8153
rect 22707 8144 22765 8150
rect 22707 8141 22719 8144
rect 22666 8113 22719 8141
rect 22666 8101 22672 8113
rect 22707 8110 22719 8113
rect 22753 8110 22765 8144
rect 22707 8104 22765 8110
rect 3411 8070 3469 8076
rect 3411 8036 3423 8070
rect 3457 8067 3469 8070
rect 3888 8067 3894 8079
rect 3457 8039 3894 8067
rect 3457 8036 3469 8039
rect 3411 8030 3469 8036
rect 3888 8027 3894 8039
rect 3946 8027 3952 8079
rect 3987 8070 4045 8076
rect 3987 8036 3999 8070
rect 4033 8067 4045 8070
rect 4563 8070 4621 8076
rect 4563 8067 4575 8070
rect 4033 8039 4575 8067
rect 4033 8036 4045 8039
rect 3987 8030 4045 8036
rect 4563 8036 4575 8039
rect 4609 8036 4621 8070
rect 4563 8030 4621 8036
rect 5235 8070 5293 8076
rect 5235 8036 5247 8070
rect 5281 8067 5293 8070
rect 5811 8070 5869 8076
rect 5811 8067 5823 8070
rect 5281 8039 5823 8067
rect 5281 8036 5293 8039
rect 5235 8030 5293 8036
rect 5811 8036 5823 8039
rect 5857 8036 5869 8070
rect 5811 8030 5869 8036
rect 6483 8070 6541 8076
rect 6483 8036 6495 8070
rect 6529 8067 6541 8070
rect 7059 8070 7117 8076
rect 7059 8067 7071 8070
rect 6529 8039 7071 8067
rect 6529 8036 6541 8039
rect 6483 8030 6541 8036
rect 7059 8036 7071 8039
rect 7105 8036 7117 8070
rect 7059 8030 7117 8036
rect 7731 8070 7789 8076
rect 7731 8036 7743 8070
rect 7777 8067 7789 8070
rect 8307 8070 8365 8076
rect 8307 8067 8319 8070
rect 7777 8039 8319 8067
rect 7777 8036 7789 8039
rect 7731 8030 7789 8036
rect 8307 8036 8319 8039
rect 8353 8036 8365 8070
rect 8307 8030 8365 8036
rect 8979 8070 9037 8076
rect 8979 8036 8991 8070
rect 9025 8067 9037 8070
rect 9555 8070 9613 8076
rect 9555 8067 9567 8070
rect 9025 8039 9567 8067
rect 9025 8036 9037 8039
rect 8979 8030 9037 8036
rect 9555 8036 9567 8039
rect 9601 8036 9613 8070
rect 9555 8030 9613 8036
rect 10227 8070 10285 8076
rect 10227 8036 10239 8070
rect 10273 8067 10285 8070
rect 10803 8070 10861 8076
rect 10803 8067 10815 8070
rect 10273 8039 10815 8067
rect 10273 8036 10285 8039
rect 10227 8030 10285 8036
rect 10803 8036 10815 8039
rect 10849 8036 10861 8070
rect 10803 8030 10861 8036
rect 11475 8070 11533 8076
rect 11475 8036 11487 8070
rect 11521 8067 11533 8070
rect 12051 8070 12109 8076
rect 12051 8067 12063 8070
rect 11521 8039 12063 8067
rect 11521 8036 11533 8039
rect 11475 8030 11533 8036
rect 12051 8036 12063 8039
rect 12097 8036 12109 8070
rect 12051 8030 12109 8036
rect 12723 8070 12781 8076
rect 12723 8036 12735 8070
rect 12769 8067 12781 8070
rect 13299 8070 13357 8076
rect 13299 8067 13311 8070
rect 12769 8039 13311 8067
rect 12769 8036 12781 8039
rect 12723 8030 12781 8036
rect 13299 8036 13311 8039
rect 13345 8036 13357 8070
rect 13299 8030 13357 8036
rect 13971 8070 14029 8076
rect 13971 8036 13983 8070
rect 14017 8067 14029 8070
rect 14547 8070 14605 8076
rect 14547 8067 14559 8070
rect 14017 8039 14559 8067
rect 14017 8036 14029 8039
rect 13971 8030 14029 8036
rect 14547 8036 14559 8039
rect 14593 8036 14605 8070
rect 14547 8030 14605 8036
rect 15219 8070 15277 8076
rect 15219 8036 15231 8070
rect 15265 8067 15277 8070
rect 15795 8070 15853 8076
rect 15795 8067 15807 8070
rect 15265 8039 15807 8067
rect 15265 8036 15277 8039
rect 15219 8030 15277 8036
rect 15795 8036 15807 8039
rect 15841 8036 15853 8070
rect 15795 8030 15853 8036
rect 16467 8070 16525 8076
rect 16467 8036 16479 8070
rect 16513 8067 16525 8070
rect 17043 8070 17101 8076
rect 17043 8067 17055 8070
rect 16513 8039 17055 8067
rect 16513 8036 16525 8039
rect 16467 8030 16525 8036
rect 17043 8036 17055 8039
rect 17089 8036 17101 8070
rect 17043 8030 17101 8036
rect 17715 8070 17773 8076
rect 17715 8036 17727 8070
rect 17761 8067 17773 8070
rect 18291 8070 18349 8076
rect 18291 8067 18303 8070
rect 17761 8039 18303 8067
rect 17761 8036 17773 8039
rect 17715 8030 17773 8036
rect 18291 8036 18303 8039
rect 18337 8036 18349 8070
rect 18291 8030 18349 8036
rect 18963 8070 19021 8076
rect 18963 8036 18975 8070
rect 19009 8067 19021 8070
rect 19539 8070 19597 8076
rect 19539 8067 19551 8070
rect 19009 8039 19551 8067
rect 19009 8036 19021 8039
rect 18963 8030 19021 8036
rect 19539 8036 19551 8039
rect 19585 8036 19597 8070
rect 19539 8030 19597 8036
rect 20211 8070 20269 8076
rect 20211 8036 20223 8070
rect 20257 8067 20269 8070
rect 20787 8070 20845 8076
rect 20787 8067 20799 8070
rect 20257 8039 20799 8067
rect 20257 8036 20269 8039
rect 20211 8030 20269 8036
rect 20787 8036 20799 8039
rect 20833 8036 20845 8070
rect 20787 8030 20845 8036
rect 21459 8070 21517 8076
rect 21459 8036 21471 8070
rect 21505 8067 21517 8070
rect 22035 8070 22093 8076
rect 22035 8067 22047 8070
rect 21505 8039 22047 8067
rect 21505 8036 21517 8039
rect 21459 8030 21517 8036
rect 22035 8036 22047 8039
rect 22081 8036 22093 8070
rect 22035 8030 22093 8036
rect 1952 7746 23264 7768
rect 1952 7694 7158 7746
rect 7210 7694 7222 7746
rect 7274 7694 7286 7746
rect 7338 7694 7350 7746
rect 7402 7694 12486 7746
rect 12538 7694 12550 7746
rect 12602 7694 12614 7746
rect 12666 7694 12678 7746
rect 12730 7694 17814 7746
rect 17866 7694 17878 7746
rect 17930 7694 17942 7746
rect 17994 7694 18006 7746
rect 18058 7694 23264 7746
rect 1952 7672 23264 7694
rect 3888 7583 3894 7635
rect 3946 7623 3952 7635
rect 3987 7626 4045 7632
rect 3987 7623 3999 7626
rect 3946 7595 3999 7623
rect 3946 7583 3952 7595
rect 3987 7592 3999 7595
rect 4033 7592 4045 7626
rect 3987 7586 4045 7592
rect 3411 7404 3469 7410
rect 3411 7370 3423 7404
rect 3457 7401 3469 7404
rect 5235 7404 5293 7410
rect 5235 7401 5247 7404
rect 3457 7373 5247 7401
rect 3457 7370 3469 7373
rect 3411 7364 3469 7370
rect 5235 7370 5247 7373
rect 5281 7370 5293 7404
rect 5235 7364 5293 7370
rect 5907 7404 5965 7410
rect 5907 7370 5919 7404
rect 5953 7401 5965 7404
rect 7731 7404 7789 7410
rect 7731 7401 7743 7404
rect 5953 7373 7743 7401
rect 5953 7370 5965 7373
rect 5907 7364 5965 7370
rect 7731 7370 7743 7373
rect 7777 7370 7789 7404
rect 8979 7404 9037 7410
rect 8979 7401 8991 7404
rect 7731 7364 7789 7370
rect 8322 7373 8991 7401
rect 4659 7330 4717 7336
rect 4659 7296 4671 7330
rect 4705 7296 4717 7330
rect 4659 7290 4717 7296
rect 7155 7330 7213 7336
rect 7155 7296 7167 7330
rect 7201 7327 7213 7330
rect 8322 7327 8350 7373
rect 8979 7370 8991 7373
rect 9025 7370 9037 7404
rect 8979 7364 9037 7370
rect 9651 7404 9709 7410
rect 9651 7370 9663 7404
rect 9697 7401 9709 7404
rect 11475 7404 11533 7410
rect 11475 7401 11487 7404
rect 9697 7373 11487 7401
rect 9697 7370 9709 7373
rect 9651 7364 9709 7370
rect 11475 7370 11487 7373
rect 11521 7370 11533 7404
rect 11475 7364 11533 7370
rect 12147 7404 12205 7410
rect 12147 7370 12159 7404
rect 12193 7401 12205 7404
rect 13971 7404 14029 7410
rect 13971 7401 13983 7404
rect 12193 7373 13983 7401
rect 12193 7370 12205 7373
rect 12147 7364 12205 7370
rect 13971 7370 13983 7373
rect 14017 7370 14029 7404
rect 13971 7364 14029 7370
rect 14547 7404 14605 7410
rect 14547 7370 14559 7404
rect 14593 7401 14605 7404
rect 16467 7404 16525 7410
rect 16467 7401 16479 7404
rect 14593 7373 16479 7401
rect 14593 7370 14605 7373
rect 14547 7364 14605 7370
rect 16467 7370 16479 7373
rect 16513 7370 16525 7404
rect 16467 7364 16525 7370
rect 17139 7404 17197 7410
rect 17139 7370 17151 7404
rect 17185 7401 17197 7404
rect 18963 7404 19021 7410
rect 18963 7401 18975 7404
rect 17185 7373 18975 7401
rect 17185 7370 17197 7373
rect 17139 7364 17197 7370
rect 18963 7370 18975 7373
rect 19009 7370 19021 7404
rect 18963 7364 19021 7370
rect 19635 7404 19693 7410
rect 19635 7370 19647 7404
rect 19681 7401 19693 7404
rect 21459 7404 21517 7410
rect 21459 7401 21471 7404
rect 19681 7373 21471 7401
rect 19681 7370 19693 7373
rect 19635 7364 19693 7370
rect 21459 7370 21471 7373
rect 21505 7370 21517 7404
rect 21459 7364 21517 7370
rect 7201 7299 8350 7327
rect 8403 7330 8461 7336
rect 7201 7296 7213 7299
rect 7155 7290 7213 7296
rect 8403 7296 8415 7330
rect 8449 7327 8461 7330
rect 10227 7330 10285 7336
rect 10227 7327 10239 7330
rect 8449 7299 10239 7327
rect 8449 7296 8461 7299
rect 8403 7290 8461 7296
rect 10227 7296 10239 7299
rect 10273 7296 10285 7330
rect 10227 7290 10285 7296
rect 10899 7330 10957 7336
rect 10899 7296 10911 7330
rect 10945 7327 10957 7330
rect 12723 7330 12781 7336
rect 12723 7327 12735 7330
rect 10945 7299 12735 7327
rect 10945 7296 10957 7299
rect 10899 7290 10957 7296
rect 12723 7296 12735 7299
rect 12769 7296 12781 7330
rect 12723 7290 12781 7296
rect 13395 7330 13453 7336
rect 13395 7296 13407 7330
rect 13441 7327 13453 7330
rect 15219 7330 15277 7336
rect 15219 7327 15231 7330
rect 13441 7299 15231 7327
rect 13441 7296 13453 7299
rect 13395 7290 13453 7296
rect 15219 7296 15231 7299
rect 15265 7296 15277 7330
rect 15219 7290 15277 7296
rect 15891 7330 15949 7336
rect 15891 7296 15903 7330
rect 15937 7327 15949 7330
rect 17715 7330 17773 7336
rect 17715 7327 17727 7330
rect 15937 7299 17727 7327
rect 15937 7296 15949 7299
rect 15891 7290 15949 7296
rect 17715 7296 17727 7299
rect 17761 7296 17773 7330
rect 17715 7290 17773 7296
rect 18387 7330 18445 7336
rect 18387 7296 18399 7330
rect 18433 7327 18445 7330
rect 20211 7330 20269 7336
rect 20211 7327 20223 7330
rect 18433 7299 20223 7327
rect 18433 7296 18445 7299
rect 18387 7290 18445 7296
rect 20211 7296 20223 7299
rect 20257 7296 20269 7330
rect 20211 7290 20269 7296
rect 20883 7330 20941 7336
rect 20883 7296 20895 7330
rect 20929 7296 20941 7330
rect 22128 7327 22134 7339
rect 22089 7299 22134 7327
rect 20883 7290 20941 7296
rect 4674 7253 4702 7290
rect 6483 7256 6541 7262
rect 6483 7253 6495 7256
rect 4674 7225 6495 7253
rect 6483 7222 6495 7225
rect 6529 7222 6541 7256
rect 20898 7253 20926 7290
rect 22128 7287 22134 7299
rect 22186 7287 22192 7339
rect 22707 7256 22765 7262
rect 22707 7253 22719 7256
rect 20898 7225 22719 7253
rect 6483 7216 6541 7222
rect 22707 7222 22719 7225
rect 22753 7222 22765 7256
rect 22707 7216 22765 7222
rect 1952 7080 23264 7102
rect 1952 7028 4494 7080
rect 4546 7028 4558 7080
rect 4610 7028 4622 7080
rect 4674 7028 4686 7080
rect 4738 7028 9822 7080
rect 9874 7028 9886 7080
rect 9938 7028 9950 7080
rect 10002 7028 10014 7080
rect 10066 7028 15150 7080
rect 15202 7028 15214 7080
rect 15266 7028 15278 7080
rect 15330 7028 15342 7080
rect 15394 7028 20478 7080
rect 20530 7028 20542 7080
rect 20594 7028 20606 7080
rect 20658 7028 20670 7080
rect 20722 7028 23264 7080
rect 1952 7006 23264 7028
rect 22128 6917 22134 6969
rect 22186 6957 22192 6969
rect 22707 6960 22765 6966
rect 22707 6957 22719 6960
rect 22186 6929 22719 6957
rect 22186 6917 22192 6929
rect 22707 6926 22719 6929
rect 22753 6926 22765 6960
rect 22707 6920 22765 6926
rect 3411 6738 3469 6744
rect 3411 6704 3423 6738
rect 3457 6735 3469 6738
rect 3888 6735 3894 6747
rect 3457 6707 3894 6735
rect 3457 6704 3469 6707
rect 3411 6698 3469 6704
rect 3888 6695 3894 6707
rect 3946 6695 3952 6747
rect 3987 6738 4045 6744
rect 3987 6704 3999 6738
rect 4033 6735 4045 6738
rect 4563 6738 4621 6744
rect 4563 6735 4575 6738
rect 4033 6707 4575 6735
rect 4033 6704 4045 6707
rect 3987 6698 4045 6704
rect 4563 6704 4575 6707
rect 4609 6704 4621 6738
rect 4563 6698 4621 6704
rect 5235 6738 5293 6744
rect 5235 6704 5247 6738
rect 5281 6735 5293 6738
rect 5811 6738 5869 6744
rect 5811 6735 5823 6738
rect 5281 6707 5823 6735
rect 5281 6704 5293 6707
rect 5235 6698 5293 6704
rect 5811 6704 5823 6707
rect 5857 6704 5869 6738
rect 5811 6698 5869 6704
rect 6483 6738 6541 6744
rect 6483 6704 6495 6738
rect 6529 6735 6541 6738
rect 7059 6738 7117 6744
rect 7059 6735 7071 6738
rect 6529 6707 7071 6735
rect 6529 6704 6541 6707
rect 6483 6698 6541 6704
rect 7059 6704 7071 6707
rect 7105 6704 7117 6738
rect 7059 6698 7117 6704
rect 7731 6738 7789 6744
rect 7731 6704 7743 6738
rect 7777 6735 7789 6738
rect 8307 6738 8365 6744
rect 8307 6735 8319 6738
rect 7777 6707 8319 6735
rect 7777 6704 7789 6707
rect 7731 6698 7789 6704
rect 8307 6704 8319 6707
rect 8353 6704 8365 6738
rect 8307 6698 8365 6704
rect 8979 6738 9037 6744
rect 8979 6704 8991 6738
rect 9025 6735 9037 6738
rect 9555 6738 9613 6744
rect 9555 6735 9567 6738
rect 9025 6707 9567 6735
rect 9025 6704 9037 6707
rect 8979 6698 9037 6704
rect 9555 6704 9567 6707
rect 9601 6704 9613 6738
rect 9555 6698 9613 6704
rect 10227 6738 10285 6744
rect 10227 6704 10239 6738
rect 10273 6735 10285 6738
rect 10803 6738 10861 6744
rect 10803 6735 10815 6738
rect 10273 6707 10815 6735
rect 10273 6704 10285 6707
rect 10227 6698 10285 6704
rect 10803 6704 10815 6707
rect 10849 6704 10861 6738
rect 10803 6698 10861 6704
rect 11475 6738 11533 6744
rect 11475 6704 11487 6738
rect 11521 6735 11533 6738
rect 12051 6738 12109 6744
rect 12051 6735 12063 6738
rect 11521 6707 12063 6735
rect 11521 6704 11533 6707
rect 11475 6698 11533 6704
rect 12051 6704 12063 6707
rect 12097 6704 12109 6738
rect 12051 6698 12109 6704
rect 12723 6738 12781 6744
rect 12723 6704 12735 6738
rect 12769 6735 12781 6738
rect 13299 6738 13357 6744
rect 13299 6735 13311 6738
rect 12769 6707 13311 6735
rect 12769 6704 12781 6707
rect 12723 6698 12781 6704
rect 13299 6704 13311 6707
rect 13345 6704 13357 6738
rect 13299 6698 13357 6704
rect 13971 6738 14029 6744
rect 13971 6704 13983 6738
rect 14017 6735 14029 6738
rect 14547 6738 14605 6744
rect 14547 6735 14559 6738
rect 14017 6707 14559 6735
rect 14017 6704 14029 6707
rect 13971 6698 14029 6704
rect 14547 6704 14559 6707
rect 14593 6704 14605 6738
rect 14547 6698 14605 6704
rect 15219 6738 15277 6744
rect 15219 6704 15231 6738
rect 15265 6735 15277 6738
rect 15795 6738 15853 6744
rect 15795 6735 15807 6738
rect 15265 6707 15807 6735
rect 15265 6704 15277 6707
rect 15219 6698 15277 6704
rect 15795 6704 15807 6707
rect 15841 6704 15853 6738
rect 15795 6698 15853 6704
rect 16467 6738 16525 6744
rect 16467 6704 16479 6738
rect 16513 6735 16525 6738
rect 17043 6738 17101 6744
rect 17043 6735 17055 6738
rect 16513 6707 17055 6735
rect 16513 6704 16525 6707
rect 16467 6698 16525 6704
rect 17043 6704 17055 6707
rect 17089 6704 17101 6738
rect 17043 6698 17101 6704
rect 17715 6738 17773 6744
rect 17715 6704 17727 6738
rect 17761 6735 17773 6738
rect 18291 6738 18349 6744
rect 18291 6735 18303 6738
rect 17761 6707 18303 6735
rect 17761 6704 17773 6707
rect 17715 6698 17773 6704
rect 18291 6704 18303 6707
rect 18337 6704 18349 6738
rect 18291 6698 18349 6704
rect 18963 6738 19021 6744
rect 18963 6704 18975 6738
rect 19009 6735 19021 6738
rect 19539 6738 19597 6744
rect 19539 6735 19551 6738
rect 19009 6707 19551 6735
rect 19009 6704 19021 6707
rect 18963 6698 19021 6704
rect 19539 6704 19551 6707
rect 19585 6704 19597 6738
rect 19539 6698 19597 6704
rect 20211 6738 20269 6744
rect 20211 6704 20223 6738
rect 20257 6735 20269 6738
rect 20787 6738 20845 6744
rect 20787 6735 20799 6738
rect 20257 6707 20799 6735
rect 20257 6704 20269 6707
rect 20211 6698 20269 6704
rect 20787 6704 20799 6707
rect 20833 6704 20845 6738
rect 20787 6698 20845 6704
rect 21459 6738 21517 6744
rect 21459 6704 21471 6738
rect 21505 6735 21517 6738
rect 22035 6738 22093 6744
rect 22035 6735 22047 6738
rect 21505 6707 22047 6735
rect 21505 6704 21517 6707
rect 21459 6698 21517 6704
rect 22035 6704 22047 6707
rect 22081 6704 22093 6738
rect 22035 6698 22093 6704
rect 1952 6414 23264 6436
rect 1952 6362 7158 6414
rect 7210 6362 7222 6414
rect 7274 6362 7286 6414
rect 7338 6362 7350 6414
rect 7402 6362 12486 6414
rect 12538 6362 12550 6414
rect 12602 6362 12614 6414
rect 12666 6362 12678 6414
rect 12730 6362 17814 6414
rect 17866 6362 17878 6414
rect 17930 6362 17942 6414
rect 17994 6362 18006 6414
rect 18058 6362 23264 6414
rect 1952 6340 23264 6362
rect 3888 6251 3894 6303
rect 3946 6291 3952 6303
rect 3987 6294 4045 6300
rect 3987 6291 3999 6294
rect 3946 6263 3999 6291
rect 3946 6251 3952 6263
rect 3987 6260 3999 6263
rect 4033 6260 4045 6294
rect 3987 6254 4045 6260
rect 21459 6146 21517 6152
rect 21459 6143 21471 6146
rect 20802 6115 21471 6143
rect 3411 6072 3469 6078
rect 3411 6038 3423 6072
rect 3457 6069 3469 6072
rect 5235 6072 5293 6078
rect 5235 6069 5247 6072
rect 3457 6041 5247 6069
rect 3457 6038 3469 6041
rect 3411 6032 3469 6038
rect 5235 6038 5247 6041
rect 5281 6038 5293 6072
rect 5235 6032 5293 6038
rect 5907 6072 5965 6078
rect 5907 6038 5919 6072
rect 5953 6069 5965 6072
rect 7731 6072 7789 6078
rect 7731 6069 7743 6072
rect 5953 6041 7743 6069
rect 5953 6038 5965 6041
rect 5907 6032 5965 6038
rect 7731 6038 7743 6041
rect 7777 6038 7789 6072
rect 8979 6072 9037 6078
rect 8979 6069 8991 6072
rect 7731 6032 7789 6038
rect 8322 6041 8991 6069
rect 4659 5998 4717 6004
rect 4659 5964 4671 5998
rect 4705 5964 4717 5998
rect 4659 5958 4717 5964
rect 7155 5998 7213 6004
rect 7155 5964 7167 5998
rect 7201 5995 7213 5998
rect 8322 5995 8350 6041
rect 8979 6038 8991 6041
rect 9025 6038 9037 6072
rect 8979 6032 9037 6038
rect 9651 6072 9709 6078
rect 9651 6038 9663 6072
rect 9697 6069 9709 6072
rect 11475 6072 11533 6078
rect 11475 6069 11487 6072
rect 9697 6041 11487 6069
rect 9697 6038 9709 6041
rect 9651 6032 9709 6038
rect 11475 6038 11487 6041
rect 11521 6038 11533 6072
rect 11475 6032 11533 6038
rect 12147 6072 12205 6078
rect 12147 6038 12159 6072
rect 12193 6069 12205 6072
rect 13971 6072 14029 6078
rect 13971 6069 13983 6072
rect 12193 6041 13983 6069
rect 12193 6038 12205 6041
rect 12147 6032 12205 6038
rect 13971 6038 13983 6041
rect 14017 6038 14029 6072
rect 13971 6032 14029 6038
rect 14547 6072 14605 6078
rect 14547 6038 14559 6072
rect 14593 6069 14605 6072
rect 16467 6072 16525 6078
rect 16467 6069 16479 6072
rect 14593 6041 16479 6069
rect 14593 6038 14605 6041
rect 14547 6032 14605 6038
rect 16467 6038 16479 6041
rect 16513 6038 16525 6072
rect 16467 6032 16525 6038
rect 18387 6072 18445 6078
rect 18387 6038 18399 6072
rect 18433 6069 18445 6072
rect 20211 6072 20269 6078
rect 20211 6069 20223 6072
rect 18433 6041 20223 6069
rect 18433 6038 18445 6041
rect 18387 6032 18445 6038
rect 20211 6038 20223 6041
rect 20257 6038 20269 6072
rect 20211 6032 20269 6038
rect 7201 5967 8350 5995
rect 8403 5998 8461 6004
rect 7201 5964 7213 5967
rect 7155 5958 7213 5964
rect 8403 5964 8415 5998
rect 8449 5995 8461 5998
rect 10227 5998 10285 6004
rect 10227 5995 10239 5998
rect 8449 5967 10239 5995
rect 8449 5964 8461 5967
rect 8403 5958 8461 5964
rect 10227 5964 10239 5967
rect 10273 5964 10285 5998
rect 10227 5958 10285 5964
rect 10899 5998 10957 6004
rect 10899 5964 10911 5998
rect 10945 5995 10957 5998
rect 12723 5998 12781 6004
rect 12723 5995 12735 5998
rect 10945 5967 12735 5995
rect 10945 5964 10957 5967
rect 10899 5958 10957 5964
rect 12723 5964 12735 5967
rect 12769 5964 12781 5998
rect 12723 5958 12781 5964
rect 13395 5998 13453 6004
rect 13395 5964 13407 5998
rect 13441 5995 13453 5998
rect 15219 5998 15277 6004
rect 15219 5995 15231 5998
rect 13441 5967 15231 5995
rect 13441 5964 13453 5967
rect 13395 5958 13453 5964
rect 15219 5964 15231 5967
rect 15265 5964 15277 5998
rect 15219 5958 15277 5964
rect 15891 5998 15949 6004
rect 15891 5964 15903 5998
rect 15937 5964 15949 5998
rect 15891 5958 15949 5964
rect 17139 5998 17197 6004
rect 17139 5964 17151 5998
rect 17185 5995 17197 5998
rect 18963 5998 19021 6004
rect 18963 5995 18975 5998
rect 17185 5967 18975 5995
rect 17185 5964 17197 5967
rect 17139 5958 17197 5964
rect 18963 5964 18975 5967
rect 19009 5964 19021 5998
rect 18963 5958 19021 5964
rect 19635 5998 19693 6004
rect 19635 5964 19647 5998
rect 19681 5995 19693 5998
rect 20802 5995 20830 6115
rect 21459 6112 21471 6115
rect 21505 6112 21517 6146
rect 21459 6106 21517 6112
rect 19681 5967 20830 5995
rect 20883 5998 20941 6004
rect 19681 5964 19693 5967
rect 19635 5958 19693 5964
rect 20883 5964 20895 5998
rect 20929 5964 20941 5998
rect 20883 5958 20941 5964
rect 22131 5998 22189 6004
rect 22131 5964 22143 5998
rect 22177 5995 22189 5998
rect 22608 5995 22614 6007
rect 22177 5967 22614 5995
rect 22177 5964 22189 5967
rect 22131 5958 22189 5964
rect 4674 5921 4702 5958
rect 6483 5924 6541 5930
rect 6483 5921 6495 5924
rect 4674 5893 6495 5921
rect 6483 5890 6495 5893
rect 6529 5890 6541 5924
rect 15906 5921 15934 5958
rect 17715 5924 17773 5930
rect 17715 5921 17727 5924
rect 15906 5893 17727 5921
rect 6483 5884 6541 5890
rect 17715 5890 17727 5893
rect 17761 5890 17773 5924
rect 20898 5921 20926 5958
rect 22608 5955 22614 5967
rect 22666 5955 22672 6007
rect 22707 5924 22765 5930
rect 22707 5921 22719 5924
rect 20898 5893 22719 5921
rect 17715 5884 17773 5890
rect 22707 5890 22719 5893
rect 22753 5890 22765 5924
rect 22707 5884 22765 5890
rect 1952 5748 23264 5770
rect 1952 5696 4494 5748
rect 4546 5696 4558 5748
rect 4610 5696 4622 5748
rect 4674 5696 4686 5748
rect 4738 5696 9822 5748
rect 9874 5696 9886 5748
rect 9938 5696 9950 5748
rect 10002 5696 10014 5748
rect 10066 5696 15150 5748
rect 15202 5696 15214 5748
rect 15266 5696 15278 5748
rect 15330 5696 15342 5748
rect 15394 5696 20478 5748
rect 20530 5696 20542 5748
rect 20594 5696 20606 5748
rect 20658 5696 20670 5748
rect 20722 5696 23264 5748
rect 1952 5674 23264 5696
rect 22608 5585 22614 5637
rect 22666 5625 22672 5637
rect 22707 5628 22765 5634
rect 22707 5625 22719 5628
rect 22666 5597 22719 5625
rect 22666 5585 22672 5597
rect 22707 5594 22719 5597
rect 22753 5594 22765 5628
rect 22707 5588 22765 5594
rect 3411 5406 3469 5412
rect 3411 5372 3423 5406
rect 3457 5403 3469 5406
rect 3888 5403 3894 5415
rect 3457 5375 3894 5403
rect 3457 5372 3469 5375
rect 3411 5366 3469 5372
rect 3888 5363 3894 5375
rect 3946 5363 3952 5415
rect 3987 5406 4045 5412
rect 3987 5372 3999 5406
rect 4033 5403 4045 5406
rect 4563 5406 4621 5412
rect 4563 5403 4575 5406
rect 4033 5375 4575 5403
rect 4033 5372 4045 5375
rect 3987 5366 4045 5372
rect 4563 5372 4575 5375
rect 4609 5372 4621 5406
rect 4563 5366 4621 5372
rect 5235 5406 5293 5412
rect 5235 5372 5247 5406
rect 5281 5403 5293 5406
rect 5811 5406 5869 5412
rect 5811 5403 5823 5406
rect 5281 5375 5823 5403
rect 5281 5372 5293 5375
rect 5235 5366 5293 5372
rect 5811 5372 5823 5375
rect 5857 5372 5869 5406
rect 5811 5366 5869 5372
rect 6483 5406 6541 5412
rect 6483 5372 6495 5406
rect 6529 5403 6541 5406
rect 7059 5406 7117 5412
rect 7059 5403 7071 5406
rect 6529 5375 7071 5403
rect 6529 5372 6541 5375
rect 6483 5366 6541 5372
rect 7059 5372 7071 5375
rect 7105 5372 7117 5406
rect 7059 5366 7117 5372
rect 7731 5406 7789 5412
rect 7731 5372 7743 5406
rect 7777 5403 7789 5406
rect 8307 5406 8365 5412
rect 8307 5403 8319 5406
rect 7777 5375 8319 5403
rect 7777 5372 7789 5375
rect 7731 5366 7789 5372
rect 8307 5372 8319 5375
rect 8353 5372 8365 5406
rect 8307 5366 8365 5372
rect 8979 5406 9037 5412
rect 8979 5372 8991 5406
rect 9025 5403 9037 5406
rect 9555 5406 9613 5412
rect 9555 5403 9567 5406
rect 9025 5375 9567 5403
rect 9025 5372 9037 5375
rect 8979 5366 9037 5372
rect 9555 5372 9567 5375
rect 9601 5372 9613 5406
rect 9555 5366 9613 5372
rect 10227 5406 10285 5412
rect 10227 5372 10239 5406
rect 10273 5403 10285 5406
rect 10803 5406 10861 5412
rect 10803 5403 10815 5406
rect 10273 5375 10815 5403
rect 10273 5372 10285 5375
rect 10227 5366 10285 5372
rect 10803 5372 10815 5375
rect 10849 5372 10861 5406
rect 10803 5366 10861 5372
rect 11475 5406 11533 5412
rect 11475 5372 11487 5406
rect 11521 5403 11533 5406
rect 12051 5406 12109 5412
rect 12051 5403 12063 5406
rect 11521 5375 12063 5403
rect 11521 5372 11533 5375
rect 11475 5366 11533 5372
rect 12051 5372 12063 5375
rect 12097 5372 12109 5406
rect 12051 5366 12109 5372
rect 12723 5406 12781 5412
rect 12723 5372 12735 5406
rect 12769 5403 12781 5406
rect 13299 5406 13357 5412
rect 13299 5403 13311 5406
rect 12769 5375 13311 5403
rect 12769 5372 12781 5375
rect 12723 5366 12781 5372
rect 13299 5372 13311 5375
rect 13345 5372 13357 5406
rect 13299 5366 13357 5372
rect 13971 5406 14029 5412
rect 13971 5372 13983 5406
rect 14017 5403 14029 5406
rect 14547 5406 14605 5412
rect 14547 5403 14559 5406
rect 14017 5375 14559 5403
rect 14017 5372 14029 5375
rect 13971 5366 14029 5372
rect 14547 5372 14559 5375
rect 14593 5372 14605 5406
rect 14547 5366 14605 5372
rect 15219 5406 15277 5412
rect 15219 5372 15231 5406
rect 15265 5403 15277 5406
rect 15795 5406 15853 5412
rect 15795 5403 15807 5406
rect 15265 5375 15807 5403
rect 15265 5372 15277 5375
rect 15219 5366 15277 5372
rect 15795 5372 15807 5375
rect 15841 5372 15853 5406
rect 15795 5366 15853 5372
rect 16467 5406 16525 5412
rect 16467 5372 16479 5406
rect 16513 5403 16525 5406
rect 17043 5406 17101 5412
rect 17043 5403 17055 5406
rect 16513 5375 17055 5403
rect 16513 5372 16525 5375
rect 16467 5366 16525 5372
rect 17043 5372 17055 5375
rect 17089 5372 17101 5406
rect 17043 5366 17101 5372
rect 17715 5406 17773 5412
rect 17715 5372 17727 5406
rect 17761 5403 17773 5406
rect 18291 5406 18349 5412
rect 18291 5403 18303 5406
rect 17761 5375 18303 5403
rect 17761 5372 17773 5375
rect 17715 5366 17773 5372
rect 18291 5372 18303 5375
rect 18337 5372 18349 5406
rect 18291 5366 18349 5372
rect 18963 5406 19021 5412
rect 18963 5372 18975 5406
rect 19009 5403 19021 5406
rect 19539 5406 19597 5412
rect 19539 5403 19551 5406
rect 19009 5375 19551 5403
rect 19009 5372 19021 5375
rect 18963 5366 19021 5372
rect 19539 5372 19551 5375
rect 19585 5372 19597 5406
rect 19539 5366 19597 5372
rect 20211 5406 20269 5412
rect 20211 5372 20223 5406
rect 20257 5403 20269 5406
rect 20787 5406 20845 5412
rect 20787 5403 20799 5406
rect 20257 5375 20799 5403
rect 20257 5372 20269 5375
rect 20211 5366 20269 5372
rect 20787 5372 20799 5375
rect 20833 5372 20845 5406
rect 20787 5366 20845 5372
rect 21459 5406 21517 5412
rect 21459 5372 21471 5406
rect 21505 5403 21517 5406
rect 22035 5406 22093 5412
rect 22035 5403 22047 5406
rect 21505 5375 22047 5403
rect 21505 5372 21517 5375
rect 21459 5366 21517 5372
rect 22035 5372 22047 5375
rect 22081 5372 22093 5406
rect 22035 5366 22093 5372
rect 1952 5082 23264 5104
rect 1952 5030 7158 5082
rect 7210 5030 7222 5082
rect 7274 5030 7286 5082
rect 7338 5030 7350 5082
rect 7402 5030 12486 5082
rect 12538 5030 12550 5082
rect 12602 5030 12614 5082
rect 12666 5030 12678 5082
rect 12730 5030 17814 5082
rect 17866 5030 17878 5082
rect 17930 5030 17942 5082
rect 17994 5030 18006 5082
rect 18058 5030 23264 5082
rect 1952 5008 23264 5030
rect 3888 4919 3894 4971
rect 3946 4959 3952 4971
rect 3987 4962 4045 4968
rect 3987 4959 3999 4962
rect 3946 4931 3999 4959
rect 3946 4919 3952 4931
rect 3987 4928 3999 4931
rect 4033 4928 4045 4962
rect 3987 4922 4045 4928
rect 4659 4740 4717 4746
rect 4659 4706 4671 4740
rect 4705 4737 4717 4740
rect 6483 4740 6541 4746
rect 6483 4737 6495 4740
rect 4705 4709 6495 4737
rect 4705 4706 4717 4709
rect 4659 4700 4717 4706
rect 6483 4706 6495 4709
rect 6529 4706 6541 4740
rect 8979 4740 9037 4746
rect 8979 4737 8991 4740
rect 6483 4700 6541 4706
rect 8322 4709 8991 4737
rect 3411 4666 3469 4672
rect 3411 4632 3423 4666
rect 3457 4663 3469 4666
rect 5235 4666 5293 4672
rect 5235 4663 5247 4666
rect 3457 4635 5247 4663
rect 3457 4632 3469 4635
rect 3411 4626 3469 4632
rect 5235 4632 5247 4635
rect 5281 4632 5293 4666
rect 5235 4626 5293 4632
rect 5907 4666 5965 4672
rect 5907 4632 5919 4666
rect 5953 4632 5965 4666
rect 5907 4626 5965 4632
rect 7155 4666 7213 4672
rect 7155 4632 7167 4666
rect 7201 4663 7213 4666
rect 8322 4663 8350 4709
rect 8979 4706 8991 4709
rect 9025 4706 9037 4740
rect 8979 4700 9037 4706
rect 9651 4740 9709 4746
rect 9651 4706 9663 4740
rect 9697 4737 9709 4740
rect 11475 4740 11533 4746
rect 11475 4737 11487 4740
rect 9697 4709 11487 4737
rect 9697 4706 9709 4709
rect 9651 4700 9709 4706
rect 11475 4706 11487 4709
rect 11521 4706 11533 4740
rect 11475 4700 11533 4706
rect 12147 4740 12205 4746
rect 12147 4706 12159 4740
rect 12193 4737 12205 4740
rect 13971 4740 14029 4746
rect 13971 4737 13983 4740
rect 12193 4709 13983 4737
rect 12193 4706 12205 4709
rect 12147 4700 12205 4706
rect 13971 4706 13983 4709
rect 14017 4706 14029 4740
rect 13971 4700 14029 4706
rect 14547 4740 14605 4746
rect 14547 4706 14559 4740
rect 14593 4737 14605 4740
rect 16467 4740 16525 4746
rect 16467 4737 16479 4740
rect 14593 4709 16479 4737
rect 14593 4706 14605 4709
rect 14547 4700 14605 4706
rect 16467 4706 16479 4709
rect 16513 4706 16525 4740
rect 16467 4700 16525 4706
rect 17139 4740 17197 4746
rect 17139 4706 17151 4740
rect 17185 4737 17197 4740
rect 18963 4740 19021 4746
rect 18963 4737 18975 4740
rect 17185 4709 18975 4737
rect 17185 4706 17197 4709
rect 17139 4700 17197 4706
rect 18963 4706 18975 4709
rect 19009 4706 19021 4740
rect 18963 4700 19021 4706
rect 19635 4740 19693 4746
rect 19635 4706 19647 4740
rect 19681 4737 19693 4740
rect 21459 4740 21517 4746
rect 21459 4737 21471 4740
rect 19681 4709 21471 4737
rect 19681 4706 19693 4709
rect 19635 4700 19693 4706
rect 21459 4706 21471 4709
rect 21505 4706 21517 4740
rect 21459 4700 21517 4706
rect 7201 4635 8350 4663
rect 8403 4666 8461 4672
rect 7201 4632 7213 4635
rect 7155 4626 7213 4632
rect 8403 4632 8415 4666
rect 8449 4663 8461 4666
rect 10227 4666 10285 4672
rect 10227 4663 10239 4666
rect 8449 4635 10239 4663
rect 8449 4632 8461 4635
rect 8403 4626 8461 4632
rect 10227 4632 10239 4635
rect 10273 4632 10285 4666
rect 10227 4626 10285 4632
rect 10899 4666 10957 4672
rect 10899 4632 10911 4666
rect 10945 4663 10957 4666
rect 12723 4666 12781 4672
rect 12723 4663 12735 4666
rect 10945 4635 12735 4663
rect 10945 4632 10957 4635
rect 10899 4626 10957 4632
rect 12723 4632 12735 4635
rect 12769 4632 12781 4666
rect 12723 4626 12781 4632
rect 13395 4666 13453 4672
rect 13395 4632 13407 4666
rect 13441 4663 13453 4666
rect 15219 4666 15277 4672
rect 15219 4663 15231 4666
rect 13441 4635 15231 4663
rect 13441 4632 13453 4635
rect 13395 4626 13453 4632
rect 15219 4632 15231 4635
rect 15265 4632 15277 4666
rect 15219 4626 15277 4632
rect 15891 4666 15949 4672
rect 15891 4632 15903 4666
rect 15937 4663 15949 4666
rect 17715 4666 17773 4672
rect 17715 4663 17727 4666
rect 15937 4635 17727 4663
rect 15937 4632 15949 4635
rect 15891 4626 15949 4632
rect 17715 4632 17727 4635
rect 17761 4632 17773 4666
rect 17715 4626 17773 4632
rect 18387 4666 18445 4672
rect 18387 4632 18399 4666
rect 18433 4663 18445 4666
rect 20211 4666 20269 4672
rect 20211 4663 20223 4666
rect 18433 4635 20223 4663
rect 18433 4632 18445 4635
rect 18387 4626 18445 4632
rect 20211 4632 20223 4635
rect 20257 4632 20269 4666
rect 20211 4626 20269 4632
rect 20883 4666 20941 4672
rect 20883 4632 20895 4666
rect 20929 4632 20941 4666
rect 20883 4626 20941 4632
rect 22131 4666 22189 4672
rect 22131 4632 22143 4666
rect 22177 4663 22189 4666
rect 22608 4663 22614 4675
rect 22177 4635 22614 4663
rect 22177 4632 22189 4635
rect 22131 4626 22189 4632
rect 5922 4589 5950 4626
rect 7731 4592 7789 4598
rect 7731 4589 7743 4592
rect 5922 4561 7743 4589
rect 7731 4558 7743 4561
rect 7777 4558 7789 4592
rect 20898 4589 20926 4626
rect 22608 4623 22614 4635
rect 22666 4623 22672 4675
rect 22707 4592 22765 4598
rect 22707 4589 22719 4592
rect 20898 4561 22719 4589
rect 7731 4552 7789 4558
rect 22707 4558 22719 4561
rect 22753 4558 22765 4592
rect 22707 4552 22765 4558
rect 1952 4416 23264 4438
rect 1952 4364 4494 4416
rect 4546 4364 4558 4416
rect 4610 4364 4622 4416
rect 4674 4364 4686 4416
rect 4738 4364 9822 4416
rect 9874 4364 9886 4416
rect 9938 4364 9950 4416
rect 10002 4364 10014 4416
rect 10066 4364 15150 4416
rect 15202 4364 15214 4416
rect 15266 4364 15278 4416
rect 15330 4364 15342 4416
rect 15394 4364 20478 4416
rect 20530 4364 20542 4416
rect 20594 4364 20606 4416
rect 20658 4364 20670 4416
rect 20722 4364 23264 4416
rect 1952 4342 23264 4364
rect 22608 4253 22614 4305
rect 22666 4293 22672 4305
rect 22707 4296 22765 4302
rect 22707 4293 22719 4296
rect 22666 4265 22719 4293
rect 22666 4253 22672 4265
rect 22707 4262 22719 4265
rect 22753 4262 22765 4296
rect 22707 4256 22765 4262
rect 3411 4074 3469 4080
rect 3411 4040 3423 4074
rect 3457 4071 3469 4074
rect 3888 4071 3894 4083
rect 3457 4043 3894 4071
rect 3457 4040 3469 4043
rect 3411 4034 3469 4040
rect 3888 4031 3894 4043
rect 3946 4031 3952 4083
rect 3987 4074 4045 4080
rect 3987 4040 3999 4074
rect 4033 4071 4045 4074
rect 4563 4074 4621 4080
rect 4563 4071 4575 4074
rect 4033 4043 4575 4071
rect 4033 4040 4045 4043
rect 3987 4034 4045 4040
rect 4563 4040 4575 4043
rect 4609 4040 4621 4074
rect 4563 4034 4621 4040
rect 5235 4074 5293 4080
rect 5235 4040 5247 4074
rect 5281 4071 5293 4074
rect 5811 4074 5869 4080
rect 5811 4071 5823 4074
rect 5281 4043 5823 4071
rect 5281 4040 5293 4043
rect 5235 4034 5293 4040
rect 5811 4040 5823 4043
rect 5857 4040 5869 4074
rect 5811 4034 5869 4040
rect 6483 4074 6541 4080
rect 6483 4040 6495 4074
rect 6529 4071 6541 4074
rect 7059 4074 7117 4080
rect 7059 4071 7071 4074
rect 6529 4043 7071 4071
rect 6529 4040 6541 4043
rect 6483 4034 6541 4040
rect 7059 4040 7071 4043
rect 7105 4040 7117 4074
rect 7059 4034 7117 4040
rect 7731 4074 7789 4080
rect 7731 4040 7743 4074
rect 7777 4071 7789 4074
rect 8307 4074 8365 4080
rect 8307 4071 8319 4074
rect 7777 4043 8319 4071
rect 7777 4040 7789 4043
rect 7731 4034 7789 4040
rect 8307 4040 8319 4043
rect 8353 4040 8365 4074
rect 8307 4034 8365 4040
rect 8979 4074 9037 4080
rect 8979 4040 8991 4074
rect 9025 4071 9037 4074
rect 9555 4074 9613 4080
rect 9555 4071 9567 4074
rect 9025 4043 9567 4071
rect 9025 4040 9037 4043
rect 8979 4034 9037 4040
rect 9555 4040 9567 4043
rect 9601 4040 9613 4074
rect 9555 4034 9613 4040
rect 10227 4074 10285 4080
rect 10227 4040 10239 4074
rect 10273 4071 10285 4074
rect 10803 4074 10861 4080
rect 10803 4071 10815 4074
rect 10273 4043 10815 4071
rect 10273 4040 10285 4043
rect 10227 4034 10285 4040
rect 10803 4040 10815 4043
rect 10849 4040 10861 4074
rect 10803 4034 10861 4040
rect 11475 4074 11533 4080
rect 11475 4040 11487 4074
rect 11521 4071 11533 4074
rect 12051 4074 12109 4080
rect 12051 4071 12063 4074
rect 11521 4043 12063 4071
rect 11521 4040 11533 4043
rect 11475 4034 11533 4040
rect 12051 4040 12063 4043
rect 12097 4040 12109 4074
rect 12051 4034 12109 4040
rect 12723 4074 12781 4080
rect 12723 4040 12735 4074
rect 12769 4071 12781 4074
rect 13299 4074 13357 4080
rect 13299 4071 13311 4074
rect 12769 4043 13311 4071
rect 12769 4040 12781 4043
rect 12723 4034 12781 4040
rect 13299 4040 13311 4043
rect 13345 4040 13357 4074
rect 13299 4034 13357 4040
rect 13971 4074 14029 4080
rect 13971 4040 13983 4074
rect 14017 4071 14029 4074
rect 14547 4074 14605 4080
rect 14547 4071 14559 4074
rect 14017 4043 14559 4071
rect 14017 4040 14029 4043
rect 13971 4034 14029 4040
rect 14547 4040 14559 4043
rect 14593 4040 14605 4074
rect 14547 4034 14605 4040
rect 15219 4074 15277 4080
rect 15219 4040 15231 4074
rect 15265 4071 15277 4074
rect 15795 4074 15853 4080
rect 15795 4071 15807 4074
rect 15265 4043 15807 4071
rect 15265 4040 15277 4043
rect 15219 4034 15277 4040
rect 15795 4040 15807 4043
rect 15841 4040 15853 4074
rect 15795 4034 15853 4040
rect 16467 4074 16525 4080
rect 16467 4040 16479 4074
rect 16513 4071 16525 4074
rect 17043 4074 17101 4080
rect 17043 4071 17055 4074
rect 16513 4043 17055 4071
rect 16513 4040 16525 4043
rect 16467 4034 16525 4040
rect 17043 4040 17055 4043
rect 17089 4040 17101 4074
rect 17043 4034 17101 4040
rect 17715 4074 17773 4080
rect 17715 4040 17727 4074
rect 17761 4071 17773 4074
rect 18291 4074 18349 4080
rect 18291 4071 18303 4074
rect 17761 4043 18303 4071
rect 17761 4040 17773 4043
rect 17715 4034 17773 4040
rect 18291 4040 18303 4043
rect 18337 4040 18349 4074
rect 18291 4034 18349 4040
rect 18963 4074 19021 4080
rect 18963 4040 18975 4074
rect 19009 4071 19021 4074
rect 19539 4074 19597 4080
rect 19539 4071 19551 4074
rect 19009 4043 19551 4071
rect 19009 4040 19021 4043
rect 18963 4034 19021 4040
rect 19539 4040 19551 4043
rect 19585 4040 19597 4074
rect 19539 4034 19597 4040
rect 20211 4074 20269 4080
rect 20211 4040 20223 4074
rect 20257 4071 20269 4074
rect 20787 4074 20845 4080
rect 20787 4071 20799 4074
rect 20257 4043 20799 4071
rect 20257 4040 20269 4043
rect 20211 4034 20269 4040
rect 20787 4040 20799 4043
rect 20833 4040 20845 4074
rect 20787 4034 20845 4040
rect 21459 4074 21517 4080
rect 21459 4040 21471 4074
rect 21505 4071 21517 4074
rect 22035 4074 22093 4080
rect 22035 4071 22047 4074
rect 21505 4043 22047 4071
rect 21505 4040 21517 4043
rect 21459 4034 21517 4040
rect 22035 4040 22047 4043
rect 22081 4040 22093 4074
rect 22035 4034 22093 4040
rect 1952 3750 23264 3772
rect 1952 3698 7158 3750
rect 7210 3698 7222 3750
rect 7274 3698 7286 3750
rect 7338 3698 7350 3750
rect 7402 3698 12486 3750
rect 12538 3698 12550 3750
rect 12602 3698 12614 3750
rect 12666 3698 12678 3750
rect 12730 3698 17814 3750
rect 17866 3698 17878 3750
rect 17930 3698 17942 3750
rect 17994 3698 18006 3750
rect 18058 3698 23264 3750
rect 1952 3676 23264 3698
rect 3888 3513 3894 3565
rect 3946 3553 3952 3565
rect 3987 3556 4045 3562
rect 3987 3553 3999 3556
rect 3946 3525 3999 3553
rect 3946 3513 3952 3525
rect 3987 3522 3999 3525
rect 4033 3522 4045 3556
rect 3987 3516 4045 3522
rect 3411 3408 3469 3414
rect 3411 3374 3423 3408
rect 3457 3405 3469 3408
rect 5235 3408 5293 3414
rect 5235 3405 5247 3408
rect 3457 3377 5247 3405
rect 3457 3374 3469 3377
rect 3411 3368 3469 3374
rect 5235 3374 5247 3377
rect 5281 3374 5293 3408
rect 5235 3368 5293 3374
rect 5907 3408 5965 3414
rect 5907 3374 5919 3408
rect 5953 3405 5965 3408
rect 7731 3408 7789 3414
rect 7731 3405 7743 3408
rect 5953 3377 7743 3405
rect 5953 3374 5965 3377
rect 5907 3368 5965 3374
rect 7731 3374 7743 3377
rect 7777 3374 7789 3408
rect 8979 3408 9037 3414
rect 8979 3405 8991 3408
rect 7731 3368 7789 3374
rect 8322 3377 8991 3405
rect 4659 3334 4717 3340
rect 4659 3300 4671 3334
rect 4705 3300 4717 3334
rect 4659 3294 4717 3300
rect 7155 3334 7213 3340
rect 7155 3300 7167 3334
rect 7201 3331 7213 3334
rect 8322 3331 8350 3377
rect 8979 3374 8991 3377
rect 9025 3374 9037 3408
rect 8979 3368 9037 3374
rect 9651 3408 9709 3414
rect 9651 3374 9663 3408
rect 9697 3405 9709 3408
rect 11475 3408 11533 3414
rect 11475 3405 11487 3408
rect 9697 3377 11487 3405
rect 9697 3374 9709 3377
rect 9651 3368 9709 3374
rect 11475 3374 11487 3377
rect 11521 3374 11533 3408
rect 11475 3368 11533 3374
rect 12147 3408 12205 3414
rect 12147 3374 12159 3408
rect 12193 3405 12205 3408
rect 13971 3408 14029 3414
rect 13971 3405 13983 3408
rect 12193 3377 13983 3405
rect 12193 3374 12205 3377
rect 12147 3368 12205 3374
rect 13971 3374 13983 3377
rect 14017 3374 14029 3408
rect 13971 3368 14029 3374
rect 14547 3408 14605 3414
rect 14547 3374 14559 3408
rect 14593 3405 14605 3408
rect 16467 3408 16525 3414
rect 16467 3405 16479 3408
rect 14593 3377 16479 3405
rect 14593 3374 14605 3377
rect 14547 3368 14605 3374
rect 16467 3374 16479 3377
rect 16513 3374 16525 3408
rect 16467 3368 16525 3374
rect 17139 3408 17197 3414
rect 17139 3374 17151 3408
rect 17185 3405 17197 3408
rect 18963 3408 19021 3414
rect 18963 3405 18975 3408
rect 17185 3377 18975 3405
rect 17185 3374 17197 3377
rect 17139 3368 17197 3374
rect 18963 3374 18975 3377
rect 19009 3374 19021 3408
rect 18963 3368 19021 3374
rect 19635 3408 19693 3414
rect 19635 3374 19647 3408
rect 19681 3405 19693 3408
rect 21459 3408 21517 3414
rect 21459 3405 21471 3408
rect 19681 3377 21471 3405
rect 19681 3374 19693 3377
rect 19635 3368 19693 3374
rect 21459 3374 21471 3377
rect 21505 3374 21517 3408
rect 21459 3368 21517 3374
rect 7201 3303 8350 3331
rect 8403 3334 8461 3340
rect 7201 3300 7213 3303
rect 7155 3294 7213 3300
rect 8403 3300 8415 3334
rect 8449 3331 8461 3334
rect 10227 3334 10285 3340
rect 10227 3331 10239 3334
rect 8449 3303 10239 3331
rect 8449 3300 8461 3303
rect 8403 3294 8461 3300
rect 10227 3300 10239 3303
rect 10273 3300 10285 3334
rect 10227 3294 10285 3300
rect 10899 3334 10957 3340
rect 10899 3300 10911 3334
rect 10945 3331 10957 3334
rect 12723 3334 12781 3340
rect 12723 3331 12735 3334
rect 10945 3303 12735 3331
rect 10945 3300 10957 3303
rect 10899 3294 10957 3300
rect 12723 3300 12735 3303
rect 12769 3300 12781 3334
rect 12723 3294 12781 3300
rect 13395 3334 13453 3340
rect 13395 3300 13407 3334
rect 13441 3331 13453 3334
rect 15219 3334 15277 3340
rect 15219 3331 15231 3334
rect 13441 3303 15231 3331
rect 13441 3300 13453 3303
rect 13395 3294 13453 3300
rect 15219 3300 15231 3303
rect 15265 3300 15277 3334
rect 15219 3294 15277 3300
rect 15891 3334 15949 3340
rect 15891 3300 15903 3334
rect 15937 3331 15949 3334
rect 17715 3334 17773 3340
rect 17715 3331 17727 3334
rect 15937 3303 17727 3331
rect 15937 3300 15949 3303
rect 15891 3294 15949 3300
rect 17715 3300 17727 3303
rect 17761 3300 17773 3334
rect 17715 3294 17773 3300
rect 18387 3334 18445 3340
rect 18387 3300 18399 3334
rect 18433 3331 18445 3334
rect 20211 3334 20269 3340
rect 20211 3331 20223 3334
rect 18433 3303 20223 3331
rect 18433 3300 18445 3303
rect 18387 3294 18445 3300
rect 20211 3300 20223 3303
rect 20257 3300 20269 3334
rect 20211 3294 20269 3300
rect 20883 3334 20941 3340
rect 20883 3300 20895 3334
rect 20929 3300 20941 3334
rect 20883 3294 20941 3300
rect 22131 3334 22189 3340
rect 22131 3300 22143 3334
rect 22177 3331 22189 3334
rect 22608 3331 22614 3343
rect 22177 3303 22614 3331
rect 22177 3300 22189 3303
rect 22131 3294 22189 3300
rect 4674 3257 4702 3294
rect 6483 3260 6541 3266
rect 6483 3257 6495 3260
rect 4674 3229 6495 3257
rect 6483 3226 6495 3229
rect 6529 3226 6541 3260
rect 20898 3257 20926 3294
rect 22608 3291 22614 3303
rect 22666 3291 22672 3343
rect 22707 3260 22765 3266
rect 22707 3257 22719 3260
rect 20898 3229 22719 3257
rect 6483 3220 6541 3226
rect 22707 3226 22719 3229
rect 22753 3226 22765 3260
rect 22707 3220 22765 3226
rect 1952 3084 23264 3106
rect 1952 3032 4494 3084
rect 4546 3032 4558 3084
rect 4610 3032 4622 3084
rect 4674 3032 4686 3084
rect 4738 3032 9822 3084
rect 9874 3032 9886 3084
rect 9938 3032 9950 3084
rect 10002 3032 10014 3084
rect 10066 3032 15150 3084
rect 15202 3032 15214 3084
rect 15266 3032 15278 3084
rect 15330 3032 15342 3084
rect 15394 3032 20478 3084
rect 20530 3032 20542 3084
rect 20594 3032 20606 3084
rect 20658 3032 20670 3084
rect 20722 3032 23264 3084
rect 1952 3010 23264 3032
rect 22608 2773 22614 2825
rect 22666 2813 22672 2825
rect 22707 2816 22765 2822
rect 22707 2813 22719 2816
rect 22666 2785 22719 2813
rect 22666 2773 22672 2785
rect 22707 2782 22719 2785
rect 22753 2782 22765 2816
rect 22707 2776 22765 2782
rect 3411 2742 3469 2748
rect 3411 2708 3423 2742
rect 3457 2739 3469 2742
rect 3888 2739 3894 2751
rect 3457 2711 3894 2739
rect 3457 2708 3469 2711
rect 3411 2702 3469 2708
rect 3888 2699 3894 2711
rect 3946 2699 3952 2751
rect 3987 2742 4045 2748
rect 3987 2708 3999 2742
rect 4033 2739 4045 2742
rect 4563 2742 4621 2748
rect 4563 2739 4575 2742
rect 4033 2711 4575 2739
rect 4033 2708 4045 2711
rect 3987 2702 4045 2708
rect 4563 2708 4575 2711
rect 4609 2708 4621 2742
rect 4563 2702 4621 2708
rect 5235 2742 5293 2748
rect 5235 2708 5247 2742
rect 5281 2739 5293 2742
rect 5811 2742 5869 2748
rect 5811 2739 5823 2742
rect 5281 2711 5823 2739
rect 5281 2708 5293 2711
rect 5235 2702 5293 2708
rect 5811 2708 5823 2711
rect 5857 2708 5869 2742
rect 5811 2702 5869 2708
rect 6483 2742 6541 2748
rect 6483 2708 6495 2742
rect 6529 2739 6541 2742
rect 7059 2742 7117 2748
rect 7059 2739 7071 2742
rect 6529 2711 7071 2739
rect 6529 2708 6541 2711
rect 6483 2702 6541 2708
rect 7059 2708 7071 2711
rect 7105 2708 7117 2742
rect 7059 2702 7117 2708
rect 7731 2742 7789 2748
rect 7731 2708 7743 2742
rect 7777 2739 7789 2742
rect 8307 2742 8365 2748
rect 8307 2739 8319 2742
rect 7777 2711 8319 2739
rect 7777 2708 7789 2711
rect 7731 2702 7789 2708
rect 8307 2708 8319 2711
rect 8353 2708 8365 2742
rect 8307 2702 8365 2708
rect 8979 2742 9037 2748
rect 8979 2708 8991 2742
rect 9025 2739 9037 2742
rect 9555 2742 9613 2748
rect 9555 2739 9567 2742
rect 9025 2711 9567 2739
rect 9025 2708 9037 2711
rect 8979 2702 9037 2708
rect 9555 2708 9567 2711
rect 9601 2708 9613 2742
rect 9555 2702 9613 2708
rect 10227 2742 10285 2748
rect 10227 2708 10239 2742
rect 10273 2739 10285 2742
rect 10803 2742 10861 2748
rect 10803 2739 10815 2742
rect 10273 2711 10815 2739
rect 10273 2708 10285 2711
rect 10227 2702 10285 2708
rect 10803 2708 10815 2711
rect 10849 2708 10861 2742
rect 10803 2702 10861 2708
rect 11475 2742 11533 2748
rect 11475 2708 11487 2742
rect 11521 2739 11533 2742
rect 12051 2742 12109 2748
rect 12051 2739 12063 2742
rect 11521 2711 12063 2739
rect 11521 2708 11533 2711
rect 11475 2702 11533 2708
rect 12051 2708 12063 2711
rect 12097 2708 12109 2742
rect 12051 2702 12109 2708
rect 12723 2742 12781 2748
rect 12723 2708 12735 2742
rect 12769 2739 12781 2742
rect 13299 2742 13357 2748
rect 13299 2739 13311 2742
rect 12769 2711 13311 2739
rect 12769 2708 12781 2711
rect 12723 2702 12781 2708
rect 13299 2708 13311 2711
rect 13345 2708 13357 2742
rect 13299 2702 13357 2708
rect 13971 2742 14029 2748
rect 13971 2708 13983 2742
rect 14017 2739 14029 2742
rect 14547 2742 14605 2748
rect 14547 2739 14559 2742
rect 14017 2711 14559 2739
rect 14017 2708 14029 2711
rect 13971 2702 14029 2708
rect 14547 2708 14559 2711
rect 14593 2708 14605 2742
rect 14547 2702 14605 2708
rect 15219 2742 15277 2748
rect 15219 2708 15231 2742
rect 15265 2739 15277 2742
rect 15795 2742 15853 2748
rect 15795 2739 15807 2742
rect 15265 2711 15807 2739
rect 15265 2708 15277 2711
rect 15219 2702 15277 2708
rect 15795 2708 15807 2711
rect 15841 2708 15853 2742
rect 15795 2702 15853 2708
rect 16467 2742 16525 2748
rect 16467 2708 16479 2742
rect 16513 2739 16525 2742
rect 17043 2742 17101 2748
rect 17043 2739 17055 2742
rect 16513 2711 17055 2739
rect 16513 2708 16525 2711
rect 16467 2702 16525 2708
rect 17043 2708 17055 2711
rect 17089 2708 17101 2742
rect 17043 2702 17101 2708
rect 17715 2742 17773 2748
rect 17715 2708 17727 2742
rect 17761 2739 17773 2742
rect 18291 2742 18349 2748
rect 18291 2739 18303 2742
rect 17761 2711 18303 2739
rect 17761 2708 17773 2711
rect 17715 2702 17773 2708
rect 18291 2708 18303 2711
rect 18337 2708 18349 2742
rect 18291 2702 18349 2708
rect 18963 2742 19021 2748
rect 18963 2708 18975 2742
rect 19009 2739 19021 2742
rect 19539 2742 19597 2748
rect 19539 2739 19551 2742
rect 19009 2711 19551 2739
rect 19009 2708 19021 2711
rect 18963 2702 19021 2708
rect 19539 2708 19551 2711
rect 19585 2708 19597 2742
rect 19539 2702 19597 2708
rect 20211 2742 20269 2748
rect 20211 2708 20223 2742
rect 20257 2739 20269 2742
rect 20787 2742 20845 2748
rect 20787 2739 20799 2742
rect 20257 2711 20799 2739
rect 20257 2708 20269 2711
rect 20211 2702 20269 2708
rect 20787 2708 20799 2711
rect 20833 2708 20845 2742
rect 20787 2702 20845 2708
rect 21459 2742 21517 2748
rect 21459 2708 21471 2742
rect 21505 2739 21517 2742
rect 22035 2742 22093 2748
rect 22035 2739 22047 2742
rect 21505 2711 22047 2739
rect 21505 2708 21517 2711
rect 21459 2702 21517 2708
rect 22035 2708 22047 2711
rect 22081 2708 22093 2742
rect 22035 2702 22093 2708
rect 1952 2418 23264 2440
rect 1952 2366 7158 2418
rect 7210 2366 7222 2418
rect 7274 2366 7286 2418
rect 7338 2366 7350 2418
rect 7402 2366 12486 2418
rect 12538 2366 12550 2418
rect 12602 2366 12614 2418
rect 12666 2366 12678 2418
rect 12730 2366 17814 2418
rect 17866 2366 17878 2418
rect 17930 2366 17942 2418
rect 17994 2366 18006 2418
rect 18058 2366 23264 2418
rect 1952 2344 23264 2366
rect 3888 2255 3894 2307
rect 3946 2295 3952 2307
rect 3987 2298 4045 2304
rect 3987 2295 3999 2298
rect 3946 2267 3999 2295
rect 3946 2255 3952 2267
rect 3987 2264 3999 2267
rect 4033 2264 4045 2298
rect 3987 2258 4045 2264
rect 11970 2045 12766 2073
rect 3315 2002 3373 2008
rect 3315 1968 3327 2002
rect 3361 1968 3373 2002
rect 3315 1962 3373 1968
rect 4659 2002 4717 2008
rect 4659 1968 4671 2002
rect 4705 1968 4717 2002
rect 4659 1962 4717 1968
rect 5907 2002 5965 2008
rect 5907 1968 5919 2002
rect 5953 1999 5965 2002
rect 7155 2002 7213 2008
rect 5953 1971 6814 1999
rect 5953 1968 5965 1971
rect 5907 1962 5965 1968
rect 3330 1851 3358 1962
rect 4674 1925 4702 1962
rect 6483 1928 6541 1934
rect 6483 1925 6495 1928
rect 4674 1897 6495 1925
rect 6483 1894 6495 1897
rect 6529 1894 6541 1928
rect 6786 1925 6814 1971
rect 7155 1968 7167 2002
rect 7201 1999 7213 2002
rect 8403 2002 8461 2008
rect 7201 1971 8350 1999
rect 7201 1968 7213 1971
rect 7155 1962 7213 1968
rect 7731 1928 7789 1934
rect 7731 1925 7743 1928
rect 6786 1897 7743 1925
rect 6483 1888 6541 1894
rect 7731 1894 7743 1897
rect 7777 1894 7789 1928
rect 7731 1888 7789 1894
rect 5235 1854 5293 1860
rect 5235 1851 5247 1854
rect 3330 1823 5247 1851
rect 5235 1820 5247 1823
rect 5281 1820 5293 1854
rect 8322 1851 8350 1971
rect 8403 1968 8415 2002
rect 8449 1968 8461 2002
rect 8403 1962 8461 1968
rect 9651 2002 9709 2008
rect 9651 1968 9663 2002
rect 9697 1999 9709 2002
rect 10899 2002 10957 2008
rect 9697 1971 10558 1999
rect 9697 1968 9709 1971
rect 9651 1962 9709 1968
rect 8418 1925 8446 1962
rect 10227 1928 10285 1934
rect 10227 1925 10239 1928
rect 8418 1897 10239 1925
rect 10227 1894 10239 1897
rect 10273 1894 10285 1928
rect 10227 1888 10285 1894
rect 8979 1854 9037 1860
rect 8979 1851 8991 1854
rect 8322 1823 8991 1851
rect 5235 1814 5293 1820
rect 8979 1820 8991 1823
rect 9025 1820 9037 1854
rect 10530 1851 10558 1971
rect 10899 1968 10911 2002
rect 10945 1999 10957 2002
rect 11970 1999 11998 2045
rect 12738 2008 12766 2045
rect 14466 2045 15262 2073
rect 10945 1971 11998 1999
rect 12051 2002 12109 2008
rect 10945 1968 10957 1971
rect 10899 1962 10957 1968
rect 12051 1968 12063 2002
rect 12097 1968 12109 2002
rect 12051 1962 12109 1968
rect 12723 2002 12781 2008
rect 12723 1968 12735 2002
rect 12769 1968 12781 2002
rect 12723 1962 12781 1968
rect 13395 2002 13453 2008
rect 13395 1968 13407 2002
rect 13441 1999 13453 2002
rect 14466 1999 14494 2045
rect 15234 2008 15262 2045
rect 13441 1971 14494 1999
rect 14547 2002 14605 2008
rect 13441 1968 13453 1971
rect 13395 1962 13453 1968
rect 14547 1968 14559 2002
rect 14593 1968 14605 2002
rect 14547 1962 14605 1968
rect 15219 2002 15277 2008
rect 15219 1968 15231 2002
rect 15265 1968 15277 2002
rect 15219 1962 15277 1968
rect 15891 2002 15949 2008
rect 15891 1968 15903 2002
rect 15937 1968 15949 2002
rect 15891 1962 15949 1968
rect 17139 2002 17197 2008
rect 17139 1968 17151 2002
rect 17185 1999 17197 2002
rect 18387 2002 18445 2008
rect 17185 1971 18046 1999
rect 17185 1968 17197 1971
rect 17139 1962 17197 1968
rect 11475 1854 11533 1860
rect 11475 1851 11487 1854
rect 10530 1823 11487 1851
rect 8979 1814 9037 1820
rect 11475 1820 11487 1823
rect 11521 1820 11533 1854
rect 12066 1851 12094 1962
rect 13971 1854 14029 1860
rect 13971 1851 13983 1854
rect 12066 1823 13983 1851
rect 11475 1814 11533 1820
rect 13971 1820 13983 1823
rect 14017 1820 14029 1854
rect 14562 1851 14590 1962
rect 15906 1925 15934 1962
rect 17715 1928 17773 1934
rect 17715 1925 17727 1928
rect 15906 1897 17727 1925
rect 17715 1894 17727 1897
rect 17761 1894 17773 1928
rect 17715 1888 17773 1894
rect 16467 1854 16525 1860
rect 16467 1851 16479 1854
rect 14562 1823 16479 1851
rect 13971 1814 14029 1820
rect 16467 1820 16479 1823
rect 16513 1820 16525 1854
rect 18018 1851 18046 1971
rect 18387 1968 18399 2002
rect 18433 1968 18445 2002
rect 18387 1962 18445 1968
rect 19635 2002 19693 2008
rect 19635 1968 19647 2002
rect 19681 1999 19693 2002
rect 20883 2002 20941 2008
rect 19681 1971 20350 1999
rect 19681 1968 19693 1971
rect 19635 1962 19693 1968
rect 18402 1925 18430 1962
rect 20211 1928 20269 1934
rect 20211 1925 20223 1928
rect 18402 1897 20223 1925
rect 20211 1894 20223 1897
rect 20257 1894 20269 1928
rect 20211 1888 20269 1894
rect 18963 1854 19021 1860
rect 18963 1851 18975 1854
rect 18018 1823 18975 1851
rect 16467 1814 16525 1820
rect 18963 1820 18975 1823
rect 19009 1820 19021 1854
rect 20322 1851 20350 1971
rect 20883 1968 20895 2002
rect 20929 1968 20941 2002
rect 22128 1999 22134 2011
rect 22089 1971 22134 1999
rect 20883 1962 20941 1968
rect 20898 1925 20926 1962
rect 22128 1959 22134 1971
rect 22186 1959 22192 2011
rect 22707 1928 22765 1934
rect 22707 1925 22719 1928
rect 20898 1897 22719 1925
rect 22707 1894 22719 1897
rect 22753 1894 22765 1928
rect 22707 1888 22765 1894
rect 21459 1854 21517 1860
rect 21459 1851 21471 1854
rect 20322 1823 21471 1851
rect 18963 1814 19021 1820
rect 21459 1820 21471 1823
rect 21505 1820 21517 1854
rect 21459 1814 21517 1820
rect 1952 1752 23264 1774
rect 1952 1700 4494 1752
rect 4546 1700 4558 1752
rect 4610 1700 4622 1752
rect 4674 1700 4686 1752
rect 4738 1700 9822 1752
rect 9874 1700 9886 1752
rect 9938 1700 9950 1752
rect 10002 1700 10014 1752
rect 10066 1700 15150 1752
rect 15202 1700 15214 1752
rect 15266 1700 15278 1752
rect 15330 1700 15342 1752
rect 15394 1700 20478 1752
rect 20530 1700 20542 1752
rect 20594 1700 20606 1752
rect 20658 1700 20670 1752
rect 20722 1700 23264 1752
rect 1952 1678 23264 1700
rect 22128 1589 22134 1641
rect 22186 1629 22192 1641
rect 22707 1632 22765 1638
rect 22707 1629 22719 1632
rect 22186 1601 22719 1629
rect 22186 1589 22192 1601
rect 22707 1598 22719 1601
rect 22753 1598 22765 1632
rect 22707 1592 22765 1598
rect 2352 1367 2358 1419
rect 2410 1407 2416 1419
rect 3024 1407 3030 1419
rect 2410 1379 3030 1407
rect 2410 1367 2416 1379
rect 3024 1367 3030 1379
rect 3082 1407 3088 1419
rect 3315 1410 3373 1416
rect 3315 1407 3327 1410
rect 3082 1379 3327 1407
rect 3082 1367 3088 1379
rect 3315 1376 3327 1379
rect 3361 1376 3373 1410
rect 3315 1370 3373 1376
rect 3987 1410 4045 1416
rect 3987 1376 3999 1410
rect 4033 1407 4045 1410
rect 4563 1410 4621 1416
rect 4563 1407 4575 1410
rect 4033 1379 4575 1407
rect 4033 1376 4045 1379
rect 3987 1370 4045 1376
rect 4563 1376 4575 1379
rect 4609 1376 4621 1410
rect 4563 1370 4621 1376
rect 5235 1410 5293 1416
rect 5235 1376 5247 1410
rect 5281 1407 5293 1410
rect 5811 1410 5869 1416
rect 5811 1407 5823 1410
rect 5281 1379 5823 1407
rect 5281 1376 5293 1379
rect 5235 1370 5293 1376
rect 5811 1376 5823 1379
rect 5857 1376 5869 1410
rect 5811 1370 5869 1376
rect 6483 1410 6541 1416
rect 6483 1376 6495 1410
rect 6529 1407 6541 1410
rect 7059 1410 7117 1416
rect 7059 1407 7071 1410
rect 6529 1379 7071 1407
rect 6529 1376 6541 1379
rect 6483 1370 6541 1376
rect 7059 1376 7071 1379
rect 7105 1376 7117 1410
rect 7059 1370 7117 1376
rect 7731 1410 7789 1416
rect 7731 1376 7743 1410
rect 7777 1407 7789 1410
rect 8307 1410 8365 1416
rect 8307 1407 8319 1410
rect 7777 1379 8319 1407
rect 7777 1376 7789 1379
rect 7731 1370 7789 1376
rect 8307 1376 8319 1379
rect 8353 1376 8365 1410
rect 8307 1370 8365 1376
rect 8979 1410 9037 1416
rect 8979 1376 8991 1410
rect 9025 1407 9037 1410
rect 9555 1410 9613 1416
rect 9555 1407 9567 1410
rect 9025 1379 9567 1407
rect 9025 1376 9037 1379
rect 8979 1370 9037 1376
rect 9555 1376 9567 1379
rect 9601 1376 9613 1410
rect 9555 1370 9613 1376
rect 10227 1410 10285 1416
rect 10227 1376 10239 1410
rect 10273 1407 10285 1410
rect 10803 1410 10861 1416
rect 10803 1407 10815 1410
rect 10273 1379 10815 1407
rect 10273 1376 10285 1379
rect 10227 1370 10285 1376
rect 10803 1376 10815 1379
rect 10849 1376 10861 1410
rect 10803 1370 10861 1376
rect 11475 1410 11533 1416
rect 11475 1376 11487 1410
rect 11521 1407 11533 1410
rect 12051 1410 12109 1416
rect 12051 1407 12063 1410
rect 11521 1379 12063 1407
rect 11521 1376 11533 1379
rect 11475 1370 11533 1376
rect 12051 1376 12063 1379
rect 12097 1376 12109 1410
rect 12051 1370 12109 1376
rect 12723 1410 12781 1416
rect 12723 1376 12735 1410
rect 12769 1407 12781 1410
rect 13299 1410 13357 1416
rect 13299 1407 13311 1410
rect 12769 1379 13311 1407
rect 12769 1376 12781 1379
rect 12723 1370 12781 1376
rect 13299 1376 13311 1379
rect 13345 1376 13357 1410
rect 13299 1370 13357 1376
rect 13971 1410 14029 1416
rect 13971 1376 13983 1410
rect 14017 1407 14029 1410
rect 14547 1410 14605 1416
rect 14547 1407 14559 1410
rect 14017 1379 14559 1407
rect 14017 1376 14029 1379
rect 13971 1370 14029 1376
rect 14547 1376 14559 1379
rect 14593 1376 14605 1410
rect 14547 1370 14605 1376
rect 15219 1410 15277 1416
rect 15219 1376 15231 1410
rect 15265 1407 15277 1410
rect 15795 1410 15853 1416
rect 15795 1407 15807 1410
rect 15265 1379 15807 1407
rect 15265 1376 15277 1379
rect 15219 1370 15277 1376
rect 15795 1376 15807 1379
rect 15841 1376 15853 1410
rect 15795 1370 15853 1376
rect 16467 1410 16525 1416
rect 16467 1376 16479 1410
rect 16513 1407 16525 1410
rect 17043 1410 17101 1416
rect 17043 1407 17055 1410
rect 16513 1379 17055 1407
rect 16513 1376 16525 1379
rect 16467 1370 16525 1376
rect 17043 1376 17055 1379
rect 17089 1376 17101 1410
rect 17043 1370 17101 1376
rect 17715 1410 17773 1416
rect 17715 1376 17727 1410
rect 17761 1407 17773 1410
rect 18291 1410 18349 1416
rect 18291 1407 18303 1410
rect 17761 1379 18303 1407
rect 17761 1376 17773 1379
rect 17715 1370 17773 1376
rect 18291 1376 18303 1379
rect 18337 1376 18349 1410
rect 18291 1370 18349 1376
rect 18963 1410 19021 1416
rect 18963 1376 18975 1410
rect 19009 1407 19021 1410
rect 19539 1410 19597 1416
rect 19539 1407 19551 1410
rect 19009 1379 19551 1407
rect 19009 1376 19021 1379
rect 18963 1370 19021 1376
rect 19539 1376 19551 1379
rect 19585 1376 19597 1410
rect 19539 1370 19597 1376
rect 20211 1410 20269 1416
rect 20211 1376 20223 1410
rect 20257 1407 20269 1410
rect 20787 1410 20845 1416
rect 20787 1407 20799 1410
rect 20257 1379 20799 1407
rect 20257 1376 20269 1379
rect 20211 1370 20269 1376
rect 20787 1376 20799 1379
rect 20833 1376 20845 1410
rect 20787 1370 20845 1376
rect 21459 1410 21517 1416
rect 21459 1376 21471 1410
rect 21505 1407 21517 1410
rect 22035 1410 22093 1416
rect 22035 1407 22047 1410
rect 21505 1379 22047 1407
rect 21505 1376 21517 1379
rect 21459 1370 21517 1376
rect 22035 1376 22047 1379
rect 22081 1376 22093 1410
rect 22035 1370 22093 1376
rect 1952 1086 23264 1108
rect 1952 1034 7158 1086
rect 7210 1034 7222 1086
rect 7274 1034 7286 1086
rect 7338 1034 7350 1086
rect 7402 1034 12486 1086
rect 12538 1034 12550 1086
rect 12602 1034 12614 1086
rect 12666 1034 12678 1086
rect 12730 1034 17814 1086
rect 17866 1034 17878 1086
rect 17930 1034 17942 1086
rect 17994 1034 18006 1086
rect 18058 1034 23264 1086
rect 1952 1012 23264 1034
<< via1 >>
rect 4494 27008 4546 27060
rect 4558 27008 4610 27060
rect 4622 27008 4674 27060
rect 4686 27008 4738 27060
rect 9822 27008 9874 27060
rect 9886 27008 9938 27060
rect 9950 27008 10002 27060
rect 10014 27008 10066 27060
rect 15150 27008 15202 27060
rect 15214 27008 15266 27060
rect 15278 27008 15330 27060
rect 15342 27008 15394 27060
rect 20478 27008 20530 27060
rect 20542 27008 20594 27060
rect 20606 27008 20658 27060
rect 20670 27008 20722 27060
rect 2742 26940 2794 26949
rect 2742 26906 2751 26940
rect 2751 26906 2785 26940
rect 2785 26906 2794 26940
rect 2742 26897 2794 26906
rect 2742 26749 2794 26801
rect 2358 26601 2410 26653
rect 7158 26342 7210 26394
rect 7222 26342 7274 26394
rect 7286 26342 7338 26394
rect 7350 26342 7402 26394
rect 12486 26342 12538 26394
rect 12550 26342 12602 26394
rect 12614 26342 12666 26394
rect 12678 26342 12730 26394
rect 17814 26342 17866 26394
rect 17878 26342 17930 26394
rect 17942 26342 17994 26394
rect 18006 26342 18058 26394
rect 2742 26274 2794 26283
rect 2742 26240 2751 26274
rect 2751 26240 2785 26274
rect 2785 26240 2794 26274
rect 2742 26231 2794 26240
rect 2454 26009 2506 26061
rect 2358 25978 2410 25987
rect 2358 25944 2367 25978
rect 2367 25944 2401 25978
rect 2401 25944 2410 25978
rect 2358 25935 2410 25944
rect 3894 25935 3946 25987
rect 4494 25676 4546 25728
rect 4558 25676 4610 25728
rect 4622 25676 4674 25728
rect 4686 25676 4738 25728
rect 9822 25676 9874 25728
rect 9886 25676 9938 25728
rect 9950 25676 10002 25728
rect 10014 25676 10066 25728
rect 15150 25676 15202 25728
rect 15214 25676 15266 25728
rect 15278 25676 15330 25728
rect 15342 25676 15394 25728
rect 20478 25676 20530 25728
rect 20542 25676 20594 25728
rect 20606 25676 20658 25728
rect 20670 25676 20722 25728
rect 3894 25565 3946 25617
rect 2358 25417 2410 25469
rect 2742 25417 2794 25469
rect 7158 25010 7210 25062
rect 7222 25010 7274 25062
rect 7286 25010 7338 25062
rect 7350 25010 7402 25062
rect 12486 25010 12538 25062
rect 12550 25010 12602 25062
rect 12614 25010 12666 25062
rect 12678 25010 12730 25062
rect 17814 25010 17866 25062
rect 17878 25010 17930 25062
rect 17942 25010 17994 25062
rect 18006 25010 18058 25062
rect 2742 24942 2794 24951
rect 2742 24908 2751 24942
rect 2751 24908 2785 24942
rect 2785 24908 2794 24942
rect 2742 24899 2794 24908
rect 2070 24720 2122 24729
rect 2070 24686 2079 24720
rect 2079 24686 2113 24720
rect 2113 24686 2122 24720
rect 2070 24677 2122 24686
rect 2742 24603 2794 24655
rect 5142 24603 5194 24655
rect 4494 24344 4546 24396
rect 4558 24344 4610 24396
rect 4622 24344 4674 24396
rect 4686 24344 4738 24396
rect 9822 24344 9874 24396
rect 9886 24344 9938 24396
rect 9950 24344 10002 24396
rect 10014 24344 10066 24396
rect 15150 24344 15202 24396
rect 15214 24344 15266 24396
rect 15278 24344 15330 24396
rect 15342 24344 15394 24396
rect 20478 24344 20530 24396
rect 20542 24344 20594 24396
rect 20606 24344 20658 24396
rect 20670 24344 20722 24396
rect 5142 24233 5194 24285
rect 2742 24011 2794 24063
rect 7158 23678 7210 23730
rect 7222 23678 7274 23730
rect 7286 23678 7338 23730
rect 7350 23678 7402 23730
rect 12486 23678 12538 23730
rect 12550 23678 12602 23730
rect 12614 23678 12666 23730
rect 12678 23678 12730 23730
rect 17814 23678 17866 23730
rect 17878 23678 17930 23730
rect 17942 23678 17994 23730
rect 18006 23678 18058 23730
rect 2742 23536 2794 23545
rect 2742 23502 2751 23536
rect 2751 23502 2785 23536
rect 2785 23502 2794 23536
rect 2742 23493 2794 23502
rect 2070 23388 2122 23397
rect 2070 23354 2079 23388
rect 2079 23354 2113 23388
rect 2113 23354 2122 23388
rect 2070 23345 2122 23354
rect 2742 23271 2794 23323
rect 7734 23197 7786 23249
rect 4494 23012 4546 23064
rect 4558 23012 4610 23064
rect 4622 23012 4674 23064
rect 4686 23012 4738 23064
rect 9822 23012 9874 23064
rect 9886 23012 9938 23064
rect 9950 23012 10002 23064
rect 10014 23012 10066 23064
rect 15150 23012 15202 23064
rect 15214 23012 15266 23064
rect 15278 23012 15330 23064
rect 15342 23012 15394 23064
rect 20478 23012 20530 23064
rect 20542 23012 20594 23064
rect 20606 23012 20658 23064
rect 20670 23012 20722 23064
rect 2742 22679 2794 22731
rect 7734 22722 7786 22731
rect 7734 22688 7743 22722
rect 7743 22688 7777 22722
rect 7777 22688 7786 22722
rect 7734 22679 7786 22688
rect 7158 22346 7210 22398
rect 7222 22346 7274 22398
rect 7286 22346 7338 22398
rect 7350 22346 7402 22398
rect 12486 22346 12538 22398
rect 12550 22346 12602 22398
rect 12614 22346 12666 22398
rect 12678 22346 12730 22398
rect 17814 22346 17866 22398
rect 17878 22346 17930 22398
rect 17942 22346 17994 22398
rect 18006 22346 18058 22398
rect 2742 22278 2794 22287
rect 2742 22244 2751 22278
rect 2751 22244 2785 22278
rect 2785 22244 2794 22278
rect 2742 22235 2794 22244
rect 2070 22056 2122 22065
rect 2070 22022 2079 22056
rect 2079 22022 2113 22056
rect 2113 22022 2122 22056
rect 2070 22013 2122 22022
rect 2742 21939 2794 21991
rect 12630 21939 12682 21991
rect 4494 21680 4546 21732
rect 4558 21680 4610 21732
rect 4622 21680 4674 21732
rect 4686 21680 4738 21732
rect 9822 21680 9874 21732
rect 9886 21680 9938 21732
rect 9950 21680 10002 21732
rect 10014 21680 10066 21732
rect 15150 21680 15202 21732
rect 15214 21680 15266 21732
rect 15278 21680 15330 21732
rect 15342 21680 15394 21732
rect 20478 21680 20530 21732
rect 20542 21680 20594 21732
rect 20606 21680 20658 21732
rect 20670 21680 20722 21732
rect 12630 21569 12682 21621
rect 2742 21347 2794 21399
rect 7158 21014 7210 21066
rect 7222 21014 7274 21066
rect 7286 21014 7338 21066
rect 7350 21014 7402 21066
rect 12486 21014 12538 21066
rect 12550 21014 12602 21066
rect 12614 21014 12666 21066
rect 12678 21014 12730 21066
rect 17814 21014 17866 21066
rect 17878 21014 17930 21066
rect 17942 21014 17994 21066
rect 18006 21014 18058 21066
rect 2742 20946 2794 20955
rect 2742 20912 2751 20946
rect 2751 20912 2785 20946
rect 2785 20912 2794 20946
rect 2742 20903 2794 20912
rect 2454 20681 2506 20733
rect 2358 20650 2410 20659
rect 2358 20616 2367 20650
rect 2367 20616 2401 20650
rect 2401 20616 2410 20650
rect 2358 20607 2410 20616
rect 22614 20607 22666 20659
rect 4494 20348 4546 20400
rect 4558 20348 4610 20400
rect 4622 20348 4674 20400
rect 4686 20348 4738 20400
rect 9822 20348 9874 20400
rect 9886 20348 9938 20400
rect 9950 20348 10002 20400
rect 10014 20348 10066 20400
rect 15150 20348 15202 20400
rect 15214 20348 15266 20400
rect 15278 20348 15330 20400
rect 15342 20348 15394 20400
rect 20478 20348 20530 20400
rect 20542 20348 20594 20400
rect 20606 20348 20658 20400
rect 20670 20348 20722 20400
rect 22614 20237 22666 20289
rect 2358 20089 2410 20141
rect 2742 20089 2794 20141
rect 7158 19682 7210 19734
rect 7222 19682 7274 19734
rect 7286 19682 7338 19734
rect 7350 19682 7402 19734
rect 12486 19682 12538 19734
rect 12550 19682 12602 19734
rect 12614 19682 12666 19734
rect 12678 19682 12730 19734
rect 17814 19682 17866 19734
rect 17878 19682 17930 19734
rect 17942 19682 17994 19734
rect 18006 19682 18058 19734
rect 2742 19614 2794 19623
rect 2742 19580 2751 19614
rect 2751 19580 2785 19614
rect 2785 19580 2794 19614
rect 2742 19571 2794 19580
rect 2070 19392 2122 19401
rect 2070 19358 2079 19392
rect 2079 19358 2113 19392
rect 2113 19358 2122 19392
rect 2070 19349 2122 19358
rect 2358 19318 2410 19327
rect 2358 19284 2367 19318
rect 2367 19284 2401 19318
rect 2401 19284 2410 19318
rect 2358 19275 2410 19284
rect 22614 19275 22666 19327
rect 4494 19016 4546 19068
rect 4558 19016 4610 19068
rect 4622 19016 4674 19068
rect 4686 19016 4738 19068
rect 9822 19016 9874 19068
rect 9886 19016 9938 19068
rect 9950 19016 10002 19068
rect 10014 19016 10066 19068
rect 15150 19016 15202 19068
rect 15214 19016 15266 19068
rect 15278 19016 15330 19068
rect 15342 19016 15394 19068
rect 20478 19016 20530 19068
rect 20542 19016 20594 19068
rect 20606 19016 20658 19068
rect 20670 19016 20722 19068
rect 22614 18831 22666 18883
rect 3894 18683 3946 18735
rect 7158 18350 7210 18402
rect 7222 18350 7274 18402
rect 7286 18350 7338 18402
rect 7350 18350 7402 18402
rect 12486 18350 12538 18402
rect 12550 18350 12602 18402
rect 12614 18350 12666 18402
rect 12678 18350 12730 18402
rect 17814 18350 17866 18402
rect 17878 18350 17930 18402
rect 17942 18350 17994 18402
rect 18006 18350 18058 18402
rect 3894 18091 3946 18143
rect 22134 17986 22186 17995
rect 22134 17952 22143 17986
rect 22143 17952 22177 17986
rect 22177 17952 22186 17986
rect 22134 17943 22186 17952
rect 4494 17684 4546 17736
rect 4558 17684 4610 17736
rect 4622 17684 4674 17736
rect 4686 17684 4738 17736
rect 9822 17684 9874 17736
rect 9886 17684 9938 17736
rect 9950 17684 10002 17736
rect 10014 17684 10066 17736
rect 15150 17684 15202 17736
rect 15214 17684 15266 17736
rect 15278 17684 15330 17736
rect 15342 17684 15394 17736
rect 20478 17684 20530 17736
rect 20542 17684 20594 17736
rect 20606 17684 20658 17736
rect 20670 17684 20722 17736
rect 22134 17573 22186 17625
rect 2358 17425 2410 17477
rect 7158 17018 7210 17070
rect 7222 17018 7274 17070
rect 7286 17018 7338 17070
rect 7350 17018 7402 17070
rect 12486 17018 12538 17070
rect 12550 17018 12602 17070
rect 12614 17018 12666 17070
rect 12678 17018 12730 17070
rect 17814 17018 17866 17070
rect 17878 17018 17930 17070
rect 17942 17018 17994 17070
rect 18006 17018 18058 17070
rect 2358 16907 2410 16959
rect 2070 16728 2122 16737
rect 2070 16694 2079 16728
rect 2079 16694 2113 16728
rect 2113 16694 2122 16728
rect 2070 16685 2122 16694
rect 2358 16654 2410 16663
rect 2358 16620 2367 16654
rect 2367 16620 2401 16654
rect 2401 16620 2410 16654
rect 2358 16611 2410 16620
rect 22614 16611 22666 16663
rect 4494 16352 4546 16404
rect 4558 16352 4610 16404
rect 4622 16352 4674 16404
rect 4686 16352 4738 16404
rect 9822 16352 9874 16404
rect 9886 16352 9938 16404
rect 9950 16352 10002 16404
rect 10014 16352 10066 16404
rect 15150 16352 15202 16404
rect 15214 16352 15266 16404
rect 15278 16352 15330 16404
rect 15342 16352 15394 16404
rect 20478 16352 20530 16404
rect 20542 16352 20594 16404
rect 20606 16352 20658 16404
rect 20670 16352 20722 16404
rect 22614 16241 22666 16293
rect 3894 16019 3946 16071
rect 7158 15686 7210 15738
rect 7222 15686 7274 15738
rect 7286 15686 7338 15738
rect 7350 15686 7402 15738
rect 12486 15686 12538 15738
rect 12550 15686 12602 15738
rect 12614 15686 12666 15738
rect 12678 15686 12730 15738
rect 17814 15686 17866 15738
rect 17878 15686 17930 15738
rect 17942 15686 17994 15738
rect 18006 15686 18058 15738
rect 3894 15575 3946 15627
rect 22614 15279 22666 15331
rect 4494 15020 4546 15072
rect 4558 15020 4610 15072
rect 4622 15020 4674 15072
rect 4686 15020 4738 15072
rect 9822 15020 9874 15072
rect 9886 15020 9938 15072
rect 9950 15020 10002 15072
rect 10014 15020 10066 15072
rect 15150 15020 15202 15072
rect 15214 15020 15266 15072
rect 15278 15020 15330 15072
rect 15342 15020 15394 15072
rect 20478 15020 20530 15072
rect 20542 15020 20594 15072
rect 20606 15020 20658 15072
rect 20670 15020 20722 15072
rect 22614 14909 22666 14961
rect 3894 14687 3946 14739
rect 7158 14354 7210 14406
rect 7222 14354 7274 14406
rect 7286 14354 7338 14406
rect 7350 14354 7402 14406
rect 12486 14354 12538 14406
rect 12550 14354 12602 14406
rect 12614 14354 12666 14406
rect 12678 14354 12730 14406
rect 17814 14354 17866 14406
rect 17878 14354 17930 14406
rect 17942 14354 17994 14406
rect 18006 14354 18058 14406
rect 3894 14243 3946 14295
rect 22614 13947 22666 13999
rect 4494 13688 4546 13740
rect 4558 13688 4610 13740
rect 4622 13688 4674 13740
rect 4686 13688 4738 13740
rect 9822 13688 9874 13740
rect 9886 13688 9938 13740
rect 9950 13688 10002 13740
rect 10014 13688 10066 13740
rect 15150 13688 15202 13740
rect 15214 13688 15266 13740
rect 15278 13688 15330 13740
rect 15342 13688 15394 13740
rect 20478 13688 20530 13740
rect 20542 13688 20594 13740
rect 20606 13688 20658 13740
rect 20670 13688 20722 13740
rect 22614 13503 22666 13555
rect 3894 13355 3946 13407
rect 7158 13022 7210 13074
rect 7222 13022 7274 13074
rect 7286 13022 7338 13074
rect 7350 13022 7402 13074
rect 12486 13022 12538 13074
rect 12550 13022 12602 13074
rect 12614 13022 12666 13074
rect 12678 13022 12730 13074
rect 17814 13022 17866 13074
rect 17878 13022 17930 13074
rect 17942 13022 17994 13074
rect 18006 13022 18058 13074
rect 3894 12911 3946 12963
rect 22134 12658 22186 12667
rect 22134 12624 22143 12658
rect 22143 12624 22177 12658
rect 22177 12624 22186 12658
rect 22134 12615 22186 12624
rect 4494 12356 4546 12408
rect 4558 12356 4610 12408
rect 4622 12356 4674 12408
rect 4686 12356 4738 12408
rect 9822 12356 9874 12408
rect 9886 12356 9938 12408
rect 9950 12356 10002 12408
rect 10014 12356 10066 12408
rect 15150 12356 15202 12408
rect 15214 12356 15266 12408
rect 15278 12356 15330 12408
rect 15342 12356 15394 12408
rect 20478 12356 20530 12408
rect 20542 12356 20594 12408
rect 20606 12356 20658 12408
rect 20670 12356 20722 12408
rect 22134 12245 22186 12297
rect 2358 12097 2410 12149
rect 7158 11690 7210 11742
rect 7222 11690 7274 11742
rect 7286 11690 7338 11742
rect 7350 11690 7402 11742
rect 12486 11690 12538 11742
rect 12550 11690 12602 11742
rect 12614 11690 12666 11742
rect 12678 11690 12730 11742
rect 17814 11690 17866 11742
rect 17878 11690 17930 11742
rect 17942 11690 17994 11742
rect 18006 11690 18058 11742
rect 2358 11579 2410 11631
rect 2070 11400 2122 11409
rect 2070 11366 2079 11400
rect 2079 11366 2113 11400
rect 2113 11366 2122 11400
rect 2070 11357 2122 11366
rect 2358 11326 2410 11335
rect 2358 11292 2367 11326
rect 2367 11292 2401 11326
rect 2401 11292 2410 11326
rect 2358 11283 2410 11292
rect 22614 11283 22666 11335
rect 4494 11024 4546 11076
rect 4558 11024 4610 11076
rect 4622 11024 4674 11076
rect 4686 11024 4738 11076
rect 9822 11024 9874 11076
rect 9886 11024 9938 11076
rect 9950 11024 10002 11076
rect 10014 11024 10066 11076
rect 15150 11024 15202 11076
rect 15214 11024 15266 11076
rect 15278 11024 15330 11076
rect 15342 11024 15394 11076
rect 20478 11024 20530 11076
rect 20542 11024 20594 11076
rect 20606 11024 20658 11076
rect 20670 11024 20722 11076
rect 22614 10913 22666 10965
rect 3894 10691 3946 10743
rect 7158 10358 7210 10410
rect 7222 10358 7274 10410
rect 7286 10358 7338 10410
rect 7350 10358 7402 10410
rect 12486 10358 12538 10410
rect 12550 10358 12602 10410
rect 12614 10358 12666 10410
rect 12678 10358 12730 10410
rect 17814 10358 17866 10410
rect 17878 10358 17930 10410
rect 17942 10358 17994 10410
rect 18006 10358 18058 10410
rect 3894 10247 3946 10299
rect 22614 9951 22666 10003
rect 4494 9692 4546 9744
rect 4558 9692 4610 9744
rect 4622 9692 4674 9744
rect 4686 9692 4738 9744
rect 9822 9692 9874 9744
rect 9886 9692 9938 9744
rect 9950 9692 10002 9744
rect 10014 9692 10066 9744
rect 15150 9692 15202 9744
rect 15214 9692 15266 9744
rect 15278 9692 15330 9744
rect 15342 9692 15394 9744
rect 20478 9692 20530 9744
rect 20542 9692 20594 9744
rect 20606 9692 20658 9744
rect 20670 9692 20722 9744
rect 22614 9581 22666 9633
rect 3894 9359 3946 9411
rect 7158 9026 7210 9078
rect 7222 9026 7274 9078
rect 7286 9026 7338 9078
rect 7350 9026 7402 9078
rect 12486 9026 12538 9078
rect 12550 9026 12602 9078
rect 12614 9026 12666 9078
rect 12678 9026 12730 9078
rect 17814 9026 17866 9078
rect 17878 9026 17930 9078
rect 17942 9026 17994 9078
rect 18006 9026 18058 9078
rect 3894 8915 3946 8967
rect 22614 8619 22666 8671
rect 4494 8360 4546 8412
rect 4558 8360 4610 8412
rect 4622 8360 4674 8412
rect 4686 8360 4738 8412
rect 9822 8360 9874 8412
rect 9886 8360 9938 8412
rect 9950 8360 10002 8412
rect 10014 8360 10066 8412
rect 15150 8360 15202 8412
rect 15214 8360 15266 8412
rect 15278 8360 15330 8412
rect 15342 8360 15394 8412
rect 20478 8360 20530 8412
rect 20542 8360 20594 8412
rect 20606 8360 20658 8412
rect 20670 8360 20722 8412
rect 22614 8101 22666 8153
rect 3894 8027 3946 8079
rect 7158 7694 7210 7746
rect 7222 7694 7274 7746
rect 7286 7694 7338 7746
rect 7350 7694 7402 7746
rect 12486 7694 12538 7746
rect 12550 7694 12602 7746
rect 12614 7694 12666 7746
rect 12678 7694 12730 7746
rect 17814 7694 17866 7746
rect 17878 7694 17930 7746
rect 17942 7694 17994 7746
rect 18006 7694 18058 7746
rect 3894 7583 3946 7635
rect 22134 7330 22186 7339
rect 22134 7296 22143 7330
rect 22143 7296 22177 7330
rect 22177 7296 22186 7330
rect 22134 7287 22186 7296
rect 4494 7028 4546 7080
rect 4558 7028 4610 7080
rect 4622 7028 4674 7080
rect 4686 7028 4738 7080
rect 9822 7028 9874 7080
rect 9886 7028 9938 7080
rect 9950 7028 10002 7080
rect 10014 7028 10066 7080
rect 15150 7028 15202 7080
rect 15214 7028 15266 7080
rect 15278 7028 15330 7080
rect 15342 7028 15394 7080
rect 20478 7028 20530 7080
rect 20542 7028 20594 7080
rect 20606 7028 20658 7080
rect 20670 7028 20722 7080
rect 22134 6917 22186 6969
rect 3894 6695 3946 6747
rect 7158 6362 7210 6414
rect 7222 6362 7274 6414
rect 7286 6362 7338 6414
rect 7350 6362 7402 6414
rect 12486 6362 12538 6414
rect 12550 6362 12602 6414
rect 12614 6362 12666 6414
rect 12678 6362 12730 6414
rect 17814 6362 17866 6414
rect 17878 6362 17930 6414
rect 17942 6362 17994 6414
rect 18006 6362 18058 6414
rect 3894 6251 3946 6303
rect 22614 5955 22666 6007
rect 4494 5696 4546 5748
rect 4558 5696 4610 5748
rect 4622 5696 4674 5748
rect 4686 5696 4738 5748
rect 9822 5696 9874 5748
rect 9886 5696 9938 5748
rect 9950 5696 10002 5748
rect 10014 5696 10066 5748
rect 15150 5696 15202 5748
rect 15214 5696 15266 5748
rect 15278 5696 15330 5748
rect 15342 5696 15394 5748
rect 20478 5696 20530 5748
rect 20542 5696 20594 5748
rect 20606 5696 20658 5748
rect 20670 5696 20722 5748
rect 22614 5585 22666 5637
rect 3894 5363 3946 5415
rect 7158 5030 7210 5082
rect 7222 5030 7274 5082
rect 7286 5030 7338 5082
rect 7350 5030 7402 5082
rect 12486 5030 12538 5082
rect 12550 5030 12602 5082
rect 12614 5030 12666 5082
rect 12678 5030 12730 5082
rect 17814 5030 17866 5082
rect 17878 5030 17930 5082
rect 17942 5030 17994 5082
rect 18006 5030 18058 5082
rect 3894 4919 3946 4971
rect 22614 4623 22666 4675
rect 4494 4364 4546 4416
rect 4558 4364 4610 4416
rect 4622 4364 4674 4416
rect 4686 4364 4738 4416
rect 9822 4364 9874 4416
rect 9886 4364 9938 4416
rect 9950 4364 10002 4416
rect 10014 4364 10066 4416
rect 15150 4364 15202 4416
rect 15214 4364 15266 4416
rect 15278 4364 15330 4416
rect 15342 4364 15394 4416
rect 20478 4364 20530 4416
rect 20542 4364 20594 4416
rect 20606 4364 20658 4416
rect 20670 4364 20722 4416
rect 22614 4253 22666 4305
rect 3894 4031 3946 4083
rect 7158 3698 7210 3750
rect 7222 3698 7274 3750
rect 7286 3698 7338 3750
rect 7350 3698 7402 3750
rect 12486 3698 12538 3750
rect 12550 3698 12602 3750
rect 12614 3698 12666 3750
rect 12678 3698 12730 3750
rect 17814 3698 17866 3750
rect 17878 3698 17930 3750
rect 17942 3698 17994 3750
rect 18006 3698 18058 3750
rect 3894 3513 3946 3565
rect 22614 3291 22666 3343
rect 4494 3032 4546 3084
rect 4558 3032 4610 3084
rect 4622 3032 4674 3084
rect 4686 3032 4738 3084
rect 9822 3032 9874 3084
rect 9886 3032 9938 3084
rect 9950 3032 10002 3084
rect 10014 3032 10066 3084
rect 15150 3032 15202 3084
rect 15214 3032 15266 3084
rect 15278 3032 15330 3084
rect 15342 3032 15394 3084
rect 20478 3032 20530 3084
rect 20542 3032 20594 3084
rect 20606 3032 20658 3084
rect 20670 3032 20722 3084
rect 22614 2773 22666 2825
rect 3894 2699 3946 2751
rect 7158 2366 7210 2418
rect 7222 2366 7274 2418
rect 7286 2366 7338 2418
rect 7350 2366 7402 2418
rect 12486 2366 12538 2418
rect 12550 2366 12602 2418
rect 12614 2366 12666 2418
rect 12678 2366 12730 2418
rect 17814 2366 17866 2418
rect 17878 2366 17930 2418
rect 17942 2366 17994 2418
rect 18006 2366 18058 2418
rect 3894 2255 3946 2307
rect 22134 2002 22186 2011
rect 22134 1968 22143 2002
rect 22143 1968 22177 2002
rect 22177 1968 22186 2002
rect 22134 1959 22186 1968
rect 4494 1700 4546 1752
rect 4558 1700 4610 1752
rect 4622 1700 4674 1752
rect 4686 1700 4738 1752
rect 9822 1700 9874 1752
rect 9886 1700 9938 1752
rect 9950 1700 10002 1752
rect 10014 1700 10066 1752
rect 15150 1700 15202 1752
rect 15214 1700 15266 1752
rect 15278 1700 15330 1752
rect 15342 1700 15394 1752
rect 20478 1700 20530 1752
rect 20542 1700 20594 1752
rect 20606 1700 20658 1752
rect 20670 1700 20722 1752
rect 22134 1589 22186 1641
rect 2358 1367 2410 1419
rect 3030 1367 3082 1419
rect 7158 1034 7210 1086
rect 7222 1034 7274 1086
rect 7286 1034 7338 1086
rect 7350 1034 7402 1086
rect 12486 1034 12538 1086
rect 12550 1034 12602 1086
rect 12614 1034 12666 1086
rect 12678 1034 12730 1086
rect 17814 1034 17866 1086
rect 17878 1034 17930 1086
rect 17942 1034 17994 1086
rect 18006 1034 18058 1086
<< metal2 >>
rect 2740 27358 2796 27367
rect 2740 27293 2796 27302
rect 2754 26955 2782 27293
rect 4468 27062 4764 27082
rect 4524 27060 4548 27062
rect 4604 27060 4628 27062
rect 4684 27060 4708 27062
rect 4546 27008 4548 27060
rect 4610 27008 4622 27060
rect 4684 27008 4686 27060
rect 4524 27006 4548 27008
rect 4604 27006 4628 27008
rect 4684 27006 4708 27008
rect 4468 26986 4764 27006
rect 9796 27062 10092 27082
rect 9852 27060 9876 27062
rect 9932 27060 9956 27062
rect 10012 27060 10036 27062
rect 9874 27008 9876 27060
rect 9938 27008 9950 27060
rect 10012 27008 10014 27060
rect 9852 27006 9876 27008
rect 9932 27006 9956 27008
rect 10012 27006 10036 27008
rect 9796 26986 10092 27006
rect 15124 27062 15420 27082
rect 15180 27060 15204 27062
rect 15260 27060 15284 27062
rect 15340 27060 15364 27062
rect 15202 27008 15204 27060
rect 15266 27008 15278 27060
rect 15340 27008 15342 27060
rect 15180 27006 15204 27008
rect 15260 27006 15284 27008
rect 15340 27006 15364 27008
rect 15124 26986 15420 27006
rect 20452 27062 20748 27082
rect 20508 27060 20532 27062
rect 20588 27060 20612 27062
rect 20668 27060 20692 27062
rect 20530 27008 20532 27060
rect 20594 27008 20606 27060
rect 20668 27008 20670 27060
rect 20508 27006 20532 27008
rect 20588 27006 20612 27008
rect 20668 27006 20692 27008
rect 20452 26986 20748 27006
rect 2742 26949 2794 26955
rect 2742 26891 2794 26897
rect 2742 26801 2794 26807
rect 2742 26743 2794 26749
rect 2358 26653 2410 26659
rect 2358 26595 2410 26601
rect 2370 26183 2398 26595
rect 2754 26289 2782 26743
rect 7132 26396 7428 26416
rect 7188 26394 7212 26396
rect 7268 26394 7292 26396
rect 7348 26394 7372 26396
rect 7210 26342 7212 26394
rect 7274 26342 7286 26394
rect 7348 26342 7350 26394
rect 7188 26340 7212 26342
rect 7268 26340 7292 26342
rect 7348 26340 7372 26342
rect 7132 26320 7428 26340
rect 12460 26396 12756 26416
rect 12516 26394 12540 26396
rect 12596 26394 12620 26396
rect 12676 26394 12700 26396
rect 12538 26342 12540 26394
rect 12602 26342 12614 26394
rect 12676 26342 12678 26394
rect 12516 26340 12540 26342
rect 12596 26340 12620 26342
rect 12676 26340 12700 26342
rect 12460 26320 12756 26340
rect 17788 26396 18084 26416
rect 17844 26394 17868 26396
rect 17924 26394 17948 26396
rect 18004 26394 18028 26396
rect 17866 26342 17868 26394
rect 17930 26342 17942 26394
rect 18004 26342 18006 26394
rect 17844 26340 17868 26342
rect 17924 26340 17948 26342
rect 18004 26340 18028 26342
rect 17788 26320 18084 26340
rect 2742 26283 2794 26289
rect 2742 26225 2794 26231
rect 2356 26174 2412 26183
rect 2356 26109 2412 26118
rect 2454 26061 2506 26067
rect 2454 26003 2506 26009
rect 2358 25987 2410 25993
rect 2358 25929 2410 25935
rect 2370 25475 2398 25929
rect 2466 25591 2494 26003
rect 3894 25987 3946 25993
rect 3894 25929 3946 25935
rect 3906 25623 3934 25929
rect 4468 25730 4764 25750
rect 4524 25728 4548 25730
rect 4604 25728 4628 25730
rect 4684 25728 4708 25730
rect 4546 25676 4548 25728
rect 4610 25676 4622 25728
rect 4684 25676 4686 25728
rect 4524 25674 4548 25676
rect 4604 25674 4628 25676
rect 4684 25674 4708 25676
rect 4468 25654 4764 25674
rect 9796 25730 10092 25750
rect 9852 25728 9876 25730
rect 9932 25728 9956 25730
rect 10012 25728 10036 25730
rect 9874 25676 9876 25728
rect 9938 25676 9950 25728
rect 10012 25676 10014 25728
rect 9852 25674 9876 25676
rect 9932 25674 9956 25676
rect 10012 25674 10036 25676
rect 9796 25654 10092 25674
rect 15124 25730 15420 25750
rect 15180 25728 15204 25730
rect 15260 25728 15284 25730
rect 15340 25728 15364 25730
rect 15202 25676 15204 25728
rect 15266 25676 15278 25728
rect 15340 25676 15342 25728
rect 15180 25674 15204 25676
rect 15260 25674 15284 25676
rect 15340 25674 15364 25676
rect 15124 25654 15420 25674
rect 20452 25730 20748 25750
rect 20508 25728 20532 25730
rect 20588 25728 20612 25730
rect 20668 25728 20692 25730
rect 20530 25676 20532 25728
rect 20594 25676 20606 25728
rect 20668 25676 20670 25728
rect 20508 25674 20532 25676
rect 20588 25674 20612 25676
rect 20668 25674 20692 25676
rect 20452 25654 20748 25674
rect 3894 25617 3946 25623
rect 2452 25582 2508 25591
rect 3894 25559 3946 25565
rect 2452 25517 2508 25526
rect 2358 25469 2410 25475
rect 2358 25411 2410 25417
rect 2742 25469 2794 25475
rect 2742 25411 2794 25417
rect 2754 24957 2782 25411
rect 7132 25064 7428 25084
rect 7188 25062 7212 25064
rect 7268 25062 7292 25064
rect 7348 25062 7372 25064
rect 7210 25010 7212 25062
rect 7274 25010 7286 25062
rect 7348 25010 7350 25062
rect 7188 25008 7212 25010
rect 7268 25008 7292 25010
rect 7348 25008 7372 25010
rect 7132 24988 7428 25008
rect 12460 25064 12756 25084
rect 12516 25062 12540 25064
rect 12596 25062 12620 25064
rect 12676 25062 12700 25064
rect 12538 25010 12540 25062
rect 12602 25010 12614 25062
rect 12676 25010 12678 25062
rect 12516 25008 12540 25010
rect 12596 25008 12620 25010
rect 12676 25008 12700 25010
rect 12460 24988 12756 25008
rect 17788 25064 18084 25084
rect 17844 25062 17868 25064
rect 17924 25062 17948 25064
rect 18004 25062 18028 25064
rect 17866 25010 17868 25062
rect 17930 25010 17942 25062
rect 18004 25010 18006 25062
rect 17844 25008 17868 25010
rect 17924 25008 17948 25010
rect 18004 25008 18028 25010
rect 17788 24988 18084 25008
rect 2742 24951 2794 24957
rect 2742 24893 2794 24899
rect 2070 24729 2122 24735
rect 2068 24694 2070 24703
rect 2122 24694 2124 24703
rect 2068 24629 2124 24638
rect 2742 24655 2794 24661
rect 2742 24597 2794 24603
rect 5142 24655 5194 24661
rect 5142 24597 5194 24603
rect 2754 24069 2782 24597
rect 4468 24398 4764 24418
rect 4524 24396 4548 24398
rect 4604 24396 4628 24398
rect 4684 24396 4708 24398
rect 4546 24344 4548 24396
rect 4610 24344 4622 24396
rect 4684 24344 4686 24396
rect 4524 24342 4548 24344
rect 4604 24342 4628 24344
rect 4684 24342 4708 24344
rect 4468 24322 4764 24342
rect 5154 24291 5182 24597
rect 9796 24398 10092 24418
rect 9852 24396 9876 24398
rect 9932 24396 9956 24398
rect 10012 24396 10036 24398
rect 9874 24344 9876 24396
rect 9938 24344 9950 24396
rect 10012 24344 10014 24396
rect 9852 24342 9876 24344
rect 9932 24342 9956 24344
rect 10012 24342 10036 24344
rect 9796 24322 10092 24342
rect 15124 24398 15420 24418
rect 15180 24396 15204 24398
rect 15260 24396 15284 24398
rect 15340 24396 15364 24398
rect 15202 24344 15204 24396
rect 15266 24344 15278 24396
rect 15340 24344 15342 24396
rect 15180 24342 15204 24344
rect 15260 24342 15284 24344
rect 15340 24342 15364 24344
rect 15124 24322 15420 24342
rect 20452 24398 20748 24418
rect 20508 24396 20532 24398
rect 20588 24396 20612 24398
rect 20668 24396 20692 24398
rect 20530 24344 20532 24396
rect 20594 24344 20606 24396
rect 20668 24344 20670 24396
rect 20508 24342 20532 24344
rect 20588 24342 20612 24344
rect 20668 24342 20692 24344
rect 20452 24322 20748 24342
rect 5142 24285 5194 24291
rect 5142 24227 5194 24233
rect 2742 24063 2794 24069
rect 2742 24005 2794 24011
rect 2754 23551 2782 24005
rect 7132 23732 7428 23752
rect 7188 23730 7212 23732
rect 7268 23730 7292 23732
rect 7348 23730 7372 23732
rect 7210 23678 7212 23730
rect 7274 23678 7286 23730
rect 7348 23678 7350 23730
rect 7188 23676 7212 23678
rect 7268 23676 7292 23678
rect 7348 23676 7372 23678
rect 7132 23656 7428 23676
rect 12460 23732 12756 23752
rect 12516 23730 12540 23732
rect 12596 23730 12620 23732
rect 12676 23730 12700 23732
rect 12538 23678 12540 23730
rect 12602 23678 12614 23730
rect 12676 23678 12678 23730
rect 12516 23676 12540 23678
rect 12596 23676 12620 23678
rect 12676 23676 12700 23678
rect 12460 23656 12756 23676
rect 17788 23732 18084 23752
rect 17844 23730 17868 23732
rect 17924 23730 17948 23732
rect 18004 23730 18028 23732
rect 17866 23678 17868 23730
rect 17930 23678 17942 23730
rect 18004 23678 18006 23730
rect 17844 23676 17868 23678
rect 17924 23676 17948 23678
rect 18004 23676 18028 23678
rect 17788 23656 18084 23676
rect 2742 23545 2794 23551
rect 2742 23487 2794 23493
rect 2070 23397 2122 23403
rect 2068 23362 2070 23371
rect 2122 23362 2124 23371
rect 2068 23297 2124 23306
rect 2742 23323 2794 23329
rect 2742 23265 2794 23271
rect 2754 22737 2782 23265
rect 7734 23249 7786 23255
rect 7734 23191 7786 23197
rect 4468 23066 4764 23086
rect 4524 23064 4548 23066
rect 4604 23064 4628 23066
rect 4684 23064 4708 23066
rect 4546 23012 4548 23064
rect 4610 23012 4622 23064
rect 4684 23012 4686 23064
rect 4524 23010 4548 23012
rect 4604 23010 4628 23012
rect 4684 23010 4708 23012
rect 4468 22990 4764 23010
rect 7746 22737 7774 23191
rect 9796 23066 10092 23086
rect 9852 23064 9876 23066
rect 9932 23064 9956 23066
rect 10012 23064 10036 23066
rect 9874 23012 9876 23064
rect 9938 23012 9950 23064
rect 10012 23012 10014 23064
rect 9852 23010 9876 23012
rect 9932 23010 9956 23012
rect 10012 23010 10036 23012
rect 9796 22990 10092 23010
rect 15124 23066 15420 23086
rect 15180 23064 15204 23066
rect 15260 23064 15284 23066
rect 15340 23064 15364 23066
rect 15202 23012 15204 23064
rect 15266 23012 15278 23064
rect 15340 23012 15342 23064
rect 15180 23010 15204 23012
rect 15260 23010 15284 23012
rect 15340 23010 15364 23012
rect 15124 22990 15420 23010
rect 20452 23066 20748 23086
rect 20508 23064 20532 23066
rect 20588 23064 20612 23066
rect 20668 23064 20692 23066
rect 20530 23012 20532 23064
rect 20594 23012 20606 23064
rect 20668 23012 20670 23064
rect 20508 23010 20532 23012
rect 20588 23010 20612 23012
rect 20668 23010 20692 23012
rect 20452 22990 20748 23010
rect 2742 22731 2794 22737
rect 2742 22673 2794 22679
rect 7734 22731 7786 22737
rect 7734 22673 7786 22679
rect 2754 22293 2782 22673
rect 7132 22400 7428 22420
rect 7188 22398 7212 22400
rect 7268 22398 7292 22400
rect 7348 22398 7372 22400
rect 7210 22346 7212 22398
rect 7274 22346 7286 22398
rect 7348 22346 7350 22398
rect 7188 22344 7212 22346
rect 7268 22344 7292 22346
rect 7348 22344 7372 22346
rect 7132 22324 7428 22344
rect 12460 22400 12756 22420
rect 12516 22398 12540 22400
rect 12596 22398 12620 22400
rect 12676 22398 12700 22400
rect 12538 22346 12540 22398
rect 12602 22346 12614 22398
rect 12676 22346 12678 22398
rect 12516 22344 12540 22346
rect 12596 22344 12620 22346
rect 12676 22344 12700 22346
rect 12460 22324 12756 22344
rect 17788 22400 18084 22420
rect 17844 22398 17868 22400
rect 17924 22398 17948 22400
rect 18004 22398 18028 22400
rect 17866 22346 17868 22398
rect 17930 22346 17942 22398
rect 18004 22346 18006 22398
rect 17844 22344 17868 22346
rect 17924 22344 17948 22346
rect 18004 22344 18028 22346
rect 17788 22324 18084 22344
rect 2742 22287 2794 22293
rect 2742 22229 2794 22235
rect 2070 22065 2122 22071
rect 2070 22007 2122 22013
rect 2082 21891 2110 22007
rect 2742 21991 2794 21997
rect 2742 21933 2794 21939
rect 12630 21991 12682 21997
rect 12630 21933 12682 21939
rect 2068 21882 2124 21891
rect 2068 21817 2124 21826
rect 2754 21405 2782 21933
rect 4468 21734 4764 21754
rect 4524 21732 4548 21734
rect 4604 21732 4628 21734
rect 4684 21732 4708 21734
rect 4546 21680 4548 21732
rect 4610 21680 4622 21732
rect 4684 21680 4686 21732
rect 4524 21678 4548 21680
rect 4604 21678 4628 21680
rect 4684 21678 4708 21680
rect 4468 21658 4764 21678
rect 9796 21734 10092 21754
rect 9852 21732 9876 21734
rect 9932 21732 9956 21734
rect 10012 21732 10036 21734
rect 9874 21680 9876 21732
rect 9938 21680 9950 21732
rect 10012 21680 10014 21732
rect 9852 21678 9876 21680
rect 9932 21678 9956 21680
rect 10012 21678 10036 21680
rect 9796 21658 10092 21678
rect 12642 21627 12670 21933
rect 15124 21734 15420 21754
rect 15180 21732 15204 21734
rect 15260 21732 15284 21734
rect 15340 21732 15364 21734
rect 15202 21680 15204 21732
rect 15266 21680 15278 21732
rect 15340 21680 15342 21732
rect 15180 21678 15204 21680
rect 15260 21678 15284 21680
rect 15340 21678 15364 21680
rect 15124 21658 15420 21678
rect 20452 21734 20748 21754
rect 20508 21732 20532 21734
rect 20588 21732 20612 21734
rect 20668 21732 20692 21734
rect 20530 21680 20532 21732
rect 20594 21680 20606 21732
rect 20668 21680 20670 21732
rect 20508 21678 20532 21680
rect 20588 21678 20612 21680
rect 20668 21678 20692 21680
rect 20452 21658 20748 21678
rect 12630 21621 12682 21627
rect 12630 21563 12682 21569
rect 2742 21399 2794 21405
rect 2742 21341 2794 21347
rect 2754 20961 2782 21341
rect 7132 21068 7428 21088
rect 7188 21066 7212 21068
rect 7268 21066 7292 21068
rect 7348 21066 7372 21068
rect 7210 21014 7212 21066
rect 7274 21014 7286 21066
rect 7348 21014 7350 21066
rect 7188 21012 7212 21014
rect 7268 21012 7292 21014
rect 7348 21012 7372 21014
rect 7132 20992 7428 21012
rect 12460 21068 12756 21088
rect 12516 21066 12540 21068
rect 12596 21066 12620 21068
rect 12676 21066 12700 21068
rect 12538 21014 12540 21066
rect 12602 21014 12614 21066
rect 12676 21014 12678 21066
rect 12516 21012 12540 21014
rect 12596 21012 12620 21014
rect 12676 21012 12700 21014
rect 12460 20992 12756 21012
rect 17788 21068 18084 21088
rect 17844 21066 17868 21068
rect 17924 21066 17948 21068
rect 18004 21066 18028 21068
rect 17866 21014 17868 21066
rect 17930 21014 17942 21066
rect 18004 21014 18006 21066
rect 17844 21012 17868 21014
rect 17924 21012 17948 21014
rect 18004 21012 18028 21014
rect 17788 20992 18084 21012
rect 2742 20955 2794 20961
rect 2742 20897 2794 20903
rect 2454 20733 2506 20739
rect 2454 20675 2506 20681
rect 2358 20659 2410 20665
rect 2358 20601 2410 20607
rect 2370 20147 2398 20601
rect 2358 20141 2410 20147
rect 2466 20115 2494 20675
rect 22614 20659 22666 20665
rect 22614 20601 22666 20607
rect 4468 20402 4764 20422
rect 4524 20400 4548 20402
rect 4604 20400 4628 20402
rect 4684 20400 4708 20402
rect 4546 20348 4548 20400
rect 4610 20348 4622 20400
rect 4684 20348 4686 20400
rect 4524 20346 4548 20348
rect 4604 20346 4628 20348
rect 4684 20346 4708 20348
rect 4468 20326 4764 20346
rect 9796 20402 10092 20422
rect 9852 20400 9876 20402
rect 9932 20400 9956 20402
rect 10012 20400 10036 20402
rect 9874 20348 9876 20400
rect 9938 20348 9950 20400
rect 10012 20348 10014 20400
rect 9852 20346 9876 20348
rect 9932 20346 9956 20348
rect 10012 20346 10036 20348
rect 9796 20326 10092 20346
rect 15124 20402 15420 20422
rect 15180 20400 15204 20402
rect 15260 20400 15284 20402
rect 15340 20400 15364 20402
rect 15202 20348 15204 20400
rect 15266 20348 15278 20400
rect 15340 20348 15342 20400
rect 15180 20346 15204 20348
rect 15260 20346 15284 20348
rect 15340 20346 15364 20348
rect 15124 20326 15420 20346
rect 20452 20402 20748 20422
rect 20508 20400 20532 20402
rect 20588 20400 20612 20402
rect 20668 20400 20692 20402
rect 20530 20348 20532 20400
rect 20594 20348 20606 20400
rect 20668 20348 20670 20400
rect 20508 20346 20532 20348
rect 20588 20346 20612 20348
rect 20668 20346 20692 20348
rect 20452 20326 20748 20346
rect 22626 20295 22654 20601
rect 22614 20289 22666 20295
rect 22614 20231 22666 20237
rect 2742 20141 2794 20147
rect 2358 20083 2410 20089
rect 2452 20106 2508 20115
rect 2742 20083 2794 20089
rect 2452 20041 2508 20050
rect 2754 19629 2782 20083
rect 7132 19736 7428 19756
rect 7188 19734 7212 19736
rect 7268 19734 7292 19736
rect 7348 19734 7372 19736
rect 7210 19682 7212 19734
rect 7274 19682 7286 19734
rect 7348 19682 7350 19734
rect 7188 19680 7212 19682
rect 7268 19680 7292 19682
rect 7348 19680 7372 19682
rect 7132 19660 7428 19680
rect 12460 19736 12756 19756
rect 12516 19734 12540 19736
rect 12596 19734 12620 19736
rect 12676 19734 12700 19736
rect 12538 19682 12540 19734
rect 12602 19682 12614 19734
rect 12676 19682 12678 19734
rect 12516 19680 12540 19682
rect 12596 19680 12620 19682
rect 12676 19680 12700 19682
rect 12460 19660 12756 19680
rect 17788 19736 18084 19756
rect 17844 19734 17868 19736
rect 17924 19734 17948 19736
rect 18004 19734 18028 19736
rect 17866 19682 17868 19734
rect 17930 19682 17942 19734
rect 18004 19682 18006 19734
rect 17844 19680 17868 19682
rect 17924 19680 17948 19682
rect 18004 19680 18028 19682
rect 17788 19660 18084 19680
rect 2742 19623 2794 19629
rect 2742 19565 2794 19571
rect 2070 19401 2122 19407
rect 2068 19366 2070 19375
rect 2122 19366 2124 19375
rect 2068 19301 2124 19310
rect 2358 19327 2410 19333
rect 2358 19269 2410 19275
rect 22614 19327 22666 19333
rect 22614 19269 22666 19275
rect 2370 17483 2398 19269
rect 4468 19070 4764 19090
rect 4524 19068 4548 19070
rect 4604 19068 4628 19070
rect 4684 19068 4708 19070
rect 4546 19016 4548 19068
rect 4610 19016 4622 19068
rect 4684 19016 4686 19068
rect 4524 19014 4548 19016
rect 4604 19014 4628 19016
rect 4684 19014 4708 19016
rect 4468 18994 4764 19014
rect 9796 19070 10092 19090
rect 9852 19068 9876 19070
rect 9932 19068 9956 19070
rect 10012 19068 10036 19070
rect 9874 19016 9876 19068
rect 9938 19016 9950 19068
rect 10012 19016 10014 19068
rect 9852 19014 9876 19016
rect 9932 19014 9956 19016
rect 10012 19014 10036 19016
rect 9796 18994 10092 19014
rect 15124 19070 15420 19090
rect 15180 19068 15204 19070
rect 15260 19068 15284 19070
rect 15340 19068 15364 19070
rect 15202 19016 15204 19068
rect 15266 19016 15278 19068
rect 15340 19016 15342 19068
rect 15180 19014 15204 19016
rect 15260 19014 15284 19016
rect 15340 19014 15364 19016
rect 15124 18994 15420 19014
rect 20452 19070 20748 19090
rect 20508 19068 20532 19070
rect 20588 19068 20612 19070
rect 20668 19068 20692 19070
rect 20530 19016 20532 19068
rect 20594 19016 20606 19068
rect 20668 19016 20670 19068
rect 20508 19014 20532 19016
rect 20588 19014 20612 19016
rect 20668 19014 20692 19016
rect 20452 18994 20748 19014
rect 22626 18889 22654 19269
rect 22614 18883 22666 18889
rect 22614 18825 22666 18831
rect 3894 18735 3946 18741
rect 3894 18677 3946 18683
rect 3906 18149 3934 18677
rect 7132 18404 7428 18424
rect 7188 18402 7212 18404
rect 7268 18402 7292 18404
rect 7348 18402 7372 18404
rect 7210 18350 7212 18402
rect 7274 18350 7286 18402
rect 7348 18350 7350 18402
rect 7188 18348 7212 18350
rect 7268 18348 7292 18350
rect 7348 18348 7372 18350
rect 7132 18328 7428 18348
rect 12460 18404 12756 18424
rect 12516 18402 12540 18404
rect 12596 18402 12620 18404
rect 12676 18402 12700 18404
rect 12538 18350 12540 18402
rect 12602 18350 12614 18402
rect 12676 18350 12678 18402
rect 12516 18348 12540 18350
rect 12596 18348 12620 18350
rect 12676 18348 12700 18350
rect 12460 18328 12756 18348
rect 17788 18404 18084 18424
rect 17844 18402 17868 18404
rect 17924 18402 17948 18404
rect 18004 18402 18028 18404
rect 17866 18350 17868 18402
rect 17930 18350 17942 18402
rect 18004 18350 18006 18402
rect 17844 18348 17868 18350
rect 17924 18348 17948 18350
rect 18004 18348 18028 18350
rect 17788 18328 18084 18348
rect 3894 18143 3946 18149
rect 3894 18085 3946 18091
rect 22134 17995 22186 18001
rect 22134 17937 22186 17943
rect 4468 17738 4764 17758
rect 4524 17736 4548 17738
rect 4604 17736 4628 17738
rect 4684 17736 4708 17738
rect 4546 17684 4548 17736
rect 4610 17684 4622 17736
rect 4684 17684 4686 17736
rect 4524 17682 4548 17684
rect 4604 17682 4628 17684
rect 4684 17682 4708 17684
rect 4468 17662 4764 17682
rect 9796 17738 10092 17758
rect 9852 17736 9876 17738
rect 9932 17736 9956 17738
rect 10012 17736 10036 17738
rect 9874 17684 9876 17736
rect 9938 17684 9950 17736
rect 10012 17684 10014 17736
rect 9852 17682 9876 17684
rect 9932 17682 9956 17684
rect 10012 17682 10036 17684
rect 9796 17662 10092 17682
rect 15124 17738 15420 17758
rect 15180 17736 15204 17738
rect 15260 17736 15284 17738
rect 15340 17736 15364 17738
rect 15202 17684 15204 17736
rect 15266 17684 15278 17736
rect 15340 17684 15342 17736
rect 15180 17682 15204 17684
rect 15260 17682 15284 17684
rect 15340 17682 15364 17684
rect 15124 17662 15420 17682
rect 20452 17738 20748 17758
rect 20508 17736 20532 17738
rect 20588 17736 20612 17738
rect 20668 17736 20692 17738
rect 20530 17684 20532 17736
rect 20594 17684 20606 17736
rect 20668 17684 20670 17736
rect 20508 17682 20532 17684
rect 20588 17682 20612 17684
rect 20668 17682 20692 17684
rect 20452 17662 20748 17682
rect 22146 17631 22174 17937
rect 22134 17625 22186 17631
rect 22134 17567 22186 17573
rect 2358 17477 2410 17483
rect 2358 17419 2410 17425
rect 2370 16965 2398 17419
rect 7132 17072 7428 17092
rect 7188 17070 7212 17072
rect 7268 17070 7292 17072
rect 7348 17070 7372 17072
rect 7210 17018 7212 17070
rect 7274 17018 7286 17070
rect 7348 17018 7350 17070
rect 7188 17016 7212 17018
rect 7268 17016 7292 17018
rect 7348 17016 7372 17018
rect 7132 16996 7428 17016
rect 12460 17072 12756 17092
rect 12516 17070 12540 17072
rect 12596 17070 12620 17072
rect 12676 17070 12700 17072
rect 12538 17018 12540 17070
rect 12602 17018 12614 17070
rect 12676 17018 12678 17070
rect 12516 17016 12540 17018
rect 12596 17016 12620 17018
rect 12676 17016 12700 17018
rect 12460 16996 12756 17016
rect 17788 17072 18084 17092
rect 17844 17070 17868 17072
rect 17924 17070 17948 17072
rect 18004 17070 18028 17072
rect 17866 17018 17868 17070
rect 17930 17018 17942 17070
rect 18004 17018 18006 17070
rect 17844 17016 17868 17018
rect 17924 17016 17948 17018
rect 18004 17016 18028 17018
rect 17788 16996 18084 17016
rect 2358 16959 2410 16965
rect 2358 16901 2410 16907
rect 2070 16737 2122 16743
rect 2070 16679 2122 16685
rect 2082 16119 2110 16679
rect 2358 16663 2410 16669
rect 2358 16605 2410 16611
rect 22614 16663 22666 16669
rect 22614 16605 22666 16611
rect 2068 16110 2124 16119
rect 2068 16045 2124 16054
rect 2370 12155 2398 16605
rect 4468 16406 4764 16426
rect 4524 16404 4548 16406
rect 4604 16404 4628 16406
rect 4684 16404 4708 16406
rect 4546 16352 4548 16404
rect 4610 16352 4622 16404
rect 4684 16352 4686 16404
rect 4524 16350 4548 16352
rect 4604 16350 4628 16352
rect 4684 16350 4708 16352
rect 4468 16330 4764 16350
rect 9796 16406 10092 16426
rect 9852 16404 9876 16406
rect 9932 16404 9956 16406
rect 10012 16404 10036 16406
rect 9874 16352 9876 16404
rect 9938 16352 9950 16404
rect 10012 16352 10014 16404
rect 9852 16350 9876 16352
rect 9932 16350 9956 16352
rect 10012 16350 10036 16352
rect 9796 16330 10092 16350
rect 15124 16406 15420 16426
rect 15180 16404 15204 16406
rect 15260 16404 15284 16406
rect 15340 16404 15364 16406
rect 15202 16352 15204 16404
rect 15266 16352 15278 16404
rect 15340 16352 15342 16404
rect 15180 16350 15204 16352
rect 15260 16350 15284 16352
rect 15340 16350 15364 16352
rect 15124 16330 15420 16350
rect 20452 16406 20748 16426
rect 20508 16404 20532 16406
rect 20588 16404 20612 16406
rect 20668 16404 20692 16406
rect 20530 16352 20532 16404
rect 20594 16352 20606 16404
rect 20668 16352 20670 16404
rect 20508 16350 20532 16352
rect 20588 16350 20612 16352
rect 20668 16350 20692 16352
rect 20452 16330 20748 16350
rect 22626 16299 22654 16605
rect 22614 16293 22666 16299
rect 22614 16235 22666 16241
rect 3894 16071 3946 16077
rect 3894 16013 3946 16019
rect 3906 15633 3934 16013
rect 7132 15740 7428 15760
rect 7188 15738 7212 15740
rect 7268 15738 7292 15740
rect 7348 15738 7372 15740
rect 7210 15686 7212 15738
rect 7274 15686 7286 15738
rect 7348 15686 7350 15738
rect 7188 15684 7212 15686
rect 7268 15684 7292 15686
rect 7348 15684 7372 15686
rect 7132 15664 7428 15684
rect 12460 15740 12756 15760
rect 12516 15738 12540 15740
rect 12596 15738 12620 15740
rect 12676 15738 12700 15740
rect 12538 15686 12540 15738
rect 12602 15686 12614 15738
rect 12676 15686 12678 15738
rect 12516 15684 12540 15686
rect 12596 15684 12620 15686
rect 12676 15684 12700 15686
rect 12460 15664 12756 15684
rect 17788 15740 18084 15760
rect 17844 15738 17868 15740
rect 17924 15738 17948 15740
rect 18004 15738 18028 15740
rect 17866 15686 17868 15738
rect 17930 15686 17942 15738
rect 18004 15686 18006 15738
rect 17844 15684 17868 15686
rect 17924 15684 17948 15686
rect 18004 15684 18028 15686
rect 17788 15664 18084 15684
rect 3894 15627 3946 15633
rect 3894 15569 3946 15575
rect 22614 15331 22666 15337
rect 22614 15273 22666 15279
rect 4468 15074 4764 15094
rect 4524 15072 4548 15074
rect 4604 15072 4628 15074
rect 4684 15072 4708 15074
rect 4546 15020 4548 15072
rect 4610 15020 4622 15072
rect 4684 15020 4686 15072
rect 4524 15018 4548 15020
rect 4604 15018 4628 15020
rect 4684 15018 4708 15020
rect 4468 14998 4764 15018
rect 9796 15074 10092 15094
rect 9852 15072 9876 15074
rect 9932 15072 9956 15074
rect 10012 15072 10036 15074
rect 9874 15020 9876 15072
rect 9938 15020 9950 15072
rect 10012 15020 10014 15072
rect 9852 15018 9876 15020
rect 9932 15018 9956 15020
rect 10012 15018 10036 15020
rect 9796 14998 10092 15018
rect 15124 15074 15420 15094
rect 15180 15072 15204 15074
rect 15260 15072 15284 15074
rect 15340 15072 15364 15074
rect 15202 15020 15204 15072
rect 15266 15020 15278 15072
rect 15340 15020 15342 15072
rect 15180 15018 15204 15020
rect 15260 15018 15284 15020
rect 15340 15018 15364 15020
rect 15124 14998 15420 15018
rect 20452 15074 20748 15094
rect 20508 15072 20532 15074
rect 20588 15072 20612 15074
rect 20668 15072 20692 15074
rect 20530 15020 20532 15072
rect 20594 15020 20606 15072
rect 20668 15020 20670 15072
rect 20508 15018 20532 15020
rect 20588 15018 20612 15020
rect 20668 15018 20692 15020
rect 20452 14998 20748 15018
rect 22626 14967 22654 15273
rect 22614 14961 22666 14967
rect 22614 14903 22666 14909
rect 3894 14739 3946 14745
rect 3894 14681 3946 14687
rect 3906 14301 3934 14681
rect 7132 14408 7428 14428
rect 7188 14406 7212 14408
rect 7268 14406 7292 14408
rect 7348 14406 7372 14408
rect 7210 14354 7212 14406
rect 7274 14354 7286 14406
rect 7348 14354 7350 14406
rect 7188 14352 7212 14354
rect 7268 14352 7292 14354
rect 7348 14352 7372 14354
rect 7132 14332 7428 14352
rect 12460 14408 12756 14428
rect 12516 14406 12540 14408
rect 12596 14406 12620 14408
rect 12676 14406 12700 14408
rect 12538 14354 12540 14406
rect 12602 14354 12614 14406
rect 12676 14354 12678 14406
rect 12516 14352 12540 14354
rect 12596 14352 12620 14354
rect 12676 14352 12700 14354
rect 12460 14332 12756 14352
rect 17788 14408 18084 14428
rect 17844 14406 17868 14408
rect 17924 14406 17948 14408
rect 18004 14406 18028 14408
rect 17866 14354 17868 14406
rect 17930 14354 17942 14406
rect 18004 14354 18006 14406
rect 17844 14352 17868 14354
rect 17924 14352 17948 14354
rect 18004 14352 18028 14354
rect 17788 14332 18084 14352
rect 3894 14295 3946 14301
rect 3894 14237 3946 14243
rect 22614 13999 22666 14005
rect 22614 13941 22666 13947
rect 4468 13742 4764 13762
rect 4524 13740 4548 13742
rect 4604 13740 4628 13742
rect 4684 13740 4708 13742
rect 4546 13688 4548 13740
rect 4610 13688 4622 13740
rect 4684 13688 4686 13740
rect 4524 13686 4548 13688
rect 4604 13686 4628 13688
rect 4684 13686 4708 13688
rect 4468 13666 4764 13686
rect 9796 13742 10092 13762
rect 9852 13740 9876 13742
rect 9932 13740 9956 13742
rect 10012 13740 10036 13742
rect 9874 13688 9876 13740
rect 9938 13688 9950 13740
rect 10012 13688 10014 13740
rect 9852 13686 9876 13688
rect 9932 13686 9956 13688
rect 10012 13686 10036 13688
rect 9796 13666 10092 13686
rect 15124 13742 15420 13762
rect 15180 13740 15204 13742
rect 15260 13740 15284 13742
rect 15340 13740 15364 13742
rect 15202 13688 15204 13740
rect 15266 13688 15278 13740
rect 15340 13688 15342 13740
rect 15180 13686 15204 13688
rect 15260 13686 15284 13688
rect 15340 13686 15364 13688
rect 15124 13666 15420 13686
rect 20452 13742 20748 13762
rect 20508 13740 20532 13742
rect 20588 13740 20612 13742
rect 20668 13740 20692 13742
rect 20530 13688 20532 13740
rect 20594 13688 20606 13740
rect 20668 13688 20670 13740
rect 20508 13686 20532 13688
rect 20588 13686 20612 13688
rect 20668 13686 20692 13688
rect 20452 13666 20748 13686
rect 22626 13561 22654 13941
rect 22614 13555 22666 13561
rect 22614 13497 22666 13503
rect 3894 13407 3946 13413
rect 3894 13349 3946 13355
rect 3906 12969 3934 13349
rect 7132 13076 7428 13096
rect 7188 13074 7212 13076
rect 7268 13074 7292 13076
rect 7348 13074 7372 13076
rect 7210 13022 7212 13074
rect 7274 13022 7286 13074
rect 7348 13022 7350 13074
rect 7188 13020 7212 13022
rect 7268 13020 7292 13022
rect 7348 13020 7372 13022
rect 7132 13000 7428 13020
rect 12460 13076 12756 13096
rect 12516 13074 12540 13076
rect 12596 13074 12620 13076
rect 12676 13074 12700 13076
rect 12538 13022 12540 13074
rect 12602 13022 12614 13074
rect 12676 13022 12678 13074
rect 12516 13020 12540 13022
rect 12596 13020 12620 13022
rect 12676 13020 12700 13022
rect 12460 13000 12756 13020
rect 17788 13076 18084 13096
rect 17844 13074 17868 13076
rect 17924 13074 17948 13076
rect 18004 13074 18028 13076
rect 17866 13022 17868 13074
rect 17930 13022 17942 13074
rect 18004 13022 18006 13074
rect 17844 13020 17868 13022
rect 17924 13020 17948 13022
rect 18004 13020 18028 13022
rect 17788 13000 18084 13020
rect 3894 12963 3946 12969
rect 3894 12905 3946 12911
rect 22134 12667 22186 12673
rect 22134 12609 22186 12615
rect 4468 12410 4764 12430
rect 4524 12408 4548 12410
rect 4604 12408 4628 12410
rect 4684 12408 4708 12410
rect 4546 12356 4548 12408
rect 4610 12356 4622 12408
rect 4684 12356 4686 12408
rect 4524 12354 4548 12356
rect 4604 12354 4628 12356
rect 4684 12354 4708 12356
rect 4468 12334 4764 12354
rect 9796 12410 10092 12430
rect 9852 12408 9876 12410
rect 9932 12408 9956 12410
rect 10012 12408 10036 12410
rect 9874 12356 9876 12408
rect 9938 12356 9950 12408
rect 10012 12356 10014 12408
rect 9852 12354 9876 12356
rect 9932 12354 9956 12356
rect 10012 12354 10036 12356
rect 9796 12334 10092 12354
rect 15124 12410 15420 12430
rect 15180 12408 15204 12410
rect 15260 12408 15284 12410
rect 15340 12408 15364 12410
rect 15202 12356 15204 12408
rect 15266 12356 15278 12408
rect 15340 12356 15342 12408
rect 15180 12354 15204 12356
rect 15260 12354 15284 12356
rect 15340 12354 15364 12356
rect 15124 12334 15420 12354
rect 20452 12410 20748 12430
rect 20508 12408 20532 12410
rect 20588 12408 20612 12410
rect 20668 12408 20692 12410
rect 20530 12356 20532 12408
rect 20594 12356 20606 12408
rect 20668 12356 20670 12408
rect 20508 12354 20532 12356
rect 20588 12354 20612 12356
rect 20668 12354 20692 12356
rect 20452 12334 20748 12354
rect 22146 12303 22174 12609
rect 22134 12297 22186 12303
rect 22134 12239 22186 12245
rect 2358 12149 2410 12155
rect 2358 12091 2410 12097
rect 2370 11637 2398 12091
rect 7132 11744 7428 11764
rect 7188 11742 7212 11744
rect 7268 11742 7292 11744
rect 7348 11742 7372 11744
rect 7210 11690 7212 11742
rect 7274 11690 7286 11742
rect 7348 11690 7350 11742
rect 7188 11688 7212 11690
rect 7268 11688 7292 11690
rect 7348 11688 7372 11690
rect 7132 11668 7428 11688
rect 12460 11744 12756 11764
rect 12516 11742 12540 11744
rect 12596 11742 12620 11744
rect 12676 11742 12700 11744
rect 12538 11690 12540 11742
rect 12602 11690 12614 11742
rect 12676 11690 12678 11742
rect 12516 11688 12540 11690
rect 12596 11688 12620 11690
rect 12676 11688 12700 11690
rect 12460 11668 12756 11688
rect 17788 11744 18084 11764
rect 17844 11742 17868 11744
rect 17924 11742 17948 11744
rect 18004 11742 18028 11744
rect 17866 11690 17868 11742
rect 17930 11690 17942 11742
rect 18004 11690 18006 11742
rect 17844 11688 17868 11690
rect 17924 11688 17948 11690
rect 18004 11688 18028 11690
rect 17788 11668 18084 11688
rect 2358 11631 2410 11637
rect 2358 11573 2410 11579
rect 2070 11409 2122 11415
rect 2070 11351 2122 11357
rect 2082 10791 2110 11351
rect 2358 11335 2410 11341
rect 2358 11277 2410 11283
rect 22614 11335 22666 11341
rect 22614 11277 22666 11283
rect 2068 10782 2124 10791
rect 2068 10717 2124 10726
rect 2370 1425 2398 11277
rect 4468 11078 4764 11098
rect 4524 11076 4548 11078
rect 4604 11076 4628 11078
rect 4684 11076 4708 11078
rect 4546 11024 4548 11076
rect 4610 11024 4622 11076
rect 4684 11024 4686 11076
rect 4524 11022 4548 11024
rect 4604 11022 4628 11024
rect 4684 11022 4708 11024
rect 4468 11002 4764 11022
rect 9796 11078 10092 11098
rect 9852 11076 9876 11078
rect 9932 11076 9956 11078
rect 10012 11076 10036 11078
rect 9874 11024 9876 11076
rect 9938 11024 9950 11076
rect 10012 11024 10014 11076
rect 9852 11022 9876 11024
rect 9932 11022 9956 11024
rect 10012 11022 10036 11024
rect 9796 11002 10092 11022
rect 15124 11078 15420 11098
rect 15180 11076 15204 11078
rect 15260 11076 15284 11078
rect 15340 11076 15364 11078
rect 15202 11024 15204 11076
rect 15266 11024 15278 11076
rect 15340 11024 15342 11076
rect 15180 11022 15204 11024
rect 15260 11022 15284 11024
rect 15340 11022 15364 11024
rect 15124 11002 15420 11022
rect 20452 11078 20748 11098
rect 20508 11076 20532 11078
rect 20588 11076 20612 11078
rect 20668 11076 20692 11078
rect 20530 11024 20532 11076
rect 20594 11024 20606 11076
rect 20668 11024 20670 11076
rect 20508 11022 20532 11024
rect 20588 11022 20612 11024
rect 20668 11022 20692 11024
rect 20452 11002 20748 11022
rect 22626 10971 22654 11277
rect 22614 10965 22666 10971
rect 22614 10907 22666 10913
rect 3894 10743 3946 10749
rect 3894 10685 3946 10691
rect 3906 10305 3934 10685
rect 7132 10412 7428 10432
rect 7188 10410 7212 10412
rect 7268 10410 7292 10412
rect 7348 10410 7372 10412
rect 7210 10358 7212 10410
rect 7274 10358 7286 10410
rect 7348 10358 7350 10410
rect 7188 10356 7212 10358
rect 7268 10356 7292 10358
rect 7348 10356 7372 10358
rect 7132 10336 7428 10356
rect 12460 10412 12756 10432
rect 12516 10410 12540 10412
rect 12596 10410 12620 10412
rect 12676 10410 12700 10412
rect 12538 10358 12540 10410
rect 12602 10358 12614 10410
rect 12676 10358 12678 10410
rect 12516 10356 12540 10358
rect 12596 10356 12620 10358
rect 12676 10356 12700 10358
rect 12460 10336 12756 10356
rect 17788 10412 18084 10432
rect 17844 10410 17868 10412
rect 17924 10410 17948 10412
rect 18004 10410 18028 10412
rect 17866 10358 17868 10410
rect 17930 10358 17942 10410
rect 18004 10358 18006 10410
rect 17844 10356 17868 10358
rect 17924 10356 17948 10358
rect 18004 10356 18028 10358
rect 17788 10336 18084 10356
rect 3894 10299 3946 10305
rect 3894 10241 3946 10247
rect 22614 10003 22666 10009
rect 22614 9945 22666 9951
rect 4468 9746 4764 9766
rect 4524 9744 4548 9746
rect 4604 9744 4628 9746
rect 4684 9744 4708 9746
rect 4546 9692 4548 9744
rect 4610 9692 4622 9744
rect 4684 9692 4686 9744
rect 4524 9690 4548 9692
rect 4604 9690 4628 9692
rect 4684 9690 4708 9692
rect 4468 9670 4764 9690
rect 9796 9746 10092 9766
rect 9852 9744 9876 9746
rect 9932 9744 9956 9746
rect 10012 9744 10036 9746
rect 9874 9692 9876 9744
rect 9938 9692 9950 9744
rect 10012 9692 10014 9744
rect 9852 9690 9876 9692
rect 9932 9690 9956 9692
rect 10012 9690 10036 9692
rect 9796 9670 10092 9690
rect 15124 9746 15420 9766
rect 15180 9744 15204 9746
rect 15260 9744 15284 9746
rect 15340 9744 15364 9746
rect 15202 9692 15204 9744
rect 15266 9692 15278 9744
rect 15340 9692 15342 9744
rect 15180 9690 15204 9692
rect 15260 9690 15284 9692
rect 15340 9690 15364 9692
rect 15124 9670 15420 9690
rect 20452 9746 20748 9766
rect 20508 9744 20532 9746
rect 20588 9744 20612 9746
rect 20668 9744 20692 9746
rect 20530 9692 20532 9744
rect 20594 9692 20606 9744
rect 20668 9692 20670 9744
rect 20508 9690 20532 9692
rect 20588 9690 20612 9692
rect 20668 9690 20692 9692
rect 20452 9670 20748 9690
rect 22626 9639 22654 9945
rect 22614 9633 22666 9639
rect 22614 9575 22666 9581
rect 3894 9411 3946 9417
rect 3894 9353 3946 9359
rect 3906 8973 3934 9353
rect 7132 9080 7428 9100
rect 7188 9078 7212 9080
rect 7268 9078 7292 9080
rect 7348 9078 7372 9080
rect 7210 9026 7212 9078
rect 7274 9026 7286 9078
rect 7348 9026 7350 9078
rect 7188 9024 7212 9026
rect 7268 9024 7292 9026
rect 7348 9024 7372 9026
rect 7132 9004 7428 9024
rect 12460 9080 12756 9100
rect 12516 9078 12540 9080
rect 12596 9078 12620 9080
rect 12676 9078 12700 9080
rect 12538 9026 12540 9078
rect 12602 9026 12614 9078
rect 12676 9026 12678 9078
rect 12516 9024 12540 9026
rect 12596 9024 12620 9026
rect 12676 9024 12700 9026
rect 12460 9004 12756 9024
rect 17788 9080 18084 9100
rect 17844 9078 17868 9080
rect 17924 9078 17948 9080
rect 18004 9078 18028 9080
rect 17866 9026 17868 9078
rect 17930 9026 17942 9078
rect 18004 9026 18006 9078
rect 17844 9024 17868 9026
rect 17924 9024 17948 9026
rect 18004 9024 18028 9026
rect 17788 9004 18084 9024
rect 3894 8967 3946 8973
rect 3894 8909 3946 8915
rect 22614 8671 22666 8677
rect 22614 8613 22666 8619
rect 4468 8414 4764 8434
rect 4524 8412 4548 8414
rect 4604 8412 4628 8414
rect 4684 8412 4708 8414
rect 4546 8360 4548 8412
rect 4610 8360 4622 8412
rect 4684 8360 4686 8412
rect 4524 8358 4548 8360
rect 4604 8358 4628 8360
rect 4684 8358 4708 8360
rect 4468 8338 4764 8358
rect 9796 8414 10092 8434
rect 9852 8412 9876 8414
rect 9932 8412 9956 8414
rect 10012 8412 10036 8414
rect 9874 8360 9876 8412
rect 9938 8360 9950 8412
rect 10012 8360 10014 8412
rect 9852 8358 9876 8360
rect 9932 8358 9956 8360
rect 10012 8358 10036 8360
rect 9796 8338 10092 8358
rect 15124 8414 15420 8434
rect 15180 8412 15204 8414
rect 15260 8412 15284 8414
rect 15340 8412 15364 8414
rect 15202 8360 15204 8412
rect 15266 8360 15278 8412
rect 15340 8360 15342 8412
rect 15180 8358 15204 8360
rect 15260 8358 15284 8360
rect 15340 8358 15364 8360
rect 15124 8338 15420 8358
rect 20452 8414 20748 8434
rect 20508 8412 20532 8414
rect 20588 8412 20612 8414
rect 20668 8412 20692 8414
rect 20530 8360 20532 8412
rect 20594 8360 20606 8412
rect 20668 8360 20670 8412
rect 20508 8358 20532 8360
rect 20588 8358 20612 8360
rect 20668 8358 20692 8360
rect 20452 8338 20748 8358
rect 22626 8159 22654 8613
rect 22614 8153 22666 8159
rect 22614 8095 22666 8101
rect 3894 8079 3946 8085
rect 3894 8021 3946 8027
rect 3906 7641 3934 8021
rect 7132 7748 7428 7768
rect 7188 7746 7212 7748
rect 7268 7746 7292 7748
rect 7348 7746 7372 7748
rect 7210 7694 7212 7746
rect 7274 7694 7286 7746
rect 7348 7694 7350 7746
rect 7188 7692 7212 7694
rect 7268 7692 7292 7694
rect 7348 7692 7372 7694
rect 7132 7672 7428 7692
rect 12460 7748 12756 7768
rect 12516 7746 12540 7748
rect 12596 7746 12620 7748
rect 12676 7746 12700 7748
rect 12538 7694 12540 7746
rect 12602 7694 12614 7746
rect 12676 7694 12678 7746
rect 12516 7692 12540 7694
rect 12596 7692 12620 7694
rect 12676 7692 12700 7694
rect 12460 7672 12756 7692
rect 17788 7748 18084 7768
rect 17844 7746 17868 7748
rect 17924 7746 17948 7748
rect 18004 7746 18028 7748
rect 17866 7694 17868 7746
rect 17930 7694 17942 7746
rect 18004 7694 18006 7746
rect 17844 7692 17868 7694
rect 17924 7692 17948 7694
rect 18004 7692 18028 7694
rect 17788 7672 18084 7692
rect 3894 7635 3946 7641
rect 3894 7577 3946 7583
rect 22134 7339 22186 7345
rect 22134 7281 22186 7287
rect 4468 7082 4764 7102
rect 4524 7080 4548 7082
rect 4604 7080 4628 7082
rect 4684 7080 4708 7082
rect 4546 7028 4548 7080
rect 4610 7028 4622 7080
rect 4684 7028 4686 7080
rect 4524 7026 4548 7028
rect 4604 7026 4628 7028
rect 4684 7026 4708 7028
rect 4468 7006 4764 7026
rect 9796 7082 10092 7102
rect 9852 7080 9876 7082
rect 9932 7080 9956 7082
rect 10012 7080 10036 7082
rect 9874 7028 9876 7080
rect 9938 7028 9950 7080
rect 10012 7028 10014 7080
rect 9852 7026 9876 7028
rect 9932 7026 9956 7028
rect 10012 7026 10036 7028
rect 9796 7006 10092 7026
rect 15124 7082 15420 7102
rect 15180 7080 15204 7082
rect 15260 7080 15284 7082
rect 15340 7080 15364 7082
rect 15202 7028 15204 7080
rect 15266 7028 15278 7080
rect 15340 7028 15342 7080
rect 15180 7026 15204 7028
rect 15260 7026 15284 7028
rect 15340 7026 15364 7028
rect 15124 7006 15420 7026
rect 20452 7082 20748 7102
rect 20508 7080 20532 7082
rect 20588 7080 20612 7082
rect 20668 7080 20692 7082
rect 20530 7028 20532 7080
rect 20594 7028 20606 7080
rect 20668 7028 20670 7080
rect 20508 7026 20532 7028
rect 20588 7026 20612 7028
rect 20668 7026 20692 7028
rect 20452 7006 20748 7026
rect 22146 6975 22174 7281
rect 22134 6969 22186 6975
rect 22134 6911 22186 6917
rect 3894 6747 3946 6753
rect 3894 6689 3946 6695
rect 3906 6309 3934 6689
rect 7132 6416 7428 6436
rect 7188 6414 7212 6416
rect 7268 6414 7292 6416
rect 7348 6414 7372 6416
rect 7210 6362 7212 6414
rect 7274 6362 7286 6414
rect 7348 6362 7350 6414
rect 7188 6360 7212 6362
rect 7268 6360 7292 6362
rect 7348 6360 7372 6362
rect 7132 6340 7428 6360
rect 12460 6416 12756 6436
rect 12516 6414 12540 6416
rect 12596 6414 12620 6416
rect 12676 6414 12700 6416
rect 12538 6362 12540 6414
rect 12602 6362 12614 6414
rect 12676 6362 12678 6414
rect 12516 6360 12540 6362
rect 12596 6360 12620 6362
rect 12676 6360 12700 6362
rect 12460 6340 12756 6360
rect 17788 6416 18084 6436
rect 17844 6414 17868 6416
rect 17924 6414 17948 6416
rect 18004 6414 18028 6416
rect 17866 6362 17868 6414
rect 17930 6362 17942 6414
rect 18004 6362 18006 6414
rect 17844 6360 17868 6362
rect 17924 6360 17948 6362
rect 18004 6360 18028 6362
rect 17788 6340 18084 6360
rect 3894 6303 3946 6309
rect 3894 6245 3946 6251
rect 22614 6007 22666 6013
rect 22614 5949 22666 5955
rect 4468 5750 4764 5770
rect 4524 5748 4548 5750
rect 4604 5748 4628 5750
rect 4684 5748 4708 5750
rect 4546 5696 4548 5748
rect 4610 5696 4622 5748
rect 4684 5696 4686 5748
rect 4524 5694 4548 5696
rect 4604 5694 4628 5696
rect 4684 5694 4708 5696
rect 4468 5674 4764 5694
rect 9796 5750 10092 5770
rect 9852 5748 9876 5750
rect 9932 5748 9956 5750
rect 10012 5748 10036 5750
rect 9874 5696 9876 5748
rect 9938 5696 9950 5748
rect 10012 5696 10014 5748
rect 9852 5694 9876 5696
rect 9932 5694 9956 5696
rect 10012 5694 10036 5696
rect 9796 5674 10092 5694
rect 15124 5750 15420 5770
rect 15180 5748 15204 5750
rect 15260 5748 15284 5750
rect 15340 5748 15364 5750
rect 15202 5696 15204 5748
rect 15266 5696 15278 5748
rect 15340 5696 15342 5748
rect 15180 5694 15204 5696
rect 15260 5694 15284 5696
rect 15340 5694 15364 5696
rect 15124 5674 15420 5694
rect 20452 5750 20748 5770
rect 20508 5748 20532 5750
rect 20588 5748 20612 5750
rect 20668 5748 20692 5750
rect 20530 5696 20532 5748
rect 20594 5696 20606 5748
rect 20668 5696 20670 5748
rect 20508 5694 20532 5696
rect 20588 5694 20612 5696
rect 20668 5694 20692 5696
rect 20452 5674 20748 5694
rect 22626 5643 22654 5949
rect 22614 5637 22666 5643
rect 22614 5579 22666 5585
rect 3894 5415 3946 5421
rect 3894 5357 3946 5363
rect 3906 4977 3934 5357
rect 7132 5084 7428 5104
rect 7188 5082 7212 5084
rect 7268 5082 7292 5084
rect 7348 5082 7372 5084
rect 7210 5030 7212 5082
rect 7274 5030 7286 5082
rect 7348 5030 7350 5082
rect 7188 5028 7212 5030
rect 7268 5028 7292 5030
rect 7348 5028 7372 5030
rect 7132 5008 7428 5028
rect 12460 5084 12756 5104
rect 12516 5082 12540 5084
rect 12596 5082 12620 5084
rect 12676 5082 12700 5084
rect 12538 5030 12540 5082
rect 12602 5030 12614 5082
rect 12676 5030 12678 5082
rect 12516 5028 12540 5030
rect 12596 5028 12620 5030
rect 12676 5028 12700 5030
rect 12460 5008 12756 5028
rect 17788 5084 18084 5104
rect 17844 5082 17868 5084
rect 17924 5082 17948 5084
rect 18004 5082 18028 5084
rect 17866 5030 17868 5082
rect 17930 5030 17942 5082
rect 18004 5030 18006 5082
rect 17844 5028 17868 5030
rect 17924 5028 17948 5030
rect 18004 5028 18028 5030
rect 17788 5008 18084 5028
rect 3894 4971 3946 4977
rect 3894 4913 3946 4919
rect 22614 4675 22666 4681
rect 22614 4617 22666 4623
rect 4468 4418 4764 4438
rect 4524 4416 4548 4418
rect 4604 4416 4628 4418
rect 4684 4416 4708 4418
rect 4546 4364 4548 4416
rect 4610 4364 4622 4416
rect 4684 4364 4686 4416
rect 4524 4362 4548 4364
rect 4604 4362 4628 4364
rect 4684 4362 4708 4364
rect 4468 4342 4764 4362
rect 9796 4418 10092 4438
rect 9852 4416 9876 4418
rect 9932 4416 9956 4418
rect 10012 4416 10036 4418
rect 9874 4364 9876 4416
rect 9938 4364 9950 4416
rect 10012 4364 10014 4416
rect 9852 4362 9876 4364
rect 9932 4362 9956 4364
rect 10012 4362 10036 4364
rect 9796 4342 10092 4362
rect 15124 4418 15420 4438
rect 15180 4416 15204 4418
rect 15260 4416 15284 4418
rect 15340 4416 15364 4418
rect 15202 4364 15204 4416
rect 15266 4364 15278 4416
rect 15340 4364 15342 4416
rect 15180 4362 15204 4364
rect 15260 4362 15284 4364
rect 15340 4362 15364 4364
rect 15124 4342 15420 4362
rect 20452 4418 20748 4438
rect 20508 4416 20532 4418
rect 20588 4416 20612 4418
rect 20668 4416 20692 4418
rect 20530 4364 20532 4416
rect 20594 4364 20606 4416
rect 20668 4364 20670 4416
rect 20508 4362 20532 4364
rect 20588 4362 20612 4364
rect 20668 4362 20692 4364
rect 20452 4342 20748 4362
rect 22626 4311 22654 4617
rect 22614 4305 22666 4311
rect 22614 4247 22666 4253
rect 3894 4083 3946 4089
rect 3894 4025 3946 4031
rect 3906 3571 3934 4025
rect 7132 3752 7428 3772
rect 7188 3750 7212 3752
rect 7268 3750 7292 3752
rect 7348 3750 7372 3752
rect 7210 3698 7212 3750
rect 7274 3698 7286 3750
rect 7348 3698 7350 3750
rect 7188 3696 7212 3698
rect 7268 3696 7292 3698
rect 7348 3696 7372 3698
rect 7132 3676 7428 3696
rect 12460 3752 12756 3772
rect 12516 3750 12540 3752
rect 12596 3750 12620 3752
rect 12676 3750 12700 3752
rect 12538 3698 12540 3750
rect 12602 3698 12614 3750
rect 12676 3698 12678 3750
rect 12516 3696 12540 3698
rect 12596 3696 12620 3698
rect 12676 3696 12700 3698
rect 12460 3676 12756 3696
rect 17788 3752 18084 3772
rect 17844 3750 17868 3752
rect 17924 3750 17948 3752
rect 18004 3750 18028 3752
rect 17866 3698 17868 3750
rect 17930 3698 17942 3750
rect 18004 3698 18006 3750
rect 17844 3696 17868 3698
rect 17924 3696 17948 3698
rect 18004 3696 18028 3698
rect 17788 3676 18084 3696
rect 3894 3565 3946 3571
rect 3894 3507 3946 3513
rect 22614 3343 22666 3349
rect 22614 3285 22666 3291
rect 4468 3086 4764 3106
rect 4524 3084 4548 3086
rect 4604 3084 4628 3086
rect 4684 3084 4708 3086
rect 4546 3032 4548 3084
rect 4610 3032 4622 3084
rect 4684 3032 4686 3084
rect 4524 3030 4548 3032
rect 4604 3030 4628 3032
rect 4684 3030 4708 3032
rect 4468 3010 4764 3030
rect 9796 3086 10092 3106
rect 9852 3084 9876 3086
rect 9932 3084 9956 3086
rect 10012 3084 10036 3086
rect 9874 3032 9876 3084
rect 9938 3032 9950 3084
rect 10012 3032 10014 3084
rect 9852 3030 9876 3032
rect 9932 3030 9956 3032
rect 10012 3030 10036 3032
rect 9796 3010 10092 3030
rect 15124 3086 15420 3106
rect 15180 3084 15204 3086
rect 15260 3084 15284 3086
rect 15340 3084 15364 3086
rect 15202 3032 15204 3084
rect 15266 3032 15278 3084
rect 15340 3032 15342 3084
rect 15180 3030 15204 3032
rect 15260 3030 15284 3032
rect 15340 3030 15364 3032
rect 15124 3010 15420 3030
rect 20452 3086 20748 3106
rect 20508 3084 20532 3086
rect 20588 3084 20612 3086
rect 20668 3084 20692 3086
rect 20530 3032 20532 3084
rect 20594 3032 20606 3084
rect 20668 3032 20670 3084
rect 20508 3030 20532 3032
rect 20588 3030 20612 3032
rect 20668 3030 20692 3032
rect 20452 3010 20748 3030
rect 22626 2831 22654 3285
rect 22614 2825 22666 2831
rect 22614 2767 22666 2773
rect 3894 2751 3946 2757
rect 3894 2693 3946 2699
rect 3906 2313 3934 2693
rect 7132 2420 7428 2440
rect 7188 2418 7212 2420
rect 7268 2418 7292 2420
rect 7348 2418 7372 2420
rect 7210 2366 7212 2418
rect 7274 2366 7286 2418
rect 7348 2366 7350 2418
rect 7188 2364 7212 2366
rect 7268 2364 7292 2366
rect 7348 2364 7372 2366
rect 7132 2344 7428 2364
rect 12460 2420 12756 2440
rect 12516 2418 12540 2420
rect 12596 2418 12620 2420
rect 12676 2418 12700 2420
rect 12538 2366 12540 2418
rect 12602 2366 12614 2418
rect 12676 2366 12678 2418
rect 12516 2364 12540 2366
rect 12596 2364 12620 2366
rect 12676 2364 12700 2366
rect 12460 2344 12756 2364
rect 17788 2420 18084 2440
rect 17844 2418 17868 2420
rect 17924 2418 17948 2420
rect 18004 2418 18028 2420
rect 17866 2366 17868 2418
rect 17930 2366 17942 2418
rect 18004 2366 18006 2418
rect 17844 2364 17868 2366
rect 17924 2364 17948 2366
rect 18004 2364 18028 2366
rect 17788 2344 18084 2364
rect 3894 2307 3946 2313
rect 3894 2249 3946 2255
rect 22134 2011 22186 2017
rect 22134 1953 22186 1959
rect 4468 1754 4764 1774
rect 4524 1752 4548 1754
rect 4604 1752 4628 1754
rect 4684 1752 4708 1754
rect 4546 1700 4548 1752
rect 4610 1700 4622 1752
rect 4684 1700 4686 1752
rect 4524 1698 4548 1700
rect 4604 1698 4628 1700
rect 4684 1698 4708 1700
rect 4468 1678 4764 1698
rect 9796 1754 10092 1774
rect 9852 1752 9876 1754
rect 9932 1752 9956 1754
rect 10012 1752 10036 1754
rect 9874 1700 9876 1752
rect 9938 1700 9950 1752
rect 10012 1700 10014 1752
rect 9852 1698 9876 1700
rect 9932 1698 9956 1700
rect 10012 1698 10036 1700
rect 9796 1678 10092 1698
rect 15124 1754 15420 1774
rect 15180 1752 15204 1754
rect 15260 1752 15284 1754
rect 15340 1752 15364 1754
rect 15202 1700 15204 1752
rect 15266 1700 15278 1752
rect 15340 1700 15342 1752
rect 15180 1698 15204 1700
rect 15260 1698 15284 1700
rect 15340 1698 15364 1700
rect 15124 1678 15420 1698
rect 20452 1754 20748 1774
rect 20508 1752 20532 1754
rect 20588 1752 20612 1754
rect 20668 1752 20692 1754
rect 20530 1700 20532 1752
rect 20594 1700 20606 1752
rect 20668 1700 20670 1752
rect 20508 1698 20532 1700
rect 20588 1698 20612 1700
rect 20668 1698 20692 1700
rect 20452 1678 20748 1698
rect 22146 1647 22174 1953
rect 22134 1641 22186 1647
rect 22134 1583 22186 1589
rect 2358 1419 2410 1425
rect 2358 1361 2410 1367
rect 3030 1419 3082 1425
rect 3030 1361 3082 1367
rect 3042 875 3070 1361
rect 7132 1088 7428 1108
rect 7188 1086 7212 1088
rect 7268 1086 7292 1088
rect 7348 1086 7372 1088
rect 7210 1034 7212 1086
rect 7274 1034 7286 1086
rect 7348 1034 7350 1086
rect 7188 1032 7212 1034
rect 7268 1032 7292 1034
rect 7348 1032 7372 1034
rect 7132 1012 7428 1032
rect 12460 1088 12756 1108
rect 12516 1086 12540 1088
rect 12596 1086 12620 1088
rect 12676 1086 12700 1088
rect 12538 1034 12540 1086
rect 12602 1034 12614 1086
rect 12676 1034 12678 1086
rect 12516 1032 12540 1034
rect 12596 1032 12620 1034
rect 12676 1032 12700 1034
rect 12460 1012 12756 1032
rect 17788 1088 18084 1108
rect 17844 1086 17868 1088
rect 17924 1086 17948 1088
rect 18004 1086 18028 1088
rect 17866 1034 17868 1086
rect 17930 1034 17942 1086
rect 18004 1034 18006 1086
rect 17844 1032 17868 1034
rect 17924 1032 17948 1034
rect 18004 1032 18028 1034
rect 17788 1012 18084 1032
rect 3028 866 3084 875
rect 3028 801 3084 810
<< via2 >>
rect 2740 27302 2796 27358
rect 4468 27060 4524 27062
rect 4548 27060 4604 27062
rect 4628 27060 4684 27062
rect 4708 27060 4764 27062
rect 4468 27008 4494 27060
rect 4494 27008 4524 27060
rect 4548 27008 4558 27060
rect 4558 27008 4604 27060
rect 4628 27008 4674 27060
rect 4674 27008 4684 27060
rect 4708 27008 4738 27060
rect 4738 27008 4764 27060
rect 4468 27006 4524 27008
rect 4548 27006 4604 27008
rect 4628 27006 4684 27008
rect 4708 27006 4764 27008
rect 9796 27060 9852 27062
rect 9876 27060 9932 27062
rect 9956 27060 10012 27062
rect 10036 27060 10092 27062
rect 9796 27008 9822 27060
rect 9822 27008 9852 27060
rect 9876 27008 9886 27060
rect 9886 27008 9932 27060
rect 9956 27008 10002 27060
rect 10002 27008 10012 27060
rect 10036 27008 10066 27060
rect 10066 27008 10092 27060
rect 9796 27006 9852 27008
rect 9876 27006 9932 27008
rect 9956 27006 10012 27008
rect 10036 27006 10092 27008
rect 15124 27060 15180 27062
rect 15204 27060 15260 27062
rect 15284 27060 15340 27062
rect 15364 27060 15420 27062
rect 15124 27008 15150 27060
rect 15150 27008 15180 27060
rect 15204 27008 15214 27060
rect 15214 27008 15260 27060
rect 15284 27008 15330 27060
rect 15330 27008 15340 27060
rect 15364 27008 15394 27060
rect 15394 27008 15420 27060
rect 15124 27006 15180 27008
rect 15204 27006 15260 27008
rect 15284 27006 15340 27008
rect 15364 27006 15420 27008
rect 20452 27060 20508 27062
rect 20532 27060 20588 27062
rect 20612 27060 20668 27062
rect 20692 27060 20748 27062
rect 20452 27008 20478 27060
rect 20478 27008 20508 27060
rect 20532 27008 20542 27060
rect 20542 27008 20588 27060
rect 20612 27008 20658 27060
rect 20658 27008 20668 27060
rect 20692 27008 20722 27060
rect 20722 27008 20748 27060
rect 20452 27006 20508 27008
rect 20532 27006 20588 27008
rect 20612 27006 20668 27008
rect 20692 27006 20748 27008
rect 7132 26394 7188 26396
rect 7212 26394 7268 26396
rect 7292 26394 7348 26396
rect 7372 26394 7428 26396
rect 7132 26342 7158 26394
rect 7158 26342 7188 26394
rect 7212 26342 7222 26394
rect 7222 26342 7268 26394
rect 7292 26342 7338 26394
rect 7338 26342 7348 26394
rect 7372 26342 7402 26394
rect 7402 26342 7428 26394
rect 7132 26340 7188 26342
rect 7212 26340 7268 26342
rect 7292 26340 7348 26342
rect 7372 26340 7428 26342
rect 12460 26394 12516 26396
rect 12540 26394 12596 26396
rect 12620 26394 12676 26396
rect 12700 26394 12756 26396
rect 12460 26342 12486 26394
rect 12486 26342 12516 26394
rect 12540 26342 12550 26394
rect 12550 26342 12596 26394
rect 12620 26342 12666 26394
rect 12666 26342 12676 26394
rect 12700 26342 12730 26394
rect 12730 26342 12756 26394
rect 12460 26340 12516 26342
rect 12540 26340 12596 26342
rect 12620 26340 12676 26342
rect 12700 26340 12756 26342
rect 17788 26394 17844 26396
rect 17868 26394 17924 26396
rect 17948 26394 18004 26396
rect 18028 26394 18084 26396
rect 17788 26342 17814 26394
rect 17814 26342 17844 26394
rect 17868 26342 17878 26394
rect 17878 26342 17924 26394
rect 17948 26342 17994 26394
rect 17994 26342 18004 26394
rect 18028 26342 18058 26394
rect 18058 26342 18084 26394
rect 17788 26340 17844 26342
rect 17868 26340 17924 26342
rect 17948 26340 18004 26342
rect 18028 26340 18084 26342
rect 2356 26118 2412 26174
rect 4468 25728 4524 25730
rect 4548 25728 4604 25730
rect 4628 25728 4684 25730
rect 4708 25728 4764 25730
rect 4468 25676 4494 25728
rect 4494 25676 4524 25728
rect 4548 25676 4558 25728
rect 4558 25676 4604 25728
rect 4628 25676 4674 25728
rect 4674 25676 4684 25728
rect 4708 25676 4738 25728
rect 4738 25676 4764 25728
rect 4468 25674 4524 25676
rect 4548 25674 4604 25676
rect 4628 25674 4684 25676
rect 4708 25674 4764 25676
rect 9796 25728 9852 25730
rect 9876 25728 9932 25730
rect 9956 25728 10012 25730
rect 10036 25728 10092 25730
rect 9796 25676 9822 25728
rect 9822 25676 9852 25728
rect 9876 25676 9886 25728
rect 9886 25676 9932 25728
rect 9956 25676 10002 25728
rect 10002 25676 10012 25728
rect 10036 25676 10066 25728
rect 10066 25676 10092 25728
rect 9796 25674 9852 25676
rect 9876 25674 9932 25676
rect 9956 25674 10012 25676
rect 10036 25674 10092 25676
rect 15124 25728 15180 25730
rect 15204 25728 15260 25730
rect 15284 25728 15340 25730
rect 15364 25728 15420 25730
rect 15124 25676 15150 25728
rect 15150 25676 15180 25728
rect 15204 25676 15214 25728
rect 15214 25676 15260 25728
rect 15284 25676 15330 25728
rect 15330 25676 15340 25728
rect 15364 25676 15394 25728
rect 15394 25676 15420 25728
rect 15124 25674 15180 25676
rect 15204 25674 15260 25676
rect 15284 25674 15340 25676
rect 15364 25674 15420 25676
rect 20452 25728 20508 25730
rect 20532 25728 20588 25730
rect 20612 25728 20668 25730
rect 20692 25728 20748 25730
rect 20452 25676 20478 25728
rect 20478 25676 20508 25728
rect 20532 25676 20542 25728
rect 20542 25676 20588 25728
rect 20612 25676 20658 25728
rect 20658 25676 20668 25728
rect 20692 25676 20722 25728
rect 20722 25676 20748 25728
rect 20452 25674 20508 25676
rect 20532 25674 20588 25676
rect 20612 25674 20668 25676
rect 20692 25674 20748 25676
rect 2452 25526 2508 25582
rect 7132 25062 7188 25064
rect 7212 25062 7268 25064
rect 7292 25062 7348 25064
rect 7372 25062 7428 25064
rect 7132 25010 7158 25062
rect 7158 25010 7188 25062
rect 7212 25010 7222 25062
rect 7222 25010 7268 25062
rect 7292 25010 7338 25062
rect 7338 25010 7348 25062
rect 7372 25010 7402 25062
rect 7402 25010 7428 25062
rect 7132 25008 7188 25010
rect 7212 25008 7268 25010
rect 7292 25008 7348 25010
rect 7372 25008 7428 25010
rect 12460 25062 12516 25064
rect 12540 25062 12596 25064
rect 12620 25062 12676 25064
rect 12700 25062 12756 25064
rect 12460 25010 12486 25062
rect 12486 25010 12516 25062
rect 12540 25010 12550 25062
rect 12550 25010 12596 25062
rect 12620 25010 12666 25062
rect 12666 25010 12676 25062
rect 12700 25010 12730 25062
rect 12730 25010 12756 25062
rect 12460 25008 12516 25010
rect 12540 25008 12596 25010
rect 12620 25008 12676 25010
rect 12700 25008 12756 25010
rect 17788 25062 17844 25064
rect 17868 25062 17924 25064
rect 17948 25062 18004 25064
rect 18028 25062 18084 25064
rect 17788 25010 17814 25062
rect 17814 25010 17844 25062
rect 17868 25010 17878 25062
rect 17878 25010 17924 25062
rect 17948 25010 17994 25062
rect 17994 25010 18004 25062
rect 18028 25010 18058 25062
rect 18058 25010 18084 25062
rect 17788 25008 17844 25010
rect 17868 25008 17924 25010
rect 17948 25008 18004 25010
rect 18028 25008 18084 25010
rect 2068 24677 2070 24694
rect 2070 24677 2122 24694
rect 2122 24677 2124 24694
rect 2068 24638 2124 24677
rect 4468 24396 4524 24398
rect 4548 24396 4604 24398
rect 4628 24396 4684 24398
rect 4708 24396 4764 24398
rect 4468 24344 4494 24396
rect 4494 24344 4524 24396
rect 4548 24344 4558 24396
rect 4558 24344 4604 24396
rect 4628 24344 4674 24396
rect 4674 24344 4684 24396
rect 4708 24344 4738 24396
rect 4738 24344 4764 24396
rect 4468 24342 4524 24344
rect 4548 24342 4604 24344
rect 4628 24342 4684 24344
rect 4708 24342 4764 24344
rect 9796 24396 9852 24398
rect 9876 24396 9932 24398
rect 9956 24396 10012 24398
rect 10036 24396 10092 24398
rect 9796 24344 9822 24396
rect 9822 24344 9852 24396
rect 9876 24344 9886 24396
rect 9886 24344 9932 24396
rect 9956 24344 10002 24396
rect 10002 24344 10012 24396
rect 10036 24344 10066 24396
rect 10066 24344 10092 24396
rect 9796 24342 9852 24344
rect 9876 24342 9932 24344
rect 9956 24342 10012 24344
rect 10036 24342 10092 24344
rect 15124 24396 15180 24398
rect 15204 24396 15260 24398
rect 15284 24396 15340 24398
rect 15364 24396 15420 24398
rect 15124 24344 15150 24396
rect 15150 24344 15180 24396
rect 15204 24344 15214 24396
rect 15214 24344 15260 24396
rect 15284 24344 15330 24396
rect 15330 24344 15340 24396
rect 15364 24344 15394 24396
rect 15394 24344 15420 24396
rect 15124 24342 15180 24344
rect 15204 24342 15260 24344
rect 15284 24342 15340 24344
rect 15364 24342 15420 24344
rect 20452 24396 20508 24398
rect 20532 24396 20588 24398
rect 20612 24396 20668 24398
rect 20692 24396 20748 24398
rect 20452 24344 20478 24396
rect 20478 24344 20508 24396
rect 20532 24344 20542 24396
rect 20542 24344 20588 24396
rect 20612 24344 20658 24396
rect 20658 24344 20668 24396
rect 20692 24344 20722 24396
rect 20722 24344 20748 24396
rect 20452 24342 20508 24344
rect 20532 24342 20588 24344
rect 20612 24342 20668 24344
rect 20692 24342 20748 24344
rect 7132 23730 7188 23732
rect 7212 23730 7268 23732
rect 7292 23730 7348 23732
rect 7372 23730 7428 23732
rect 7132 23678 7158 23730
rect 7158 23678 7188 23730
rect 7212 23678 7222 23730
rect 7222 23678 7268 23730
rect 7292 23678 7338 23730
rect 7338 23678 7348 23730
rect 7372 23678 7402 23730
rect 7402 23678 7428 23730
rect 7132 23676 7188 23678
rect 7212 23676 7268 23678
rect 7292 23676 7348 23678
rect 7372 23676 7428 23678
rect 12460 23730 12516 23732
rect 12540 23730 12596 23732
rect 12620 23730 12676 23732
rect 12700 23730 12756 23732
rect 12460 23678 12486 23730
rect 12486 23678 12516 23730
rect 12540 23678 12550 23730
rect 12550 23678 12596 23730
rect 12620 23678 12666 23730
rect 12666 23678 12676 23730
rect 12700 23678 12730 23730
rect 12730 23678 12756 23730
rect 12460 23676 12516 23678
rect 12540 23676 12596 23678
rect 12620 23676 12676 23678
rect 12700 23676 12756 23678
rect 17788 23730 17844 23732
rect 17868 23730 17924 23732
rect 17948 23730 18004 23732
rect 18028 23730 18084 23732
rect 17788 23678 17814 23730
rect 17814 23678 17844 23730
rect 17868 23678 17878 23730
rect 17878 23678 17924 23730
rect 17948 23678 17994 23730
rect 17994 23678 18004 23730
rect 18028 23678 18058 23730
rect 18058 23678 18084 23730
rect 17788 23676 17844 23678
rect 17868 23676 17924 23678
rect 17948 23676 18004 23678
rect 18028 23676 18084 23678
rect 2068 23345 2070 23362
rect 2070 23345 2122 23362
rect 2122 23345 2124 23362
rect 2068 23306 2124 23345
rect 4468 23064 4524 23066
rect 4548 23064 4604 23066
rect 4628 23064 4684 23066
rect 4708 23064 4764 23066
rect 4468 23012 4494 23064
rect 4494 23012 4524 23064
rect 4548 23012 4558 23064
rect 4558 23012 4604 23064
rect 4628 23012 4674 23064
rect 4674 23012 4684 23064
rect 4708 23012 4738 23064
rect 4738 23012 4764 23064
rect 4468 23010 4524 23012
rect 4548 23010 4604 23012
rect 4628 23010 4684 23012
rect 4708 23010 4764 23012
rect 9796 23064 9852 23066
rect 9876 23064 9932 23066
rect 9956 23064 10012 23066
rect 10036 23064 10092 23066
rect 9796 23012 9822 23064
rect 9822 23012 9852 23064
rect 9876 23012 9886 23064
rect 9886 23012 9932 23064
rect 9956 23012 10002 23064
rect 10002 23012 10012 23064
rect 10036 23012 10066 23064
rect 10066 23012 10092 23064
rect 9796 23010 9852 23012
rect 9876 23010 9932 23012
rect 9956 23010 10012 23012
rect 10036 23010 10092 23012
rect 15124 23064 15180 23066
rect 15204 23064 15260 23066
rect 15284 23064 15340 23066
rect 15364 23064 15420 23066
rect 15124 23012 15150 23064
rect 15150 23012 15180 23064
rect 15204 23012 15214 23064
rect 15214 23012 15260 23064
rect 15284 23012 15330 23064
rect 15330 23012 15340 23064
rect 15364 23012 15394 23064
rect 15394 23012 15420 23064
rect 15124 23010 15180 23012
rect 15204 23010 15260 23012
rect 15284 23010 15340 23012
rect 15364 23010 15420 23012
rect 20452 23064 20508 23066
rect 20532 23064 20588 23066
rect 20612 23064 20668 23066
rect 20692 23064 20748 23066
rect 20452 23012 20478 23064
rect 20478 23012 20508 23064
rect 20532 23012 20542 23064
rect 20542 23012 20588 23064
rect 20612 23012 20658 23064
rect 20658 23012 20668 23064
rect 20692 23012 20722 23064
rect 20722 23012 20748 23064
rect 20452 23010 20508 23012
rect 20532 23010 20588 23012
rect 20612 23010 20668 23012
rect 20692 23010 20748 23012
rect 7132 22398 7188 22400
rect 7212 22398 7268 22400
rect 7292 22398 7348 22400
rect 7372 22398 7428 22400
rect 7132 22346 7158 22398
rect 7158 22346 7188 22398
rect 7212 22346 7222 22398
rect 7222 22346 7268 22398
rect 7292 22346 7338 22398
rect 7338 22346 7348 22398
rect 7372 22346 7402 22398
rect 7402 22346 7428 22398
rect 7132 22344 7188 22346
rect 7212 22344 7268 22346
rect 7292 22344 7348 22346
rect 7372 22344 7428 22346
rect 12460 22398 12516 22400
rect 12540 22398 12596 22400
rect 12620 22398 12676 22400
rect 12700 22398 12756 22400
rect 12460 22346 12486 22398
rect 12486 22346 12516 22398
rect 12540 22346 12550 22398
rect 12550 22346 12596 22398
rect 12620 22346 12666 22398
rect 12666 22346 12676 22398
rect 12700 22346 12730 22398
rect 12730 22346 12756 22398
rect 12460 22344 12516 22346
rect 12540 22344 12596 22346
rect 12620 22344 12676 22346
rect 12700 22344 12756 22346
rect 17788 22398 17844 22400
rect 17868 22398 17924 22400
rect 17948 22398 18004 22400
rect 18028 22398 18084 22400
rect 17788 22346 17814 22398
rect 17814 22346 17844 22398
rect 17868 22346 17878 22398
rect 17878 22346 17924 22398
rect 17948 22346 17994 22398
rect 17994 22346 18004 22398
rect 18028 22346 18058 22398
rect 18058 22346 18084 22398
rect 17788 22344 17844 22346
rect 17868 22344 17924 22346
rect 17948 22344 18004 22346
rect 18028 22344 18084 22346
rect 2068 21826 2124 21882
rect 4468 21732 4524 21734
rect 4548 21732 4604 21734
rect 4628 21732 4684 21734
rect 4708 21732 4764 21734
rect 4468 21680 4494 21732
rect 4494 21680 4524 21732
rect 4548 21680 4558 21732
rect 4558 21680 4604 21732
rect 4628 21680 4674 21732
rect 4674 21680 4684 21732
rect 4708 21680 4738 21732
rect 4738 21680 4764 21732
rect 4468 21678 4524 21680
rect 4548 21678 4604 21680
rect 4628 21678 4684 21680
rect 4708 21678 4764 21680
rect 9796 21732 9852 21734
rect 9876 21732 9932 21734
rect 9956 21732 10012 21734
rect 10036 21732 10092 21734
rect 9796 21680 9822 21732
rect 9822 21680 9852 21732
rect 9876 21680 9886 21732
rect 9886 21680 9932 21732
rect 9956 21680 10002 21732
rect 10002 21680 10012 21732
rect 10036 21680 10066 21732
rect 10066 21680 10092 21732
rect 9796 21678 9852 21680
rect 9876 21678 9932 21680
rect 9956 21678 10012 21680
rect 10036 21678 10092 21680
rect 15124 21732 15180 21734
rect 15204 21732 15260 21734
rect 15284 21732 15340 21734
rect 15364 21732 15420 21734
rect 15124 21680 15150 21732
rect 15150 21680 15180 21732
rect 15204 21680 15214 21732
rect 15214 21680 15260 21732
rect 15284 21680 15330 21732
rect 15330 21680 15340 21732
rect 15364 21680 15394 21732
rect 15394 21680 15420 21732
rect 15124 21678 15180 21680
rect 15204 21678 15260 21680
rect 15284 21678 15340 21680
rect 15364 21678 15420 21680
rect 20452 21732 20508 21734
rect 20532 21732 20588 21734
rect 20612 21732 20668 21734
rect 20692 21732 20748 21734
rect 20452 21680 20478 21732
rect 20478 21680 20508 21732
rect 20532 21680 20542 21732
rect 20542 21680 20588 21732
rect 20612 21680 20658 21732
rect 20658 21680 20668 21732
rect 20692 21680 20722 21732
rect 20722 21680 20748 21732
rect 20452 21678 20508 21680
rect 20532 21678 20588 21680
rect 20612 21678 20668 21680
rect 20692 21678 20748 21680
rect 7132 21066 7188 21068
rect 7212 21066 7268 21068
rect 7292 21066 7348 21068
rect 7372 21066 7428 21068
rect 7132 21014 7158 21066
rect 7158 21014 7188 21066
rect 7212 21014 7222 21066
rect 7222 21014 7268 21066
rect 7292 21014 7338 21066
rect 7338 21014 7348 21066
rect 7372 21014 7402 21066
rect 7402 21014 7428 21066
rect 7132 21012 7188 21014
rect 7212 21012 7268 21014
rect 7292 21012 7348 21014
rect 7372 21012 7428 21014
rect 12460 21066 12516 21068
rect 12540 21066 12596 21068
rect 12620 21066 12676 21068
rect 12700 21066 12756 21068
rect 12460 21014 12486 21066
rect 12486 21014 12516 21066
rect 12540 21014 12550 21066
rect 12550 21014 12596 21066
rect 12620 21014 12666 21066
rect 12666 21014 12676 21066
rect 12700 21014 12730 21066
rect 12730 21014 12756 21066
rect 12460 21012 12516 21014
rect 12540 21012 12596 21014
rect 12620 21012 12676 21014
rect 12700 21012 12756 21014
rect 17788 21066 17844 21068
rect 17868 21066 17924 21068
rect 17948 21066 18004 21068
rect 18028 21066 18084 21068
rect 17788 21014 17814 21066
rect 17814 21014 17844 21066
rect 17868 21014 17878 21066
rect 17878 21014 17924 21066
rect 17948 21014 17994 21066
rect 17994 21014 18004 21066
rect 18028 21014 18058 21066
rect 18058 21014 18084 21066
rect 17788 21012 17844 21014
rect 17868 21012 17924 21014
rect 17948 21012 18004 21014
rect 18028 21012 18084 21014
rect 4468 20400 4524 20402
rect 4548 20400 4604 20402
rect 4628 20400 4684 20402
rect 4708 20400 4764 20402
rect 4468 20348 4494 20400
rect 4494 20348 4524 20400
rect 4548 20348 4558 20400
rect 4558 20348 4604 20400
rect 4628 20348 4674 20400
rect 4674 20348 4684 20400
rect 4708 20348 4738 20400
rect 4738 20348 4764 20400
rect 4468 20346 4524 20348
rect 4548 20346 4604 20348
rect 4628 20346 4684 20348
rect 4708 20346 4764 20348
rect 9796 20400 9852 20402
rect 9876 20400 9932 20402
rect 9956 20400 10012 20402
rect 10036 20400 10092 20402
rect 9796 20348 9822 20400
rect 9822 20348 9852 20400
rect 9876 20348 9886 20400
rect 9886 20348 9932 20400
rect 9956 20348 10002 20400
rect 10002 20348 10012 20400
rect 10036 20348 10066 20400
rect 10066 20348 10092 20400
rect 9796 20346 9852 20348
rect 9876 20346 9932 20348
rect 9956 20346 10012 20348
rect 10036 20346 10092 20348
rect 15124 20400 15180 20402
rect 15204 20400 15260 20402
rect 15284 20400 15340 20402
rect 15364 20400 15420 20402
rect 15124 20348 15150 20400
rect 15150 20348 15180 20400
rect 15204 20348 15214 20400
rect 15214 20348 15260 20400
rect 15284 20348 15330 20400
rect 15330 20348 15340 20400
rect 15364 20348 15394 20400
rect 15394 20348 15420 20400
rect 15124 20346 15180 20348
rect 15204 20346 15260 20348
rect 15284 20346 15340 20348
rect 15364 20346 15420 20348
rect 20452 20400 20508 20402
rect 20532 20400 20588 20402
rect 20612 20400 20668 20402
rect 20692 20400 20748 20402
rect 20452 20348 20478 20400
rect 20478 20348 20508 20400
rect 20532 20348 20542 20400
rect 20542 20348 20588 20400
rect 20612 20348 20658 20400
rect 20658 20348 20668 20400
rect 20692 20348 20722 20400
rect 20722 20348 20748 20400
rect 20452 20346 20508 20348
rect 20532 20346 20588 20348
rect 20612 20346 20668 20348
rect 20692 20346 20748 20348
rect 2452 20050 2508 20106
rect 7132 19734 7188 19736
rect 7212 19734 7268 19736
rect 7292 19734 7348 19736
rect 7372 19734 7428 19736
rect 7132 19682 7158 19734
rect 7158 19682 7188 19734
rect 7212 19682 7222 19734
rect 7222 19682 7268 19734
rect 7292 19682 7338 19734
rect 7338 19682 7348 19734
rect 7372 19682 7402 19734
rect 7402 19682 7428 19734
rect 7132 19680 7188 19682
rect 7212 19680 7268 19682
rect 7292 19680 7348 19682
rect 7372 19680 7428 19682
rect 12460 19734 12516 19736
rect 12540 19734 12596 19736
rect 12620 19734 12676 19736
rect 12700 19734 12756 19736
rect 12460 19682 12486 19734
rect 12486 19682 12516 19734
rect 12540 19682 12550 19734
rect 12550 19682 12596 19734
rect 12620 19682 12666 19734
rect 12666 19682 12676 19734
rect 12700 19682 12730 19734
rect 12730 19682 12756 19734
rect 12460 19680 12516 19682
rect 12540 19680 12596 19682
rect 12620 19680 12676 19682
rect 12700 19680 12756 19682
rect 17788 19734 17844 19736
rect 17868 19734 17924 19736
rect 17948 19734 18004 19736
rect 18028 19734 18084 19736
rect 17788 19682 17814 19734
rect 17814 19682 17844 19734
rect 17868 19682 17878 19734
rect 17878 19682 17924 19734
rect 17948 19682 17994 19734
rect 17994 19682 18004 19734
rect 18028 19682 18058 19734
rect 18058 19682 18084 19734
rect 17788 19680 17844 19682
rect 17868 19680 17924 19682
rect 17948 19680 18004 19682
rect 18028 19680 18084 19682
rect 2068 19349 2070 19366
rect 2070 19349 2122 19366
rect 2122 19349 2124 19366
rect 2068 19310 2124 19349
rect 4468 19068 4524 19070
rect 4548 19068 4604 19070
rect 4628 19068 4684 19070
rect 4708 19068 4764 19070
rect 4468 19016 4494 19068
rect 4494 19016 4524 19068
rect 4548 19016 4558 19068
rect 4558 19016 4604 19068
rect 4628 19016 4674 19068
rect 4674 19016 4684 19068
rect 4708 19016 4738 19068
rect 4738 19016 4764 19068
rect 4468 19014 4524 19016
rect 4548 19014 4604 19016
rect 4628 19014 4684 19016
rect 4708 19014 4764 19016
rect 9796 19068 9852 19070
rect 9876 19068 9932 19070
rect 9956 19068 10012 19070
rect 10036 19068 10092 19070
rect 9796 19016 9822 19068
rect 9822 19016 9852 19068
rect 9876 19016 9886 19068
rect 9886 19016 9932 19068
rect 9956 19016 10002 19068
rect 10002 19016 10012 19068
rect 10036 19016 10066 19068
rect 10066 19016 10092 19068
rect 9796 19014 9852 19016
rect 9876 19014 9932 19016
rect 9956 19014 10012 19016
rect 10036 19014 10092 19016
rect 15124 19068 15180 19070
rect 15204 19068 15260 19070
rect 15284 19068 15340 19070
rect 15364 19068 15420 19070
rect 15124 19016 15150 19068
rect 15150 19016 15180 19068
rect 15204 19016 15214 19068
rect 15214 19016 15260 19068
rect 15284 19016 15330 19068
rect 15330 19016 15340 19068
rect 15364 19016 15394 19068
rect 15394 19016 15420 19068
rect 15124 19014 15180 19016
rect 15204 19014 15260 19016
rect 15284 19014 15340 19016
rect 15364 19014 15420 19016
rect 20452 19068 20508 19070
rect 20532 19068 20588 19070
rect 20612 19068 20668 19070
rect 20692 19068 20748 19070
rect 20452 19016 20478 19068
rect 20478 19016 20508 19068
rect 20532 19016 20542 19068
rect 20542 19016 20588 19068
rect 20612 19016 20658 19068
rect 20658 19016 20668 19068
rect 20692 19016 20722 19068
rect 20722 19016 20748 19068
rect 20452 19014 20508 19016
rect 20532 19014 20588 19016
rect 20612 19014 20668 19016
rect 20692 19014 20748 19016
rect 7132 18402 7188 18404
rect 7212 18402 7268 18404
rect 7292 18402 7348 18404
rect 7372 18402 7428 18404
rect 7132 18350 7158 18402
rect 7158 18350 7188 18402
rect 7212 18350 7222 18402
rect 7222 18350 7268 18402
rect 7292 18350 7338 18402
rect 7338 18350 7348 18402
rect 7372 18350 7402 18402
rect 7402 18350 7428 18402
rect 7132 18348 7188 18350
rect 7212 18348 7268 18350
rect 7292 18348 7348 18350
rect 7372 18348 7428 18350
rect 12460 18402 12516 18404
rect 12540 18402 12596 18404
rect 12620 18402 12676 18404
rect 12700 18402 12756 18404
rect 12460 18350 12486 18402
rect 12486 18350 12516 18402
rect 12540 18350 12550 18402
rect 12550 18350 12596 18402
rect 12620 18350 12666 18402
rect 12666 18350 12676 18402
rect 12700 18350 12730 18402
rect 12730 18350 12756 18402
rect 12460 18348 12516 18350
rect 12540 18348 12596 18350
rect 12620 18348 12676 18350
rect 12700 18348 12756 18350
rect 17788 18402 17844 18404
rect 17868 18402 17924 18404
rect 17948 18402 18004 18404
rect 18028 18402 18084 18404
rect 17788 18350 17814 18402
rect 17814 18350 17844 18402
rect 17868 18350 17878 18402
rect 17878 18350 17924 18402
rect 17948 18350 17994 18402
rect 17994 18350 18004 18402
rect 18028 18350 18058 18402
rect 18058 18350 18084 18402
rect 17788 18348 17844 18350
rect 17868 18348 17924 18350
rect 17948 18348 18004 18350
rect 18028 18348 18084 18350
rect 4468 17736 4524 17738
rect 4548 17736 4604 17738
rect 4628 17736 4684 17738
rect 4708 17736 4764 17738
rect 4468 17684 4494 17736
rect 4494 17684 4524 17736
rect 4548 17684 4558 17736
rect 4558 17684 4604 17736
rect 4628 17684 4674 17736
rect 4674 17684 4684 17736
rect 4708 17684 4738 17736
rect 4738 17684 4764 17736
rect 4468 17682 4524 17684
rect 4548 17682 4604 17684
rect 4628 17682 4684 17684
rect 4708 17682 4764 17684
rect 9796 17736 9852 17738
rect 9876 17736 9932 17738
rect 9956 17736 10012 17738
rect 10036 17736 10092 17738
rect 9796 17684 9822 17736
rect 9822 17684 9852 17736
rect 9876 17684 9886 17736
rect 9886 17684 9932 17736
rect 9956 17684 10002 17736
rect 10002 17684 10012 17736
rect 10036 17684 10066 17736
rect 10066 17684 10092 17736
rect 9796 17682 9852 17684
rect 9876 17682 9932 17684
rect 9956 17682 10012 17684
rect 10036 17682 10092 17684
rect 15124 17736 15180 17738
rect 15204 17736 15260 17738
rect 15284 17736 15340 17738
rect 15364 17736 15420 17738
rect 15124 17684 15150 17736
rect 15150 17684 15180 17736
rect 15204 17684 15214 17736
rect 15214 17684 15260 17736
rect 15284 17684 15330 17736
rect 15330 17684 15340 17736
rect 15364 17684 15394 17736
rect 15394 17684 15420 17736
rect 15124 17682 15180 17684
rect 15204 17682 15260 17684
rect 15284 17682 15340 17684
rect 15364 17682 15420 17684
rect 20452 17736 20508 17738
rect 20532 17736 20588 17738
rect 20612 17736 20668 17738
rect 20692 17736 20748 17738
rect 20452 17684 20478 17736
rect 20478 17684 20508 17736
rect 20532 17684 20542 17736
rect 20542 17684 20588 17736
rect 20612 17684 20658 17736
rect 20658 17684 20668 17736
rect 20692 17684 20722 17736
rect 20722 17684 20748 17736
rect 20452 17682 20508 17684
rect 20532 17682 20588 17684
rect 20612 17682 20668 17684
rect 20692 17682 20748 17684
rect 7132 17070 7188 17072
rect 7212 17070 7268 17072
rect 7292 17070 7348 17072
rect 7372 17070 7428 17072
rect 7132 17018 7158 17070
rect 7158 17018 7188 17070
rect 7212 17018 7222 17070
rect 7222 17018 7268 17070
rect 7292 17018 7338 17070
rect 7338 17018 7348 17070
rect 7372 17018 7402 17070
rect 7402 17018 7428 17070
rect 7132 17016 7188 17018
rect 7212 17016 7268 17018
rect 7292 17016 7348 17018
rect 7372 17016 7428 17018
rect 12460 17070 12516 17072
rect 12540 17070 12596 17072
rect 12620 17070 12676 17072
rect 12700 17070 12756 17072
rect 12460 17018 12486 17070
rect 12486 17018 12516 17070
rect 12540 17018 12550 17070
rect 12550 17018 12596 17070
rect 12620 17018 12666 17070
rect 12666 17018 12676 17070
rect 12700 17018 12730 17070
rect 12730 17018 12756 17070
rect 12460 17016 12516 17018
rect 12540 17016 12596 17018
rect 12620 17016 12676 17018
rect 12700 17016 12756 17018
rect 17788 17070 17844 17072
rect 17868 17070 17924 17072
rect 17948 17070 18004 17072
rect 18028 17070 18084 17072
rect 17788 17018 17814 17070
rect 17814 17018 17844 17070
rect 17868 17018 17878 17070
rect 17878 17018 17924 17070
rect 17948 17018 17994 17070
rect 17994 17018 18004 17070
rect 18028 17018 18058 17070
rect 18058 17018 18084 17070
rect 17788 17016 17844 17018
rect 17868 17016 17924 17018
rect 17948 17016 18004 17018
rect 18028 17016 18084 17018
rect 2068 16054 2124 16110
rect 4468 16404 4524 16406
rect 4548 16404 4604 16406
rect 4628 16404 4684 16406
rect 4708 16404 4764 16406
rect 4468 16352 4494 16404
rect 4494 16352 4524 16404
rect 4548 16352 4558 16404
rect 4558 16352 4604 16404
rect 4628 16352 4674 16404
rect 4674 16352 4684 16404
rect 4708 16352 4738 16404
rect 4738 16352 4764 16404
rect 4468 16350 4524 16352
rect 4548 16350 4604 16352
rect 4628 16350 4684 16352
rect 4708 16350 4764 16352
rect 9796 16404 9852 16406
rect 9876 16404 9932 16406
rect 9956 16404 10012 16406
rect 10036 16404 10092 16406
rect 9796 16352 9822 16404
rect 9822 16352 9852 16404
rect 9876 16352 9886 16404
rect 9886 16352 9932 16404
rect 9956 16352 10002 16404
rect 10002 16352 10012 16404
rect 10036 16352 10066 16404
rect 10066 16352 10092 16404
rect 9796 16350 9852 16352
rect 9876 16350 9932 16352
rect 9956 16350 10012 16352
rect 10036 16350 10092 16352
rect 15124 16404 15180 16406
rect 15204 16404 15260 16406
rect 15284 16404 15340 16406
rect 15364 16404 15420 16406
rect 15124 16352 15150 16404
rect 15150 16352 15180 16404
rect 15204 16352 15214 16404
rect 15214 16352 15260 16404
rect 15284 16352 15330 16404
rect 15330 16352 15340 16404
rect 15364 16352 15394 16404
rect 15394 16352 15420 16404
rect 15124 16350 15180 16352
rect 15204 16350 15260 16352
rect 15284 16350 15340 16352
rect 15364 16350 15420 16352
rect 20452 16404 20508 16406
rect 20532 16404 20588 16406
rect 20612 16404 20668 16406
rect 20692 16404 20748 16406
rect 20452 16352 20478 16404
rect 20478 16352 20508 16404
rect 20532 16352 20542 16404
rect 20542 16352 20588 16404
rect 20612 16352 20658 16404
rect 20658 16352 20668 16404
rect 20692 16352 20722 16404
rect 20722 16352 20748 16404
rect 20452 16350 20508 16352
rect 20532 16350 20588 16352
rect 20612 16350 20668 16352
rect 20692 16350 20748 16352
rect 7132 15738 7188 15740
rect 7212 15738 7268 15740
rect 7292 15738 7348 15740
rect 7372 15738 7428 15740
rect 7132 15686 7158 15738
rect 7158 15686 7188 15738
rect 7212 15686 7222 15738
rect 7222 15686 7268 15738
rect 7292 15686 7338 15738
rect 7338 15686 7348 15738
rect 7372 15686 7402 15738
rect 7402 15686 7428 15738
rect 7132 15684 7188 15686
rect 7212 15684 7268 15686
rect 7292 15684 7348 15686
rect 7372 15684 7428 15686
rect 12460 15738 12516 15740
rect 12540 15738 12596 15740
rect 12620 15738 12676 15740
rect 12700 15738 12756 15740
rect 12460 15686 12486 15738
rect 12486 15686 12516 15738
rect 12540 15686 12550 15738
rect 12550 15686 12596 15738
rect 12620 15686 12666 15738
rect 12666 15686 12676 15738
rect 12700 15686 12730 15738
rect 12730 15686 12756 15738
rect 12460 15684 12516 15686
rect 12540 15684 12596 15686
rect 12620 15684 12676 15686
rect 12700 15684 12756 15686
rect 17788 15738 17844 15740
rect 17868 15738 17924 15740
rect 17948 15738 18004 15740
rect 18028 15738 18084 15740
rect 17788 15686 17814 15738
rect 17814 15686 17844 15738
rect 17868 15686 17878 15738
rect 17878 15686 17924 15738
rect 17948 15686 17994 15738
rect 17994 15686 18004 15738
rect 18028 15686 18058 15738
rect 18058 15686 18084 15738
rect 17788 15684 17844 15686
rect 17868 15684 17924 15686
rect 17948 15684 18004 15686
rect 18028 15684 18084 15686
rect 4468 15072 4524 15074
rect 4548 15072 4604 15074
rect 4628 15072 4684 15074
rect 4708 15072 4764 15074
rect 4468 15020 4494 15072
rect 4494 15020 4524 15072
rect 4548 15020 4558 15072
rect 4558 15020 4604 15072
rect 4628 15020 4674 15072
rect 4674 15020 4684 15072
rect 4708 15020 4738 15072
rect 4738 15020 4764 15072
rect 4468 15018 4524 15020
rect 4548 15018 4604 15020
rect 4628 15018 4684 15020
rect 4708 15018 4764 15020
rect 9796 15072 9852 15074
rect 9876 15072 9932 15074
rect 9956 15072 10012 15074
rect 10036 15072 10092 15074
rect 9796 15020 9822 15072
rect 9822 15020 9852 15072
rect 9876 15020 9886 15072
rect 9886 15020 9932 15072
rect 9956 15020 10002 15072
rect 10002 15020 10012 15072
rect 10036 15020 10066 15072
rect 10066 15020 10092 15072
rect 9796 15018 9852 15020
rect 9876 15018 9932 15020
rect 9956 15018 10012 15020
rect 10036 15018 10092 15020
rect 15124 15072 15180 15074
rect 15204 15072 15260 15074
rect 15284 15072 15340 15074
rect 15364 15072 15420 15074
rect 15124 15020 15150 15072
rect 15150 15020 15180 15072
rect 15204 15020 15214 15072
rect 15214 15020 15260 15072
rect 15284 15020 15330 15072
rect 15330 15020 15340 15072
rect 15364 15020 15394 15072
rect 15394 15020 15420 15072
rect 15124 15018 15180 15020
rect 15204 15018 15260 15020
rect 15284 15018 15340 15020
rect 15364 15018 15420 15020
rect 20452 15072 20508 15074
rect 20532 15072 20588 15074
rect 20612 15072 20668 15074
rect 20692 15072 20748 15074
rect 20452 15020 20478 15072
rect 20478 15020 20508 15072
rect 20532 15020 20542 15072
rect 20542 15020 20588 15072
rect 20612 15020 20658 15072
rect 20658 15020 20668 15072
rect 20692 15020 20722 15072
rect 20722 15020 20748 15072
rect 20452 15018 20508 15020
rect 20532 15018 20588 15020
rect 20612 15018 20668 15020
rect 20692 15018 20748 15020
rect 7132 14406 7188 14408
rect 7212 14406 7268 14408
rect 7292 14406 7348 14408
rect 7372 14406 7428 14408
rect 7132 14354 7158 14406
rect 7158 14354 7188 14406
rect 7212 14354 7222 14406
rect 7222 14354 7268 14406
rect 7292 14354 7338 14406
rect 7338 14354 7348 14406
rect 7372 14354 7402 14406
rect 7402 14354 7428 14406
rect 7132 14352 7188 14354
rect 7212 14352 7268 14354
rect 7292 14352 7348 14354
rect 7372 14352 7428 14354
rect 12460 14406 12516 14408
rect 12540 14406 12596 14408
rect 12620 14406 12676 14408
rect 12700 14406 12756 14408
rect 12460 14354 12486 14406
rect 12486 14354 12516 14406
rect 12540 14354 12550 14406
rect 12550 14354 12596 14406
rect 12620 14354 12666 14406
rect 12666 14354 12676 14406
rect 12700 14354 12730 14406
rect 12730 14354 12756 14406
rect 12460 14352 12516 14354
rect 12540 14352 12596 14354
rect 12620 14352 12676 14354
rect 12700 14352 12756 14354
rect 17788 14406 17844 14408
rect 17868 14406 17924 14408
rect 17948 14406 18004 14408
rect 18028 14406 18084 14408
rect 17788 14354 17814 14406
rect 17814 14354 17844 14406
rect 17868 14354 17878 14406
rect 17878 14354 17924 14406
rect 17948 14354 17994 14406
rect 17994 14354 18004 14406
rect 18028 14354 18058 14406
rect 18058 14354 18084 14406
rect 17788 14352 17844 14354
rect 17868 14352 17924 14354
rect 17948 14352 18004 14354
rect 18028 14352 18084 14354
rect 4468 13740 4524 13742
rect 4548 13740 4604 13742
rect 4628 13740 4684 13742
rect 4708 13740 4764 13742
rect 4468 13688 4494 13740
rect 4494 13688 4524 13740
rect 4548 13688 4558 13740
rect 4558 13688 4604 13740
rect 4628 13688 4674 13740
rect 4674 13688 4684 13740
rect 4708 13688 4738 13740
rect 4738 13688 4764 13740
rect 4468 13686 4524 13688
rect 4548 13686 4604 13688
rect 4628 13686 4684 13688
rect 4708 13686 4764 13688
rect 9796 13740 9852 13742
rect 9876 13740 9932 13742
rect 9956 13740 10012 13742
rect 10036 13740 10092 13742
rect 9796 13688 9822 13740
rect 9822 13688 9852 13740
rect 9876 13688 9886 13740
rect 9886 13688 9932 13740
rect 9956 13688 10002 13740
rect 10002 13688 10012 13740
rect 10036 13688 10066 13740
rect 10066 13688 10092 13740
rect 9796 13686 9852 13688
rect 9876 13686 9932 13688
rect 9956 13686 10012 13688
rect 10036 13686 10092 13688
rect 15124 13740 15180 13742
rect 15204 13740 15260 13742
rect 15284 13740 15340 13742
rect 15364 13740 15420 13742
rect 15124 13688 15150 13740
rect 15150 13688 15180 13740
rect 15204 13688 15214 13740
rect 15214 13688 15260 13740
rect 15284 13688 15330 13740
rect 15330 13688 15340 13740
rect 15364 13688 15394 13740
rect 15394 13688 15420 13740
rect 15124 13686 15180 13688
rect 15204 13686 15260 13688
rect 15284 13686 15340 13688
rect 15364 13686 15420 13688
rect 20452 13740 20508 13742
rect 20532 13740 20588 13742
rect 20612 13740 20668 13742
rect 20692 13740 20748 13742
rect 20452 13688 20478 13740
rect 20478 13688 20508 13740
rect 20532 13688 20542 13740
rect 20542 13688 20588 13740
rect 20612 13688 20658 13740
rect 20658 13688 20668 13740
rect 20692 13688 20722 13740
rect 20722 13688 20748 13740
rect 20452 13686 20508 13688
rect 20532 13686 20588 13688
rect 20612 13686 20668 13688
rect 20692 13686 20748 13688
rect 7132 13074 7188 13076
rect 7212 13074 7268 13076
rect 7292 13074 7348 13076
rect 7372 13074 7428 13076
rect 7132 13022 7158 13074
rect 7158 13022 7188 13074
rect 7212 13022 7222 13074
rect 7222 13022 7268 13074
rect 7292 13022 7338 13074
rect 7338 13022 7348 13074
rect 7372 13022 7402 13074
rect 7402 13022 7428 13074
rect 7132 13020 7188 13022
rect 7212 13020 7268 13022
rect 7292 13020 7348 13022
rect 7372 13020 7428 13022
rect 12460 13074 12516 13076
rect 12540 13074 12596 13076
rect 12620 13074 12676 13076
rect 12700 13074 12756 13076
rect 12460 13022 12486 13074
rect 12486 13022 12516 13074
rect 12540 13022 12550 13074
rect 12550 13022 12596 13074
rect 12620 13022 12666 13074
rect 12666 13022 12676 13074
rect 12700 13022 12730 13074
rect 12730 13022 12756 13074
rect 12460 13020 12516 13022
rect 12540 13020 12596 13022
rect 12620 13020 12676 13022
rect 12700 13020 12756 13022
rect 17788 13074 17844 13076
rect 17868 13074 17924 13076
rect 17948 13074 18004 13076
rect 18028 13074 18084 13076
rect 17788 13022 17814 13074
rect 17814 13022 17844 13074
rect 17868 13022 17878 13074
rect 17878 13022 17924 13074
rect 17948 13022 17994 13074
rect 17994 13022 18004 13074
rect 18028 13022 18058 13074
rect 18058 13022 18084 13074
rect 17788 13020 17844 13022
rect 17868 13020 17924 13022
rect 17948 13020 18004 13022
rect 18028 13020 18084 13022
rect 4468 12408 4524 12410
rect 4548 12408 4604 12410
rect 4628 12408 4684 12410
rect 4708 12408 4764 12410
rect 4468 12356 4494 12408
rect 4494 12356 4524 12408
rect 4548 12356 4558 12408
rect 4558 12356 4604 12408
rect 4628 12356 4674 12408
rect 4674 12356 4684 12408
rect 4708 12356 4738 12408
rect 4738 12356 4764 12408
rect 4468 12354 4524 12356
rect 4548 12354 4604 12356
rect 4628 12354 4684 12356
rect 4708 12354 4764 12356
rect 9796 12408 9852 12410
rect 9876 12408 9932 12410
rect 9956 12408 10012 12410
rect 10036 12408 10092 12410
rect 9796 12356 9822 12408
rect 9822 12356 9852 12408
rect 9876 12356 9886 12408
rect 9886 12356 9932 12408
rect 9956 12356 10002 12408
rect 10002 12356 10012 12408
rect 10036 12356 10066 12408
rect 10066 12356 10092 12408
rect 9796 12354 9852 12356
rect 9876 12354 9932 12356
rect 9956 12354 10012 12356
rect 10036 12354 10092 12356
rect 15124 12408 15180 12410
rect 15204 12408 15260 12410
rect 15284 12408 15340 12410
rect 15364 12408 15420 12410
rect 15124 12356 15150 12408
rect 15150 12356 15180 12408
rect 15204 12356 15214 12408
rect 15214 12356 15260 12408
rect 15284 12356 15330 12408
rect 15330 12356 15340 12408
rect 15364 12356 15394 12408
rect 15394 12356 15420 12408
rect 15124 12354 15180 12356
rect 15204 12354 15260 12356
rect 15284 12354 15340 12356
rect 15364 12354 15420 12356
rect 20452 12408 20508 12410
rect 20532 12408 20588 12410
rect 20612 12408 20668 12410
rect 20692 12408 20748 12410
rect 20452 12356 20478 12408
rect 20478 12356 20508 12408
rect 20532 12356 20542 12408
rect 20542 12356 20588 12408
rect 20612 12356 20658 12408
rect 20658 12356 20668 12408
rect 20692 12356 20722 12408
rect 20722 12356 20748 12408
rect 20452 12354 20508 12356
rect 20532 12354 20588 12356
rect 20612 12354 20668 12356
rect 20692 12354 20748 12356
rect 7132 11742 7188 11744
rect 7212 11742 7268 11744
rect 7292 11742 7348 11744
rect 7372 11742 7428 11744
rect 7132 11690 7158 11742
rect 7158 11690 7188 11742
rect 7212 11690 7222 11742
rect 7222 11690 7268 11742
rect 7292 11690 7338 11742
rect 7338 11690 7348 11742
rect 7372 11690 7402 11742
rect 7402 11690 7428 11742
rect 7132 11688 7188 11690
rect 7212 11688 7268 11690
rect 7292 11688 7348 11690
rect 7372 11688 7428 11690
rect 12460 11742 12516 11744
rect 12540 11742 12596 11744
rect 12620 11742 12676 11744
rect 12700 11742 12756 11744
rect 12460 11690 12486 11742
rect 12486 11690 12516 11742
rect 12540 11690 12550 11742
rect 12550 11690 12596 11742
rect 12620 11690 12666 11742
rect 12666 11690 12676 11742
rect 12700 11690 12730 11742
rect 12730 11690 12756 11742
rect 12460 11688 12516 11690
rect 12540 11688 12596 11690
rect 12620 11688 12676 11690
rect 12700 11688 12756 11690
rect 17788 11742 17844 11744
rect 17868 11742 17924 11744
rect 17948 11742 18004 11744
rect 18028 11742 18084 11744
rect 17788 11690 17814 11742
rect 17814 11690 17844 11742
rect 17868 11690 17878 11742
rect 17878 11690 17924 11742
rect 17948 11690 17994 11742
rect 17994 11690 18004 11742
rect 18028 11690 18058 11742
rect 18058 11690 18084 11742
rect 17788 11688 17844 11690
rect 17868 11688 17924 11690
rect 17948 11688 18004 11690
rect 18028 11688 18084 11690
rect 2068 10726 2124 10782
rect 4468 11076 4524 11078
rect 4548 11076 4604 11078
rect 4628 11076 4684 11078
rect 4708 11076 4764 11078
rect 4468 11024 4494 11076
rect 4494 11024 4524 11076
rect 4548 11024 4558 11076
rect 4558 11024 4604 11076
rect 4628 11024 4674 11076
rect 4674 11024 4684 11076
rect 4708 11024 4738 11076
rect 4738 11024 4764 11076
rect 4468 11022 4524 11024
rect 4548 11022 4604 11024
rect 4628 11022 4684 11024
rect 4708 11022 4764 11024
rect 9796 11076 9852 11078
rect 9876 11076 9932 11078
rect 9956 11076 10012 11078
rect 10036 11076 10092 11078
rect 9796 11024 9822 11076
rect 9822 11024 9852 11076
rect 9876 11024 9886 11076
rect 9886 11024 9932 11076
rect 9956 11024 10002 11076
rect 10002 11024 10012 11076
rect 10036 11024 10066 11076
rect 10066 11024 10092 11076
rect 9796 11022 9852 11024
rect 9876 11022 9932 11024
rect 9956 11022 10012 11024
rect 10036 11022 10092 11024
rect 15124 11076 15180 11078
rect 15204 11076 15260 11078
rect 15284 11076 15340 11078
rect 15364 11076 15420 11078
rect 15124 11024 15150 11076
rect 15150 11024 15180 11076
rect 15204 11024 15214 11076
rect 15214 11024 15260 11076
rect 15284 11024 15330 11076
rect 15330 11024 15340 11076
rect 15364 11024 15394 11076
rect 15394 11024 15420 11076
rect 15124 11022 15180 11024
rect 15204 11022 15260 11024
rect 15284 11022 15340 11024
rect 15364 11022 15420 11024
rect 20452 11076 20508 11078
rect 20532 11076 20588 11078
rect 20612 11076 20668 11078
rect 20692 11076 20748 11078
rect 20452 11024 20478 11076
rect 20478 11024 20508 11076
rect 20532 11024 20542 11076
rect 20542 11024 20588 11076
rect 20612 11024 20658 11076
rect 20658 11024 20668 11076
rect 20692 11024 20722 11076
rect 20722 11024 20748 11076
rect 20452 11022 20508 11024
rect 20532 11022 20588 11024
rect 20612 11022 20668 11024
rect 20692 11022 20748 11024
rect 7132 10410 7188 10412
rect 7212 10410 7268 10412
rect 7292 10410 7348 10412
rect 7372 10410 7428 10412
rect 7132 10358 7158 10410
rect 7158 10358 7188 10410
rect 7212 10358 7222 10410
rect 7222 10358 7268 10410
rect 7292 10358 7338 10410
rect 7338 10358 7348 10410
rect 7372 10358 7402 10410
rect 7402 10358 7428 10410
rect 7132 10356 7188 10358
rect 7212 10356 7268 10358
rect 7292 10356 7348 10358
rect 7372 10356 7428 10358
rect 12460 10410 12516 10412
rect 12540 10410 12596 10412
rect 12620 10410 12676 10412
rect 12700 10410 12756 10412
rect 12460 10358 12486 10410
rect 12486 10358 12516 10410
rect 12540 10358 12550 10410
rect 12550 10358 12596 10410
rect 12620 10358 12666 10410
rect 12666 10358 12676 10410
rect 12700 10358 12730 10410
rect 12730 10358 12756 10410
rect 12460 10356 12516 10358
rect 12540 10356 12596 10358
rect 12620 10356 12676 10358
rect 12700 10356 12756 10358
rect 17788 10410 17844 10412
rect 17868 10410 17924 10412
rect 17948 10410 18004 10412
rect 18028 10410 18084 10412
rect 17788 10358 17814 10410
rect 17814 10358 17844 10410
rect 17868 10358 17878 10410
rect 17878 10358 17924 10410
rect 17948 10358 17994 10410
rect 17994 10358 18004 10410
rect 18028 10358 18058 10410
rect 18058 10358 18084 10410
rect 17788 10356 17844 10358
rect 17868 10356 17924 10358
rect 17948 10356 18004 10358
rect 18028 10356 18084 10358
rect 4468 9744 4524 9746
rect 4548 9744 4604 9746
rect 4628 9744 4684 9746
rect 4708 9744 4764 9746
rect 4468 9692 4494 9744
rect 4494 9692 4524 9744
rect 4548 9692 4558 9744
rect 4558 9692 4604 9744
rect 4628 9692 4674 9744
rect 4674 9692 4684 9744
rect 4708 9692 4738 9744
rect 4738 9692 4764 9744
rect 4468 9690 4524 9692
rect 4548 9690 4604 9692
rect 4628 9690 4684 9692
rect 4708 9690 4764 9692
rect 9796 9744 9852 9746
rect 9876 9744 9932 9746
rect 9956 9744 10012 9746
rect 10036 9744 10092 9746
rect 9796 9692 9822 9744
rect 9822 9692 9852 9744
rect 9876 9692 9886 9744
rect 9886 9692 9932 9744
rect 9956 9692 10002 9744
rect 10002 9692 10012 9744
rect 10036 9692 10066 9744
rect 10066 9692 10092 9744
rect 9796 9690 9852 9692
rect 9876 9690 9932 9692
rect 9956 9690 10012 9692
rect 10036 9690 10092 9692
rect 15124 9744 15180 9746
rect 15204 9744 15260 9746
rect 15284 9744 15340 9746
rect 15364 9744 15420 9746
rect 15124 9692 15150 9744
rect 15150 9692 15180 9744
rect 15204 9692 15214 9744
rect 15214 9692 15260 9744
rect 15284 9692 15330 9744
rect 15330 9692 15340 9744
rect 15364 9692 15394 9744
rect 15394 9692 15420 9744
rect 15124 9690 15180 9692
rect 15204 9690 15260 9692
rect 15284 9690 15340 9692
rect 15364 9690 15420 9692
rect 20452 9744 20508 9746
rect 20532 9744 20588 9746
rect 20612 9744 20668 9746
rect 20692 9744 20748 9746
rect 20452 9692 20478 9744
rect 20478 9692 20508 9744
rect 20532 9692 20542 9744
rect 20542 9692 20588 9744
rect 20612 9692 20658 9744
rect 20658 9692 20668 9744
rect 20692 9692 20722 9744
rect 20722 9692 20748 9744
rect 20452 9690 20508 9692
rect 20532 9690 20588 9692
rect 20612 9690 20668 9692
rect 20692 9690 20748 9692
rect 7132 9078 7188 9080
rect 7212 9078 7268 9080
rect 7292 9078 7348 9080
rect 7372 9078 7428 9080
rect 7132 9026 7158 9078
rect 7158 9026 7188 9078
rect 7212 9026 7222 9078
rect 7222 9026 7268 9078
rect 7292 9026 7338 9078
rect 7338 9026 7348 9078
rect 7372 9026 7402 9078
rect 7402 9026 7428 9078
rect 7132 9024 7188 9026
rect 7212 9024 7268 9026
rect 7292 9024 7348 9026
rect 7372 9024 7428 9026
rect 12460 9078 12516 9080
rect 12540 9078 12596 9080
rect 12620 9078 12676 9080
rect 12700 9078 12756 9080
rect 12460 9026 12486 9078
rect 12486 9026 12516 9078
rect 12540 9026 12550 9078
rect 12550 9026 12596 9078
rect 12620 9026 12666 9078
rect 12666 9026 12676 9078
rect 12700 9026 12730 9078
rect 12730 9026 12756 9078
rect 12460 9024 12516 9026
rect 12540 9024 12596 9026
rect 12620 9024 12676 9026
rect 12700 9024 12756 9026
rect 17788 9078 17844 9080
rect 17868 9078 17924 9080
rect 17948 9078 18004 9080
rect 18028 9078 18084 9080
rect 17788 9026 17814 9078
rect 17814 9026 17844 9078
rect 17868 9026 17878 9078
rect 17878 9026 17924 9078
rect 17948 9026 17994 9078
rect 17994 9026 18004 9078
rect 18028 9026 18058 9078
rect 18058 9026 18084 9078
rect 17788 9024 17844 9026
rect 17868 9024 17924 9026
rect 17948 9024 18004 9026
rect 18028 9024 18084 9026
rect 4468 8412 4524 8414
rect 4548 8412 4604 8414
rect 4628 8412 4684 8414
rect 4708 8412 4764 8414
rect 4468 8360 4494 8412
rect 4494 8360 4524 8412
rect 4548 8360 4558 8412
rect 4558 8360 4604 8412
rect 4628 8360 4674 8412
rect 4674 8360 4684 8412
rect 4708 8360 4738 8412
rect 4738 8360 4764 8412
rect 4468 8358 4524 8360
rect 4548 8358 4604 8360
rect 4628 8358 4684 8360
rect 4708 8358 4764 8360
rect 9796 8412 9852 8414
rect 9876 8412 9932 8414
rect 9956 8412 10012 8414
rect 10036 8412 10092 8414
rect 9796 8360 9822 8412
rect 9822 8360 9852 8412
rect 9876 8360 9886 8412
rect 9886 8360 9932 8412
rect 9956 8360 10002 8412
rect 10002 8360 10012 8412
rect 10036 8360 10066 8412
rect 10066 8360 10092 8412
rect 9796 8358 9852 8360
rect 9876 8358 9932 8360
rect 9956 8358 10012 8360
rect 10036 8358 10092 8360
rect 15124 8412 15180 8414
rect 15204 8412 15260 8414
rect 15284 8412 15340 8414
rect 15364 8412 15420 8414
rect 15124 8360 15150 8412
rect 15150 8360 15180 8412
rect 15204 8360 15214 8412
rect 15214 8360 15260 8412
rect 15284 8360 15330 8412
rect 15330 8360 15340 8412
rect 15364 8360 15394 8412
rect 15394 8360 15420 8412
rect 15124 8358 15180 8360
rect 15204 8358 15260 8360
rect 15284 8358 15340 8360
rect 15364 8358 15420 8360
rect 20452 8412 20508 8414
rect 20532 8412 20588 8414
rect 20612 8412 20668 8414
rect 20692 8412 20748 8414
rect 20452 8360 20478 8412
rect 20478 8360 20508 8412
rect 20532 8360 20542 8412
rect 20542 8360 20588 8412
rect 20612 8360 20658 8412
rect 20658 8360 20668 8412
rect 20692 8360 20722 8412
rect 20722 8360 20748 8412
rect 20452 8358 20508 8360
rect 20532 8358 20588 8360
rect 20612 8358 20668 8360
rect 20692 8358 20748 8360
rect 7132 7746 7188 7748
rect 7212 7746 7268 7748
rect 7292 7746 7348 7748
rect 7372 7746 7428 7748
rect 7132 7694 7158 7746
rect 7158 7694 7188 7746
rect 7212 7694 7222 7746
rect 7222 7694 7268 7746
rect 7292 7694 7338 7746
rect 7338 7694 7348 7746
rect 7372 7694 7402 7746
rect 7402 7694 7428 7746
rect 7132 7692 7188 7694
rect 7212 7692 7268 7694
rect 7292 7692 7348 7694
rect 7372 7692 7428 7694
rect 12460 7746 12516 7748
rect 12540 7746 12596 7748
rect 12620 7746 12676 7748
rect 12700 7746 12756 7748
rect 12460 7694 12486 7746
rect 12486 7694 12516 7746
rect 12540 7694 12550 7746
rect 12550 7694 12596 7746
rect 12620 7694 12666 7746
rect 12666 7694 12676 7746
rect 12700 7694 12730 7746
rect 12730 7694 12756 7746
rect 12460 7692 12516 7694
rect 12540 7692 12596 7694
rect 12620 7692 12676 7694
rect 12700 7692 12756 7694
rect 17788 7746 17844 7748
rect 17868 7746 17924 7748
rect 17948 7746 18004 7748
rect 18028 7746 18084 7748
rect 17788 7694 17814 7746
rect 17814 7694 17844 7746
rect 17868 7694 17878 7746
rect 17878 7694 17924 7746
rect 17948 7694 17994 7746
rect 17994 7694 18004 7746
rect 18028 7694 18058 7746
rect 18058 7694 18084 7746
rect 17788 7692 17844 7694
rect 17868 7692 17924 7694
rect 17948 7692 18004 7694
rect 18028 7692 18084 7694
rect 4468 7080 4524 7082
rect 4548 7080 4604 7082
rect 4628 7080 4684 7082
rect 4708 7080 4764 7082
rect 4468 7028 4494 7080
rect 4494 7028 4524 7080
rect 4548 7028 4558 7080
rect 4558 7028 4604 7080
rect 4628 7028 4674 7080
rect 4674 7028 4684 7080
rect 4708 7028 4738 7080
rect 4738 7028 4764 7080
rect 4468 7026 4524 7028
rect 4548 7026 4604 7028
rect 4628 7026 4684 7028
rect 4708 7026 4764 7028
rect 9796 7080 9852 7082
rect 9876 7080 9932 7082
rect 9956 7080 10012 7082
rect 10036 7080 10092 7082
rect 9796 7028 9822 7080
rect 9822 7028 9852 7080
rect 9876 7028 9886 7080
rect 9886 7028 9932 7080
rect 9956 7028 10002 7080
rect 10002 7028 10012 7080
rect 10036 7028 10066 7080
rect 10066 7028 10092 7080
rect 9796 7026 9852 7028
rect 9876 7026 9932 7028
rect 9956 7026 10012 7028
rect 10036 7026 10092 7028
rect 15124 7080 15180 7082
rect 15204 7080 15260 7082
rect 15284 7080 15340 7082
rect 15364 7080 15420 7082
rect 15124 7028 15150 7080
rect 15150 7028 15180 7080
rect 15204 7028 15214 7080
rect 15214 7028 15260 7080
rect 15284 7028 15330 7080
rect 15330 7028 15340 7080
rect 15364 7028 15394 7080
rect 15394 7028 15420 7080
rect 15124 7026 15180 7028
rect 15204 7026 15260 7028
rect 15284 7026 15340 7028
rect 15364 7026 15420 7028
rect 20452 7080 20508 7082
rect 20532 7080 20588 7082
rect 20612 7080 20668 7082
rect 20692 7080 20748 7082
rect 20452 7028 20478 7080
rect 20478 7028 20508 7080
rect 20532 7028 20542 7080
rect 20542 7028 20588 7080
rect 20612 7028 20658 7080
rect 20658 7028 20668 7080
rect 20692 7028 20722 7080
rect 20722 7028 20748 7080
rect 20452 7026 20508 7028
rect 20532 7026 20588 7028
rect 20612 7026 20668 7028
rect 20692 7026 20748 7028
rect 7132 6414 7188 6416
rect 7212 6414 7268 6416
rect 7292 6414 7348 6416
rect 7372 6414 7428 6416
rect 7132 6362 7158 6414
rect 7158 6362 7188 6414
rect 7212 6362 7222 6414
rect 7222 6362 7268 6414
rect 7292 6362 7338 6414
rect 7338 6362 7348 6414
rect 7372 6362 7402 6414
rect 7402 6362 7428 6414
rect 7132 6360 7188 6362
rect 7212 6360 7268 6362
rect 7292 6360 7348 6362
rect 7372 6360 7428 6362
rect 12460 6414 12516 6416
rect 12540 6414 12596 6416
rect 12620 6414 12676 6416
rect 12700 6414 12756 6416
rect 12460 6362 12486 6414
rect 12486 6362 12516 6414
rect 12540 6362 12550 6414
rect 12550 6362 12596 6414
rect 12620 6362 12666 6414
rect 12666 6362 12676 6414
rect 12700 6362 12730 6414
rect 12730 6362 12756 6414
rect 12460 6360 12516 6362
rect 12540 6360 12596 6362
rect 12620 6360 12676 6362
rect 12700 6360 12756 6362
rect 17788 6414 17844 6416
rect 17868 6414 17924 6416
rect 17948 6414 18004 6416
rect 18028 6414 18084 6416
rect 17788 6362 17814 6414
rect 17814 6362 17844 6414
rect 17868 6362 17878 6414
rect 17878 6362 17924 6414
rect 17948 6362 17994 6414
rect 17994 6362 18004 6414
rect 18028 6362 18058 6414
rect 18058 6362 18084 6414
rect 17788 6360 17844 6362
rect 17868 6360 17924 6362
rect 17948 6360 18004 6362
rect 18028 6360 18084 6362
rect 4468 5748 4524 5750
rect 4548 5748 4604 5750
rect 4628 5748 4684 5750
rect 4708 5748 4764 5750
rect 4468 5696 4494 5748
rect 4494 5696 4524 5748
rect 4548 5696 4558 5748
rect 4558 5696 4604 5748
rect 4628 5696 4674 5748
rect 4674 5696 4684 5748
rect 4708 5696 4738 5748
rect 4738 5696 4764 5748
rect 4468 5694 4524 5696
rect 4548 5694 4604 5696
rect 4628 5694 4684 5696
rect 4708 5694 4764 5696
rect 9796 5748 9852 5750
rect 9876 5748 9932 5750
rect 9956 5748 10012 5750
rect 10036 5748 10092 5750
rect 9796 5696 9822 5748
rect 9822 5696 9852 5748
rect 9876 5696 9886 5748
rect 9886 5696 9932 5748
rect 9956 5696 10002 5748
rect 10002 5696 10012 5748
rect 10036 5696 10066 5748
rect 10066 5696 10092 5748
rect 9796 5694 9852 5696
rect 9876 5694 9932 5696
rect 9956 5694 10012 5696
rect 10036 5694 10092 5696
rect 15124 5748 15180 5750
rect 15204 5748 15260 5750
rect 15284 5748 15340 5750
rect 15364 5748 15420 5750
rect 15124 5696 15150 5748
rect 15150 5696 15180 5748
rect 15204 5696 15214 5748
rect 15214 5696 15260 5748
rect 15284 5696 15330 5748
rect 15330 5696 15340 5748
rect 15364 5696 15394 5748
rect 15394 5696 15420 5748
rect 15124 5694 15180 5696
rect 15204 5694 15260 5696
rect 15284 5694 15340 5696
rect 15364 5694 15420 5696
rect 20452 5748 20508 5750
rect 20532 5748 20588 5750
rect 20612 5748 20668 5750
rect 20692 5748 20748 5750
rect 20452 5696 20478 5748
rect 20478 5696 20508 5748
rect 20532 5696 20542 5748
rect 20542 5696 20588 5748
rect 20612 5696 20658 5748
rect 20658 5696 20668 5748
rect 20692 5696 20722 5748
rect 20722 5696 20748 5748
rect 20452 5694 20508 5696
rect 20532 5694 20588 5696
rect 20612 5694 20668 5696
rect 20692 5694 20748 5696
rect 7132 5082 7188 5084
rect 7212 5082 7268 5084
rect 7292 5082 7348 5084
rect 7372 5082 7428 5084
rect 7132 5030 7158 5082
rect 7158 5030 7188 5082
rect 7212 5030 7222 5082
rect 7222 5030 7268 5082
rect 7292 5030 7338 5082
rect 7338 5030 7348 5082
rect 7372 5030 7402 5082
rect 7402 5030 7428 5082
rect 7132 5028 7188 5030
rect 7212 5028 7268 5030
rect 7292 5028 7348 5030
rect 7372 5028 7428 5030
rect 12460 5082 12516 5084
rect 12540 5082 12596 5084
rect 12620 5082 12676 5084
rect 12700 5082 12756 5084
rect 12460 5030 12486 5082
rect 12486 5030 12516 5082
rect 12540 5030 12550 5082
rect 12550 5030 12596 5082
rect 12620 5030 12666 5082
rect 12666 5030 12676 5082
rect 12700 5030 12730 5082
rect 12730 5030 12756 5082
rect 12460 5028 12516 5030
rect 12540 5028 12596 5030
rect 12620 5028 12676 5030
rect 12700 5028 12756 5030
rect 17788 5082 17844 5084
rect 17868 5082 17924 5084
rect 17948 5082 18004 5084
rect 18028 5082 18084 5084
rect 17788 5030 17814 5082
rect 17814 5030 17844 5082
rect 17868 5030 17878 5082
rect 17878 5030 17924 5082
rect 17948 5030 17994 5082
rect 17994 5030 18004 5082
rect 18028 5030 18058 5082
rect 18058 5030 18084 5082
rect 17788 5028 17844 5030
rect 17868 5028 17924 5030
rect 17948 5028 18004 5030
rect 18028 5028 18084 5030
rect 4468 4416 4524 4418
rect 4548 4416 4604 4418
rect 4628 4416 4684 4418
rect 4708 4416 4764 4418
rect 4468 4364 4494 4416
rect 4494 4364 4524 4416
rect 4548 4364 4558 4416
rect 4558 4364 4604 4416
rect 4628 4364 4674 4416
rect 4674 4364 4684 4416
rect 4708 4364 4738 4416
rect 4738 4364 4764 4416
rect 4468 4362 4524 4364
rect 4548 4362 4604 4364
rect 4628 4362 4684 4364
rect 4708 4362 4764 4364
rect 9796 4416 9852 4418
rect 9876 4416 9932 4418
rect 9956 4416 10012 4418
rect 10036 4416 10092 4418
rect 9796 4364 9822 4416
rect 9822 4364 9852 4416
rect 9876 4364 9886 4416
rect 9886 4364 9932 4416
rect 9956 4364 10002 4416
rect 10002 4364 10012 4416
rect 10036 4364 10066 4416
rect 10066 4364 10092 4416
rect 9796 4362 9852 4364
rect 9876 4362 9932 4364
rect 9956 4362 10012 4364
rect 10036 4362 10092 4364
rect 15124 4416 15180 4418
rect 15204 4416 15260 4418
rect 15284 4416 15340 4418
rect 15364 4416 15420 4418
rect 15124 4364 15150 4416
rect 15150 4364 15180 4416
rect 15204 4364 15214 4416
rect 15214 4364 15260 4416
rect 15284 4364 15330 4416
rect 15330 4364 15340 4416
rect 15364 4364 15394 4416
rect 15394 4364 15420 4416
rect 15124 4362 15180 4364
rect 15204 4362 15260 4364
rect 15284 4362 15340 4364
rect 15364 4362 15420 4364
rect 20452 4416 20508 4418
rect 20532 4416 20588 4418
rect 20612 4416 20668 4418
rect 20692 4416 20748 4418
rect 20452 4364 20478 4416
rect 20478 4364 20508 4416
rect 20532 4364 20542 4416
rect 20542 4364 20588 4416
rect 20612 4364 20658 4416
rect 20658 4364 20668 4416
rect 20692 4364 20722 4416
rect 20722 4364 20748 4416
rect 20452 4362 20508 4364
rect 20532 4362 20588 4364
rect 20612 4362 20668 4364
rect 20692 4362 20748 4364
rect 7132 3750 7188 3752
rect 7212 3750 7268 3752
rect 7292 3750 7348 3752
rect 7372 3750 7428 3752
rect 7132 3698 7158 3750
rect 7158 3698 7188 3750
rect 7212 3698 7222 3750
rect 7222 3698 7268 3750
rect 7292 3698 7338 3750
rect 7338 3698 7348 3750
rect 7372 3698 7402 3750
rect 7402 3698 7428 3750
rect 7132 3696 7188 3698
rect 7212 3696 7268 3698
rect 7292 3696 7348 3698
rect 7372 3696 7428 3698
rect 12460 3750 12516 3752
rect 12540 3750 12596 3752
rect 12620 3750 12676 3752
rect 12700 3750 12756 3752
rect 12460 3698 12486 3750
rect 12486 3698 12516 3750
rect 12540 3698 12550 3750
rect 12550 3698 12596 3750
rect 12620 3698 12666 3750
rect 12666 3698 12676 3750
rect 12700 3698 12730 3750
rect 12730 3698 12756 3750
rect 12460 3696 12516 3698
rect 12540 3696 12596 3698
rect 12620 3696 12676 3698
rect 12700 3696 12756 3698
rect 17788 3750 17844 3752
rect 17868 3750 17924 3752
rect 17948 3750 18004 3752
rect 18028 3750 18084 3752
rect 17788 3698 17814 3750
rect 17814 3698 17844 3750
rect 17868 3698 17878 3750
rect 17878 3698 17924 3750
rect 17948 3698 17994 3750
rect 17994 3698 18004 3750
rect 18028 3698 18058 3750
rect 18058 3698 18084 3750
rect 17788 3696 17844 3698
rect 17868 3696 17924 3698
rect 17948 3696 18004 3698
rect 18028 3696 18084 3698
rect 4468 3084 4524 3086
rect 4548 3084 4604 3086
rect 4628 3084 4684 3086
rect 4708 3084 4764 3086
rect 4468 3032 4494 3084
rect 4494 3032 4524 3084
rect 4548 3032 4558 3084
rect 4558 3032 4604 3084
rect 4628 3032 4674 3084
rect 4674 3032 4684 3084
rect 4708 3032 4738 3084
rect 4738 3032 4764 3084
rect 4468 3030 4524 3032
rect 4548 3030 4604 3032
rect 4628 3030 4684 3032
rect 4708 3030 4764 3032
rect 9796 3084 9852 3086
rect 9876 3084 9932 3086
rect 9956 3084 10012 3086
rect 10036 3084 10092 3086
rect 9796 3032 9822 3084
rect 9822 3032 9852 3084
rect 9876 3032 9886 3084
rect 9886 3032 9932 3084
rect 9956 3032 10002 3084
rect 10002 3032 10012 3084
rect 10036 3032 10066 3084
rect 10066 3032 10092 3084
rect 9796 3030 9852 3032
rect 9876 3030 9932 3032
rect 9956 3030 10012 3032
rect 10036 3030 10092 3032
rect 15124 3084 15180 3086
rect 15204 3084 15260 3086
rect 15284 3084 15340 3086
rect 15364 3084 15420 3086
rect 15124 3032 15150 3084
rect 15150 3032 15180 3084
rect 15204 3032 15214 3084
rect 15214 3032 15260 3084
rect 15284 3032 15330 3084
rect 15330 3032 15340 3084
rect 15364 3032 15394 3084
rect 15394 3032 15420 3084
rect 15124 3030 15180 3032
rect 15204 3030 15260 3032
rect 15284 3030 15340 3032
rect 15364 3030 15420 3032
rect 20452 3084 20508 3086
rect 20532 3084 20588 3086
rect 20612 3084 20668 3086
rect 20692 3084 20748 3086
rect 20452 3032 20478 3084
rect 20478 3032 20508 3084
rect 20532 3032 20542 3084
rect 20542 3032 20588 3084
rect 20612 3032 20658 3084
rect 20658 3032 20668 3084
rect 20692 3032 20722 3084
rect 20722 3032 20748 3084
rect 20452 3030 20508 3032
rect 20532 3030 20588 3032
rect 20612 3030 20668 3032
rect 20692 3030 20748 3032
rect 7132 2418 7188 2420
rect 7212 2418 7268 2420
rect 7292 2418 7348 2420
rect 7372 2418 7428 2420
rect 7132 2366 7158 2418
rect 7158 2366 7188 2418
rect 7212 2366 7222 2418
rect 7222 2366 7268 2418
rect 7292 2366 7338 2418
rect 7338 2366 7348 2418
rect 7372 2366 7402 2418
rect 7402 2366 7428 2418
rect 7132 2364 7188 2366
rect 7212 2364 7268 2366
rect 7292 2364 7348 2366
rect 7372 2364 7428 2366
rect 12460 2418 12516 2420
rect 12540 2418 12596 2420
rect 12620 2418 12676 2420
rect 12700 2418 12756 2420
rect 12460 2366 12486 2418
rect 12486 2366 12516 2418
rect 12540 2366 12550 2418
rect 12550 2366 12596 2418
rect 12620 2366 12666 2418
rect 12666 2366 12676 2418
rect 12700 2366 12730 2418
rect 12730 2366 12756 2418
rect 12460 2364 12516 2366
rect 12540 2364 12596 2366
rect 12620 2364 12676 2366
rect 12700 2364 12756 2366
rect 17788 2418 17844 2420
rect 17868 2418 17924 2420
rect 17948 2418 18004 2420
rect 18028 2418 18084 2420
rect 17788 2366 17814 2418
rect 17814 2366 17844 2418
rect 17868 2366 17878 2418
rect 17878 2366 17924 2418
rect 17948 2366 17994 2418
rect 17994 2366 18004 2418
rect 18028 2366 18058 2418
rect 18058 2366 18084 2418
rect 17788 2364 17844 2366
rect 17868 2364 17924 2366
rect 17948 2364 18004 2366
rect 18028 2364 18084 2366
rect 4468 1752 4524 1754
rect 4548 1752 4604 1754
rect 4628 1752 4684 1754
rect 4708 1752 4764 1754
rect 4468 1700 4494 1752
rect 4494 1700 4524 1752
rect 4548 1700 4558 1752
rect 4558 1700 4604 1752
rect 4628 1700 4674 1752
rect 4674 1700 4684 1752
rect 4708 1700 4738 1752
rect 4738 1700 4764 1752
rect 4468 1698 4524 1700
rect 4548 1698 4604 1700
rect 4628 1698 4684 1700
rect 4708 1698 4764 1700
rect 9796 1752 9852 1754
rect 9876 1752 9932 1754
rect 9956 1752 10012 1754
rect 10036 1752 10092 1754
rect 9796 1700 9822 1752
rect 9822 1700 9852 1752
rect 9876 1700 9886 1752
rect 9886 1700 9932 1752
rect 9956 1700 10002 1752
rect 10002 1700 10012 1752
rect 10036 1700 10066 1752
rect 10066 1700 10092 1752
rect 9796 1698 9852 1700
rect 9876 1698 9932 1700
rect 9956 1698 10012 1700
rect 10036 1698 10092 1700
rect 15124 1752 15180 1754
rect 15204 1752 15260 1754
rect 15284 1752 15340 1754
rect 15364 1752 15420 1754
rect 15124 1700 15150 1752
rect 15150 1700 15180 1752
rect 15204 1700 15214 1752
rect 15214 1700 15260 1752
rect 15284 1700 15330 1752
rect 15330 1700 15340 1752
rect 15364 1700 15394 1752
rect 15394 1700 15420 1752
rect 15124 1698 15180 1700
rect 15204 1698 15260 1700
rect 15284 1698 15340 1700
rect 15364 1698 15420 1700
rect 20452 1752 20508 1754
rect 20532 1752 20588 1754
rect 20612 1752 20668 1754
rect 20692 1752 20748 1754
rect 20452 1700 20478 1752
rect 20478 1700 20508 1752
rect 20532 1700 20542 1752
rect 20542 1700 20588 1752
rect 20612 1700 20658 1752
rect 20658 1700 20668 1752
rect 20692 1700 20722 1752
rect 20722 1700 20748 1752
rect 20452 1698 20508 1700
rect 20532 1698 20588 1700
rect 20612 1698 20668 1700
rect 20692 1698 20748 1700
rect 7132 1086 7188 1088
rect 7212 1086 7268 1088
rect 7292 1086 7348 1088
rect 7372 1086 7428 1088
rect 7132 1034 7158 1086
rect 7158 1034 7188 1086
rect 7212 1034 7222 1086
rect 7222 1034 7268 1086
rect 7292 1034 7338 1086
rect 7338 1034 7348 1086
rect 7372 1034 7402 1086
rect 7402 1034 7428 1086
rect 7132 1032 7188 1034
rect 7212 1032 7268 1034
rect 7292 1032 7348 1034
rect 7372 1032 7428 1034
rect 12460 1086 12516 1088
rect 12540 1086 12596 1088
rect 12620 1086 12676 1088
rect 12700 1086 12756 1088
rect 12460 1034 12486 1086
rect 12486 1034 12516 1086
rect 12540 1034 12550 1086
rect 12550 1034 12596 1086
rect 12620 1034 12666 1086
rect 12666 1034 12676 1086
rect 12700 1034 12730 1086
rect 12730 1034 12756 1086
rect 12460 1032 12516 1034
rect 12540 1032 12596 1034
rect 12620 1032 12676 1034
rect 12700 1032 12756 1034
rect 17788 1086 17844 1088
rect 17868 1086 17924 1088
rect 17948 1086 18004 1088
rect 18028 1086 18084 1088
rect 17788 1034 17814 1086
rect 17814 1034 17844 1086
rect 17868 1034 17878 1086
rect 17878 1034 17924 1086
rect 17948 1034 17994 1086
rect 17994 1034 18004 1086
rect 18028 1034 18058 1086
rect 18058 1034 18084 1086
rect 17788 1032 17844 1034
rect 17868 1032 17924 1034
rect 17948 1032 18004 1034
rect 18028 1032 18084 1034
rect 3028 810 3084 866
<< metal3 >>
rect 2735 27360 2801 27363
rect 830 27358 2801 27360
rect 830 27302 2740 27358
rect 2796 27302 2801 27358
rect 830 27300 2801 27302
rect 830 27192 890 27300
rect 2735 27297 2801 27300
rect 800 26936 920 27192
rect 4456 27066 4776 27067
rect 4456 27002 4464 27066
rect 4528 27002 4544 27066
rect 4608 27002 4624 27066
rect 4688 27002 4704 27066
rect 4768 27002 4776 27066
rect 4456 27001 4776 27002
rect 9784 27066 10104 27067
rect 9784 27002 9792 27066
rect 9856 27002 9872 27066
rect 9936 27002 9952 27066
rect 10016 27002 10032 27066
rect 10096 27002 10104 27066
rect 9784 27001 10104 27002
rect 15112 27066 15432 27067
rect 15112 27002 15120 27066
rect 15184 27002 15200 27066
rect 15264 27002 15280 27066
rect 15344 27002 15360 27066
rect 15424 27002 15432 27066
rect 15112 27001 15432 27002
rect 20440 27066 20760 27067
rect 20440 27002 20448 27066
rect 20512 27002 20528 27066
rect 20592 27002 20608 27066
rect 20672 27002 20688 27066
rect 20752 27002 20760 27066
rect 20440 27001 20760 27002
rect 800 26256 920 26512
rect 7120 26400 7440 26401
rect 7120 26336 7128 26400
rect 7192 26336 7208 26400
rect 7272 26336 7288 26400
rect 7352 26336 7368 26400
rect 7432 26336 7440 26400
rect 7120 26335 7440 26336
rect 12448 26400 12768 26401
rect 12448 26336 12456 26400
rect 12520 26336 12536 26400
rect 12600 26336 12616 26400
rect 12680 26336 12696 26400
rect 12760 26336 12768 26400
rect 12448 26335 12768 26336
rect 17776 26400 18096 26401
rect 17776 26336 17784 26400
rect 17848 26336 17864 26400
rect 17928 26336 17944 26400
rect 18008 26336 18024 26400
rect 18088 26336 18096 26400
rect 17776 26335 18096 26336
rect 830 26176 890 26256
rect 2351 26176 2417 26179
rect 830 26174 2417 26176
rect 830 26118 2356 26174
rect 2412 26118 2417 26174
rect 830 26116 2417 26118
rect 2351 26113 2417 26116
rect 800 25584 920 25832
rect 4456 25734 4776 25735
rect 4456 25670 4464 25734
rect 4528 25670 4544 25734
rect 4608 25670 4624 25734
rect 4688 25670 4704 25734
rect 4768 25670 4776 25734
rect 4456 25669 4776 25670
rect 9784 25734 10104 25735
rect 9784 25670 9792 25734
rect 9856 25670 9872 25734
rect 9936 25670 9952 25734
rect 10016 25670 10032 25734
rect 10096 25670 10104 25734
rect 9784 25669 10104 25670
rect 15112 25734 15432 25735
rect 15112 25670 15120 25734
rect 15184 25670 15200 25734
rect 15264 25670 15280 25734
rect 15344 25670 15360 25734
rect 15424 25670 15432 25734
rect 15112 25669 15432 25670
rect 20440 25734 20760 25735
rect 20440 25670 20448 25734
rect 20512 25670 20528 25734
rect 20592 25670 20608 25734
rect 20672 25670 20688 25734
rect 20752 25670 20760 25734
rect 20440 25669 20760 25670
rect 2447 25584 2513 25587
rect 800 25582 2513 25584
rect 800 25576 2452 25582
rect 830 25526 2452 25576
rect 2508 25526 2513 25582
rect 830 25524 2513 25526
rect 2447 25521 2513 25524
rect 7120 25068 7440 25069
rect 7120 25004 7128 25068
rect 7192 25004 7208 25068
rect 7272 25004 7288 25068
rect 7352 25004 7368 25068
rect 7432 25004 7440 25068
rect 7120 25003 7440 25004
rect 12448 25068 12768 25069
rect 12448 25004 12456 25068
rect 12520 25004 12536 25068
rect 12600 25004 12616 25068
rect 12680 25004 12696 25068
rect 12760 25004 12768 25068
rect 12448 25003 12768 25004
rect 17776 25068 18096 25069
rect 17776 25004 17784 25068
rect 17848 25004 17864 25068
rect 17928 25004 17944 25068
rect 18008 25004 18024 25068
rect 18088 25004 18096 25068
rect 17776 25003 18096 25004
rect 2063 24696 2129 24699
rect 830 24694 2129 24696
rect 830 24638 2068 24694
rect 2124 24638 2129 24694
rect 830 24636 2129 24638
rect 830 24472 890 24636
rect 2063 24633 2129 24636
rect 800 24216 920 24472
rect 4456 24402 4776 24403
rect 4456 24338 4464 24402
rect 4528 24338 4544 24402
rect 4608 24338 4624 24402
rect 4688 24338 4704 24402
rect 4768 24338 4776 24402
rect 4456 24337 4776 24338
rect 9784 24402 10104 24403
rect 9784 24338 9792 24402
rect 9856 24338 9872 24402
rect 9936 24338 9952 24402
rect 10016 24338 10032 24402
rect 10096 24338 10104 24402
rect 9784 24337 10104 24338
rect 15112 24402 15432 24403
rect 15112 24338 15120 24402
rect 15184 24338 15200 24402
rect 15264 24338 15280 24402
rect 15344 24338 15360 24402
rect 15424 24338 15432 24402
rect 15112 24337 15432 24338
rect 20440 24402 20760 24403
rect 20440 24338 20448 24402
rect 20512 24338 20528 24402
rect 20592 24338 20608 24402
rect 20672 24338 20688 24402
rect 20752 24338 20760 24402
rect 20440 24337 20760 24338
rect 7120 23736 7440 23737
rect 7120 23672 7128 23736
rect 7192 23672 7208 23736
rect 7272 23672 7288 23736
rect 7352 23672 7368 23736
rect 7432 23672 7440 23736
rect 7120 23671 7440 23672
rect 12448 23736 12768 23737
rect 12448 23672 12456 23736
rect 12520 23672 12536 23736
rect 12600 23672 12616 23736
rect 12680 23672 12696 23736
rect 12760 23672 12768 23736
rect 12448 23671 12768 23672
rect 17776 23736 18096 23737
rect 17776 23672 17784 23736
rect 17848 23672 17864 23736
rect 17928 23672 17944 23736
rect 18008 23672 18024 23736
rect 18088 23672 18096 23736
rect 17776 23671 18096 23672
rect 2063 23364 2129 23367
rect 830 23362 2129 23364
rect 830 23306 2068 23362
rect 2124 23306 2129 23362
rect 830 23304 2129 23306
rect 830 23112 890 23304
rect 2063 23301 2129 23304
rect 800 22856 920 23112
rect 4456 23070 4776 23071
rect 4456 23006 4464 23070
rect 4528 23006 4544 23070
rect 4608 23006 4624 23070
rect 4688 23006 4704 23070
rect 4768 23006 4776 23070
rect 4456 23005 4776 23006
rect 9784 23070 10104 23071
rect 9784 23006 9792 23070
rect 9856 23006 9872 23070
rect 9936 23006 9952 23070
rect 10016 23006 10032 23070
rect 10096 23006 10104 23070
rect 9784 23005 10104 23006
rect 15112 23070 15432 23071
rect 15112 23006 15120 23070
rect 15184 23006 15200 23070
rect 15264 23006 15280 23070
rect 15344 23006 15360 23070
rect 15424 23006 15432 23070
rect 15112 23005 15432 23006
rect 20440 23070 20760 23071
rect 20440 23006 20448 23070
rect 20512 23006 20528 23070
rect 20592 23006 20608 23070
rect 20672 23006 20688 23070
rect 20752 23006 20760 23070
rect 20440 23005 20760 23006
rect 7120 22404 7440 22405
rect 7120 22340 7128 22404
rect 7192 22340 7208 22404
rect 7272 22340 7288 22404
rect 7352 22340 7368 22404
rect 7432 22340 7440 22404
rect 7120 22339 7440 22340
rect 12448 22404 12768 22405
rect 12448 22340 12456 22404
rect 12520 22340 12536 22404
rect 12600 22340 12616 22404
rect 12680 22340 12696 22404
rect 12760 22340 12768 22404
rect 12448 22339 12768 22340
rect 17776 22404 18096 22405
rect 17776 22340 17784 22404
rect 17848 22340 17864 22404
rect 17928 22340 17944 22404
rect 18008 22340 18024 22404
rect 18088 22340 18096 22404
rect 17776 22339 18096 22340
rect 830 21972 1118 22032
rect 830 21888 890 21972
rect 800 21632 920 21888
rect 1058 21884 1118 21972
rect 2063 21884 2129 21887
rect 1058 21882 2129 21884
rect 1058 21826 2068 21882
rect 2124 21826 2129 21882
rect 1058 21824 2129 21826
rect 2063 21821 2129 21824
rect 4456 21738 4776 21739
rect 4456 21674 4464 21738
rect 4528 21674 4544 21738
rect 4608 21674 4624 21738
rect 4688 21674 4704 21738
rect 4768 21674 4776 21738
rect 4456 21673 4776 21674
rect 9784 21738 10104 21739
rect 9784 21674 9792 21738
rect 9856 21674 9872 21738
rect 9936 21674 9952 21738
rect 10016 21674 10032 21738
rect 10096 21674 10104 21738
rect 9784 21673 10104 21674
rect 15112 21738 15432 21739
rect 15112 21674 15120 21738
rect 15184 21674 15200 21738
rect 15264 21674 15280 21738
rect 15344 21674 15360 21738
rect 15424 21674 15432 21738
rect 15112 21673 15432 21674
rect 20440 21738 20760 21739
rect 20440 21674 20448 21738
rect 20512 21674 20528 21738
rect 20592 21674 20608 21738
rect 20672 21674 20688 21738
rect 20752 21674 20760 21738
rect 20440 21673 20760 21674
rect 7120 21072 7440 21073
rect 7120 21008 7128 21072
rect 7192 21008 7208 21072
rect 7272 21008 7288 21072
rect 7352 21008 7368 21072
rect 7432 21008 7440 21072
rect 7120 21007 7440 21008
rect 12448 21072 12768 21073
rect 12448 21008 12456 21072
rect 12520 21008 12536 21072
rect 12600 21008 12616 21072
rect 12680 21008 12696 21072
rect 12760 21008 12768 21072
rect 12448 21007 12768 21008
rect 17776 21072 18096 21073
rect 17776 21008 17784 21072
rect 17848 21008 17864 21072
rect 17928 21008 17944 21072
rect 18008 21008 18024 21072
rect 18088 21008 18096 21072
rect 17776 21007 18096 21008
rect 800 20272 920 20528
rect 4456 20406 4776 20407
rect 4456 20342 4464 20406
rect 4528 20342 4544 20406
rect 4608 20342 4624 20406
rect 4688 20342 4704 20406
rect 4768 20342 4776 20406
rect 4456 20341 4776 20342
rect 9784 20406 10104 20407
rect 9784 20342 9792 20406
rect 9856 20342 9872 20406
rect 9936 20342 9952 20406
rect 10016 20342 10032 20406
rect 10096 20342 10104 20406
rect 9784 20341 10104 20342
rect 15112 20406 15432 20407
rect 15112 20342 15120 20406
rect 15184 20342 15200 20406
rect 15264 20342 15280 20406
rect 15344 20342 15360 20406
rect 15424 20342 15432 20406
rect 15112 20341 15432 20342
rect 20440 20406 20760 20407
rect 20440 20342 20448 20406
rect 20512 20342 20528 20406
rect 20592 20342 20608 20406
rect 20672 20342 20688 20406
rect 20752 20342 20760 20406
rect 20440 20341 20760 20342
rect 830 20108 890 20272
rect 2447 20108 2513 20111
rect 830 20106 2513 20108
rect 830 20050 2452 20106
rect 2508 20050 2513 20106
rect 830 20048 2513 20050
rect 2447 20045 2513 20048
rect 7120 19740 7440 19741
rect 7120 19676 7128 19740
rect 7192 19676 7208 19740
rect 7272 19676 7288 19740
rect 7352 19676 7368 19740
rect 7432 19676 7440 19740
rect 7120 19675 7440 19676
rect 12448 19740 12768 19741
rect 12448 19676 12456 19740
rect 12520 19676 12536 19740
rect 12600 19676 12616 19740
rect 12680 19676 12696 19740
rect 12760 19676 12768 19740
rect 12448 19675 12768 19676
rect 17776 19740 18096 19741
rect 17776 19676 17784 19740
rect 17848 19676 17864 19740
rect 17928 19676 17944 19740
rect 18008 19676 18024 19740
rect 18088 19676 18096 19740
rect 17776 19675 18096 19676
rect 2063 19368 2129 19371
rect 830 19366 2129 19368
rect 830 19310 2068 19366
rect 2124 19310 2129 19366
rect 830 19308 2129 19310
rect 830 19168 890 19308
rect 2063 19305 2129 19308
rect 800 18912 920 19168
rect 4456 19074 4776 19075
rect 4456 19010 4464 19074
rect 4528 19010 4544 19074
rect 4608 19010 4624 19074
rect 4688 19010 4704 19074
rect 4768 19010 4776 19074
rect 4456 19009 4776 19010
rect 9784 19074 10104 19075
rect 9784 19010 9792 19074
rect 9856 19010 9872 19074
rect 9936 19010 9952 19074
rect 10016 19010 10032 19074
rect 10096 19010 10104 19074
rect 9784 19009 10104 19010
rect 15112 19074 15432 19075
rect 15112 19010 15120 19074
rect 15184 19010 15200 19074
rect 15264 19010 15280 19074
rect 15344 19010 15360 19074
rect 15424 19010 15432 19074
rect 15112 19009 15432 19010
rect 20440 19074 20760 19075
rect 20440 19010 20448 19074
rect 20512 19010 20528 19074
rect 20592 19010 20608 19074
rect 20672 19010 20688 19074
rect 20752 19010 20760 19074
rect 20440 19009 20760 19010
rect 7120 18408 7440 18409
rect 7120 18344 7128 18408
rect 7192 18344 7208 18408
rect 7272 18344 7288 18408
rect 7352 18344 7368 18408
rect 7432 18344 7440 18408
rect 7120 18343 7440 18344
rect 12448 18408 12768 18409
rect 12448 18344 12456 18408
rect 12520 18344 12536 18408
rect 12600 18344 12616 18408
rect 12680 18344 12696 18408
rect 12760 18344 12768 18408
rect 12448 18343 12768 18344
rect 17776 18408 18096 18409
rect 17776 18344 17784 18408
rect 17848 18344 17864 18408
rect 17928 18344 17944 18408
rect 18008 18344 18024 18408
rect 18088 18344 18096 18408
rect 17776 18343 18096 18344
rect 4456 17742 4776 17743
rect 4456 17678 4464 17742
rect 4528 17678 4544 17742
rect 4608 17678 4624 17742
rect 4688 17678 4704 17742
rect 4768 17678 4776 17742
rect 4456 17677 4776 17678
rect 9784 17742 10104 17743
rect 9784 17678 9792 17742
rect 9856 17678 9872 17742
rect 9936 17678 9952 17742
rect 10016 17678 10032 17742
rect 10096 17678 10104 17742
rect 9784 17677 10104 17678
rect 15112 17742 15432 17743
rect 15112 17678 15120 17742
rect 15184 17678 15200 17742
rect 15264 17678 15280 17742
rect 15344 17678 15360 17742
rect 15424 17678 15432 17742
rect 15112 17677 15432 17678
rect 20440 17742 20760 17743
rect 20440 17678 20448 17742
rect 20512 17678 20528 17742
rect 20592 17678 20608 17742
rect 20672 17678 20688 17742
rect 20752 17678 20760 17742
rect 20440 17677 20760 17678
rect 7120 17076 7440 17077
rect 7120 17012 7128 17076
rect 7192 17012 7208 17076
rect 7272 17012 7288 17076
rect 7352 17012 7368 17076
rect 7432 17012 7440 17076
rect 7120 17011 7440 17012
rect 12448 17076 12768 17077
rect 12448 17012 12456 17076
rect 12520 17012 12536 17076
rect 12600 17012 12616 17076
rect 12680 17012 12696 17076
rect 12760 17012 12768 17076
rect 12448 17011 12768 17012
rect 17776 17076 18096 17077
rect 17776 17012 17784 17076
rect 17848 17012 17864 17076
rect 17928 17012 17944 17076
rect 18008 17012 18024 17076
rect 18088 17012 18096 17076
rect 17776 17011 18096 17012
rect 800 16192 920 16448
rect 4456 16410 4776 16411
rect 4456 16346 4464 16410
rect 4528 16346 4544 16410
rect 4608 16346 4624 16410
rect 4688 16346 4704 16410
rect 4768 16346 4776 16410
rect 4456 16345 4776 16346
rect 9784 16410 10104 16411
rect 9784 16346 9792 16410
rect 9856 16346 9872 16410
rect 9936 16346 9952 16410
rect 10016 16346 10032 16410
rect 10096 16346 10104 16410
rect 9784 16345 10104 16346
rect 15112 16410 15432 16411
rect 15112 16346 15120 16410
rect 15184 16346 15200 16410
rect 15264 16346 15280 16410
rect 15344 16346 15360 16410
rect 15424 16346 15432 16410
rect 15112 16345 15432 16346
rect 20440 16410 20760 16411
rect 20440 16346 20448 16410
rect 20512 16346 20528 16410
rect 20592 16346 20608 16410
rect 20672 16346 20688 16410
rect 20752 16346 20760 16410
rect 20440 16345 20760 16346
rect 830 16112 890 16192
rect 2063 16112 2129 16115
rect 830 16110 2129 16112
rect 830 16054 2068 16110
rect 2124 16054 2129 16110
rect 830 16052 2129 16054
rect 2063 16049 2129 16052
rect 7120 15744 7440 15745
rect 7120 15680 7128 15744
rect 7192 15680 7208 15744
rect 7272 15680 7288 15744
rect 7352 15680 7368 15744
rect 7432 15680 7440 15744
rect 7120 15679 7440 15680
rect 12448 15744 12768 15745
rect 12448 15680 12456 15744
rect 12520 15680 12536 15744
rect 12600 15680 12616 15744
rect 12680 15680 12696 15744
rect 12760 15680 12768 15744
rect 12448 15679 12768 15680
rect 17776 15744 18096 15745
rect 17776 15680 17784 15744
rect 17848 15680 17864 15744
rect 17928 15680 17944 15744
rect 18008 15680 18024 15744
rect 18088 15680 18096 15744
rect 17776 15679 18096 15680
rect 4456 15078 4776 15079
rect 4456 15014 4464 15078
rect 4528 15014 4544 15078
rect 4608 15014 4624 15078
rect 4688 15014 4704 15078
rect 4768 15014 4776 15078
rect 4456 15013 4776 15014
rect 9784 15078 10104 15079
rect 9784 15014 9792 15078
rect 9856 15014 9872 15078
rect 9936 15014 9952 15078
rect 10016 15014 10032 15078
rect 10096 15014 10104 15078
rect 9784 15013 10104 15014
rect 15112 15078 15432 15079
rect 15112 15014 15120 15078
rect 15184 15014 15200 15078
rect 15264 15014 15280 15078
rect 15344 15014 15360 15078
rect 15424 15014 15432 15078
rect 15112 15013 15432 15014
rect 20440 15078 20760 15079
rect 20440 15014 20448 15078
rect 20512 15014 20528 15078
rect 20592 15014 20608 15078
rect 20672 15014 20688 15078
rect 20752 15014 20760 15078
rect 20440 15013 20760 15014
rect 7120 14412 7440 14413
rect 7120 14348 7128 14412
rect 7192 14348 7208 14412
rect 7272 14348 7288 14412
rect 7352 14348 7368 14412
rect 7432 14348 7440 14412
rect 7120 14347 7440 14348
rect 12448 14412 12768 14413
rect 12448 14348 12456 14412
rect 12520 14348 12536 14412
rect 12600 14348 12616 14412
rect 12680 14348 12696 14412
rect 12760 14348 12768 14412
rect 12448 14347 12768 14348
rect 17776 14412 18096 14413
rect 17776 14348 17784 14412
rect 17848 14348 17864 14412
rect 17928 14348 17944 14412
rect 18008 14348 18024 14412
rect 18088 14348 18096 14412
rect 17776 14347 18096 14348
rect 4456 13746 4776 13747
rect 4456 13682 4464 13746
rect 4528 13682 4544 13746
rect 4608 13682 4624 13746
rect 4688 13682 4704 13746
rect 4768 13682 4776 13746
rect 4456 13681 4776 13682
rect 9784 13746 10104 13747
rect 9784 13682 9792 13746
rect 9856 13682 9872 13746
rect 9936 13682 9952 13746
rect 10016 13682 10032 13746
rect 10096 13682 10104 13746
rect 9784 13681 10104 13682
rect 15112 13746 15432 13747
rect 15112 13682 15120 13746
rect 15184 13682 15200 13746
rect 15264 13682 15280 13746
rect 15344 13682 15360 13746
rect 15424 13682 15432 13746
rect 15112 13681 15432 13682
rect 20440 13746 20760 13747
rect 20440 13682 20448 13746
rect 20512 13682 20528 13746
rect 20592 13682 20608 13746
rect 20672 13682 20688 13746
rect 20752 13682 20760 13746
rect 20440 13681 20760 13682
rect 7120 13080 7440 13081
rect 7120 13016 7128 13080
rect 7192 13016 7208 13080
rect 7272 13016 7288 13080
rect 7352 13016 7368 13080
rect 7432 13016 7440 13080
rect 7120 13015 7440 13016
rect 12448 13080 12768 13081
rect 12448 13016 12456 13080
rect 12520 13016 12536 13080
rect 12600 13016 12616 13080
rect 12680 13016 12696 13080
rect 12760 13016 12768 13080
rect 12448 13015 12768 13016
rect 17776 13080 18096 13081
rect 17776 13016 17784 13080
rect 17848 13016 17864 13080
rect 17928 13016 17944 13080
rect 18008 13016 18024 13080
rect 18088 13016 18096 13080
rect 17776 13015 18096 13016
rect 4456 12414 4776 12415
rect 4456 12350 4464 12414
rect 4528 12350 4544 12414
rect 4608 12350 4624 12414
rect 4688 12350 4704 12414
rect 4768 12350 4776 12414
rect 4456 12349 4776 12350
rect 9784 12414 10104 12415
rect 9784 12350 9792 12414
rect 9856 12350 9872 12414
rect 9936 12350 9952 12414
rect 10016 12350 10032 12414
rect 10096 12350 10104 12414
rect 9784 12349 10104 12350
rect 15112 12414 15432 12415
rect 15112 12350 15120 12414
rect 15184 12350 15200 12414
rect 15264 12350 15280 12414
rect 15344 12350 15360 12414
rect 15424 12350 15432 12414
rect 15112 12349 15432 12350
rect 20440 12414 20760 12415
rect 20440 12350 20448 12414
rect 20512 12350 20528 12414
rect 20592 12350 20608 12414
rect 20672 12350 20688 12414
rect 20752 12350 20760 12414
rect 20440 12349 20760 12350
rect 7120 11748 7440 11749
rect 7120 11684 7128 11748
rect 7192 11684 7208 11748
rect 7272 11684 7288 11748
rect 7352 11684 7368 11748
rect 7432 11684 7440 11748
rect 7120 11683 7440 11684
rect 12448 11748 12768 11749
rect 12448 11684 12456 11748
rect 12520 11684 12536 11748
rect 12600 11684 12616 11748
rect 12680 11684 12696 11748
rect 12760 11684 12768 11748
rect 12448 11683 12768 11684
rect 17776 11748 18096 11749
rect 17776 11684 17784 11748
rect 17848 11684 17864 11748
rect 17928 11684 17944 11748
rect 18008 11684 18024 11748
rect 18088 11684 18096 11748
rect 17776 11683 18096 11684
rect 800 10888 920 11144
rect 4456 11082 4776 11083
rect 4456 11018 4464 11082
rect 4528 11018 4544 11082
rect 4608 11018 4624 11082
rect 4688 11018 4704 11082
rect 4768 11018 4776 11082
rect 4456 11017 4776 11018
rect 9784 11082 10104 11083
rect 9784 11018 9792 11082
rect 9856 11018 9872 11082
rect 9936 11018 9952 11082
rect 10016 11018 10032 11082
rect 10096 11018 10104 11082
rect 9784 11017 10104 11018
rect 15112 11082 15432 11083
rect 15112 11018 15120 11082
rect 15184 11018 15200 11082
rect 15264 11018 15280 11082
rect 15344 11018 15360 11082
rect 15424 11018 15432 11082
rect 15112 11017 15432 11018
rect 20440 11082 20760 11083
rect 20440 11018 20448 11082
rect 20512 11018 20528 11082
rect 20592 11018 20608 11082
rect 20672 11018 20688 11082
rect 20752 11018 20760 11082
rect 20440 11017 20760 11018
rect 830 10784 890 10888
rect 2063 10784 2129 10787
rect 830 10782 2129 10784
rect 830 10726 2068 10782
rect 2124 10726 2129 10782
rect 830 10724 2129 10726
rect 2063 10721 2129 10724
rect 7120 10416 7440 10417
rect 7120 10352 7128 10416
rect 7192 10352 7208 10416
rect 7272 10352 7288 10416
rect 7352 10352 7368 10416
rect 7432 10352 7440 10416
rect 7120 10351 7440 10352
rect 12448 10416 12768 10417
rect 12448 10352 12456 10416
rect 12520 10352 12536 10416
rect 12600 10352 12616 10416
rect 12680 10352 12696 10416
rect 12760 10352 12768 10416
rect 12448 10351 12768 10352
rect 17776 10416 18096 10417
rect 17776 10352 17784 10416
rect 17848 10352 17864 10416
rect 17928 10352 17944 10416
rect 18008 10352 18024 10416
rect 18088 10352 18096 10416
rect 17776 10351 18096 10352
rect 4456 9750 4776 9751
rect 4456 9686 4464 9750
rect 4528 9686 4544 9750
rect 4608 9686 4624 9750
rect 4688 9686 4704 9750
rect 4768 9686 4776 9750
rect 4456 9685 4776 9686
rect 9784 9750 10104 9751
rect 9784 9686 9792 9750
rect 9856 9686 9872 9750
rect 9936 9686 9952 9750
rect 10016 9686 10032 9750
rect 10096 9686 10104 9750
rect 9784 9685 10104 9686
rect 15112 9750 15432 9751
rect 15112 9686 15120 9750
rect 15184 9686 15200 9750
rect 15264 9686 15280 9750
rect 15344 9686 15360 9750
rect 15424 9686 15432 9750
rect 15112 9685 15432 9686
rect 20440 9750 20760 9751
rect 20440 9686 20448 9750
rect 20512 9686 20528 9750
rect 20592 9686 20608 9750
rect 20672 9686 20688 9750
rect 20752 9686 20760 9750
rect 20440 9685 20760 9686
rect 7120 9084 7440 9085
rect 7120 9020 7128 9084
rect 7192 9020 7208 9084
rect 7272 9020 7288 9084
rect 7352 9020 7368 9084
rect 7432 9020 7440 9084
rect 7120 9019 7440 9020
rect 12448 9084 12768 9085
rect 12448 9020 12456 9084
rect 12520 9020 12536 9084
rect 12600 9020 12616 9084
rect 12680 9020 12696 9084
rect 12760 9020 12768 9084
rect 12448 9019 12768 9020
rect 17776 9084 18096 9085
rect 17776 9020 17784 9084
rect 17848 9020 17864 9084
rect 17928 9020 17944 9084
rect 18008 9020 18024 9084
rect 18088 9020 18096 9084
rect 17776 9019 18096 9020
rect 4456 8418 4776 8419
rect 4456 8354 4464 8418
rect 4528 8354 4544 8418
rect 4608 8354 4624 8418
rect 4688 8354 4704 8418
rect 4768 8354 4776 8418
rect 4456 8353 4776 8354
rect 9784 8418 10104 8419
rect 9784 8354 9792 8418
rect 9856 8354 9872 8418
rect 9936 8354 9952 8418
rect 10016 8354 10032 8418
rect 10096 8354 10104 8418
rect 9784 8353 10104 8354
rect 15112 8418 15432 8419
rect 15112 8354 15120 8418
rect 15184 8354 15200 8418
rect 15264 8354 15280 8418
rect 15344 8354 15360 8418
rect 15424 8354 15432 8418
rect 15112 8353 15432 8354
rect 20440 8418 20760 8419
rect 20440 8354 20448 8418
rect 20512 8354 20528 8418
rect 20592 8354 20608 8418
rect 20672 8354 20688 8418
rect 20752 8354 20760 8418
rect 20440 8353 20760 8354
rect 7120 7752 7440 7753
rect 7120 7688 7128 7752
rect 7192 7688 7208 7752
rect 7272 7688 7288 7752
rect 7352 7688 7368 7752
rect 7432 7688 7440 7752
rect 7120 7687 7440 7688
rect 12448 7752 12768 7753
rect 12448 7688 12456 7752
rect 12520 7688 12536 7752
rect 12600 7688 12616 7752
rect 12680 7688 12696 7752
rect 12760 7688 12768 7752
rect 12448 7687 12768 7688
rect 17776 7752 18096 7753
rect 17776 7688 17784 7752
rect 17848 7688 17864 7752
rect 17928 7688 17944 7752
rect 18008 7688 18024 7752
rect 18088 7688 18096 7752
rect 17776 7687 18096 7688
rect 4456 7086 4776 7087
rect 4456 7022 4464 7086
rect 4528 7022 4544 7086
rect 4608 7022 4624 7086
rect 4688 7022 4704 7086
rect 4768 7022 4776 7086
rect 4456 7021 4776 7022
rect 9784 7086 10104 7087
rect 9784 7022 9792 7086
rect 9856 7022 9872 7086
rect 9936 7022 9952 7086
rect 10016 7022 10032 7086
rect 10096 7022 10104 7086
rect 9784 7021 10104 7022
rect 15112 7086 15432 7087
rect 15112 7022 15120 7086
rect 15184 7022 15200 7086
rect 15264 7022 15280 7086
rect 15344 7022 15360 7086
rect 15424 7022 15432 7086
rect 15112 7021 15432 7022
rect 20440 7086 20760 7087
rect 20440 7022 20448 7086
rect 20512 7022 20528 7086
rect 20592 7022 20608 7086
rect 20672 7022 20688 7086
rect 20752 7022 20760 7086
rect 20440 7021 20760 7022
rect 7120 6420 7440 6421
rect 7120 6356 7128 6420
rect 7192 6356 7208 6420
rect 7272 6356 7288 6420
rect 7352 6356 7368 6420
rect 7432 6356 7440 6420
rect 7120 6355 7440 6356
rect 12448 6420 12768 6421
rect 12448 6356 12456 6420
rect 12520 6356 12536 6420
rect 12600 6356 12616 6420
rect 12680 6356 12696 6420
rect 12760 6356 12768 6420
rect 12448 6355 12768 6356
rect 17776 6420 18096 6421
rect 17776 6356 17784 6420
rect 17848 6356 17864 6420
rect 17928 6356 17944 6420
rect 18008 6356 18024 6420
rect 18088 6356 18096 6420
rect 17776 6355 18096 6356
rect 4456 5754 4776 5755
rect 4456 5690 4464 5754
rect 4528 5690 4544 5754
rect 4608 5690 4624 5754
rect 4688 5690 4704 5754
rect 4768 5690 4776 5754
rect 4456 5689 4776 5690
rect 9784 5754 10104 5755
rect 9784 5690 9792 5754
rect 9856 5690 9872 5754
rect 9936 5690 9952 5754
rect 10016 5690 10032 5754
rect 10096 5690 10104 5754
rect 9784 5689 10104 5690
rect 15112 5754 15432 5755
rect 15112 5690 15120 5754
rect 15184 5690 15200 5754
rect 15264 5690 15280 5754
rect 15344 5690 15360 5754
rect 15424 5690 15432 5754
rect 15112 5689 15432 5690
rect 20440 5754 20760 5755
rect 20440 5690 20448 5754
rect 20512 5690 20528 5754
rect 20592 5690 20608 5754
rect 20672 5690 20688 5754
rect 20752 5690 20760 5754
rect 20440 5689 20760 5690
rect 7120 5088 7440 5089
rect 7120 5024 7128 5088
rect 7192 5024 7208 5088
rect 7272 5024 7288 5088
rect 7352 5024 7368 5088
rect 7432 5024 7440 5088
rect 7120 5023 7440 5024
rect 12448 5088 12768 5089
rect 12448 5024 12456 5088
rect 12520 5024 12536 5088
rect 12600 5024 12616 5088
rect 12680 5024 12696 5088
rect 12760 5024 12768 5088
rect 12448 5023 12768 5024
rect 17776 5088 18096 5089
rect 17776 5024 17784 5088
rect 17848 5024 17864 5088
rect 17928 5024 17944 5088
rect 18008 5024 18024 5088
rect 18088 5024 18096 5088
rect 17776 5023 18096 5024
rect 4456 4422 4776 4423
rect 4456 4358 4464 4422
rect 4528 4358 4544 4422
rect 4608 4358 4624 4422
rect 4688 4358 4704 4422
rect 4768 4358 4776 4422
rect 4456 4357 4776 4358
rect 9784 4422 10104 4423
rect 9784 4358 9792 4422
rect 9856 4358 9872 4422
rect 9936 4358 9952 4422
rect 10016 4358 10032 4422
rect 10096 4358 10104 4422
rect 9784 4357 10104 4358
rect 15112 4422 15432 4423
rect 15112 4358 15120 4422
rect 15184 4358 15200 4422
rect 15264 4358 15280 4422
rect 15344 4358 15360 4422
rect 15424 4358 15432 4422
rect 15112 4357 15432 4358
rect 20440 4422 20760 4423
rect 20440 4358 20448 4422
rect 20512 4358 20528 4422
rect 20592 4358 20608 4422
rect 20672 4358 20688 4422
rect 20752 4358 20760 4422
rect 20440 4357 20760 4358
rect 7120 3756 7440 3757
rect 7120 3692 7128 3756
rect 7192 3692 7208 3756
rect 7272 3692 7288 3756
rect 7352 3692 7368 3756
rect 7432 3692 7440 3756
rect 7120 3691 7440 3692
rect 12448 3756 12768 3757
rect 12448 3692 12456 3756
rect 12520 3692 12536 3756
rect 12600 3692 12616 3756
rect 12680 3692 12696 3756
rect 12760 3692 12768 3756
rect 12448 3691 12768 3692
rect 17776 3756 18096 3757
rect 17776 3692 17784 3756
rect 17848 3692 17864 3756
rect 17928 3692 17944 3756
rect 18008 3692 18024 3756
rect 18088 3692 18096 3756
rect 17776 3691 18096 3692
rect 4456 3090 4776 3091
rect 4456 3026 4464 3090
rect 4528 3026 4544 3090
rect 4608 3026 4624 3090
rect 4688 3026 4704 3090
rect 4768 3026 4776 3090
rect 4456 3025 4776 3026
rect 9784 3090 10104 3091
rect 9784 3026 9792 3090
rect 9856 3026 9872 3090
rect 9936 3026 9952 3090
rect 10016 3026 10032 3090
rect 10096 3026 10104 3090
rect 9784 3025 10104 3026
rect 15112 3090 15432 3091
rect 15112 3026 15120 3090
rect 15184 3026 15200 3090
rect 15264 3026 15280 3090
rect 15344 3026 15360 3090
rect 15424 3026 15432 3090
rect 15112 3025 15432 3026
rect 20440 3090 20760 3091
rect 20440 3026 20448 3090
rect 20512 3026 20528 3090
rect 20592 3026 20608 3090
rect 20672 3026 20688 3090
rect 20752 3026 20760 3090
rect 20440 3025 20760 3026
rect 7120 2424 7440 2425
rect 7120 2360 7128 2424
rect 7192 2360 7208 2424
rect 7272 2360 7288 2424
rect 7352 2360 7368 2424
rect 7432 2360 7440 2424
rect 7120 2359 7440 2360
rect 12448 2424 12768 2425
rect 12448 2360 12456 2424
rect 12520 2360 12536 2424
rect 12600 2360 12616 2424
rect 12680 2360 12696 2424
rect 12760 2360 12768 2424
rect 12448 2359 12768 2360
rect 17776 2424 18096 2425
rect 17776 2360 17784 2424
rect 17848 2360 17864 2424
rect 17928 2360 17944 2424
rect 18008 2360 18024 2424
rect 18088 2360 18096 2424
rect 17776 2359 18096 2360
rect 4456 1758 4776 1759
rect 4456 1694 4464 1758
rect 4528 1694 4544 1758
rect 4608 1694 4624 1758
rect 4688 1694 4704 1758
rect 4768 1694 4776 1758
rect 4456 1693 4776 1694
rect 9784 1758 10104 1759
rect 9784 1694 9792 1758
rect 9856 1694 9872 1758
rect 9936 1694 9952 1758
rect 10016 1694 10032 1758
rect 10096 1694 10104 1758
rect 9784 1693 10104 1694
rect 15112 1758 15432 1759
rect 15112 1694 15120 1758
rect 15184 1694 15200 1758
rect 15264 1694 15280 1758
rect 15344 1694 15360 1758
rect 15424 1694 15432 1758
rect 15112 1693 15432 1694
rect 20440 1758 20760 1759
rect 20440 1694 20448 1758
rect 20512 1694 20528 1758
rect 20592 1694 20608 1758
rect 20672 1694 20688 1758
rect 20752 1694 20760 1758
rect 20440 1693 20760 1694
rect 800 960 920 1216
rect 7120 1092 7440 1093
rect 7120 1028 7128 1092
rect 7192 1028 7208 1092
rect 7272 1028 7288 1092
rect 7352 1028 7368 1092
rect 7432 1028 7440 1092
rect 7120 1027 7440 1028
rect 12448 1092 12768 1093
rect 12448 1028 12456 1092
rect 12520 1028 12536 1092
rect 12600 1028 12616 1092
rect 12680 1028 12696 1092
rect 12760 1028 12768 1092
rect 12448 1027 12768 1028
rect 17776 1092 18096 1093
rect 17776 1028 17784 1092
rect 17848 1028 17864 1092
rect 17928 1028 17944 1092
rect 18008 1028 18024 1092
rect 18088 1028 18096 1092
rect 17776 1027 18096 1028
rect 830 868 890 960
rect 3023 868 3089 871
rect 830 866 3089 868
rect 830 810 3028 866
rect 3084 810 3089 866
rect 830 808 3089 810
rect 3023 805 3089 808
<< via3 >>
rect 4464 27062 4528 27066
rect 4464 27006 4468 27062
rect 4468 27006 4524 27062
rect 4524 27006 4528 27062
rect 4464 27002 4528 27006
rect 4544 27062 4608 27066
rect 4544 27006 4548 27062
rect 4548 27006 4604 27062
rect 4604 27006 4608 27062
rect 4544 27002 4608 27006
rect 4624 27062 4688 27066
rect 4624 27006 4628 27062
rect 4628 27006 4684 27062
rect 4684 27006 4688 27062
rect 4624 27002 4688 27006
rect 4704 27062 4768 27066
rect 4704 27006 4708 27062
rect 4708 27006 4764 27062
rect 4764 27006 4768 27062
rect 4704 27002 4768 27006
rect 9792 27062 9856 27066
rect 9792 27006 9796 27062
rect 9796 27006 9852 27062
rect 9852 27006 9856 27062
rect 9792 27002 9856 27006
rect 9872 27062 9936 27066
rect 9872 27006 9876 27062
rect 9876 27006 9932 27062
rect 9932 27006 9936 27062
rect 9872 27002 9936 27006
rect 9952 27062 10016 27066
rect 9952 27006 9956 27062
rect 9956 27006 10012 27062
rect 10012 27006 10016 27062
rect 9952 27002 10016 27006
rect 10032 27062 10096 27066
rect 10032 27006 10036 27062
rect 10036 27006 10092 27062
rect 10092 27006 10096 27062
rect 10032 27002 10096 27006
rect 15120 27062 15184 27066
rect 15120 27006 15124 27062
rect 15124 27006 15180 27062
rect 15180 27006 15184 27062
rect 15120 27002 15184 27006
rect 15200 27062 15264 27066
rect 15200 27006 15204 27062
rect 15204 27006 15260 27062
rect 15260 27006 15264 27062
rect 15200 27002 15264 27006
rect 15280 27062 15344 27066
rect 15280 27006 15284 27062
rect 15284 27006 15340 27062
rect 15340 27006 15344 27062
rect 15280 27002 15344 27006
rect 15360 27062 15424 27066
rect 15360 27006 15364 27062
rect 15364 27006 15420 27062
rect 15420 27006 15424 27062
rect 15360 27002 15424 27006
rect 20448 27062 20512 27066
rect 20448 27006 20452 27062
rect 20452 27006 20508 27062
rect 20508 27006 20512 27062
rect 20448 27002 20512 27006
rect 20528 27062 20592 27066
rect 20528 27006 20532 27062
rect 20532 27006 20588 27062
rect 20588 27006 20592 27062
rect 20528 27002 20592 27006
rect 20608 27062 20672 27066
rect 20608 27006 20612 27062
rect 20612 27006 20668 27062
rect 20668 27006 20672 27062
rect 20608 27002 20672 27006
rect 20688 27062 20752 27066
rect 20688 27006 20692 27062
rect 20692 27006 20748 27062
rect 20748 27006 20752 27062
rect 20688 27002 20752 27006
rect 7128 26396 7192 26400
rect 7128 26340 7132 26396
rect 7132 26340 7188 26396
rect 7188 26340 7192 26396
rect 7128 26336 7192 26340
rect 7208 26396 7272 26400
rect 7208 26340 7212 26396
rect 7212 26340 7268 26396
rect 7268 26340 7272 26396
rect 7208 26336 7272 26340
rect 7288 26396 7352 26400
rect 7288 26340 7292 26396
rect 7292 26340 7348 26396
rect 7348 26340 7352 26396
rect 7288 26336 7352 26340
rect 7368 26396 7432 26400
rect 7368 26340 7372 26396
rect 7372 26340 7428 26396
rect 7428 26340 7432 26396
rect 7368 26336 7432 26340
rect 12456 26396 12520 26400
rect 12456 26340 12460 26396
rect 12460 26340 12516 26396
rect 12516 26340 12520 26396
rect 12456 26336 12520 26340
rect 12536 26396 12600 26400
rect 12536 26340 12540 26396
rect 12540 26340 12596 26396
rect 12596 26340 12600 26396
rect 12536 26336 12600 26340
rect 12616 26396 12680 26400
rect 12616 26340 12620 26396
rect 12620 26340 12676 26396
rect 12676 26340 12680 26396
rect 12616 26336 12680 26340
rect 12696 26396 12760 26400
rect 12696 26340 12700 26396
rect 12700 26340 12756 26396
rect 12756 26340 12760 26396
rect 12696 26336 12760 26340
rect 17784 26396 17848 26400
rect 17784 26340 17788 26396
rect 17788 26340 17844 26396
rect 17844 26340 17848 26396
rect 17784 26336 17848 26340
rect 17864 26396 17928 26400
rect 17864 26340 17868 26396
rect 17868 26340 17924 26396
rect 17924 26340 17928 26396
rect 17864 26336 17928 26340
rect 17944 26396 18008 26400
rect 17944 26340 17948 26396
rect 17948 26340 18004 26396
rect 18004 26340 18008 26396
rect 17944 26336 18008 26340
rect 18024 26396 18088 26400
rect 18024 26340 18028 26396
rect 18028 26340 18084 26396
rect 18084 26340 18088 26396
rect 18024 26336 18088 26340
rect 4464 25730 4528 25734
rect 4464 25674 4468 25730
rect 4468 25674 4524 25730
rect 4524 25674 4528 25730
rect 4464 25670 4528 25674
rect 4544 25730 4608 25734
rect 4544 25674 4548 25730
rect 4548 25674 4604 25730
rect 4604 25674 4608 25730
rect 4544 25670 4608 25674
rect 4624 25730 4688 25734
rect 4624 25674 4628 25730
rect 4628 25674 4684 25730
rect 4684 25674 4688 25730
rect 4624 25670 4688 25674
rect 4704 25730 4768 25734
rect 4704 25674 4708 25730
rect 4708 25674 4764 25730
rect 4764 25674 4768 25730
rect 4704 25670 4768 25674
rect 9792 25730 9856 25734
rect 9792 25674 9796 25730
rect 9796 25674 9852 25730
rect 9852 25674 9856 25730
rect 9792 25670 9856 25674
rect 9872 25730 9936 25734
rect 9872 25674 9876 25730
rect 9876 25674 9932 25730
rect 9932 25674 9936 25730
rect 9872 25670 9936 25674
rect 9952 25730 10016 25734
rect 9952 25674 9956 25730
rect 9956 25674 10012 25730
rect 10012 25674 10016 25730
rect 9952 25670 10016 25674
rect 10032 25730 10096 25734
rect 10032 25674 10036 25730
rect 10036 25674 10092 25730
rect 10092 25674 10096 25730
rect 10032 25670 10096 25674
rect 15120 25730 15184 25734
rect 15120 25674 15124 25730
rect 15124 25674 15180 25730
rect 15180 25674 15184 25730
rect 15120 25670 15184 25674
rect 15200 25730 15264 25734
rect 15200 25674 15204 25730
rect 15204 25674 15260 25730
rect 15260 25674 15264 25730
rect 15200 25670 15264 25674
rect 15280 25730 15344 25734
rect 15280 25674 15284 25730
rect 15284 25674 15340 25730
rect 15340 25674 15344 25730
rect 15280 25670 15344 25674
rect 15360 25730 15424 25734
rect 15360 25674 15364 25730
rect 15364 25674 15420 25730
rect 15420 25674 15424 25730
rect 15360 25670 15424 25674
rect 20448 25730 20512 25734
rect 20448 25674 20452 25730
rect 20452 25674 20508 25730
rect 20508 25674 20512 25730
rect 20448 25670 20512 25674
rect 20528 25730 20592 25734
rect 20528 25674 20532 25730
rect 20532 25674 20588 25730
rect 20588 25674 20592 25730
rect 20528 25670 20592 25674
rect 20608 25730 20672 25734
rect 20608 25674 20612 25730
rect 20612 25674 20668 25730
rect 20668 25674 20672 25730
rect 20608 25670 20672 25674
rect 20688 25730 20752 25734
rect 20688 25674 20692 25730
rect 20692 25674 20748 25730
rect 20748 25674 20752 25730
rect 20688 25670 20752 25674
rect 7128 25064 7192 25068
rect 7128 25008 7132 25064
rect 7132 25008 7188 25064
rect 7188 25008 7192 25064
rect 7128 25004 7192 25008
rect 7208 25064 7272 25068
rect 7208 25008 7212 25064
rect 7212 25008 7268 25064
rect 7268 25008 7272 25064
rect 7208 25004 7272 25008
rect 7288 25064 7352 25068
rect 7288 25008 7292 25064
rect 7292 25008 7348 25064
rect 7348 25008 7352 25064
rect 7288 25004 7352 25008
rect 7368 25064 7432 25068
rect 7368 25008 7372 25064
rect 7372 25008 7428 25064
rect 7428 25008 7432 25064
rect 7368 25004 7432 25008
rect 12456 25064 12520 25068
rect 12456 25008 12460 25064
rect 12460 25008 12516 25064
rect 12516 25008 12520 25064
rect 12456 25004 12520 25008
rect 12536 25064 12600 25068
rect 12536 25008 12540 25064
rect 12540 25008 12596 25064
rect 12596 25008 12600 25064
rect 12536 25004 12600 25008
rect 12616 25064 12680 25068
rect 12616 25008 12620 25064
rect 12620 25008 12676 25064
rect 12676 25008 12680 25064
rect 12616 25004 12680 25008
rect 12696 25064 12760 25068
rect 12696 25008 12700 25064
rect 12700 25008 12756 25064
rect 12756 25008 12760 25064
rect 12696 25004 12760 25008
rect 17784 25064 17848 25068
rect 17784 25008 17788 25064
rect 17788 25008 17844 25064
rect 17844 25008 17848 25064
rect 17784 25004 17848 25008
rect 17864 25064 17928 25068
rect 17864 25008 17868 25064
rect 17868 25008 17924 25064
rect 17924 25008 17928 25064
rect 17864 25004 17928 25008
rect 17944 25064 18008 25068
rect 17944 25008 17948 25064
rect 17948 25008 18004 25064
rect 18004 25008 18008 25064
rect 17944 25004 18008 25008
rect 18024 25064 18088 25068
rect 18024 25008 18028 25064
rect 18028 25008 18084 25064
rect 18084 25008 18088 25064
rect 18024 25004 18088 25008
rect 4464 24398 4528 24402
rect 4464 24342 4468 24398
rect 4468 24342 4524 24398
rect 4524 24342 4528 24398
rect 4464 24338 4528 24342
rect 4544 24398 4608 24402
rect 4544 24342 4548 24398
rect 4548 24342 4604 24398
rect 4604 24342 4608 24398
rect 4544 24338 4608 24342
rect 4624 24398 4688 24402
rect 4624 24342 4628 24398
rect 4628 24342 4684 24398
rect 4684 24342 4688 24398
rect 4624 24338 4688 24342
rect 4704 24398 4768 24402
rect 4704 24342 4708 24398
rect 4708 24342 4764 24398
rect 4764 24342 4768 24398
rect 4704 24338 4768 24342
rect 9792 24398 9856 24402
rect 9792 24342 9796 24398
rect 9796 24342 9852 24398
rect 9852 24342 9856 24398
rect 9792 24338 9856 24342
rect 9872 24398 9936 24402
rect 9872 24342 9876 24398
rect 9876 24342 9932 24398
rect 9932 24342 9936 24398
rect 9872 24338 9936 24342
rect 9952 24398 10016 24402
rect 9952 24342 9956 24398
rect 9956 24342 10012 24398
rect 10012 24342 10016 24398
rect 9952 24338 10016 24342
rect 10032 24398 10096 24402
rect 10032 24342 10036 24398
rect 10036 24342 10092 24398
rect 10092 24342 10096 24398
rect 10032 24338 10096 24342
rect 15120 24398 15184 24402
rect 15120 24342 15124 24398
rect 15124 24342 15180 24398
rect 15180 24342 15184 24398
rect 15120 24338 15184 24342
rect 15200 24398 15264 24402
rect 15200 24342 15204 24398
rect 15204 24342 15260 24398
rect 15260 24342 15264 24398
rect 15200 24338 15264 24342
rect 15280 24398 15344 24402
rect 15280 24342 15284 24398
rect 15284 24342 15340 24398
rect 15340 24342 15344 24398
rect 15280 24338 15344 24342
rect 15360 24398 15424 24402
rect 15360 24342 15364 24398
rect 15364 24342 15420 24398
rect 15420 24342 15424 24398
rect 15360 24338 15424 24342
rect 20448 24398 20512 24402
rect 20448 24342 20452 24398
rect 20452 24342 20508 24398
rect 20508 24342 20512 24398
rect 20448 24338 20512 24342
rect 20528 24398 20592 24402
rect 20528 24342 20532 24398
rect 20532 24342 20588 24398
rect 20588 24342 20592 24398
rect 20528 24338 20592 24342
rect 20608 24398 20672 24402
rect 20608 24342 20612 24398
rect 20612 24342 20668 24398
rect 20668 24342 20672 24398
rect 20608 24338 20672 24342
rect 20688 24398 20752 24402
rect 20688 24342 20692 24398
rect 20692 24342 20748 24398
rect 20748 24342 20752 24398
rect 20688 24338 20752 24342
rect 7128 23732 7192 23736
rect 7128 23676 7132 23732
rect 7132 23676 7188 23732
rect 7188 23676 7192 23732
rect 7128 23672 7192 23676
rect 7208 23732 7272 23736
rect 7208 23676 7212 23732
rect 7212 23676 7268 23732
rect 7268 23676 7272 23732
rect 7208 23672 7272 23676
rect 7288 23732 7352 23736
rect 7288 23676 7292 23732
rect 7292 23676 7348 23732
rect 7348 23676 7352 23732
rect 7288 23672 7352 23676
rect 7368 23732 7432 23736
rect 7368 23676 7372 23732
rect 7372 23676 7428 23732
rect 7428 23676 7432 23732
rect 7368 23672 7432 23676
rect 12456 23732 12520 23736
rect 12456 23676 12460 23732
rect 12460 23676 12516 23732
rect 12516 23676 12520 23732
rect 12456 23672 12520 23676
rect 12536 23732 12600 23736
rect 12536 23676 12540 23732
rect 12540 23676 12596 23732
rect 12596 23676 12600 23732
rect 12536 23672 12600 23676
rect 12616 23732 12680 23736
rect 12616 23676 12620 23732
rect 12620 23676 12676 23732
rect 12676 23676 12680 23732
rect 12616 23672 12680 23676
rect 12696 23732 12760 23736
rect 12696 23676 12700 23732
rect 12700 23676 12756 23732
rect 12756 23676 12760 23732
rect 12696 23672 12760 23676
rect 17784 23732 17848 23736
rect 17784 23676 17788 23732
rect 17788 23676 17844 23732
rect 17844 23676 17848 23732
rect 17784 23672 17848 23676
rect 17864 23732 17928 23736
rect 17864 23676 17868 23732
rect 17868 23676 17924 23732
rect 17924 23676 17928 23732
rect 17864 23672 17928 23676
rect 17944 23732 18008 23736
rect 17944 23676 17948 23732
rect 17948 23676 18004 23732
rect 18004 23676 18008 23732
rect 17944 23672 18008 23676
rect 18024 23732 18088 23736
rect 18024 23676 18028 23732
rect 18028 23676 18084 23732
rect 18084 23676 18088 23732
rect 18024 23672 18088 23676
rect 4464 23066 4528 23070
rect 4464 23010 4468 23066
rect 4468 23010 4524 23066
rect 4524 23010 4528 23066
rect 4464 23006 4528 23010
rect 4544 23066 4608 23070
rect 4544 23010 4548 23066
rect 4548 23010 4604 23066
rect 4604 23010 4608 23066
rect 4544 23006 4608 23010
rect 4624 23066 4688 23070
rect 4624 23010 4628 23066
rect 4628 23010 4684 23066
rect 4684 23010 4688 23066
rect 4624 23006 4688 23010
rect 4704 23066 4768 23070
rect 4704 23010 4708 23066
rect 4708 23010 4764 23066
rect 4764 23010 4768 23066
rect 4704 23006 4768 23010
rect 9792 23066 9856 23070
rect 9792 23010 9796 23066
rect 9796 23010 9852 23066
rect 9852 23010 9856 23066
rect 9792 23006 9856 23010
rect 9872 23066 9936 23070
rect 9872 23010 9876 23066
rect 9876 23010 9932 23066
rect 9932 23010 9936 23066
rect 9872 23006 9936 23010
rect 9952 23066 10016 23070
rect 9952 23010 9956 23066
rect 9956 23010 10012 23066
rect 10012 23010 10016 23066
rect 9952 23006 10016 23010
rect 10032 23066 10096 23070
rect 10032 23010 10036 23066
rect 10036 23010 10092 23066
rect 10092 23010 10096 23066
rect 10032 23006 10096 23010
rect 15120 23066 15184 23070
rect 15120 23010 15124 23066
rect 15124 23010 15180 23066
rect 15180 23010 15184 23066
rect 15120 23006 15184 23010
rect 15200 23066 15264 23070
rect 15200 23010 15204 23066
rect 15204 23010 15260 23066
rect 15260 23010 15264 23066
rect 15200 23006 15264 23010
rect 15280 23066 15344 23070
rect 15280 23010 15284 23066
rect 15284 23010 15340 23066
rect 15340 23010 15344 23066
rect 15280 23006 15344 23010
rect 15360 23066 15424 23070
rect 15360 23010 15364 23066
rect 15364 23010 15420 23066
rect 15420 23010 15424 23066
rect 15360 23006 15424 23010
rect 20448 23066 20512 23070
rect 20448 23010 20452 23066
rect 20452 23010 20508 23066
rect 20508 23010 20512 23066
rect 20448 23006 20512 23010
rect 20528 23066 20592 23070
rect 20528 23010 20532 23066
rect 20532 23010 20588 23066
rect 20588 23010 20592 23066
rect 20528 23006 20592 23010
rect 20608 23066 20672 23070
rect 20608 23010 20612 23066
rect 20612 23010 20668 23066
rect 20668 23010 20672 23066
rect 20608 23006 20672 23010
rect 20688 23066 20752 23070
rect 20688 23010 20692 23066
rect 20692 23010 20748 23066
rect 20748 23010 20752 23066
rect 20688 23006 20752 23010
rect 7128 22400 7192 22404
rect 7128 22344 7132 22400
rect 7132 22344 7188 22400
rect 7188 22344 7192 22400
rect 7128 22340 7192 22344
rect 7208 22400 7272 22404
rect 7208 22344 7212 22400
rect 7212 22344 7268 22400
rect 7268 22344 7272 22400
rect 7208 22340 7272 22344
rect 7288 22400 7352 22404
rect 7288 22344 7292 22400
rect 7292 22344 7348 22400
rect 7348 22344 7352 22400
rect 7288 22340 7352 22344
rect 7368 22400 7432 22404
rect 7368 22344 7372 22400
rect 7372 22344 7428 22400
rect 7428 22344 7432 22400
rect 7368 22340 7432 22344
rect 12456 22400 12520 22404
rect 12456 22344 12460 22400
rect 12460 22344 12516 22400
rect 12516 22344 12520 22400
rect 12456 22340 12520 22344
rect 12536 22400 12600 22404
rect 12536 22344 12540 22400
rect 12540 22344 12596 22400
rect 12596 22344 12600 22400
rect 12536 22340 12600 22344
rect 12616 22400 12680 22404
rect 12616 22344 12620 22400
rect 12620 22344 12676 22400
rect 12676 22344 12680 22400
rect 12616 22340 12680 22344
rect 12696 22400 12760 22404
rect 12696 22344 12700 22400
rect 12700 22344 12756 22400
rect 12756 22344 12760 22400
rect 12696 22340 12760 22344
rect 17784 22400 17848 22404
rect 17784 22344 17788 22400
rect 17788 22344 17844 22400
rect 17844 22344 17848 22400
rect 17784 22340 17848 22344
rect 17864 22400 17928 22404
rect 17864 22344 17868 22400
rect 17868 22344 17924 22400
rect 17924 22344 17928 22400
rect 17864 22340 17928 22344
rect 17944 22400 18008 22404
rect 17944 22344 17948 22400
rect 17948 22344 18004 22400
rect 18004 22344 18008 22400
rect 17944 22340 18008 22344
rect 18024 22400 18088 22404
rect 18024 22344 18028 22400
rect 18028 22344 18084 22400
rect 18084 22344 18088 22400
rect 18024 22340 18088 22344
rect 4464 21734 4528 21738
rect 4464 21678 4468 21734
rect 4468 21678 4524 21734
rect 4524 21678 4528 21734
rect 4464 21674 4528 21678
rect 4544 21734 4608 21738
rect 4544 21678 4548 21734
rect 4548 21678 4604 21734
rect 4604 21678 4608 21734
rect 4544 21674 4608 21678
rect 4624 21734 4688 21738
rect 4624 21678 4628 21734
rect 4628 21678 4684 21734
rect 4684 21678 4688 21734
rect 4624 21674 4688 21678
rect 4704 21734 4768 21738
rect 4704 21678 4708 21734
rect 4708 21678 4764 21734
rect 4764 21678 4768 21734
rect 4704 21674 4768 21678
rect 9792 21734 9856 21738
rect 9792 21678 9796 21734
rect 9796 21678 9852 21734
rect 9852 21678 9856 21734
rect 9792 21674 9856 21678
rect 9872 21734 9936 21738
rect 9872 21678 9876 21734
rect 9876 21678 9932 21734
rect 9932 21678 9936 21734
rect 9872 21674 9936 21678
rect 9952 21734 10016 21738
rect 9952 21678 9956 21734
rect 9956 21678 10012 21734
rect 10012 21678 10016 21734
rect 9952 21674 10016 21678
rect 10032 21734 10096 21738
rect 10032 21678 10036 21734
rect 10036 21678 10092 21734
rect 10092 21678 10096 21734
rect 10032 21674 10096 21678
rect 15120 21734 15184 21738
rect 15120 21678 15124 21734
rect 15124 21678 15180 21734
rect 15180 21678 15184 21734
rect 15120 21674 15184 21678
rect 15200 21734 15264 21738
rect 15200 21678 15204 21734
rect 15204 21678 15260 21734
rect 15260 21678 15264 21734
rect 15200 21674 15264 21678
rect 15280 21734 15344 21738
rect 15280 21678 15284 21734
rect 15284 21678 15340 21734
rect 15340 21678 15344 21734
rect 15280 21674 15344 21678
rect 15360 21734 15424 21738
rect 15360 21678 15364 21734
rect 15364 21678 15420 21734
rect 15420 21678 15424 21734
rect 15360 21674 15424 21678
rect 20448 21734 20512 21738
rect 20448 21678 20452 21734
rect 20452 21678 20508 21734
rect 20508 21678 20512 21734
rect 20448 21674 20512 21678
rect 20528 21734 20592 21738
rect 20528 21678 20532 21734
rect 20532 21678 20588 21734
rect 20588 21678 20592 21734
rect 20528 21674 20592 21678
rect 20608 21734 20672 21738
rect 20608 21678 20612 21734
rect 20612 21678 20668 21734
rect 20668 21678 20672 21734
rect 20608 21674 20672 21678
rect 20688 21734 20752 21738
rect 20688 21678 20692 21734
rect 20692 21678 20748 21734
rect 20748 21678 20752 21734
rect 20688 21674 20752 21678
rect 7128 21068 7192 21072
rect 7128 21012 7132 21068
rect 7132 21012 7188 21068
rect 7188 21012 7192 21068
rect 7128 21008 7192 21012
rect 7208 21068 7272 21072
rect 7208 21012 7212 21068
rect 7212 21012 7268 21068
rect 7268 21012 7272 21068
rect 7208 21008 7272 21012
rect 7288 21068 7352 21072
rect 7288 21012 7292 21068
rect 7292 21012 7348 21068
rect 7348 21012 7352 21068
rect 7288 21008 7352 21012
rect 7368 21068 7432 21072
rect 7368 21012 7372 21068
rect 7372 21012 7428 21068
rect 7428 21012 7432 21068
rect 7368 21008 7432 21012
rect 12456 21068 12520 21072
rect 12456 21012 12460 21068
rect 12460 21012 12516 21068
rect 12516 21012 12520 21068
rect 12456 21008 12520 21012
rect 12536 21068 12600 21072
rect 12536 21012 12540 21068
rect 12540 21012 12596 21068
rect 12596 21012 12600 21068
rect 12536 21008 12600 21012
rect 12616 21068 12680 21072
rect 12616 21012 12620 21068
rect 12620 21012 12676 21068
rect 12676 21012 12680 21068
rect 12616 21008 12680 21012
rect 12696 21068 12760 21072
rect 12696 21012 12700 21068
rect 12700 21012 12756 21068
rect 12756 21012 12760 21068
rect 12696 21008 12760 21012
rect 17784 21068 17848 21072
rect 17784 21012 17788 21068
rect 17788 21012 17844 21068
rect 17844 21012 17848 21068
rect 17784 21008 17848 21012
rect 17864 21068 17928 21072
rect 17864 21012 17868 21068
rect 17868 21012 17924 21068
rect 17924 21012 17928 21068
rect 17864 21008 17928 21012
rect 17944 21068 18008 21072
rect 17944 21012 17948 21068
rect 17948 21012 18004 21068
rect 18004 21012 18008 21068
rect 17944 21008 18008 21012
rect 18024 21068 18088 21072
rect 18024 21012 18028 21068
rect 18028 21012 18084 21068
rect 18084 21012 18088 21068
rect 18024 21008 18088 21012
rect 4464 20402 4528 20406
rect 4464 20346 4468 20402
rect 4468 20346 4524 20402
rect 4524 20346 4528 20402
rect 4464 20342 4528 20346
rect 4544 20402 4608 20406
rect 4544 20346 4548 20402
rect 4548 20346 4604 20402
rect 4604 20346 4608 20402
rect 4544 20342 4608 20346
rect 4624 20402 4688 20406
rect 4624 20346 4628 20402
rect 4628 20346 4684 20402
rect 4684 20346 4688 20402
rect 4624 20342 4688 20346
rect 4704 20402 4768 20406
rect 4704 20346 4708 20402
rect 4708 20346 4764 20402
rect 4764 20346 4768 20402
rect 4704 20342 4768 20346
rect 9792 20402 9856 20406
rect 9792 20346 9796 20402
rect 9796 20346 9852 20402
rect 9852 20346 9856 20402
rect 9792 20342 9856 20346
rect 9872 20402 9936 20406
rect 9872 20346 9876 20402
rect 9876 20346 9932 20402
rect 9932 20346 9936 20402
rect 9872 20342 9936 20346
rect 9952 20402 10016 20406
rect 9952 20346 9956 20402
rect 9956 20346 10012 20402
rect 10012 20346 10016 20402
rect 9952 20342 10016 20346
rect 10032 20402 10096 20406
rect 10032 20346 10036 20402
rect 10036 20346 10092 20402
rect 10092 20346 10096 20402
rect 10032 20342 10096 20346
rect 15120 20402 15184 20406
rect 15120 20346 15124 20402
rect 15124 20346 15180 20402
rect 15180 20346 15184 20402
rect 15120 20342 15184 20346
rect 15200 20402 15264 20406
rect 15200 20346 15204 20402
rect 15204 20346 15260 20402
rect 15260 20346 15264 20402
rect 15200 20342 15264 20346
rect 15280 20402 15344 20406
rect 15280 20346 15284 20402
rect 15284 20346 15340 20402
rect 15340 20346 15344 20402
rect 15280 20342 15344 20346
rect 15360 20402 15424 20406
rect 15360 20346 15364 20402
rect 15364 20346 15420 20402
rect 15420 20346 15424 20402
rect 15360 20342 15424 20346
rect 20448 20402 20512 20406
rect 20448 20346 20452 20402
rect 20452 20346 20508 20402
rect 20508 20346 20512 20402
rect 20448 20342 20512 20346
rect 20528 20402 20592 20406
rect 20528 20346 20532 20402
rect 20532 20346 20588 20402
rect 20588 20346 20592 20402
rect 20528 20342 20592 20346
rect 20608 20402 20672 20406
rect 20608 20346 20612 20402
rect 20612 20346 20668 20402
rect 20668 20346 20672 20402
rect 20608 20342 20672 20346
rect 20688 20402 20752 20406
rect 20688 20346 20692 20402
rect 20692 20346 20748 20402
rect 20748 20346 20752 20402
rect 20688 20342 20752 20346
rect 7128 19736 7192 19740
rect 7128 19680 7132 19736
rect 7132 19680 7188 19736
rect 7188 19680 7192 19736
rect 7128 19676 7192 19680
rect 7208 19736 7272 19740
rect 7208 19680 7212 19736
rect 7212 19680 7268 19736
rect 7268 19680 7272 19736
rect 7208 19676 7272 19680
rect 7288 19736 7352 19740
rect 7288 19680 7292 19736
rect 7292 19680 7348 19736
rect 7348 19680 7352 19736
rect 7288 19676 7352 19680
rect 7368 19736 7432 19740
rect 7368 19680 7372 19736
rect 7372 19680 7428 19736
rect 7428 19680 7432 19736
rect 7368 19676 7432 19680
rect 12456 19736 12520 19740
rect 12456 19680 12460 19736
rect 12460 19680 12516 19736
rect 12516 19680 12520 19736
rect 12456 19676 12520 19680
rect 12536 19736 12600 19740
rect 12536 19680 12540 19736
rect 12540 19680 12596 19736
rect 12596 19680 12600 19736
rect 12536 19676 12600 19680
rect 12616 19736 12680 19740
rect 12616 19680 12620 19736
rect 12620 19680 12676 19736
rect 12676 19680 12680 19736
rect 12616 19676 12680 19680
rect 12696 19736 12760 19740
rect 12696 19680 12700 19736
rect 12700 19680 12756 19736
rect 12756 19680 12760 19736
rect 12696 19676 12760 19680
rect 17784 19736 17848 19740
rect 17784 19680 17788 19736
rect 17788 19680 17844 19736
rect 17844 19680 17848 19736
rect 17784 19676 17848 19680
rect 17864 19736 17928 19740
rect 17864 19680 17868 19736
rect 17868 19680 17924 19736
rect 17924 19680 17928 19736
rect 17864 19676 17928 19680
rect 17944 19736 18008 19740
rect 17944 19680 17948 19736
rect 17948 19680 18004 19736
rect 18004 19680 18008 19736
rect 17944 19676 18008 19680
rect 18024 19736 18088 19740
rect 18024 19680 18028 19736
rect 18028 19680 18084 19736
rect 18084 19680 18088 19736
rect 18024 19676 18088 19680
rect 4464 19070 4528 19074
rect 4464 19014 4468 19070
rect 4468 19014 4524 19070
rect 4524 19014 4528 19070
rect 4464 19010 4528 19014
rect 4544 19070 4608 19074
rect 4544 19014 4548 19070
rect 4548 19014 4604 19070
rect 4604 19014 4608 19070
rect 4544 19010 4608 19014
rect 4624 19070 4688 19074
rect 4624 19014 4628 19070
rect 4628 19014 4684 19070
rect 4684 19014 4688 19070
rect 4624 19010 4688 19014
rect 4704 19070 4768 19074
rect 4704 19014 4708 19070
rect 4708 19014 4764 19070
rect 4764 19014 4768 19070
rect 4704 19010 4768 19014
rect 9792 19070 9856 19074
rect 9792 19014 9796 19070
rect 9796 19014 9852 19070
rect 9852 19014 9856 19070
rect 9792 19010 9856 19014
rect 9872 19070 9936 19074
rect 9872 19014 9876 19070
rect 9876 19014 9932 19070
rect 9932 19014 9936 19070
rect 9872 19010 9936 19014
rect 9952 19070 10016 19074
rect 9952 19014 9956 19070
rect 9956 19014 10012 19070
rect 10012 19014 10016 19070
rect 9952 19010 10016 19014
rect 10032 19070 10096 19074
rect 10032 19014 10036 19070
rect 10036 19014 10092 19070
rect 10092 19014 10096 19070
rect 10032 19010 10096 19014
rect 15120 19070 15184 19074
rect 15120 19014 15124 19070
rect 15124 19014 15180 19070
rect 15180 19014 15184 19070
rect 15120 19010 15184 19014
rect 15200 19070 15264 19074
rect 15200 19014 15204 19070
rect 15204 19014 15260 19070
rect 15260 19014 15264 19070
rect 15200 19010 15264 19014
rect 15280 19070 15344 19074
rect 15280 19014 15284 19070
rect 15284 19014 15340 19070
rect 15340 19014 15344 19070
rect 15280 19010 15344 19014
rect 15360 19070 15424 19074
rect 15360 19014 15364 19070
rect 15364 19014 15420 19070
rect 15420 19014 15424 19070
rect 15360 19010 15424 19014
rect 20448 19070 20512 19074
rect 20448 19014 20452 19070
rect 20452 19014 20508 19070
rect 20508 19014 20512 19070
rect 20448 19010 20512 19014
rect 20528 19070 20592 19074
rect 20528 19014 20532 19070
rect 20532 19014 20588 19070
rect 20588 19014 20592 19070
rect 20528 19010 20592 19014
rect 20608 19070 20672 19074
rect 20608 19014 20612 19070
rect 20612 19014 20668 19070
rect 20668 19014 20672 19070
rect 20608 19010 20672 19014
rect 20688 19070 20752 19074
rect 20688 19014 20692 19070
rect 20692 19014 20748 19070
rect 20748 19014 20752 19070
rect 20688 19010 20752 19014
rect 7128 18404 7192 18408
rect 7128 18348 7132 18404
rect 7132 18348 7188 18404
rect 7188 18348 7192 18404
rect 7128 18344 7192 18348
rect 7208 18404 7272 18408
rect 7208 18348 7212 18404
rect 7212 18348 7268 18404
rect 7268 18348 7272 18404
rect 7208 18344 7272 18348
rect 7288 18404 7352 18408
rect 7288 18348 7292 18404
rect 7292 18348 7348 18404
rect 7348 18348 7352 18404
rect 7288 18344 7352 18348
rect 7368 18404 7432 18408
rect 7368 18348 7372 18404
rect 7372 18348 7428 18404
rect 7428 18348 7432 18404
rect 7368 18344 7432 18348
rect 12456 18404 12520 18408
rect 12456 18348 12460 18404
rect 12460 18348 12516 18404
rect 12516 18348 12520 18404
rect 12456 18344 12520 18348
rect 12536 18404 12600 18408
rect 12536 18348 12540 18404
rect 12540 18348 12596 18404
rect 12596 18348 12600 18404
rect 12536 18344 12600 18348
rect 12616 18404 12680 18408
rect 12616 18348 12620 18404
rect 12620 18348 12676 18404
rect 12676 18348 12680 18404
rect 12616 18344 12680 18348
rect 12696 18404 12760 18408
rect 12696 18348 12700 18404
rect 12700 18348 12756 18404
rect 12756 18348 12760 18404
rect 12696 18344 12760 18348
rect 17784 18404 17848 18408
rect 17784 18348 17788 18404
rect 17788 18348 17844 18404
rect 17844 18348 17848 18404
rect 17784 18344 17848 18348
rect 17864 18404 17928 18408
rect 17864 18348 17868 18404
rect 17868 18348 17924 18404
rect 17924 18348 17928 18404
rect 17864 18344 17928 18348
rect 17944 18404 18008 18408
rect 17944 18348 17948 18404
rect 17948 18348 18004 18404
rect 18004 18348 18008 18404
rect 17944 18344 18008 18348
rect 18024 18404 18088 18408
rect 18024 18348 18028 18404
rect 18028 18348 18084 18404
rect 18084 18348 18088 18404
rect 18024 18344 18088 18348
rect 4464 17738 4528 17742
rect 4464 17682 4468 17738
rect 4468 17682 4524 17738
rect 4524 17682 4528 17738
rect 4464 17678 4528 17682
rect 4544 17738 4608 17742
rect 4544 17682 4548 17738
rect 4548 17682 4604 17738
rect 4604 17682 4608 17738
rect 4544 17678 4608 17682
rect 4624 17738 4688 17742
rect 4624 17682 4628 17738
rect 4628 17682 4684 17738
rect 4684 17682 4688 17738
rect 4624 17678 4688 17682
rect 4704 17738 4768 17742
rect 4704 17682 4708 17738
rect 4708 17682 4764 17738
rect 4764 17682 4768 17738
rect 4704 17678 4768 17682
rect 9792 17738 9856 17742
rect 9792 17682 9796 17738
rect 9796 17682 9852 17738
rect 9852 17682 9856 17738
rect 9792 17678 9856 17682
rect 9872 17738 9936 17742
rect 9872 17682 9876 17738
rect 9876 17682 9932 17738
rect 9932 17682 9936 17738
rect 9872 17678 9936 17682
rect 9952 17738 10016 17742
rect 9952 17682 9956 17738
rect 9956 17682 10012 17738
rect 10012 17682 10016 17738
rect 9952 17678 10016 17682
rect 10032 17738 10096 17742
rect 10032 17682 10036 17738
rect 10036 17682 10092 17738
rect 10092 17682 10096 17738
rect 10032 17678 10096 17682
rect 15120 17738 15184 17742
rect 15120 17682 15124 17738
rect 15124 17682 15180 17738
rect 15180 17682 15184 17738
rect 15120 17678 15184 17682
rect 15200 17738 15264 17742
rect 15200 17682 15204 17738
rect 15204 17682 15260 17738
rect 15260 17682 15264 17738
rect 15200 17678 15264 17682
rect 15280 17738 15344 17742
rect 15280 17682 15284 17738
rect 15284 17682 15340 17738
rect 15340 17682 15344 17738
rect 15280 17678 15344 17682
rect 15360 17738 15424 17742
rect 15360 17682 15364 17738
rect 15364 17682 15420 17738
rect 15420 17682 15424 17738
rect 15360 17678 15424 17682
rect 20448 17738 20512 17742
rect 20448 17682 20452 17738
rect 20452 17682 20508 17738
rect 20508 17682 20512 17738
rect 20448 17678 20512 17682
rect 20528 17738 20592 17742
rect 20528 17682 20532 17738
rect 20532 17682 20588 17738
rect 20588 17682 20592 17738
rect 20528 17678 20592 17682
rect 20608 17738 20672 17742
rect 20608 17682 20612 17738
rect 20612 17682 20668 17738
rect 20668 17682 20672 17738
rect 20608 17678 20672 17682
rect 20688 17738 20752 17742
rect 20688 17682 20692 17738
rect 20692 17682 20748 17738
rect 20748 17682 20752 17738
rect 20688 17678 20752 17682
rect 7128 17072 7192 17076
rect 7128 17016 7132 17072
rect 7132 17016 7188 17072
rect 7188 17016 7192 17072
rect 7128 17012 7192 17016
rect 7208 17072 7272 17076
rect 7208 17016 7212 17072
rect 7212 17016 7268 17072
rect 7268 17016 7272 17072
rect 7208 17012 7272 17016
rect 7288 17072 7352 17076
rect 7288 17016 7292 17072
rect 7292 17016 7348 17072
rect 7348 17016 7352 17072
rect 7288 17012 7352 17016
rect 7368 17072 7432 17076
rect 7368 17016 7372 17072
rect 7372 17016 7428 17072
rect 7428 17016 7432 17072
rect 7368 17012 7432 17016
rect 12456 17072 12520 17076
rect 12456 17016 12460 17072
rect 12460 17016 12516 17072
rect 12516 17016 12520 17072
rect 12456 17012 12520 17016
rect 12536 17072 12600 17076
rect 12536 17016 12540 17072
rect 12540 17016 12596 17072
rect 12596 17016 12600 17072
rect 12536 17012 12600 17016
rect 12616 17072 12680 17076
rect 12616 17016 12620 17072
rect 12620 17016 12676 17072
rect 12676 17016 12680 17072
rect 12616 17012 12680 17016
rect 12696 17072 12760 17076
rect 12696 17016 12700 17072
rect 12700 17016 12756 17072
rect 12756 17016 12760 17072
rect 12696 17012 12760 17016
rect 17784 17072 17848 17076
rect 17784 17016 17788 17072
rect 17788 17016 17844 17072
rect 17844 17016 17848 17072
rect 17784 17012 17848 17016
rect 17864 17072 17928 17076
rect 17864 17016 17868 17072
rect 17868 17016 17924 17072
rect 17924 17016 17928 17072
rect 17864 17012 17928 17016
rect 17944 17072 18008 17076
rect 17944 17016 17948 17072
rect 17948 17016 18004 17072
rect 18004 17016 18008 17072
rect 17944 17012 18008 17016
rect 18024 17072 18088 17076
rect 18024 17016 18028 17072
rect 18028 17016 18084 17072
rect 18084 17016 18088 17072
rect 18024 17012 18088 17016
rect 4464 16406 4528 16410
rect 4464 16350 4468 16406
rect 4468 16350 4524 16406
rect 4524 16350 4528 16406
rect 4464 16346 4528 16350
rect 4544 16406 4608 16410
rect 4544 16350 4548 16406
rect 4548 16350 4604 16406
rect 4604 16350 4608 16406
rect 4544 16346 4608 16350
rect 4624 16406 4688 16410
rect 4624 16350 4628 16406
rect 4628 16350 4684 16406
rect 4684 16350 4688 16406
rect 4624 16346 4688 16350
rect 4704 16406 4768 16410
rect 4704 16350 4708 16406
rect 4708 16350 4764 16406
rect 4764 16350 4768 16406
rect 4704 16346 4768 16350
rect 9792 16406 9856 16410
rect 9792 16350 9796 16406
rect 9796 16350 9852 16406
rect 9852 16350 9856 16406
rect 9792 16346 9856 16350
rect 9872 16406 9936 16410
rect 9872 16350 9876 16406
rect 9876 16350 9932 16406
rect 9932 16350 9936 16406
rect 9872 16346 9936 16350
rect 9952 16406 10016 16410
rect 9952 16350 9956 16406
rect 9956 16350 10012 16406
rect 10012 16350 10016 16406
rect 9952 16346 10016 16350
rect 10032 16406 10096 16410
rect 10032 16350 10036 16406
rect 10036 16350 10092 16406
rect 10092 16350 10096 16406
rect 10032 16346 10096 16350
rect 15120 16406 15184 16410
rect 15120 16350 15124 16406
rect 15124 16350 15180 16406
rect 15180 16350 15184 16406
rect 15120 16346 15184 16350
rect 15200 16406 15264 16410
rect 15200 16350 15204 16406
rect 15204 16350 15260 16406
rect 15260 16350 15264 16406
rect 15200 16346 15264 16350
rect 15280 16406 15344 16410
rect 15280 16350 15284 16406
rect 15284 16350 15340 16406
rect 15340 16350 15344 16406
rect 15280 16346 15344 16350
rect 15360 16406 15424 16410
rect 15360 16350 15364 16406
rect 15364 16350 15420 16406
rect 15420 16350 15424 16406
rect 15360 16346 15424 16350
rect 20448 16406 20512 16410
rect 20448 16350 20452 16406
rect 20452 16350 20508 16406
rect 20508 16350 20512 16406
rect 20448 16346 20512 16350
rect 20528 16406 20592 16410
rect 20528 16350 20532 16406
rect 20532 16350 20588 16406
rect 20588 16350 20592 16406
rect 20528 16346 20592 16350
rect 20608 16406 20672 16410
rect 20608 16350 20612 16406
rect 20612 16350 20668 16406
rect 20668 16350 20672 16406
rect 20608 16346 20672 16350
rect 20688 16406 20752 16410
rect 20688 16350 20692 16406
rect 20692 16350 20748 16406
rect 20748 16350 20752 16406
rect 20688 16346 20752 16350
rect 7128 15740 7192 15744
rect 7128 15684 7132 15740
rect 7132 15684 7188 15740
rect 7188 15684 7192 15740
rect 7128 15680 7192 15684
rect 7208 15740 7272 15744
rect 7208 15684 7212 15740
rect 7212 15684 7268 15740
rect 7268 15684 7272 15740
rect 7208 15680 7272 15684
rect 7288 15740 7352 15744
rect 7288 15684 7292 15740
rect 7292 15684 7348 15740
rect 7348 15684 7352 15740
rect 7288 15680 7352 15684
rect 7368 15740 7432 15744
rect 7368 15684 7372 15740
rect 7372 15684 7428 15740
rect 7428 15684 7432 15740
rect 7368 15680 7432 15684
rect 12456 15740 12520 15744
rect 12456 15684 12460 15740
rect 12460 15684 12516 15740
rect 12516 15684 12520 15740
rect 12456 15680 12520 15684
rect 12536 15740 12600 15744
rect 12536 15684 12540 15740
rect 12540 15684 12596 15740
rect 12596 15684 12600 15740
rect 12536 15680 12600 15684
rect 12616 15740 12680 15744
rect 12616 15684 12620 15740
rect 12620 15684 12676 15740
rect 12676 15684 12680 15740
rect 12616 15680 12680 15684
rect 12696 15740 12760 15744
rect 12696 15684 12700 15740
rect 12700 15684 12756 15740
rect 12756 15684 12760 15740
rect 12696 15680 12760 15684
rect 17784 15740 17848 15744
rect 17784 15684 17788 15740
rect 17788 15684 17844 15740
rect 17844 15684 17848 15740
rect 17784 15680 17848 15684
rect 17864 15740 17928 15744
rect 17864 15684 17868 15740
rect 17868 15684 17924 15740
rect 17924 15684 17928 15740
rect 17864 15680 17928 15684
rect 17944 15740 18008 15744
rect 17944 15684 17948 15740
rect 17948 15684 18004 15740
rect 18004 15684 18008 15740
rect 17944 15680 18008 15684
rect 18024 15740 18088 15744
rect 18024 15684 18028 15740
rect 18028 15684 18084 15740
rect 18084 15684 18088 15740
rect 18024 15680 18088 15684
rect 4464 15074 4528 15078
rect 4464 15018 4468 15074
rect 4468 15018 4524 15074
rect 4524 15018 4528 15074
rect 4464 15014 4528 15018
rect 4544 15074 4608 15078
rect 4544 15018 4548 15074
rect 4548 15018 4604 15074
rect 4604 15018 4608 15074
rect 4544 15014 4608 15018
rect 4624 15074 4688 15078
rect 4624 15018 4628 15074
rect 4628 15018 4684 15074
rect 4684 15018 4688 15074
rect 4624 15014 4688 15018
rect 4704 15074 4768 15078
rect 4704 15018 4708 15074
rect 4708 15018 4764 15074
rect 4764 15018 4768 15074
rect 4704 15014 4768 15018
rect 9792 15074 9856 15078
rect 9792 15018 9796 15074
rect 9796 15018 9852 15074
rect 9852 15018 9856 15074
rect 9792 15014 9856 15018
rect 9872 15074 9936 15078
rect 9872 15018 9876 15074
rect 9876 15018 9932 15074
rect 9932 15018 9936 15074
rect 9872 15014 9936 15018
rect 9952 15074 10016 15078
rect 9952 15018 9956 15074
rect 9956 15018 10012 15074
rect 10012 15018 10016 15074
rect 9952 15014 10016 15018
rect 10032 15074 10096 15078
rect 10032 15018 10036 15074
rect 10036 15018 10092 15074
rect 10092 15018 10096 15074
rect 10032 15014 10096 15018
rect 15120 15074 15184 15078
rect 15120 15018 15124 15074
rect 15124 15018 15180 15074
rect 15180 15018 15184 15074
rect 15120 15014 15184 15018
rect 15200 15074 15264 15078
rect 15200 15018 15204 15074
rect 15204 15018 15260 15074
rect 15260 15018 15264 15074
rect 15200 15014 15264 15018
rect 15280 15074 15344 15078
rect 15280 15018 15284 15074
rect 15284 15018 15340 15074
rect 15340 15018 15344 15074
rect 15280 15014 15344 15018
rect 15360 15074 15424 15078
rect 15360 15018 15364 15074
rect 15364 15018 15420 15074
rect 15420 15018 15424 15074
rect 15360 15014 15424 15018
rect 20448 15074 20512 15078
rect 20448 15018 20452 15074
rect 20452 15018 20508 15074
rect 20508 15018 20512 15074
rect 20448 15014 20512 15018
rect 20528 15074 20592 15078
rect 20528 15018 20532 15074
rect 20532 15018 20588 15074
rect 20588 15018 20592 15074
rect 20528 15014 20592 15018
rect 20608 15074 20672 15078
rect 20608 15018 20612 15074
rect 20612 15018 20668 15074
rect 20668 15018 20672 15074
rect 20608 15014 20672 15018
rect 20688 15074 20752 15078
rect 20688 15018 20692 15074
rect 20692 15018 20748 15074
rect 20748 15018 20752 15074
rect 20688 15014 20752 15018
rect 7128 14408 7192 14412
rect 7128 14352 7132 14408
rect 7132 14352 7188 14408
rect 7188 14352 7192 14408
rect 7128 14348 7192 14352
rect 7208 14408 7272 14412
rect 7208 14352 7212 14408
rect 7212 14352 7268 14408
rect 7268 14352 7272 14408
rect 7208 14348 7272 14352
rect 7288 14408 7352 14412
rect 7288 14352 7292 14408
rect 7292 14352 7348 14408
rect 7348 14352 7352 14408
rect 7288 14348 7352 14352
rect 7368 14408 7432 14412
rect 7368 14352 7372 14408
rect 7372 14352 7428 14408
rect 7428 14352 7432 14408
rect 7368 14348 7432 14352
rect 12456 14408 12520 14412
rect 12456 14352 12460 14408
rect 12460 14352 12516 14408
rect 12516 14352 12520 14408
rect 12456 14348 12520 14352
rect 12536 14408 12600 14412
rect 12536 14352 12540 14408
rect 12540 14352 12596 14408
rect 12596 14352 12600 14408
rect 12536 14348 12600 14352
rect 12616 14408 12680 14412
rect 12616 14352 12620 14408
rect 12620 14352 12676 14408
rect 12676 14352 12680 14408
rect 12616 14348 12680 14352
rect 12696 14408 12760 14412
rect 12696 14352 12700 14408
rect 12700 14352 12756 14408
rect 12756 14352 12760 14408
rect 12696 14348 12760 14352
rect 17784 14408 17848 14412
rect 17784 14352 17788 14408
rect 17788 14352 17844 14408
rect 17844 14352 17848 14408
rect 17784 14348 17848 14352
rect 17864 14408 17928 14412
rect 17864 14352 17868 14408
rect 17868 14352 17924 14408
rect 17924 14352 17928 14408
rect 17864 14348 17928 14352
rect 17944 14408 18008 14412
rect 17944 14352 17948 14408
rect 17948 14352 18004 14408
rect 18004 14352 18008 14408
rect 17944 14348 18008 14352
rect 18024 14408 18088 14412
rect 18024 14352 18028 14408
rect 18028 14352 18084 14408
rect 18084 14352 18088 14408
rect 18024 14348 18088 14352
rect 4464 13742 4528 13746
rect 4464 13686 4468 13742
rect 4468 13686 4524 13742
rect 4524 13686 4528 13742
rect 4464 13682 4528 13686
rect 4544 13742 4608 13746
rect 4544 13686 4548 13742
rect 4548 13686 4604 13742
rect 4604 13686 4608 13742
rect 4544 13682 4608 13686
rect 4624 13742 4688 13746
rect 4624 13686 4628 13742
rect 4628 13686 4684 13742
rect 4684 13686 4688 13742
rect 4624 13682 4688 13686
rect 4704 13742 4768 13746
rect 4704 13686 4708 13742
rect 4708 13686 4764 13742
rect 4764 13686 4768 13742
rect 4704 13682 4768 13686
rect 9792 13742 9856 13746
rect 9792 13686 9796 13742
rect 9796 13686 9852 13742
rect 9852 13686 9856 13742
rect 9792 13682 9856 13686
rect 9872 13742 9936 13746
rect 9872 13686 9876 13742
rect 9876 13686 9932 13742
rect 9932 13686 9936 13742
rect 9872 13682 9936 13686
rect 9952 13742 10016 13746
rect 9952 13686 9956 13742
rect 9956 13686 10012 13742
rect 10012 13686 10016 13742
rect 9952 13682 10016 13686
rect 10032 13742 10096 13746
rect 10032 13686 10036 13742
rect 10036 13686 10092 13742
rect 10092 13686 10096 13742
rect 10032 13682 10096 13686
rect 15120 13742 15184 13746
rect 15120 13686 15124 13742
rect 15124 13686 15180 13742
rect 15180 13686 15184 13742
rect 15120 13682 15184 13686
rect 15200 13742 15264 13746
rect 15200 13686 15204 13742
rect 15204 13686 15260 13742
rect 15260 13686 15264 13742
rect 15200 13682 15264 13686
rect 15280 13742 15344 13746
rect 15280 13686 15284 13742
rect 15284 13686 15340 13742
rect 15340 13686 15344 13742
rect 15280 13682 15344 13686
rect 15360 13742 15424 13746
rect 15360 13686 15364 13742
rect 15364 13686 15420 13742
rect 15420 13686 15424 13742
rect 15360 13682 15424 13686
rect 20448 13742 20512 13746
rect 20448 13686 20452 13742
rect 20452 13686 20508 13742
rect 20508 13686 20512 13742
rect 20448 13682 20512 13686
rect 20528 13742 20592 13746
rect 20528 13686 20532 13742
rect 20532 13686 20588 13742
rect 20588 13686 20592 13742
rect 20528 13682 20592 13686
rect 20608 13742 20672 13746
rect 20608 13686 20612 13742
rect 20612 13686 20668 13742
rect 20668 13686 20672 13742
rect 20608 13682 20672 13686
rect 20688 13742 20752 13746
rect 20688 13686 20692 13742
rect 20692 13686 20748 13742
rect 20748 13686 20752 13742
rect 20688 13682 20752 13686
rect 7128 13076 7192 13080
rect 7128 13020 7132 13076
rect 7132 13020 7188 13076
rect 7188 13020 7192 13076
rect 7128 13016 7192 13020
rect 7208 13076 7272 13080
rect 7208 13020 7212 13076
rect 7212 13020 7268 13076
rect 7268 13020 7272 13076
rect 7208 13016 7272 13020
rect 7288 13076 7352 13080
rect 7288 13020 7292 13076
rect 7292 13020 7348 13076
rect 7348 13020 7352 13076
rect 7288 13016 7352 13020
rect 7368 13076 7432 13080
rect 7368 13020 7372 13076
rect 7372 13020 7428 13076
rect 7428 13020 7432 13076
rect 7368 13016 7432 13020
rect 12456 13076 12520 13080
rect 12456 13020 12460 13076
rect 12460 13020 12516 13076
rect 12516 13020 12520 13076
rect 12456 13016 12520 13020
rect 12536 13076 12600 13080
rect 12536 13020 12540 13076
rect 12540 13020 12596 13076
rect 12596 13020 12600 13076
rect 12536 13016 12600 13020
rect 12616 13076 12680 13080
rect 12616 13020 12620 13076
rect 12620 13020 12676 13076
rect 12676 13020 12680 13076
rect 12616 13016 12680 13020
rect 12696 13076 12760 13080
rect 12696 13020 12700 13076
rect 12700 13020 12756 13076
rect 12756 13020 12760 13076
rect 12696 13016 12760 13020
rect 17784 13076 17848 13080
rect 17784 13020 17788 13076
rect 17788 13020 17844 13076
rect 17844 13020 17848 13076
rect 17784 13016 17848 13020
rect 17864 13076 17928 13080
rect 17864 13020 17868 13076
rect 17868 13020 17924 13076
rect 17924 13020 17928 13076
rect 17864 13016 17928 13020
rect 17944 13076 18008 13080
rect 17944 13020 17948 13076
rect 17948 13020 18004 13076
rect 18004 13020 18008 13076
rect 17944 13016 18008 13020
rect 18024 13076 18088 13080
rect 18024 13020 18028 13076
rect 18028 13020 18084 13076
rect 18084 13020 18088 13076
rect 18024 13016 18088 13020
rect 4464 12410 4528 12414
rect 4464 12354 4468 12410
rect 4468 12354 4524 12410
rect 4524 12354 4528 12410
rect 4464 12350 4528 12354
rect 4544 12410 4608 12414
rect 4544 12354 4548 12410
rect 4548 12354 4604 12410
rect 4604 12354 4608 12410
rect 4544 12350 4608 12354
rect 4624 12410 4688 12414
rect 4624 12354 4628 12410
rect 4628 12354 4684 12410
rect 4684 12354 4688 12410
rect 4624 12350 4688 12354
rect 4704 12410 4768 12414
rect 4704 12354 4708 12410
rect 4708 12354 4764 12410
rect 4764 12354 4768 12410
rect 4704 12350 4768 12354
rect 9792 12410 9856 12414
rect 9792 12354 9796 12410
rect 9796 12354 9852 12410
rect 9852 12354 9856 12410
rect 9792 12350 9856 12354
rect 9872 12410 9936 12414
rect 9872 12354 9876 12410
rect 9876 12354 9932 12410
rect 9932 12354 9936 12410
rect 9872 12350 9936 12354
rect 9952 12410 10016 12414
rect 9952 12354 9956 12410
rect 9956 12354 10012 12410
rect 10012 12354 10016 12410
rect 9952 12350 10016 12354
rect 10032 12410 10096 12414
rect 10032 12354 10036 12410
rect 10036 12354 10092 12410
rect 10092 12354 10096 12410
rect 10032 12350 10096 12354
rect 15120 12410 15184 12414
rect 15120 12354 15124 12410
rect 15124 12354 15180 12410
rect 15180 12354 15184 12410
rect 15120 12350 15184 12354
rect 15200 12410 15264 12414
rect 15200 12354 15204 12410
rect 15204 12354 15260 12410
rect 15260 12354 15264 12410
rect 15200 12350 15264 12354
rect 15280 12410 15344 12414
rect 15280 12354 15284 12410
rect 15284 12354 15340 12410
rect 15340 12354 15344 12410
rect 15280 12350 15344 12354
rect 15360 12410 15424 12414
rect 15360 12354 15364 12410
rect 15364 12354 15420 12410
rect 15420 12354 15424 12410
rect 15360 12350 15424 12354
rect 20448 12410 20512 12414
rect 20448 12354 20452 12410
rect 20452 12354 20508 12410
rect 20508 12354 20512 12410
rect 20448 12350 20512 12354
rect 20528 12410 20592 12414
rect 20528 12354 20532 12410
rect 20532 12354 20588 12410
rect 20588 12354 20592 12410
rect 20528 12350 20592 12354
rect 20608 12410 20672 12414
rect 20608 12354 20612 12410
rect 20612 12354 20668 12410
rect 20668 12354 20672 12410
rect 20608 12350 20672 12354
rect 20688 12410 20752 12414
rect 20688 12354 20692 12410
rect 20692 12354 20748 12410
rect 20748 12354 20752 12410
rect 20688 12350 20752 12354
rect 7128 11744 7192 11748
rect 7128 11688 7132 11744
rect 7132 11688 7188 11744
rect 7188 11688 7192 11744
rect 7128 11684 7192 11688
rect 7208 11744 7272 11748
rect 7208 11688 7212 11744
rect 7212 11688 7268 11744
rect 7268 11688 7272 11744
rect 7208 11684 7272 11688
rect 7288 11744 7352 11748
rect 7288 11688 7292 11744
rect 7292 11688 7348 11744
rect 7348 11688 7352 11744
rect 7288 11684 7352 11688
rect 7368 11744 7432 11748
rect 7368 11688 7372 11744
rect 7372 11688 7428 11744
rect 7428 11688 7432 11744
rect 7368 11684 7432 11688
rect 12456 11744 12520 11748
rect 12456 11688 12460 11744
rect 12460 11688 12516 11744
rect 12516 11688 12520 11744
rect 12456 11684 12520 11688
rect 12536 11744 12600 11748
rect 12536 11688 12540 11744
rect 12540 11688 12596 11744
rect 12596 11688 12600 11744
rect 12536 11684 12600 11688
rect 12616 11744 12680 11748
rect 12616 11688 12620 11744
rect 12620 11688 12676 11744
rect 12676 11688 12680 11744
rect 12616 11684 12680 11688
rect 12696 11744 12760 11748
rect 12696 11688 12700 11744
rect 12700 11688 12756 11744
rect 12756 11688 12760 11744
rect 12696 11684 12760 11688
rect 17784 11744 17848 11748
rect 17784 11688 17788 11744
rect 17788 11688 17844 11744
rect 17844 11688 17848 11744
rect 17784 11684 17848 11688
rect 17864 11744 17928 11748
rect 17864 11688 17868 11744
rect 17868 11688 17924 11744
rect 17924 11688 17928 11744
rect 17864 11684 17928 11688
rect 17944 11744 18008 11748
rect 17944 11688 17948 11744
rect 17948 11688 18004 11744
rect 18004 11688 18008 11744
rect 17944 11684 18008 11688
rect 18024 11744 18088 11748
rect 18024 11688 18028 11744
rect 18028 11688 18084 11744
rect 18084 11688 18088 11744
rect 18024 11684 18088 11688
rect 4464 11078 4528 11082
rect 4464 11022 4468 11078
rect 4468 11022 4524 11078
rect 4524 11022 4528 11078
rect 4464 11018 4528 11022
rect 4544 11078 4608 11082
rect 4544 11022 4548 11078
rect 4548 11022 4604 11078
rect 4604 11022 4608 11078
rect 4544 11018 4608 11022
rect 4624 11078 4688 11082
rect 4624 11022 4628 11078
rect 4628 11022 4684 11078
rect 4684 11022 4688 11078
rect 4624 11018 4688 11022
rect 4704 11078 4768 11082
rect 4704 11022 4708 11078
rect 4708 11022 4764 11078
rect 4764 11022 4768 11078
rect 4704 11018 4768 11022
rect 9792 11078 9856 11082
rect 9792 11022 9796 11078
rect 9796 11022 9852 11078
rect 9852 11022 9856 11078
rect 9792 11018 9856 11022
rect 9872 11078 9936 11082
rect 9872 11022 9876 11078
rect 9876 11022 9932 11078
rect 9932 11022 9936 11078
rect 9872 11018 9936 11022
rect 9952 11078 10016 11082
rect 9952 11022 9956 11078
rect 9956 11022 10012 11078
rect 10012 11022 10016 11078
rect 9952 11018 10016 11022
rect 10032 11078 10096 11082
rect 10032 11022 10036 11078
rect 10036 11022 10092 11078
rect 10092 11022 10096 11078
rect 10032 11018 10096 11022
rect 15120 11078 15184 11082
rect 15120 11022 15124 11078
rect 15124 11022 15180 11078
rect 15180 11022 15184 11078
rect 15120 11018 15184 11022
rect 15200 11078 15264 11082
rect 15200 11022 15204 11078
rect 15204 11022 15260 11078
rect 15260 11022 15264 11078
rect 15200 11018 15264 11022
rect 15280 11078 15344 11082
rect 15280 11022 15284 11078
rect 15284 11022 15340 11078
rect 15340 11022 15344 11078
rect 15280 11018 15344 11022
rect 15360 11078 15424 11082
rect 15360 11022 15364 11078
rect 15364 11022 15420 11078
rect 15420 11022 15424 11078
rect 15360 11018 15424 11022
rect 20448 11078 20512 11082
rect 20448 11022 20452 11078
rect 20452 11022 20508 11078
rect 20508 11022 20512 11078
rect 20448 11018 20512 11022
rect 20528 11078 20592 11082
rect 20528 11022 20532 11078
rect 20532 11022 20588 11078
rect 20588 11022 20592 11078
rect 20528 11018 20592 11022
rect 20608 11078 20672 11082
rect 20608 11022 20612 11078
rect 20612 11022 20668 11078
rect 20668 11022 20672 11078
rect 20608 11018 20672 11022
rect 20688 11078 20752 11082
rect 20688 11022 20692 11078
rect 20692 11022 20748 11078
rect 20748 11022 20752 11078
rect 20688 11018 20752 11022
rect 7128 10412 7192 10416
rect 7128 10356 7132 10412
rect 7132 10356 7188 10412
rect 7188 10356 7192 10412
rect 7128 10352 7192 10356
rect 7208 10412 7272 10416
rect 7208 10356 7212 10412
rect 7212 10356 7268 10412
rect 7268 10356 7272 10412
rect 7208 10352 7272 10356
rect 7288 10412 7352 10416
rect 7288 10356 7292 10412
rect 7292 10356 7348 10412
rect 7348 10356 7352 10412
rect 7288 10352 7352 10356
rect 7368 10412 7432 10416
rect 7368 10356 7372 10412
rect 7372 10356 7428 10412
rect 7428 10356 7432 10412
rect 7368 10352 7432 10356
rect 12456 10412 12520 10416
rect 12456 10356 12460 10412
rect 12460 10356 12516 10412
rect 12516 10356 12520 10412
rect 12456 10352 12520 10356
rect 12536 10412 12600 10416
rect 12536 10356 12540 10412
rect 12540 10356 12596 10412
rect 12596 10356 12600 10412
rect 12536 10352 12600 10356
rect 12616 10412 12680 10416
rect 12616 10356 12620 10412
rect 12620 10356 12676 10412
rect 12676 10356 12680 10412
rect 12616 10352 12680 10356
rect 12696 10412 12760 10416
rect 12696 10356 12700 10412
rect 12700 10356 12756 10412
rect 12756 10356 12760 10412
rect 12696 10352 12760 10356
rect 17784 10412 17848 10416
rect 17784 10356 17788 10412
rect 17788 10356 17844 10412
rect 17844 10356 17848 10412
rect 17784 10352 17848 10356
rect 17864 10412 17928 10416
rect 17864 10356 17868 10412
rect 17868 10356 17924 10412
rect 17924 10356 17928 10412
rect 17864 10352 17928 10356
rect 17944 10412 18008 10416
rect 17944 10356 17948 10412
rect 17948 10356 18004 10412
rect 18004 10356 18008 10412
rect 17944 10352 18008 10356
rect 18024 10412 18088 10416
rect 18024 10356 18028 10412
rect 18028 10356 18084 10412
rect 18084 10356 18088 10412
rect 18024 10352 18088 10356
rect 4464 9746 4528 9750
rect 4464 9690 4468 9746
rect 4468 9690 4524 9746
rect 4524 9690 4528 9746
rect 4464 9686 4528 9690
rect 4544 9746 4608 9750
rect 4544 9690 4548 9746
rect 4548 9690 4604 9746
rect 4604 9690 4608 9746
rect 4544 9686 4608 9690
rect 4624 9746 4688 9750
rect 4624 9690 4628 9746
rect 4628 9690 4684 9746
rect 4684 9690 4688 9746
rect 4624 9686 4688 9690
rect 4704 9746 4768 9750
rect 4704 9690 4708 9746
rect 4708 9690 4764 9746
rect 4764 9690 4768 9746
rect 4704 9686 4768 9690
rect 9792 9746 9856 9750
rect 9792 9690 9796 9746
rect 9796 9690 9852 9746
rect 9852 9690 9856 9746
rect 9792 9686 9856 9690
rect 9872 9746 9936 9750
rect 9872 9690 9876 9746
rect 9876 9690 9932 9746
rect 9932 9690 9936 9746
rect 9872 9686 9936 9690
rect 9952 9746 10016 9750
rect 9952 9690 9956 9746
rect 9956 9690 10012 9746
rect 10012 9690 10016 9746
rect 9952 9686 10016 9690
rect 10032 9746 10096 9750
rect 10032 9690 10036 9746
rect 10036 9690 10092 9746
rect 10092 9690 10096 9746
rect 10032 9686 10096 9690
rect 15120 9746 15184 9750
rect 15120 9690 15124 9746
rect 15124 9690 15180 9746
rect 15180 9690 15184 9746
rect 15120 9686 15184 9690
rect 15200 9746 15264 9750
rect 15200 9690 15204 9746
rect 15204 9690 15260 9746
rect 15260 9690 15264 9746
rect 15200 9686 15264 9690
rect 15280 9746 15344 9750
rect 15280 9690 15284 9746
rect 15284 9690 15340 9746
rect 15340 9690 15344 9746
rect 15280 9686 15344 9690
rect 15360 9746 15424 9750
rect 15360 9690 15364 9746
rect 15364 9690 15420 9746
rect 15420 9690 15424 9746
rect 15360 9686 15424 9690
rect 20448 9746 20512 9750
rect 20448 9690 20452 9746
rect 20452 9690 20508 9746
rect 20508 9690 20512 9746
rect 20448 9686 20512 9690
rect 20528 9746 20592 9750
rect 20528 9690 20532 9746
rect 20532 9690 20588 9746
rect 20588 9690 20592 9746
rect 20528 9686 20592 9690
rect 20608 9746 20672 9750
rect 20608 9690 20612 9746
rect 20612 9690 20668 9746
rect 20668 9690 20672 9746
rect 20608 9686 20672 9690
rect 20688 9746 20752 9750
rect 20688 9690 20692 9746
rect 20692 9690 20748 9746
rect 20748 9690 20752 9746
rect 20688 9686 20752 9690
rect 7128 9080 7192 9084
rect 7128 9024 7132 9080
rect 7132 9024 7188 9080
rect 7188 9024 7192 9080
rect 7128 9020 7192 9024
rect 7208 9080 7272 9084
rect 7208 9024 7212 9080
rect 7212 9024 7268 9080
rect 7268 9024 7272 9080
rect 7208 9020 7272 9024
rect 7288 9080 7352 9084
rect 7288 9024 7292 9080
rect 7292 9024 7348 9080
rect 7348 9024 7352 9080
rect 7288 9020 7352 9024
rect 7368 9080 7432 9084
rect 7368 9024 7372 9080
rect 7372 9024 7428 9080
rect 7428 9024 7432 9080
rect 7368 9020 7432 9024
rect 12456 9080 12520 9084
rect 12456 9024 12460 9080
rect 12460 9024 12516 9080
rect 12516 9024 12520 9080
rect 12456 9020 12520 9024
rect 12536 9080 12600 9084
rect 12536 9024 12540 9080
rect 12540 9024 12596 9080
rect 12596 9024 12600 9080
rect 12536 9020 12600 9024
rect 12616 9080 12680 9084
rect 12616 9024 12620 9080
rect 12620 9024 12676 9080
rect 12676 9024 12680 9080
rect 12616 9020 12680 9024
rect 12696 9080 12760 9084
rect 12696 9024 12700 9080
rect 12700 9024 12756 9080
rect 12756 9024 12760 9080
rect 12696 9020 12760 9024
rect 17784 9080 17848 9084
rect 17784 9024 17788 9080
rect 17788 9024 17844 9080
rect 17844 9024 17848 9080
rect 17784 9020 17848 9024
rect 17864 9080 17928 9084
rect 17864 9024 17868 9080
rect 17868 9024 17924 9080
rect 17924 9024 17928 9080
rect 17864 9020 17928 9024
rect 17944 9080 18008 9084
rect 17944 9024 17948 9080
rect 17948 9024 18004 9080
rect 18004 9024 18008 9080
rect 17944 9020 18008 9024
rect 18024 9080 18088 9084
rect 18024 9024 18028 9080
rect 18028 9024 18084 9080
rect 18084 9024 18088 9080
rect 18024 9020 18088 9024
rect 4464 8414 4528 8418
rect 4464 8358 4468 8414
rect 4468 8358 4524 8414
rect 4524 8358 4528 8414
rect 4464 8354 4528 8358
rect 4544 8414 4608 8418
rect 4544 8358 4548 8414
rect 4548 8358 4604 8414
rect 4604 8358 4608 8414
rect 4544 8354 4608 8358
rect 4624 8414 4688 8418
rect 4624 8358 4628 8414
rect 4628 8358 4684 8414
rect 4684 8358 4688 8414
rect 4624 8354 4688 8358
rect 4704 8414 4768 8418
rect 4704 8358 4708 8414
rect 4708 8358 4764 8414
rect 4764 8358 4768 8414
rect 4704 8354 4768 8358
rect 9792 8414 9856 8418
rect 9792 8358 9796 8414
rect 9796 8358 9852 8414
rect 9852 8358 9856 8414
rect 9792 8354 9856 8358
rect 9872 8414 9936 8418
rect 9872 8358 9876 8414
rect 9876 8358 9932 8414
rect 9932 8358 9936 8414
rect 9872 8354 9936 8358
rect 9952 8414 10016 8418
rect 9952 8358 9956 8414
rect 9956 8358 10012 8414
rect 10012 8358 10016 8414
rect 9952 8354 10016 8358
rect 10032 8414 10096 8418
rect 10032 8358 10036 8414
rect 10036 8358 10092 8414
rect 10092 8358 10096 8414
rect 10032 8354 10096 8358
rect 15120 8414 15184 8418
rect 15120 8358 15124 8414
rect 15124 8358 15180 8414
rect 15180 8358 15184 8414
rect 15120 8354 15184 8358
rect 15200 8414 15264 8418
rect 15200 8358 15204 8414
rect 15204 8358 15260 8414
rect 15260 8358 15264 8414
rect 15200 8354 15264 8358
rect 15280 8414 15344 8418
rect 15280 8358 15284 8414
rect 15284 8358 15340 8414
rect 15340 8358 15344 8414
rect 15280 8354 15344 8358
rect 15360 8414 15424 8418
rect 15360 8358 15364 8414
rect 15364 8358 15420 8414
rect 15420 8358 15424 8414
rect 15360 8354 15424 8358
rect 20448 8414 20512 8418
rect 20448 8358 20452 8414
rect 20452 8358 20508 8414
rect 20508 8358 20512 8414
rect 20448 8354 20512 8358
rect 20528 8414 20592 8418
rect 20528 8358 20532 8414
rect 20532 8358 20588 8414
rect 20588 8358 20592 8414
rect 20528 8354 20592 8358
rect 20608 8414 20672 8418
rect 20608 8358 20612 8414
rect 20612 8358 20668 8414
rect 20668 8358 20672 8414
rect 20608 8354 20672 8358
rect 20688 8414 20752 8418
rect 20688 8358 20692 8414
rect 20692 8358 20748 8414
rect 20748 8358 20752 8414
rect 20688 8354 20752 8358
rect 7128 7748 7192 7752
rect 7128 7692 7132 7748
rect 7132 7692 7188 7748
rect 7188 7692 7192 7748
rect 7128 7688 7192 7692
rect 7208 7748 7272 7752
rect 7208 7692 7212 7748
rect 7212 7692 7268 7748
rect 7268 7692 7272 7748
rect 7208 7688 7272 7692
rect 7288 7748 7352 7752
rect 7288 7692 7292 7748
rect 7292 7692 7348 7748
rect 7348 7692 7352 7748
rect 7288 7688 7352 7692
rect 7368 7748 7432 7752
rect 7368 7692 7372 7748
rect 7372 7692 7428 7748
rect 7428 7692 7432 7748
rect 7368 7688 7432 7692
rect 12456 7748 12520 7752
rect 12456 7692 12460 7748
rect 12460 7692 12516 7748
rect 12516 7692 12520 7748
rect 12456 7688 12520 7692
rect 12536 7748 12600 7752
rect 12536 7692 12540 7748
rect 12540 7692 12596 7748
rect 12596 7692 12600 7748
rect 12536 7688 12600 7692
rect 12616 7748 12680 7752
rect 12616 7692 12620 7748
rect 12620 7692 12676 7748
rect 12676 7692 12680 7748
rect 12616 7688 12680 7692
rect 12696 7748 12760 7752
rect 12696 7692 12700 7748
rect 12700 7692 12756 7748
rect 12756 7692 12760 7748
rect 12696 7688 12760 7692
rect 17784 7748 17848 7752
rect 17784 7692 17788 7748
rect 17788 7692 17844 7748
rect 17844 7692 17848 7748
rect 17784 7688 17848 7692
rect 17864 7748 17928 7752
rect 17864 7692 17868 7748
rect 17868 7692 17924 7748
rect 17924 7692 17928 7748
rect 17864 7688 17928 7692
rect 17944 7748 18008 7752
rect 17944 7692 17948 7748
rect 17948 7692 18004 7748
rect 18004 7692 18008 7748
rect 17944 7688 18008 7692
rect 18024 7748 18088 7752
rect 18024 7692 18028 7748
rect 18028 7692 18084 7748
rect 18084 7692 18088 7748
rect 18024 7688 18088 7692
rect 4464 7082 4528 7086
rect 4464 7026 4468 7082
rect 4468 7026 4524 7082
rect 4524 7026 4528 7082
rect 4464 7022 4528 7026
rect 4544 7082 4608 7086
rect 4544 7026 4548 7082
rect 4548 7026 4604 7082
rect 4604 7026 4608 7082
rect 4544 7022 4608 7026
rect 4624 7082 4688 7086
rect 4624 7026 4628 7082
rect 4628 7026 4684 7082
rect 4684 7026 4688 7082
rect 4624 7022 4688 7026
rect 4704 7082 4768 7086
rect 4704 7026 4708 7082
rect 4708 7026 4764 7082
rect 4764 7026 4768 7082
rect 4704 7022 4768 7026
rect 9792 7082 9856 7086
rect 9792 7026 9796 7082
rect 9796 7026 9852 7082
rect 9852 7026 9856 7082
rect 9792 7022 9856 7026
rect 9872 7082 9936 7086
rect 9872 7026 9876 7082
rect 9876 7026 9932 7082
rect 9932 7026 9936 7082
rect 9872 7022 9936 7026
rect 9952 7082 10016 7086
rect 9952 7026 9956 7082
rect 9956 7026 10012 7082
rect 10012 7026 10016 7082
rect 9952 7022 10016 7026
rect 10032 7082 10096 7086
rect 10032 7026 10036 7082
rect 10036 7026 10092 7082
rect 10092 7026 10096 7082
rect 10032 7022 10096 7026
rect 15120 7082 15184 7086
rect 15120 7026 15124 7082
rect 15124 7026 15180 7082
rect 15180 7026 15184 7082
rect 15120 7022 15184 7026
rect 15200 7082 15264 7086
rect 15200 7026 15204 7082
rect 15204 7026 15260 7082
rect 15260 7026 15264 7082
rect 15200 7022 15264 7026
rect 15280 7082 15344 7086
rect 15280 7026 15284 7082
rect 15284 7026 15340 7082
rect 15340 7026 15344 7082
rect 15280 7022 15344 7026
rect 15360 7082 15424 7086
rect 15360 7026 15364 7082
rect 15364 7026 15420 7082
rect 15420 7026 15424 7082
rect 15360 7022 15424 7026
rect 20448 7082 20512 7086
rect 20448 7026 20452 7082
rect 20452 7026 20508 7082
rect 20508 7026 20512 7082
rect 20448 7022 20512 7026
rect 20528 7082 20592 7086
rect 20528 7026 20532 7082
rect 20532 7026 20588 7082
rect 20588 7026 20592 7082
rect 20528 7022 20592 7026
rect 20608 7082 20672 7086
rect 20608 7026 20612 7082
rect 20612 7026 20668 7082
rect 20668 7026 20672 7082
rect 20608 7022 20672 7026
rect 20688 7082 20752 7086
rect 20688 7026 20692 7082
rect 20692 7026 20748 7082
rect 20748 7026 20752 7082
rect 20688 7022 20752 7026
rect 7128 6416 7192 6420
rect 7128 6360 7132 6416
rect 7132 6360 7188 6416
rect 7188 6360 7192 6416
rect 7128 6356 7192 6360
rect 7208 6416 7272 6420
rect 7208 6360 7212 6416
rect 7212 6360 7268 6416
rect 7268 6360 7272 6416
rect 7208 6356 7272 6360
rect 7288 6416 7352 6420
rect 7288 6360 7292 6416
rect 7292 6360 7348 6416
rect 7348 6360 7352 6416
rect 7288 6356 7352 6360
rect 7368 6416 7432 6420
rect 7368 6360 7372 6416
rect 7372 6360 7428 6416
rect 7428 6360 7432 6416
rect 7368 6356 7432 6360
rect 12456 6416 12520 6420
rect 12456 6360 12460 6416
rect 12460 6360 12516 6416
rect 12516 6360 12520 6416
rect 12456 6356 12520 6360
rect 12536 6416 12600 6420
rect 12536 6360 12540 6416
rect 12540 6360 12596 6416
rect 12596 6360 12600 6416
rect 12536 6356 12600 6360
rect 12616 6416 12680 6420
rect 12616 6360 12620 6416
rect 12620 6360 12676 6416
rect 12676 6360 12680 6416
rect 12616 6356 12680 6360
rect 12696 6416 12760 6420
rect 12696 6360 12700 6416
rect 12700 6360 12756 6416
rect 12756 6360 12760 6416
rect 12696 6356 12760 6360
rect 17784 6416 17848 6420
rect 17784 6360 17788 6416
rect 17788 6360 17844 6416
rect 17844 6360 17848 6416
rect 17784 6356 17848 6360
rect 17864 6416 17928 6420
rect 17864 6360 17868 6416
rect 17868 6360 17924 6416
rect 17924 6360 17928 6416
rect 17864 6356 17928 6360
rect 17944 6416 18008 6420
rect 17944 6360 17948 6416
rect 17948 6360 18004 6416
rect 18004 6360 18008 6416
rect 17944 6356 18008 6360
rect 18024 6416 18088 6420
rect 18024 6360 18028 6416
rect 18028 6360 18084 6416
rect 18084 6360 18088 6416
rect 18024 6356 18088 6360
rect 4464 5750 4528 5754
rect 4464 5694 4468 5750
rect 4468 5694 4524 5750
rect 4524 5694 4528 5750
rect 4464 5690 4528 5694
rect 4544 5750 4608 5754
rect 4544 5694 4548 5750
rect 4548 5694 4604 5750
rect 4604 5694 4608 5750
rect 4544 5690 4608 5694
rect 4624 5750 4688 5754
rect 4624 5694 4628 5750
rect 4628 5694 4684 5750
rect 4684 5694 4688 5750
rect 4624 5690 4688 5694
rect 4704 5750 4768 5754
rect 4704 5694 4708 5750
rect 4708 5694 4764 5750
rect 4764 5694 4768 5750
rect 4704 5690 4768 5694
rect 9792 5750 9856 5754
rect 9792 5694 9796 5750
rect 9796 5694 9852 5750
rect 9852 5694 9856 5750
rect 9792 5690 9856 5694
rect 9872 5750 9936 5754
rect 9872 5694 9876 5750
rect 9876 5694 9932 5750
rect 9932 5694 9936 5750
rect 9872 5690 9936 5694
rect 9952 5750 10016 5754
rect 9952 5694 9956 5750
rect 9956 5694 10012 5750
rect 10012 5694 10016 5750
rect 9952 5690 10016 5694
rect 10032 5750 10096 5754
rect 10032 5694 10036 5750
rect 10036 5694 10092 5750
rect 10092 5694 10096 5750
rect 10032 5690 10096 5694
rect 15120 5750 15184 5754
rect 15120 5694 15124 5750
rect 15124 5694 15180 5750
rect 15180 5694 15184 5750
rect 15120 5690 15184 5694
rect 15200 5750 15264 5754
rect 15200 5694 15204 5750
rect 15204 5694 15260 5750
rect 15260 5694 15264 5750
rect 15200 5690 15264 5694
rect 15280 5750 15344 5754
rect 15280 5694 15284 5750
rect 15284 5694 15340 5750
rect 15340 5694 15344 5750
rect 15280 5690 15344 5694
rect 15360 5750 15424 5754
rect 15360 5694 15364 5750
rect 15364 5694 15420 5750
rect 15420 5694 15424 5750
rect 15360 5690 15424 5694
rect 20448 5750 20512 5754
rect 20448 5694 20452 5750
rect 20452 5694 20508 5750
rect 20508 5694 20512 5750
rect 20448 5690 20512 5694
rect 20528 5750 20592 5754
rect 20528 5694 20532 5750
rect 20532 5694 20588 5750
rect 20588 5694 20592 5750
rect 20528 5690 20592 5694
rect 20608 5750 20672 5754
rect 20608 5694 20612 5750
rect 20612 5694 20668 5750
rect 20668 5694 20672 5750
rect 20608 5690 20672 5694
rect 20688 5750 20752 5754
rect 20688 5694 20692 5750
rect 20692 5694 20748 5750
rect 20748 5694 20752 5750
rect 20688 5690 20752 5694
rect 7128 5084 7192 5088
rect 7128 5028 7132 5084
rect 7132 5028 7188 5084
rect 7188 5028 7192 5084
rect 7128 5024 7192 5028
rect 7208 5084 7272 5088
rect 7208 5028 7212 5084
rect 7212 5028 7268 5084
rect 7268 5028 7272 5084
rect 7208 5024 7272 5028
rect 7288 5084 7352 5088
rect 7288 5028 7292 5084
rect 7292 5028 7348 5084
rect 7348 5028 7352 5084
rect 7288 5024 7352 5028
rect 7368 5084 7432 5088
rect 7368 5028 7372 5084
rect 7372 5028 7428 5084
rect 7428 5028 7432 5084
rect 7368 5024 7432 5028
rect 12456 5084 12520 5088
rect 12456 5028 12460 5084
rect 12460 5028 12516 5084
rect 12516 5028 12520 5084
rect 12456 5024 12520 5028
rect 12536 5084 12600 5088
rect 12536 5028 12540 5084
rect 12540 5028 12596 5084
rect 12596 5028 12600 5084
rect 12536 5024 12600 5028
rect 12616 5084 12680 5088
rect 12616 5028 12620 5084
rect 12620 5028 12676 5084
rect 12676 5028 12680 5084
rect 12616 5024 12680 5028
rect 12696 5084 12760 5088
rect 12696 5028 12700 5084
rect 12700 5028 12756 5084
rect 12756 5028 12760 5084
rect 12696 5024 12760 5028
rect 17784 5084 17848 5088
rect 17784 5028 17788 5084
rect 17788 5028 17844 5084
rect 17844 5028 17848 5084
rect 17784 5024 17848 5028
rect 17864 5084 17928 5088
rect 17864 5028 17868 5084
rect 17868 5028 17924 5084
rect 17924 5028 17928 5084
rect 17864 5024 17928 5028
rect 17944 5084 18008 5088
rect 17944 5028 17948 5084
rect 17948 5028 18004 5084
rect 18004 5028 18008 5084
rect 17944 5024 18008 5028
rect 18024 5084 18088 5088
rect 18024 5028 18028 5084
rect 18028 5028 18084 5084
rect 18084 5028 18088 5084
rect 18024 5024 18088 5028
rect 4464 4418 4528 4422
rect 4464 4362 4468 4418
rect 4468 4362 4524 4418
rect 4524 4362 4528 4418
rect 4464 4358 4528 4362
rect 4544 4418 4608 4422
rect 4544 4362 4548 4418
rect 4548 4362 4604 4418
rect 4604 4362 4608 4418
rect 4544 4358 4608 4362
rect 4624 4418 4688 4422
rect 4624 4362 4628 4418
rect 4628 4362 4684 4418
rect 4684 4362 4688 4418
rect 4624 4358 4688 4362
rect 4704 4418 4768 4422
rect 4704 4362 4708 4418
rect 4708 4362 4764 4418
rect 4764 4362 4768 4418
rect 4704 4358 4768 4362
rect 9792 4418 9856 4422
rect 9792 4362 9796 4418
rect 9796 4362 9852 4418
rect 9852 4362 9856 4418
rect 9792 4358 9856 4362
rect 9872 4418 9936 4422
rect 9872 4362 9876 4418
rect 9876 4362 9932 4418
rect 9932 4362 9936 4418
rect 9872 4358 9936 4362
rect 9952 4418 10016 4422
rect 9952 4362 9956 4418
rect 9956 4362 10012 4418
rect 10012 4362 10016 4418
rect 9952 4358 10016 4362
rect 10032 4418 10096 4422
rect 10032 4362 10036 4418
rect 10036 4362 10092 4418
rect 10092 4362 10096 4418
rect 10032 4358 10096 4362
rect 15120 4418 15184 4422
rect 15120 4362 15124 4418
rect 15124 4362 15180 4418
rect 15180 4362 15184 4418
rect 15120 4358 15184 4362
rect 15200 4418 15264 4422
rect 15200 4362 15204 4418
rect 15204 4362 15260 4418
rect 15260 4362 15264 4418
rect 15200 4358 15264 4362
rect 15280 4418 15344 4422
rect 15280 4362 15284 4418
rect 15284 4362 15340 4418
rect 15340 4362 15344 4418
rect 15280 4358 15344 4362
rect 15360 4418 15424 4422
rect 15360 4362 15364 4418
rect 15364 4362 15420 4418
rect 15420 4362 15424 4418
rect 15360 4358 15424 4362
rect 20448 4418 20512 4422
rect 20448 4362 20452 4418
rect 20452 4362 20508 4418
rect 20508 4362 20512 4418
rect 20448 4358 20512 4362
rect 20528 4418 20592 4422
rect 20528 4362 20532 4418
rect 20532 4362 20588 4418
rect 20588 4362 20592 4418
rect 20528 4358 20592 4362
rect 20608 4418 20672 4422
rect 20608 4362 20612 4418
rect 20612 4362 20668 4418
rect 20668 4362 20672 4418
rect 20608 4358 20672 4362
rect 20688 4418 20752 4422
rect 20688 4362 20692 4418
rect 20692 4362 20748 4418
rect 20748 4362 20752 4418
rect 20688 4358 20752 4362
rect 7128 3752 7192 3756
rect 7128 3696 7132 3752
rect 7132 3696 7188 3752
rect 7188 3696 7192 3752
rect 7128 3692 7192 3696
rect 7208 3752 7272 3756
rect 7208 3696 7212 3752
rect 7212 3696 7268 3752
rect 7268 3696 7272 3752
rect 7208 3692 7272 3696
rect 7288 3752 7352 3756
rect 7288 3696 7292 3752
rect 7292 3696 7348 3752
rect 7348 3696 7352 3752
rect 7288 3692 7352 3696
rect 7368 3752 7432 3756
rect 7368 3696 7372 3752
rect 7372 3696 7428 3752
rect 7428 3696 7432 3752
rect 7368 3692 7432 3696
rect 12456 3752 12520 3756
rect 12456 3696 12460 3752
rect 12460 3696 12516 3752
rect 12516 3696 12520 3752
rect 12456 3692 12520 3696
rect 12536 3752 12600 3756
rect 12536 3696 12540 3752
rect 12540 3696 12596 3752
rect 12596 3696 12600 3752
rect 12536 3692 12600 3696
rect 12616 3752 12680 3756
rect 12616 3696 12620 3752
rect 12620 3696 12676 3752
rect 12676 3696 12680 3752
rect 12616 3692 12680 3696
rect 12696 3752 12760 3756
rect 12696 3696 12700 3752
rect 12700 3696 12756 3752
rect 12756 3696 12760 3752
rect 12696 3692 12760 3696
rect 17784 3752 17848 3756
rect 17784 3696 17788 3752
rect 17788 3696 17844 3752
rect 17844 3696 17848 3752
rect 17784 3692 17848 3696
rect 17864 3752 17928 3756
rect 17864 3696 17868 3752
rect 17868 3696 17924 3752
rect 17924 3696 17928 3752
rect 17864 3692 17928 3696
rect 17944 3752 18008 3756
rect 17944 3696 17948 3752
rect 17948 3696 18004 3752
rect 18004 3696 18008 3752
rect 17944 3692 18008 3696
rect 18024 3752 18088 3756
rect 18024 3696 18028 3752
rect 18028 3696 18084 3752
rect 18084 3696 18088 3752
rect 18024 3692 18088 3696
rect 4464 3086 4528 3090
rect 4464 3030 4468 3086
rect 4468 3030 4524 3086
rect 4524 3030 4528 3086
rect 4464 3026 4528 3030
rect 4544 3086 4608 3090
rect 4544 3030 4548 3086
rect 4548 3030 4604 3086
rect 4604 3030 4608 3086
rect 4544 3026 4608 3030
rect 4624 3086 4688 3090
rect 4624 3030 4628 3086
rect 4628 3030 4684 3086
rect 4684 3030 4688 3086
rect 4624 3026 4688 3030
rect 4704 3086 4768 3090
rect 4704 3030 4708 3086
rect 4708 3030 4764 3086
rect 4764 3030 4768 3086
rect 4704 3026 4768 3030
rect 9792 3086 9856 3090
rect 9792 3030 9796 3086
rect 9796 3030 9852 3086
rect 9852 3030 9856 3086
rect 9792 3026 9856 3030
rect 9872 3086 9936 3090
rect 9872 3030 9876 3086
rect 9876 3030 9932 3086
rect 9932 3030 9936 3086
rect 9872 3026 9936 3030
rect 9952 3086 10016 3090
rect 9952 3030 9956 3086
rect 9956 3030 10012 3086
rect 10012 3030 10016 3086
rect 9952 3026 10016 3030
rect 10032 3086 10096 3090
rect 10032 3030 10036 3086
rect 10036 3030 10092 3086
rect 10092 3030 10096 3086
rect 10032 3026 10096 3030
rect 15120 3086 15184 3090
rect 15120 3030 15124 3086
rect 15124 3030 15180 3086
rect 15180 3030 15184 3086
rect 15120 3026 15184 3030
rect 15200 3086 15264 3090
rect 15200 3030 15204 3086
rect 15204 3030 15260 3086
rect 15260 3030 15264 3086
rect 15200 3026 15264 3030
rect 15280 3086 15344 3090
rect 15280 3030 15284 3086
rect 15284 3030 15340 3086
rect 15340 3030 15344 3086
rect 15280 3026 15344 3030
rect 15360 3086 15424 3090
rect 15360 3030 15364 3086
rect 15364 3030 15420 3086
rect 15420 3030 15424 3086
rect 15360 3026 15424 3030
rect 20448 3086 20512 3090
rect 20448 3030 20452 3086
rect 20452 3030 20508 3086
rect 20508 3030 20512 3086
rect 20448 3026 20512 3030
rect 20528 3086 20592 3090
rect 20528 3030 20532 3086
rect 20532 3030 20588 3086
rect 20588 3030 20592 3086
rect 20528 3026 20592 3030
rect 20608 3086 20672 3090
rect 20608 3030 20612 3086
rect 20612 3030 20668 3086
rect 20668 3030 20672 3086
rect 20608 3026 20672 3030
rect 20688 3086 20752 3090
rect 20688 3030 20692 3086
rect 20692 3030 20748 3086
rect 20748 3030 20752 3086
rect 20688 3026 20752 3030
rect 7128 2420 7192 2424
rect 7128 2364 7132 2420
rect 7132 2364 7188 2420
rect 7188 2364 7192 2420
rect 7128 2360 7192 2364
rect 7208 2420 7272 2424
rect 7208 2364 7212 2420
rect 7212 2364 7268 2420
rect 7268 2364 7272 2420
rect 7208 2360 7272 2364
rect 7288 2420 7352 2424
rect 7288 2364 7292 2420
rect 7292 2364 7348 2420
rect 7348 2364 7352 2420
rect 7288 2360 7352 2364
rect 7368 2420 7432 2424
rect 7368 2364 7372 2420
rect 7372 2364 7428 2420
rect 7428 2364 7432 2420
rect 7368 2360 7432 2364
rect 12456 2420 12520 2424
rect 12456 2364 12460 2420
rect 12460 2364 12516 2420
rect 12516 2364 12520 2420
rect 12456 2360 12520 2364
rect 12536 2420 12600 2424
rect 12536 2364 12540 2420
rect 12540 2364 12596 2420
rect 12596 2364 12600 2420
rect 12536 2360 12600 2364
rect 12616 2420 12680 2424
rect 12616 2364 12620 2420
rect 12620 2364 12676 2420
rect 12676 2364 12680 2420
rect 12616 2360 12680 2364
rect 12696 2420 12760 2424
rect 12696 2364 12700 2420
rect 12700 2364 12756 2420
rect 12756 2364 12760 2420
rect 12696 2360 12760 2364
rect 17784 2420 17848 2424
rect 17784 2364 17788 2420
rect 17788 2364 17844 2420
rect 17844 2364 17848 2420
rect 17784 2360 17848 2364
rect 17864 2420 17928 2424
rect 17864 2364 17868 2420
rect 17868 2364 17924 2420
rect 17924 2364 17928 2420
rect 17864 2360 17928 2364
rect 17944 2420 18008 2424
rect 17944 2364 17948 2420
rect 17948 2364 18004 2420
rect 18004 2364 18008 2420
rect 17944 2360 18008 2364
rect 18024 2420 18088 2424
rect 18024 2364 18028 2420
rect 18028 2364 18084 2420
rect 18084 2364 18088 2420
rect 18024 2360 18088 2364
rect 4464 1754 4528 1758
rect 4464 1698 4468 1754
rect 4468 1698 4524 1754
rect 4524 1698 4528 1754
rect 4464 1694 4528 1698
rect 4544 1754 4608 1758
rect 4544 1698 4548 1754
rect 4548 1698 4604 1754
rect 4604 1698 4608 1754
rect 4544 1694 4608 1698
rect 4624 1754 4688 1758
rect 4624 1698 4628 1754
rect 4628 1698 4684 1754
rect 4684 1698 4688 1754
rect 4624 1694 4688 1698
rect 4704 1754 4768 1758
rect 4704 1698 4708 1754
rect 4708 1698 4764 1754
rect 4764 1698 4768 1754
rect 4704 1694 4768 1698
rect 9792 1754 9856 1758
rect 9792 1698 9796 1754
rect 9796 1698 9852 1754
rect 9852 1698 9856 1754
rect 9792 1694 9856 1698
rect 9872 1754 9936 1758
rect 9872 1698 9876 1754
rect 9876 1698 9932 1754
rect 9932 1698 9936 1754
rect 9872 1694 9936 1698
rect 9952 1754 10016 1758
rect 9952 1698 9956 1754
rect 9956 1698 10012 1754
rect 10012 1698 10016 1754
rect 9952 1694 10016 1698
rect 10032 1754 10096 1758
rect 10032 1698 10036 1754
rect 10036 1698 10092 1754
rect 10092 1698 10096 1754
rect 10032 1694 10096 1698
rect 15120 1754 15184 1758
rect 15120 1698 15124 1754
rect 15124 1698 15180 1754
rect 15180 1698 15184 1754
rect 15120 1694 15184 1698
rect 15200 1754 15264 1758
rect 15200 1698 15204 1754
rect 15204 1698 15260 1754
rect 15260 1698 15264 1754
rect 15200 1694 15264 1698
rect 15280 1754 15344 1758
rect 15280 1698 15284 1754
rect 15284 1698 15340 1754
rect 15340 1698 15344 1754
rect 15280 1694 15344 1698
rect 15360 1754 15424 1758
rect 15360 1698 15364 1754
rect 15364 1698 15420 1754
rect 15420 1698 15424 1754
rect 15360 1694 15424 1698
rect 20448 1754 20512 1758
rect 20448 1698 20452 1754
rect 20452 1698 20508 1754
rect 20508 1698 20512 1754
rect 20448 1694 20512 1698
rect 20528 1754 20592 1758
rect 20528 1698 20532 1754
rect 20532 1698 20588 1754
rect 20588 1698 20592 1754
rect 20528 1694 20592 1698
rect 20608 1754 20672 1758
rect 20608 1698 20612 1754
rect 20612 1698 20668 1754
rect 20668 1698 20672 1754
rect 20608 1694 20672 1698
rect 20688 1754 20752 1758
rect 20688 1698 20692 1754
rect 20692 1698 20748 1754
rect 20748 1698 20752 1754
rect 20688 1694 20752 1698
rect 7128 1088 7192 1092
rect 7128 1032 7132 1088
rect 7132 1032 7188 1088
rect 7188 1032 7192 1088
rect 7128 1028 7192 1032
rect 7208 1088 7272 1092
rect 7208 1032 7212 1088
rect 7212 1032 7268 1088
rect 7268 1032 7272 1088
rect 7208 1028 7272 1032
rect 7288 1088 7352 1092
rect 7288 1032 7292 1088
rect 7292 1032 7348 1088
rect 7348 1032 7352 1088
rect 7288 1028 7352 1032
rect 7368 1088 7432 1092
rect 7368 1032 7372 1088
rect 7372 1032 7428 1088
rect 7428 1032 7432 1088
rect 7368 1028 7432 1032
rect 12456 1088 12520 1092
rect 12456 1032 12460 1088
rect 12460 1032 12516 1088
rect 12516 1032 12520 1088
rect 12456 1028 12520 1032
rect 12536 1088 12600 1092
rect 12536 1032 12540 1088
rect 12540 1032 12596 1088
rect 12596 1032 12600 1088
rect 12536 1028 12600 1032
rect 12616 1088 12680 1092
rect 12616 1032 12620 1088
rect 12620 1032 12676 1088
rect 12676 1032 12680 1088
rect 12616 1028 12680 1032
rect 12696 1088 12760 1092
rect 12696 1032 12700 1088
rect 12700 1032 12756 1088
rect 12756 1032 12760 1088
rect 12696 1028 12760 1032
rect 17784 1088 17848 1092
rect 17784 1032 17788 1088
rect 17788 1032 17844 1088
rect 17844 1032 17848 1088
rect 17784 1028 17848 1032
rect 17864 1088 17928 1092
rect 17864 1032 17868 1088
rect 17868 1032 17924 1088
rect 17924 1032 17928 1088
rect 17864 1028 17928 1032
rect 17944 1088 18008 1092
rect 17944 1032 17948 1088
rect 17948 1032 18004 1088
rect 18004 1032 18008 1088
rect 17944 1028 18008 1032
rect 18024 1088 18088 1092
rect 18024 1032 18028 1088
rect 18028 1032 18084 1088
rect 18084 1032 18088 1088
rect 18024 1028 18088 1032
<< metal4 >>
rect 4456 27066 4776 27082
rect 4456 27002 4464 27066
rect 4528 27002 4544 27066
rect 4608 27002 4624 27066
rect 4688 27002 4704 27066
rect 4768 27002 4776 27066
rect 4456 25734 4776 27002
rect 4456 25670 4464 25734
rect 4528 25670 4544 25734
rect 4608 25670 4624 25734
rect 4688 25670 4704 25734
rect 4768 25670 4776 25734
rect 4456 24402 4776 25670
rect 4456 24338 4464 24402
rect 4528 24338 4544 24402
rect 4608 24338 4624 24402
rect 4688 24338 4704 24402
rect 4768 24338 4776 24402
rect 4456 23070 4776 24338
rect 4456 23006 4464 23070
rect 4528 23006 4544 23070
rect 4608 23006 4624 23070
rect 4688 23006 4704 23070
rect 4768 23006 4776 23070
rect 4456 21738 4776 23006
rect 4456 21674 4464 21738
rect 4528 21674 4544 21738
rect 4608 21674 4624 21738
rect 4688 21674 4704 21738
rect 4768 21674 4776 21738
rect 4456 20970 4776 21674
rect 4456 20734 4498 20970
rect 4734 20734 4776 20970
rect 4456 20406 4776 20734
rect 4456 20342 4464 20406
rect 4528 20342 4544 20406
rect 4608 20342 4624 20406
rect 4688 20342 4704 20406
rect 4768 20342 4776 20406
rect 4456 19074 4776 20342
rect 4456 19010 4464 19074
rect 4528 19010 4544 19074
rect 4608 19010 4624 19074
rect 4688 19010 4704 19074
rect 4768 19010 4776 19074
rect 4456 17742 4776 19010
rect 4456 17678 4464 17742
rect 4528 17678 4544 17742
rect 4608 17678 4624 17742
rect 4688 17678 4704 17742
rect 4768 17678 4776 17742
rect 4456 16410 4776 17678
rect 4456 16346 4464 16410
rect 4528 16346 4544 16410
rect 4608 16346 4624 16410
rect 4688 16346 4704 16410
rect 4768 16346 4776 16410
rect 4456 15078 4776 16346
rect 4456 15014 4464 15078
rect 4528 15014 4544 15078
rect 4608 15014 4624 15078
rect 4688 15014 4704 15078
rect 4768 15014 4776 15078
rect 4456 13746 4776 15014
rect 4456 13682 4464 13746
rect 4528 13682 4544 13746
rect 4608 13682 4624 13746
rect 4688 13682 4704 13746
rect 4768 13682 4776 13746
rect 4456 12414 4776 13682
rect 4456 12350 4464 12414
rect 4528 12350 4544 12414
rect 4608 12350 4624 12414
rect 4688 12350 4704 12414
rect 4768 12350 4776 12414
rect 4456 11082 4776 12350
rect 4456 11018 4464 11082
rect 4528 11018 4544 11082
rect 4608 11018 4624 11082
rect 4688 11018 4704 11082
rect 4768 11018 4776 11082
rect 4456 9750 4776 11018
rect 4456 9686 4464 9750
rect 4528 9686 4544 9750
rect 4608 9686 4624 9750
rect 4688 9686 4704 9750
rect 4768 9686 4776 9750
rect 4456 8418 4776 9686
rect 4456 8354 4464 8418
rect 4528 8354 4544 8418
rect 4608 8354 4624 8418
rect 4688 8354 4704 8418
rect 4768 8354 4776 8418
rect 4456 7086 4776 8354
rect 4456 7022 4464 7086
rect 4528 7022 4544 7086
rect 4608 7022 4624 7086
rect 4688 7022 4704 7086
rect 4768 7022 4776 7086
rect 4456 5754 4776 7022
rect 4456 5690 4464 5754
rect 4528 5690 4544 5754
rect 4608 5690 4624 5754
rect 4688 5690 4704 5754
rect 4768 5690 4776 5754
rect 4456 4422 4776 5690
rect 4456 4358 4464 4422
rect 4528 4358 4544 4422
rect 4608 4358 4624 4422
rect 4688 4358 4704 4422
rect 4768 4358 4776 4422
rect 4456 3090 4776 4358
rect 4456 3026 4464 3090
rect 4528 3026 4544 3090
rect 4608 3026 4624 3090
rect 4688 3026 4704 3090
rect 4768 3026 4776 3090
rect 4456 1758 4776 3026
rect 4456 1694 4464 1758
rect 4528 1694 4544 1758
rect 4608 1694 4624 1758
rect 4688 1694 4704 1758
rect 4768 1694 4776 1758
rect 4456 1012 4776 1694
rect 7120 26400 7440 27082
rect 7120 26336 7128 26400
rect 7192 26336 7208 26400
rect 7272 26336 7288 26400
rect 7352 26336 7368 26400
rect 7432 26336 7440 26400
rect 7120 25068 7440 26336
rect 7120 25004 7128 25068
rect 7192 25004 7208 25068
rect 7272 25004 7288 25068
rect 7352 25004 7368 25068
rect 7432 25004 7440 25068
rect 7120 23736 7440 25004
rect 7120 23672 7128 23736
rect 7192 23672 7208 23736
rect 7272 23672 7288 23736
rect 7352 23672 7368 23736
rect 7432 23672 7440 23736
rect 7120 22404 7440 23672
rect 7120 22340 7128 22404
rect 7192 22340 7208 22404
rect 7272 22340 7288 22404
rect 7352 22340 7368 22404
rect 7432 22340 7440 22404
rect 7120 21072 7440 22340
rect 7120 21008 7128 21072
rect 7192 21008 7208 21072
rect 7272 21008 7288 21072
rect 7352 21008 7368 21072
rect 7432 21008 7440 21072
rect 7120 19740 7440 21008
rect 7120 19676 7128 19740
rect 7192 19676 7208 19740
rect 7272 19676 7288 19740
rect 7352 19676 7368 19740
rect 7432 19676 7440 19740
rect 7120 18408 7440 19676
rect 7120 18344 7128 18408
rect 7192 18344 7208 18408
rect 7272 18344 7288 18408
rect 7352 18344 7368 18408
rect 7432 18344 7440 18408
rect 7120 17076 7440 18344
rect 7120 17012 7128 17076
rect 7192 17012 7208 17076
rect 7272 17012 7288 17076
rect 7352 17012 7368 17076
rect 7432 17012 7440 17076
rect 7120 15744 7440 17012
rect 7120 15680 7128 15744
rect 7192 15680 7208 15744
rect 7272 15680 7288 15744
rect 7352 15680 7368 15744
rect 7432 15680 7440 15744
rect 7120 14412 7440 15680
rect 7120 14348 7128 14412
rect 7192 14348 7208 14412
rect 7272 14348 7288 14412
rect 7352 14348 7368 14412
rect 7432 14348 7440 14412
rect 7120 13080 7440 14348
rect 7120 13016 7128 13080
rect 7192 13016 7208 13080
rect 7272 13016 7288 13080
rect 7352 13016 7368 13080
rect 7432 13016 7440 13080
rect 7120 11748 7440 13016
rect 7120 11684 7128 11748
rect 7192 11684 7208 11748
rect 7272 11684 7288 11748
rect 7352 11684 7368 11748
rect 7432 11684 7440 11748
rect 7120 10416 7440 11684
rect 7120 10352 7128 10416
rect 7192 10352 7208 10416
rect 7272 10352 7288 10416
rect 7352 10352 7368 10416
rect 7432 10352 7440 10416
rect 7120 9084 7440 10352
rect 7120 9020 7128 9084
rect 7192 9020 7208 9084
rect 7272 9020 7288 9084
rect 7352 9020 7368 9084
rect 7432 9020 7440 9084
rect 7120 7752 7440 9020
rect 7120 7688 7128 7752
rect 7192 7688 7208 7752
rect 7272 7688 7288 7752
rect 7352 7688 7368 7752
rect 7432 7688 7440 7752
rect 7120 6420 7440 7688
rect 7120 6356 7128 6420
rect 7192 6356 7208 6420
rect 7272 6356 7288 6420
rect 7352 6356 7368 6420
rect 7432 6356 7440 6420
rect 7120 5088 7440 6356
rect 7120 5024 7128 5088
rect 7192 5024 7208 5088
rect 7272 5024 7288 5088
rect 7352 5024 7368 5088
rect 7432 5024 7440 5088
rect 7120 3756 7440 5024
rect 7120 3692 7128 3756
rect 7192 3692 7208 3756
rect 7272 3692 7288 3756
rect 7352 3692 7368 3756
rect 7432 3692 7440 3756
rect 7120 2970 7440 3692
rect 7120 2734 7162 2970
rect 7398 2734 7440 2970
rect 7120 2424 7440 2734
rect 7120 2360 7128 2424
rect 7192 2360 7208 2424
rect 7272 2360 7288 2424
rect 7352 2360 7368 2424
rect 7432 2360 7440 2424
rect 7120 1092 7440 2360
rect 7120 1028 7128 1092
rect 7192 1028 7208 1092
rect 7272 1028 7288 1092
rect 7352 1028 7368 1092
rect 7432 1028 7440 1092
rect 7120 1012 7440 1028
rect 9784 27066 10104 27082
rect 9784 27002 9792 27066
rect 9856 27002 9872 27066
rect 9936 27002 9952 27066
rect 10016 27002 10032 27066
rect 10096 27002 10104 27066
rect 9784 25734 10104 27002
rect 9784 25670 9792 25734
rect 9856 25670 9872 25734
rect 9936 25670 9952 25734
rect 10016 25670 10032 25734
rect 10096 25670 10104 25734
rect 9784 24402 10104 25670
rect 9784 24338 9792 24402
rect 9856 24338 9872 24402
rect 9936 24338 9952 24402
rect 10016 24338 10032 24402
rect 10096 24338 10104 24402
rect 9784 23070 10104 24338
rect 9784 23006 9792 23070
rect 9856 23006 9872 23070
rect 9936 23006 9952 23070
rect 10016 23006 10032 23070
rect 10096 23006 10104 23070
rect 9784 21738 10104 23006
rect 9784 21674 9792 21738
rect 9856 21674 9872 21738
rect 9936 21674 9952 21738
rect 10016 21674 10032 21738
rect 10096 21674 10104 21738
rect 9784 20970 10104 21674
rect 9784 20734 9826 20970
rect 10062 20734 10104 20970
rect 9784 20406 10104 20734
rect 9784 20342 9792 20406
rect 9856 20342 9872 20406
rect 9936 20342 9952 20406
rect 10016 20342 10032 20406
rect 10096 20342 10104 20406
rect 9784 19074 10104 20342
rect 9784 19010 9792 19074
rect 9856 19010 9872 19074
rect 9936 19010 9952 19074
rect 10016 19010 10032 19074
rect 10096 19010 10104 19074
rect 9784 17742 10104 19010
rect 9784 17678 9792 17742
rect 9856 17678 9872 17742
rect 9936 17678 9952 17742
rect 10016 17678 10032 17742
rect 10096 17678 10104 17742
rect 9784 16410 10104 17678
rect 9784 16346 9792 16410
rect 9856 16346 9872 16410
rect 9936 16346 9952 16410
rect 10016 16346 10032 16410
rect 10096 16346 10104 16410
rect 9784 15078 10104 16346
rect 9784 15014 9792 15078
rect 9856 15014 9872 15078
rect 9936 15014 9952 15078
rect 10016 15014 10032 15078
rect 10096 15014 10104 15078
rect 9784 13746 10104 15014
rect 9784 13682 9792 13746
rect 9856 13682 9872 13746
rect 9936 13682 9952 13746
rect 10016 13682 10032 13746
rect 10096 13682 10104 13746
rect 9784 12414 10104 13682
rect 9784 12350 9792 12414
rect 9856 12350 9872 12414
rect 9936 12350 9952 12414
rect 10016 12350 10032 12414
rect 10096 12350 10104 12414
rect 9784 11082 10104 12350
rect 9784 11018 9792 11082
rect 9856 11018 9872 11082
rect 9936 11018 9952 11082
rect 10016 11018 10032 11082
rect 10096 11018 10104 11082
rect 9784 9750 10104 11018
rect 9784 9686 9792 9750
rect 9856 9686 9872 9750
rect 9936 9686 9952 9750
rect 10016 9686 10032 9750
rect 10096 9686 10104 9750
rect 9784 8418 10104 9686
rect 9784 8354 9792 8418
rect 9856 8354 9872 8418
rect 9936 8354 9952 8418
rect 10016 8354 10032 8418
rect 10096 8354 10104 8418
rect 9784 7086 10104 8354
rect 9784 7022 9792 7086
rect 9856 7022 9872 7086
rect 9936 7022 9952 7086
rect 10016 7022 10032 7086
rect 10096 7022 10104 7086
rect 9784 5754 10104 7022
rect 9784 5690 9792 5754
rect 9856 5690 9872 5754
rect 9936 5690 9952 5754
rect 10016 5690 10032 5754
rect 10096 5690 10104 5754
rect 9784 4422 10104 5690
rect 9784 4358 9792 4422
rect 9856 4358 9872 4422
rect 9936 4358 9952 4422
rect 10016 4358 10032 4422
rect 10096 4358 10104 4422
rect 9784 3090 10104 4358
rect 9784 3026 9792 3090
rect 9856 3026 9872 3090
rect 9936 3026 9952 3090
rect 10016 3026 10032 3090
rect 10096 3026 10104 3090
rect 9784 1758 10104 3026
rect 9784 1694 9792 1758
rect 9856 1694 9872 1758
rect 9936 1694 9952 1758
rect 10016 1694 10032 1758
rect 10096 1694 10104 1758
rect 9784 1012 10104 1694
rect 12448 26400 12768 27082
rect 12448 26336 12456 26400
rect 12520 26336 12536 26400
rect 12600 26336 12616 26400
rect 12680 26336 12696 26400
rect 12760 26336 12768 26400
rect 12448 25068 12768 26336
rect 12448 25004 12456 25068
rect 12520 25004 12536 25068
rect 12600 25004 12616 25068
rect 12680 25004 12696 25068
rect 12760 25004 12768 25068
rect 12448 23736 12768 25004
rect 12448 23672 12456 23736
rect 12520 23672 12536 23736
rect 12600 23672 12616 23736
rect 12680 23672 12696 23736
rect 12760 23672 12768 23736
rect 12448 22404 12768 23672
rect 12448 22340 12456 22404
rect 12520 22340 12536 22404
rect 12600 22340 12616 22404
rect 12680 22340 12696 22404
rect 12760 22340 12768 22404
rect 12448 21072 12768 22340
rect 12448 21008 12456 21072
rect 12520 21008 12536 21072
rect 12600 21008 12616 21072
rect 12680 21008 12696 21072
rect 12760 21008 12768 21072
rect 12448 19740 12768 21008
rect 12448 19676 12456 19740
rect 12520 19676 12536 19740
rect 12600 19676 12616 19740
rect 12680 19676 12696 19740
rect 12760 19676 12768 19740
rect 12448 18408 12768 19676
rect 12448 18344 12456 18408
rect 12520 18344 12536 18408
rect 12600 18344 12616 18408
rect 12680 18344 12696 18408
rect 12760 18344 12768 18408
rect 12448 17076 12768 18344
rect 12448 17012 12456 17076
rect 12520 17012 12536 17076
rect 12600 17012 12616 17076
rect 12680 17012 12696 17076
rect 12760 17012 12768 17076
rect 12448 15744 12768 17012
rect 12448 15680 12456 15744
rect 12520 15680 12536 15744
rect 12600 15680 12616 15744
rect 12680 15680 12696 15744
rect 12760 15680 12768 15744
rect 12448 14412 12768 15680
rect 12448 14348 12456 14412
rect 12520 14348 12536 14412
rect 12600 14348 12616 14412
rect 12680 14348 12696 14412
rect 12760 14348 12768 14412
rect 12448 13080 12768 14348
rect 12448 13016 12456 13080
rect 12520 13016 12536 13080
rect 12600 13016 12616 13080
rect 12680 13016 12696 13080
rect 12760 13016 12768 13080
rect 12448 11748 12768 13016
rect 12448 11684 12456 11748
rect 12520 11684 12536 11748
rect 12600 11684 12616 11748
rect 12680 11684 12696 11748
rect 12760 11684 12768 11748
rect 12448 10416 12768 11684
rect 12448 10352 12456 10416
rect 12520 10352 12536 10416
rect 12600 10352 12616 10416
rect 12680 10352 12696 10416
rect 12760 10352 12768 10416
rect 12448 9084 12768 10352
rect 12448 9020 12456 9084
rect 12520 9020 12536 9084
rect 12600 9020 12616 9084
rect 12680 9020 12696 9084
rect 12760 9020 12768 9084
rect 12448 7752 12768 9020
rect 12448 7688 12456 7752
rect 12520 7688 12536 7752
rect 12600 7688 12616 7752
rect 12680 7688 12696 7752
rect 12760 7688 12768 7752
rect 12448 6420 12768 7688
rect 12448 6356 12456 6420
rect 12520 6356 12536 6420
rect 12600 6356 12616 6420
rect 12680 6356 12696 6420
rect 12760 6356 12768 6420
rect 12448 5088 12768 6356
rect 12448 5024 12456 5088
rect 12520 5024 12536 5088
rect 12600 5024 12616 5088
rect 12680 5024 12696 5088
rect 12760 5024 12768 5088
rect 12448 3756 12768 5024
rect 12448 3692 12456 3756
rect 12520 3692 12536 3756
rect 12600 3692 12616 3756
rect 12680 3692 12696 3756
rect 12760 3692 12768 3756
rect 12448 2970 12768 3692
rect 12448 2734 12490 2970
rect 12726 2734 12768 2970
rect 12448 2424 12768 2734
rect 12448 2360 12456 2424
rect 12520 2360 12536 2424
rect 12600 2360 12616 2424
rect 12680 2360 12696 2424
rect 12760 2360 12768 2424
rect 12448 1092 12768 2360
rect 12448 1028 12456 1092
rect 12520 1028 12536 1092
rect 12600 1028 12616 1092
rect 12680 1028 12696 1092
rect 12760 1028 12768 1092
rect 12448 1012 12768 1028
rect 15112 27066 15432 27082
rect 15112 27002 15120 27066
rect 15184 27002 15200 27066
rect 15264 27002 15280 27066
rect 15344 27002 15360 27066
rect 15424 27002 15432 27066
rect 15112 25734 15432 27002
rect 15112 25670 15120 25734
rect 15184 25670 15200 25734
rect 15264 25670 15280 25734
rect 15344 25670 15360 25734
rect 15424 25670 15432 25734
rect 15112 24402 15432 25670
rect 15112 24338 15120 24402
rect 15184 24338 15200 24402
rect 15264 24338 15280 24402
rect 15344 24338 15360 24402
rect 15424 24338 15432 24402
rect 15112 23070 15432 24338
rect 15112 23006 15120 23070
rect 15184 23006 15200 23070
rect 15264 23006 15280 23070
rect 15344 23006 15360 23070
rect 15424 23006 15432 23070
rect 15112 21738 15432 23006
rect 15112 21674 15120 21738
rect 15184 21674 15200 21738
rect 15264 21674 15280 21738
rect 15344 21674 15360 21738
rect 15424 21674 15432 21738
rect 15112 20970 15432 21674
rect 15112 20734 15154 20970
rect 15390 20734 15432 20970
rect 15112 20406 15432 20734
rect 15112 20342 15120 20406
rect 15184 20342 15200 20406
rect 15264 20342 15280 20406
rect 15344 20342 15360 20406
rect 15424 20342 15432 20406
rect 15112 19074 15432 20342
rect 15112 19010 15120 19074
rect 15184 19010 15200 19074
rect 15264 19010 15280 19074
rect 15344 19010 15360 19074
rect 15424 19010 15432 19074
rect 15112 17742 15432 19010
rect 15112 17678 15120 17742
rect 15184 17678 15200 17742
rect 15264 17678 15280 17742
rect 15344 17678 15360 17742
rect 15424 17678 15432 17742
rect 15112 16410 15432 17678
rect 15112 16346 15120 16410
rect 15184 16346 15200 16410
rect 15264 16346 15280 16410
rect 15344 16346 15360 16410
rect 15424 16346 15432 16410
rect 15112 15078 15432 16346
rect 15112 15014 15120 15078
rect 15184 15014 15200 15078
rect 15264 15014 15280 15078
rect 15344 15014 15360 15078
rect 15424 15014 15432 15078
rect 15112 13746 15432 15014
rect 15112 13682 15120 13746
rect 15184 13682 15200 13746
rect 15264 13682 15280 13746
rect 15344 13682 15360 13746
rect 15424 13682 15432 13746
rect 15112 12414 15432 13682
rect 15112 12350 15120 12414
rect 15184 12350 15200 12414
rect 15264 12350 15280 12414
rect 15344 12350 15360 12414
rect 15424 12350 15432 12414
rect 15112 11082 15432 12350
rect 15112 11018 15120 11082
rect 15184 11018 15200 11082
rect 15264 11018 15280 11082
rect 15344 11018 15360 11082
rect 15424 11018 15432 11082
rect 15112 9750 15432 11018
rect 15112 9686 15120 9750
rect 15184 9686 15200 9750
rect 15264 9686 15280 9750
rect 15344 9686 15360 9750
rect 15424 9686 15432 9750
rect 15112 8418 15432 9686
rect 15112 8354 15120 8418
rect 15184 8354 15200 8418
rect 15264 8354 15280 8418
rect 15344 8354 15360 8418
rect 15424 8354 15432 8418
rect 15112 7086 15432 8354
rect 15112 7022 15120 7086
rect 15184 7022 15200 7086
rect 15264 7022 15280 7086
rect 15344 7022 15360 7086
rect 15424 7022 15432 7086
rect 15112 5754 15432 7022
rect 15112 5690 15120 5754
rect 15184 5690 15200 5754
rect 15264 5690 15280 5754
rect 15344 5690 15360 5754
rect 15424 5690 15432 5754
rect 15112 4422 15432 5690
rect 15112 4358 15120 4422
rect 15184 4358 15200 4422
rect 15264 4358 15280 4422
rect 15344 4358 15360 4422
rect 15424 4358 15432 4422
rect 15112 3090 15432 4358
rect 15112 3026 15120 3090
rect 15184 3026 15200 3090
rect 15264 3026 15280 3090
rect 15344 3026 15360 3090
rect 15424 3026 15432 3090
rect 15112 1758 15432 3026
rect 15112 1694 15120 1758
rect 15184 1694 15200 1758
rect 15264 1694 15280 1758
rect 15344 1694 15360 1758
rect 15424 1694 15432 1758
rect 15112 1012 15432 1694
rect 17776 26400 18096 27082
rect 17776 26336 17784 26400
rect 17848 26336 17864 26400
rect 17928 26336 17944 26400
rect 18008 26336 18024 26400
rect 18088 26336 18096 26400
rect 17776 25068 18096 26336
rect 17776 25004 17784 25068
rect 17848 25004 17864 25068
rect 17928 25004 17944 25068
rect 18008 25004 18024 25068
rect 18088 25004 18096 25068
rect 17776 23736 18096 25004
rect 17776 23672 17784 23736
rect 17848 23672 17864 23736
rect 17928 23672 17944 23736
rect 18008 23672 18024 23736
rect 18088 23672 18096 23736
rect 17776 22404 18096 23672
rect 17776 22340 17784 22404
rect 17848 22340 17864 22404
rect 17928 22340 17944 22404
rect 18008 22340 18024 22404
rect 18088 22340 18096 22404
rect 17776 21072 18096 22340
rect 17776 21008 17784 21072
rect 17848 21008 17864 21072
rect 17928 21008 17944 21072
rect 18008 21008 18024 21072
rect 18088 21008 18096 21072
rect 17776 19740 18096 21008
rect 17776 19676 17784 19740
rect 17848 19676 17864 19740
rect 17928 19676 17944 19740
rect 18008 19676 18024 19740
rect 18088 19676 18096 19740
rect 17776 18408 18096 19676
rect 17776 18344 17784 18408
rect 17848 18344 17864 18408
rect 17928 18344 17944 18408
rect 18008 18344 18024 18408
rect 18088 18344 18096 18408
rect 17776 17076 18096 18344
rect 17776 17012 17784 17076
rect 17848 17012 17864 17076
rect 17928 17012 17944 17076
rect 18008 17012 18024 17076
rect 18088 17012 18096 17076
rect 17776 15744 18096 17012
rect 17776 15680 17784 15744
rect 17848 15680 17864 15744
rect 17928 15680 17944 15744
rect 18008 15680 18024 15744
rect 18088 15680 18096 15744
rect 17776 14412 18096 15680
rect 17776 14348 17784 14412
rect 17848 14348 17864 14412
rect 17928 14348 17944 14412
rect 18008 14348 18024 14412
rect 18088 14348 18096 14412
rect 17776 13080 18096 14348
rect 17776 13016 17784 13080
rect 17848 13016 17864 13080
rect 17928 13016 17944 13080
rect 18008 13016 18024 13080
rect 18088 13016 18096 13080
rect 17776 11748 18096 13016
rect 17776 11684 17784 11748
rect 17848 11684 17864 11748
rect 17928 11684 17944 11748
rect 18008 11684 18024 11748
rect 18088 11684 18096 11748
rect 17776 10416 18096 11684
rect 17776 10352 17784 10416
rect 17848 10352 17864 10416
rect 17928 10352 17944 10416
rect 18008 10352 18024 10416
rect 18088 10352 18096 10416
rect 17776 9084 18096 10352
rect 17776 9020 17784 9084
rect 17848 9020 17864 9084
rect 17928 9020 17944 9084
rect 18008 9020 18024 9084
rect 18088 9020 18096 9084
rect 17776 7752 18096 9020
rect 17776 7688 17784 7752
rect 17848 7688 17864 7752
rect 17928 7688 17944 7752
rect 18008 7688 18024 7752
rect 18088 7688 18096 7752
rect 17776 6420 18096 7688
rect 17776 6356 17784 6420
rect 17848 6356 17864 6420
rect 17928 6356 17944 6420
rect 18008 6356 18024 6420
rect 18088 6356 18096 6420
rect 17776 5088 18096 6356
rect 17776 5024 17784 5088
rect 17848 5024 17864 5088
rect 17928 5024 17944 5088
rect 18008 5024 18024 5088
rect 18088 5024 18096 5088
rect 17776 3756 18096 5024
rect 17776 3692 17784 3756
rect 17848 3692 17864 3756
rect 17928 3692 17944 3756
rect 18008 3692 18024 3756
rect 18088 3692 18096 3756
rect 17776 2970 18096 3692
rect 17776 2734 17818 2970
rect 18054 2734 18096 2970
rect 17776 2424 18096 2734
rect 17776 2360 17784 2424
rect 17848 2360 17864 2424
rect 17928 2360 17944 2424
rect 18008 2360 18024 2424
rect 18088 2360 18096 2424
rect 17776 1092 18096 2360
rect 17776 1028 17784 1092
rect 17848 1028 17864 1092
rect 17928 1028 17944 1092
rect 18008 1028 18024 1092
rect 18088 1028 18096 1092
rect 17776 1012 18096 1028
rect 20440 27066 20760 27082
rect 20440 27002 20448 27066
rect 20512 27002 20528 27066
rect 20592 27002 20608 27066
rect 20672 27002 20688 27066
rect 20752 27002 20760 27066
rect 20440 25734 20760 27002
rect 20440 25670 20448 25734
rect 20512 25670 20528 25734
rect 20592 25670 20608 25734
rect 20672 25670 20688 25734
rect 20752 25670 20760 25734
rect 20440 24402 20760 25670
rect 20440 24338 20448 24402
rect 20512 24338 20528 24402
rect 20592 24338 20608 24402
rect 20672 24338 20688 24402
rect 20752 24338 20760 24402
rect 20440 23070 20760 24338
rect 20440 23006 20448 23070
rect 20512 23006 20528 23070
rect 20592 23006 20608 23070
rect 20672 23006 20688 23070
rect 20752 23006 20760 23070
rect 20440 21738 20760 23006
rect 20440 21674 20448 21738
rect 20512 21674 20528 21738
rect 20592 21674 20608 21738
rect 20672 21674 20688 21738
rect 20752 21674 20760 21738
rect 20440 20970 20760 21674
rect 20440 20734 20482 20970
rect 20718 20734 20760 20970
rect 20440 20406 20760 20734
rect 20440 20342 20448 20406
rect 20512 20342 20528 20406
rect 20592 20342 20608 20406
rect 20672 20342 20688 20406
rect 20752 20342 20760 20406
rect 20440 19074 20760 20342
rect 20440 19010 20448 19074
rect 20512 19010 20528 19074
rect 20592 19010 20608 19074
rect 20672 19010 20688 19074
rect 20752 19010 20760 19074
rect 20440 17742 20760 19010
rect 20440 17678 20448 17742
rect 20512 17678 20528 17742
rect 20592 17678 20608 17742
rect 20672 17678 20688 17742
rect 20752 17678 20760 17742
rect 20440 16410 20760 17678
rect 20440 16346 20448 16410
rect 20512 16346 20528 16410
rect 20592 16346 20608 16410
rect 20672 16346 20688 16410
rect 20752 16346 20760 16410
rect 20440 15078 20760 16346
rect 20440 15014 20448 15078
rect 20512 15014 20528 15078
rect 20592 15014 20608 15078
rect 20672 15014 20688 15078
rect 20752 15014 20760 15078
rect 20440 13746 20760 15014
rect 20440 13682 20448 13746
rect 20512 13682 20528 13746
rect 20592 13682 20608 13746
rect 20672 13682 20688 13746
rect 20752 13682 20760 13746
rect 20440 12414 20760 13682
rect 20440 12350 20448 12414
rect 20512 12350 20528 12414
rect 20592 12350 20608 12414
rect 20672 12350 20688 12414
rect 20752 12350 20760 12414
rect 20440 11082 20760 12350
rect 20440 11018 20448 11082
rect 20512 11018 20528 11082
rect 20592 11018 20608 11082
rect 20672 11018 20688 11082
rect 20752 11018 20760 11082
rect 20440 9750 20760 11018
rect 20440 9686 20448 9750
rect 20512 9686 20528 9750
rect 20592 9686 20608 9750
rect 20672 9686 20688 9750
rect 20752 9686 20760 9750
rect 20440 8418 20760 9686
rect 20440 8354 20448 8418
rect 20512 8354 20528 8418
rect 20592 8354 20608 8418
rect 20672 8354 20688 8418
rect 20752 8354 20760 8418
rect 20440 7086 20760 8354
rect 20440 7022 20448 7086
rect 20512 7022 20528 7086
rect 20592 7022 20608 7086
rect 20672 7022 20688 7086
rect 20752 7022 20760 7086
rect 20440 5754 20760 7022
rect 20440 5690 20448 5754
rect 20512 5690 20528 5754
rect 20592 5690 20608 5754
rect 20672 5690 20688 5754
rect 20752 5690 20760 5754
rect 20440 4422 20760 5690
rect 20440 4358 20448 4422
rect 20512 4358 20528 4422
rect 20592 4358 20608 4422
rect 20672 4358 20688 4422
rect 20752 4358 20760 4422
rect 20440 3090 20760 4358
rect 20440 3026 20448 3090
rect 20512 3026 20528 3090
rect 20592 3026 20608 3090
rect 20672 3026 20688 3090
rect 20752 3026 20760 3090
rect 20440 1758 20760 3026
rect 20440 1694 20448 1758
rect 20512 1694 20528 1758
rect 20592 1694 20608 1758
rect 20672 1694 20688 1758
rect 20752 1694 20760 1758
rect 20440 1012 20760 1694
<< via4 >>
rect 4498 20734 4734 20970
rect 7162 2734 7398 2970
rect 9826 20734 10062 20970
rect 12490 2734 12726 2970
rect 15154 20734 15390 20970
rect 17818 2734 18054 2970
rect 20482 20734 20718 20970
<< metal5 >>
rect 1952 20970 23264 21012
rect 1952 20734 4498 20970
rect 4734 20734 9826 20970
rect 10062 20734 15154 20970
rect 15390 20734 20482 20970
rect 20718 20734 23264 20970
rect 1952 20692 23264 20734
rect 1952 2970 23264 3012
rect 1952 2734 7162 2970
rect 7398 2734 12490 2970
rect 12726 2734 17818 2970
rect 18054 2734 23264 2970
rect 1952 2692 23264 2734
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap1_0 $PDKPATH/libs.ref/sky130_fd_sc_ms/mag
timestamp 1607194124
transform 1 0 2816 0 1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_3 $PDKPATH/libs.ref/sky130_fd_sc_ms/mag
timestamp 1607194124
transform 1 0 2048 0 1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_2
timestamp 1607194124
transform 1 0 1952 0 1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap0_0
timestamp 1607194124
transform 1 0 2816 0 -1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_1
timestamp 1607194124
transform 1 0 2048 0 -1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_0
timestamp 1607194124
transform 1 0 1952 0 -1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_31 $PDKPATH/libs.ref/sky130_fd_sc_ms/mag
timestamp 1607194124
transform 1 0 3296 0 1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap1_0 $PDKPATH/libs.ref/sky130_fd_sc_ms/mag
timestamp 1607194124
transform 1 0 2912 0 1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_0
timestamp 1607194124
transform 1 0 3296 0 -1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap0_0
timestamp 1607194124
transform 1 0 2912 0 -1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_30
timestamp 1607194124
transform 1 0 4544 0 1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap1_1
timestamp 1607194124
transform 1 0 4160 0 1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap1_1
timestamp 1607194124
transform 1 0 4064 0 1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_1
timestamp 1607194124
transform 1 0 4544 0 -1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap0_1
timestamp 1607194124
transform 1 0 4160 0 -1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap0_1
timestamp 1607194124
transform 1 0 4064 0 -1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap1_2
timestamp 1607194124
transform 1 0 5408 0 1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap1_2
timestamp 1607194124
transform 1 0 5312 0 1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap0_2
timestamp 1607194124
transform 1 0 5408 0 -1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap0_2
timestamp 1607194124
transform 1 0 5312 0 -1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap1_3
timestamp 1607194124
transform 1 0 6656 0 1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap1_3
timestamp 1607194124
transform 1 0 6560 0 1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_29
timestamp 1607194124
transform 1 0 5792 0 1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap0_3
timestamp 1607194124
transform 1 0 6656 0 -1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap0_3
timestamp 1607194124
transform 1 0 6560 0 -1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_2
timestamp 1607194124
transform 1 0 5792 0 -1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_28
timestamp 1607194124
transform 1 0 7040 0 1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_3
timestamp 1607194124
transform 1 0 7040 0 -1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_27
timestamp 1607194124
transform 1 0 8288 0 1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap1_4
timestamp 1607194124
transform 1 0 7904 0 1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap1_4
timestamp 1607194124
transform 1 0 7808 0 1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_4
timestamp 1607194124
transform 1 0 8288 0 -1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap0_4
timestamp 1607194124
transform 1 0 7904 0 -1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap0_4
timestamp 1607194124
transform 1 0 7808 0 -1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap1_5
timestamp 1607194124
transform 1 0 9152 0 1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap1_5
timestamp 1607194124
transform 1 0 9056 0 1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap0_5
timestamp 1607194124
transform 1 0 9152 0 -1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap0_5
timestamp 1607194124
transform 1 0 9056 0 -1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap1_6
timestamp 1607194124
transform 1 0 10400 0 1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap1_6
timestamp 1607194124
transform 1 0 10304 0 1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_26
timestamp 1607194124
transform 1 0 9536 0 1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap0_6
timestamp 1607194124
transform 1 0 10400 0 -1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap0_6
timestamp 1607194124
transform 1 0 10304 0 -1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_5
timestamp 1607194124
transform 1 0 9536 0 -1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_25
timestamp 1607194124
transform 1 0 10784 0 1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_6
timestamp 1607194124
transform 1 0 10784 0 -1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_24
timestamp 1607194124
transform 1 0 12032 0 1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap1_7
timestamp 1607194124
transform 1 0 11648 0 1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap1_7
timestamp 1607194124
transform 1 0 11552 0 1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_7
timestamp 1607194124
transform 1 0 12032 0 -1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap0_7
timestamp 1607194124
transform 1 0 11648 0 -1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap0_7
timestamp 1607194124
transform 1 0 11552 0 -1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap1_8
timestamp 1607194124
transform 1 0 12896 0 1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap1_8
timestamp 1607194124
transform 1 0 12800 0 1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap0_8
timestamp 1607194124
transform 1 0 12896 0 -1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap0_8
timestamp 1607194124
transform 1 0 12800 0 -1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap1_9
timestamp 1607194124
transform 1 0 14144 0 1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap1_9
timestamp 1607194124
transform 1 0 14048 0 1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_23
timestamp 1607194124
transform 1 0 13280 0 1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap0_9
timestamp 1607194124
transform 1 0 14144 0 -1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap0_9
timestamp 1607194124
transform 1 0 14048 0 -1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_8
timestamp 1607194124
transform 1 0 13280 0 -1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_22
timestamp 1607194124
transform 1 0 14528 0 1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_9
timestamp 1607194124
transform 1 0 14528 0 -1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_21
timestamp 1607194124
transform 1 0 15776 0 1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap1_10
timestamp 1607194124
transform 1 0 15392 0 1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap1_10
timestamp 1607194124
transform 1 0 15296 0 1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_10
timestamp 1607194124
transform 1 0 15776 0 -1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap0_10
timestamp 1607194124
transform 1 0 15392 0 -1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap0_10
timestamp 1607194124
transform 1 0 15296 0 -1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap1_11
timestamp 1607194124
transform 1 0 16640 0 1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap1_11
timestamp 1607194124
transform 1 0 16544 0 1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap0_11
timestamp 1607194124
transform 1 0 16640 0 -1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap0_11
timestamp 1607194124
transform 1 0 16544 0 -1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap1_12
timestamp 1607194124
transform 1 0 17888 0 1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap1_12
timestamp 1607194124
transform 1 0 17792 0 1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_20
timestamp 1607194124
transform 1 0 17024 0 1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap0_12
timestamp 1607194124
transform 1 0 17888 0 -1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap0_12
timestamp 1607194124
transform 1 0 17792 0 -1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_11
timestamp 1607194124
transform 1 0 17024 0 -1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_19
timestamp 1607194124
transform 1 0 18272 0 1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_12
timestamp 1607194124
transform 1 0 18272 0 -1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_18
timestamp 1607194124
transform 1 0 19520 0 1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap1_13
timestamp 1607194124
transform 1 0 19136 0 1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap1_13
timestamp 1607194124
transform 1 0 19040 0 1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_13
timestamp 1607194124
transform 1 0 19520 0 -1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap0_13
timestamp 1607194124
transform 1 0 19136 0 -1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap0_13
timestamp 1607194124
transform 1 0 19040 0 -1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_17
timestamp 1607194124
transform 1 0 20768 0 1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap1_14
timestamp 1607194124
transform 1 0 20384 0 1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap1_14
timestamp 1607194124
transform 1 0 20288 0 1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_14
timestamp 1607194124
transform 1 0 20768 0 -1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap0_14
timestamp 1607194124
transform 1 0 20384 0 -1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap0_14
timestamp 1607194124
transform 1 0 20288 0 -1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap1_15
timestamp 1607194124
transform 1 0 21632 0 1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap1_15
timestamp 1607194124
transform 1 0 21536 0 1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap0_15
timestamp 1607194124
transform 1 0 21632 0 -1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap0_15
timestamp 1607194124
transform 1 0 21536 0 -1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_16
timestamp 1607194124
transform 1 0 22016 0 1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_15
timestamp 1607194124
transform 1 0 22016 0 -1 1726
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap1_16
timestamp 1607194124
transform 1 0 22880 0 1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap1_16
timestamp 1607194124
transform 1 0 22784 0 1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap0_16
timestamp 1607194124
transform 1 0 22880 0 -1 1726
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap0_16
timestamp 1607194124
transform 1 0 22784 0 -1 1726
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap2_0
timestamp 1607194124
transform 1 0 2816 0 -1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_5
timestamp 1607194124
transform 1 0 2048 0 -1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_4
timestamp 1607194124
transform 1 0 1952 0 -1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_32
timestamp 1607194124
transform 1 0 3296 0 -1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap2_0
timestamp 1607194124
transform 1 0 2912 0 -1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_33
timestamp 1607194124
transform 1 0 4544 0 -1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap2_1
timestamp 1607194124
transform 1 0 4160 0 -1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap2_1
timestamp 1607194124
transform 1 0 4064 0 -1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap2_2
timestamp 1607194124
transform 1 0 5408 0 -1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap2_2
timestamp 1607194124
transform 1 0 5312 0 -1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap2_3
timestamp 1607194124
transform 1 0 6656 0 -1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap2_3
timestamp 1607194124
transform 1 0 6560 0 -1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_34
timestamp 1607194124
transform 1 0 5792 0 -1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_35
timestamp 1607194124
transform 1 0 7040 0 -1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_36
timestamp 1607194124
transform 1 0 8288 0 -1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap2_4
timestamp 1607194124
transform 1 0 7904 0 -1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap2_4
timestamp 1607194124
transform 1 0 7808 0 -1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap2_5
timestamp 1607194124
transform 1 0 9152 0 -1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap2_5
timestamp 1607194124
transform 1 0 9056 0 -1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap2_6
timestamp 1607194124
transform 1 0 10400 0 -1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap2_6
timestamp 1607194124
transform 1 0 10304 0 -1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_37
timestamp 1607194124
transform 1 0 9536 0 -1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_38
timestamp 1607194124
transform 1 0 10784 0 -1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_39
timestamp 1607194124
transform 1 0 12032 0 -1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap2_7
timestamp 1607194124
transform 1 0 11648 0 -1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap2_7
timestamp 1607194124
transform 1 0 11552 0 -1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap2_8
timestamp 1607194124
transform 1 0 12896 0 -1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap2_8
timestamp 1607194124
transform 1 0 12800 0 -1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap2_9
timestamp 1607194124
transform 1 0 14144 0 -1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap2_9
timestamp 1607194124
transform 1 0 14048 0 -1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_40
timestamp 1607194124
transform 1 0 13280 0 -1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_41
timestamp 1607194124
transform 1 0 14528 0 -1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_42
timestamp 1607194124
transform 1 0 15776 0 -1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap2_10
timestamp 1607194124
transform 1 0 15392 0 -1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap2_10
timestamp 1607194124
transform 1 0 15296 0 -1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap2_11
timestamp 1607194124
transform 1 0 16640 0 -1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap2_11
timestamp 1607194124
transform 1 0 16544 0 -1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap2_12
timestamp 1607194124
transform 1 0 17888 0 -1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap2_12
timestamp 1607194124
transform 1 0 17792 0 -1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_43
timestamp 1607194124
transform 1 0 17024 0 -1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_44
timestamp 1607194124
transform 1 0 18272 0 -1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_45
timestamp 1607194124
transform 1 0 19520 0 -1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap2_13
timestamp 1607194124
transform 1 0 19136 0 -1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap2_13
timestamp 1607194124
transform 1 0 19040 0 -1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_46
timestamp 1607194124
transform 1 0 20768 0 -1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap2_14
timestamp 1607194124
transform 1 0 20384 0 -1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap2_14
timestamp 1607194124
transform 1 0 20288 0 -1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap2_15
timestamp 1607194124
transform 1 0 21632 0 -1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap2_15
timestamp 1607194124
transform 1 0 21536 0 -1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_47
timestamp 1607194124
transform 1 0 22016 0 -1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap2_16
timestamp 1607194124
transform 1 0 22880 0 -1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap2_16
timestamp 1607194124
transform 1 0 22784 0 -1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap3_0
timestamp 1607194124
transform 1 0 2816 0 1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_7
timestamp 1607194124
transform 1 0 2048 0 1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_6
timestamp 1607194124
transform 1 0 1952 0 1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_63
timestamp 1607194124
transform 1 0 3296 0 1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap3_0
timestamp 1607194124
transform 1 0 2912 0 1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_62
timestamp 1607194124
transform 1 0 4544 0 1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap3_1
timestamp 1607194124
transform 1 0 4160 0 1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap3_1
timestamp 1607194124
transform 1 0 4064 0 1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap3_2
timestamp 1607194124
transform 1 0 5408 0 1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap3_2
timestamp 1607194124
transform 1 0 5312 0 1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap3_3
timestamp 1607194124
transform 1 0 6656 0 1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap3_3
timestamp 1607194124
transform 1 0 6560 0 1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_61
timestamp 1607194124
transform 1 0 5792 0 1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_60
timestamp 1607194124
transform 1 0 7040 0 1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_59
timestamp 1607194124
transform 1 0 8288 0 1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap3_4
timestamp 1607194124
transform 1 0 7904 0 1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap3_4
timestamp 1607194124
transform 1 0 7808 0 1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap3_5
timestamp 1607194124
transform 1 0 9152 0 1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap3_5
timestamp 1607194124
transform 1 0 9056 0 1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap3_6
timestamp 1607194124
transform 1 0 10400 0 1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap3_6
timestamp 1607194124
transform 1 0 10304 0 1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_58
timestamp 1607194124
transform 1 0 9536 0 1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_57
timestamp 1607194124
transform 1 0 10784 0 1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_56
timestamp 1607194124
transform 1 0 12032 0 1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap3_7
timestamp 1607194124
transform 1 0 11648 0 1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap3_7
timestamp 1607194124
transform 1 0 11552 0 1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap3_8
timestamp 1607194124
transform 1 0 12896 0 1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap3_8
timestamp 1607194124
transform 1 0 12800 0 1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap3_9
timestamp 1607194124
transform 1 0 14144 0 1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap3_9
timestamp 1607194124
transform 1 0 14048 0 1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_55
timestamp 1607194124
transform 1 0 13280 0 1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_54
timestamp 1607194124
transform 1 0 14528 0 1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_53
timestamp 1607194124
transform 1 0 15776 0 1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap3_10
timestamp 1607194124
transform 1 0 15392 0 1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap3_10
timestamp 1607194124
transform 1 0 15296 0 1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap3_11
timestamp 1607194124
transform 1 0 16640 0 1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap3_11
timestamp 1607194124
transform 1 0 16544 0 1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap3_12
timestamp 1607194124
transform 1 0 17888 0 1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap3_12
timestamp 1607194124
transform 1 0 17792 0 1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_52
timestamp 1607194124
transform 1 0 17024 0 1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_51
timestamp 1607194124
transform 1 0 18272 0 1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_50
timestamp 1607194124
transform 1 0 19520 0 1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap3_13
timestamp 1607194124
transform 1 0 19136 0 1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap3_13
timestamp 1607194124
transform 1 0 19040 0 1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_49
timestamp 1607194124
transform 1 0 20768 0 1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap3_14
timestamp 1607194124
transform 1 0 20384 0 1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap3_14
timestamp 1607194124
transform 1 0 20288 0 1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap3_15
timestamp 1607194124
transform 1 0 21632 0 1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap3_15
timestamp 1607194124
transform 1 0 21536 0 1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_48
timestamp 1607194124
transform 1 0 22016 0 1 3058
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap3_16
timestamp 1607194124
transform 1 0 22880 0 1 3058
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap3_16
timestamp 1607194124
transform 1 0 22784 0 1 3058
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap4_0
timestamp 1607194124
transform 1 0 2816 0 -1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_9
timestamp 1607194124
transform 1 0 2048 0 -1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_8
timestamp 1607194124
transform 1 0 1952 0 -1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_64
timestamp 1607194124
transform 1 0 3296 0 -1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap4_0
timestamp 1607194124
transform 1 0 2912 0 -1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_65
timestamp 1607194124
transform 1 0 4544 0 -1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap4_1
timestamp 1607194124
transform 1 0 4160 0 -1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap4_1
timestamp 1607194124
transform 1 0 4064 0 -1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap4_2
timestamp 1607194124
transform 1 0 5408 0 -1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap4_2
timestamp 1607194124
transform 1 0 5312 0 -1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap4_3
timestamp 1607194124
transform 1 0 6656 0 -1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap4_3
timestamp 1607194124
transform 1 0 6560 0 -1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_66
timestamp 1607194124
transform 1 0 5792 0 -1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_67
timestamp 1607194124
transform 1 0 7040 0 -1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_68
timestamp 1607194124
transform 1 0 8288 0 -1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap4_4
timestamp 1607194124
transform 1 0 7904 0 -1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap4_4
timestamp 1607194124
transform 1 0 7808 0 -1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap4_5
timestamp 1607194124
transform 1 0 9152 0 -1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap4_5
timestamp 1607194124
transform 1 0 9056 0 -1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap4_6
timestamp 1607194124
transform 1 0 10400 0 -1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap4_6
timestamp 1607194124
transform 1 0 10304 0 -1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_69
timestamp 1607194124
transform 1 0 9536 0 -1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_70
timestamp 1607194124
transform 1 0 10784 0 -1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_71
timestamp 1607194124
transform 1 0 12032 0 -1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap4_7
timestamp 1607194124
transform 1 0 11648 0 -1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap4_7
timestamp 1607194124
transform 1 0 11552 0 -1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap4_8
timestamp 1607194124
transform 1 0 12896 0 -1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap4_8
timestamp 1607194124
transform 1 0 12800 0 -1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap4_9
timestamp 1607194124
transform 1 0 14144 0 -1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap4_9
timestamp 1607194124
transform 1 0 14048 0 -1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_72
timestamp 1607194124
transform 1 0 13280 0 -1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_73
timestamp 1607194124
transform 1 0 14528 0 -1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_74
timestamp 1607194124
transform 1 0 15776 0 -1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap4_10
timestamp 1607194124
transform 1 0 15392 0 -1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap4_10
timestamp 1607194124
transform 1 0 15296 0 -1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap4_11
timestamp 1607194124
transform 1 0 16640 0 -1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap4_11
timestamp 1607194124
transform 1 0 16544 0 -1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap4_12
timestamp 1607194124
transform 1 0 17888 0 -1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap4_12
timestamp 1607194124
transform 1 0 17792 0 -1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_75
timestamp 1607194124
transform 1 0 17024 0 -1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_76
timestamp 1607194124
transform 1 0 18272 0 -1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_77
timestamp 1607194124
transform 1 0 19520 0 -1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap4_13
timestamp 1607194124
transform 1 0 19136 0 -1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap4_13
timestamp 1607194124
transform 1 0 19040 0 -1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_78
timestamp 1607194124
transform 1 0 20768 0 -1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap4_14
timestamp 1607194124
transform 1 0 20384 0 -1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap4_14
timestamp 1607194124
transform 1 0 20288 0 -1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap4_15
timestamp 1607194124
transform 1 0 21632 0 -1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap4_15
timestamp 1607194124
transform 1 0 21536 0 -1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_79
timestamp 1607194124
transform 1 0 22016 0 -1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap4_16
timestamp 1607194124
transform 1 0 22880 0 -1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap4_16
timestamp 1607194124
transform 1 0 22784 0 -1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap5_0
timestamp 1607194124
transform 1 0 2816 0 1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_11
timestamp 1607194124
transform 1 0 2048 0 1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_10
timestamp 1607194124
transform 1 0 1952 0 1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_95
timestamp 1607194124
transform 1 0 3296 0 1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap5_0
timestamp 1607194124
transform 1 0 2912 0 1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_94
timestamp 1607194124
transform 1 0 4544 0 1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap5_1
timestamp 1607194124
transform 1 0 4160 0 1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap5_1
timestamp 1607194124
transform 1 0 4064 0 1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap5_2
timestamp 1607194124
transform 1 0 5408 0 1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap5_2
timestamp 1607194124
transform 1 0 5312 0 1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap5_3
timestamp 1607194124
transform 1 0 6656 0 1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap5_3
timestamp 1607194124
transform 1 0 6560 0 1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_93
timestamp 1607194124
transform 1 0 5792 0 1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_92
timestamp 1607194124
transform 1 0 7040 0 1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_91
timestamp 1607194124
transform 1 0 8288 0 1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap5_4
timestamp 1607194124
transform 1 0 7904 0 1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap5_4
timestamp 1607194124
transform 1 0 7808 0 1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap5_5
timestamp 1607194124
transform 1 0 9152 0 1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap5_5
timestamp 1607194124
transform 1 0 9056 0 1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap5_6
timestamp 1607194124
transform 1 0 10400 0 1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap5_6
timestamp 1607194124
transform 1 0 10304 0 1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_90
timestamp 1607194124
transform 1 0 9536 0 1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_89
timestamp 1607194124
transform 1 0 10784 0 1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_88
timestamp 1607194124
transform 1 0 12032 0 1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap5_7
timestamp 1607194124
transform 1 0 11648 0 1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap5_7
timestamp 1607194124
transform 1 0 11552 0 1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap5_8
timestamp 1607194124
transform 1 0 12896 0 1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap5_8
timestamp 1607194124
transform 1 0 12800 0 1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap5_9
timestamp 1607194124
transform 1 0 14144 0 1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap5_9
timestamp 1607194124
transform 1 0 14048 0 1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_87
timestamp 1607194124
transform 1 0 13280 0 1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_86
timestamp 1607194124
transform 1 0 14528 0 1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_85
timestamp 1607194124
transform 1 0 15776 0 1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap5_10
timestamp 1607194124
transform 1 0 15392 0 1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap5_10
timestamp 1607194124
transform 1 0 15296 0 1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap5_11
timestamp 1607194124
transform 1 0 16640 0 1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap5_11
timestamp 1607194124
transform 1 0 16544 0 1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap5_12
timestamp 1607194124
transform 1 0 17888 0 1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap5_12
timestamp 1607194124
transform 1 0 17792 0 1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_84
timestamp 1607194124
transform 1 0 17024 0 1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_83
timestamp 1607194124
transform 1 0 18272 0 1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_82
timestamp 1607194124
transform 1 0 19520 0 1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap5_13
timestamp 1607194124
transform 1 0 19136 0 1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap5_13
timestamp 1607194124
transform 1 0 19040 0 1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_81
timestamp 1607194124
transform 1 0 20768 0 1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap5_14
timestamp 1607194124
transform 1 0 20384 0 1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap5_14
timestamp 1607194124
transform 1 0 20288 0 1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap5_15
timestamp 1607194124
transform 1 0 21632 0 1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap5_15
timestamp 1607194124
transform 1 0 21536 0 1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_80
timestamp 1607194124
transform 1 0 22016 0 1 4390
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap5_16
timestamp 1607194124
transform 1 0 22880 0 1 4390
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap5_16
timestamp 1607194124
transform 1 0 22784 0 1 4390
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap6_0
timestamp 1607194124
transform 1 0 2816 0 -1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_13
timestamp 1607194124
transform 1 0 2048 0 -1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_12
timestamp 1607194124
transform 1 0 1952 0 -1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_96
timestamp 1607194124
transform 1 0 3296 0 -1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap6_0
timestamp 1607194124
transform 1 0 2912 0 -1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_97
timestamp 1607194124
transform 1 0 4544 0 -1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap6_1
timestamp 1607194124
transform 1 0 4160 0 -1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap6_1
timestamp 1607194124
transform 1 0 4064 0 -1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap6_2
timestamp 1607194124
transform 1 0 5408 0 -1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap6_2
timestamp 1607194124
transform 1 0 5312 0 -1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap6_3
timestamp 1607194124
transform 1 0 6656 0 -1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap6_3
timestamp 1607194124
transform 1 0 6560 0 -1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_98
timestamp 1607194124
transform 1 0 5792 0 -1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_99
timestamp 1607194124
transform 1 0 7040 0 -1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_100
timestamp 1607194124
transform 1 0 8288 0 -1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap6_4
timestamp 1607194124
transform 1 0 7904 0 -1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap6_4
timestamp 1607194124
transform 1 0 7808 0 -1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap6_5
timestamp 1607194124
transform 1 0 9152 0 -1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap6_5
timestamp 1607194124
transform 1 0 9056 0 -1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap6_6
timestamp 1607194124
transform 1 0 10400 0 -1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap6_6
timestamp 1607194124
transform 1 0 10304 0 -1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_101
timestamp 1607194124
transform 1 0 9536 0 -1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_102
timestamp 1607194124
transform 1 0 10784 0 -1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_103
timestamp 1607194124
transform 1 0 12032 0 -1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap6_7
timestamp 1607194124
transform 1 0 11648 0 -1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap6_7
timestamp 1607194124
transform 1 0 11552 0 -1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap6_8
timestamp 1607194124
transform 1 0 12896 0 -1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap6_8
timestamp 1607194124
transform 1 0 12800 0 -1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap6_9
timestamp 1607194124
transform 1 0 14144 0 -1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap6_9
timestamp 1607194124
transform 1 0 14048 0 -1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_104
timestamp 1607194124
transform 1 0 13280 0 -1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_105
timestamp 1607194124
transform 1 0 14528 0 -1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_106
timestamp 1607194124
transform 1 0 15776 0 -1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap6_10
timestamp 1607194124
transform 1 0 15392 0 -1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap6_10
timestamp 1607194124
transform 1 0 15296 0 -1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap6_11
timestamp 1607194124
transform 1 0 16640 0 -1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap6_11
timestamp 1607194124
transform 1 0 16544 0 -1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap6_12
timestamp 1607194124
transform 1 0 17888 0 -1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap6_12
timestamp 1607194124
transform 1 0 17792 0 -1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_107
timestamp 1607194124
transform 1 0 17024 0 -1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_108
timestamp 1607194124
transform 1 0 18272 0 -1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_109
timestamp 1607194124
transform 1 0 19520 0 -1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap6_13
timestamp 1607194124
transform 1 0 19136 0 -1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap6_13
timestamp 1607194124
transform 1 0 19040 0 -1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_110
timestamp 1607194124
transform 1 0 20768 0 -1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap6_14
timestamp 1607194124
transform 1 0 20384 0 -1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap6_14
timestamp 1607194124
transform 1 0 20288 0 -1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap6_15
timestamp 1607194124
transform 1 0 21632 0 -1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap6_15
timestamp 1607194124
transform 1 0 21536 0 -1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_111
timestamp 1607194124
transform 1 0 22016 0 -1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap6_16
timestamp 1607194124
transform 1 0 22880 0 -1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap6_16
timestamp 1607194124
transform 1 0 22784 0 -1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap8_0
timestamp 1607194124
transform 1 0 2816 0 -1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_17
timestamp 1607194124
transform 1 0 2048 0 -1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_16
timestamp 1607194124
transform 1 0 1952 0 -1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap7_0
timestamp 1607194124
transform 1 0 2816 0 1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_15
timestamp 1607194124
transform 1 0 2048 0 1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_14
timestamp 1607194124
transform 1 0 1952 0 1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_128
timestamp 1607194124
transform 1 0 3296 0 -1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap8_0
timestamp 1607194124
transform 1 0 2912 0 -1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_127
timestamp 1607194124
transform 1 0 3296 0 1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap7_0
timestamp 1607194124
transform 1 0 2912 0 1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_129
timestamp 1607194124
transform 1 0 4544 0 -1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap8_1
timestamp 1607194124
transform 1 0 4160 0 -1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap8_1
timestamp 1607194124
transform 1 0 4064 0 -1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_126
timestamp 1607194124
transform 1 0 4544 0 1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap7_1
timestamp 1607194124
transform 1 0 4160 0 1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap7_1
timestamp 1607194124
transform 1 0 4064 0 1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap8_2
timestamp 1607194124
transform 1 0 5408 0 -1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap8_2
timestamp 1607194124
transform 1 0 5312 0 -1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap7_2
timestamp 1607194124
transform 1 0 5408 0 1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap7_2
timestamp 1607194124
transform 1 0 5312 0 1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap8_3
timestamp 1607194124
transform 1 0 6656 0 -1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap8_3
timestamp 1607194124
transform 1 0 6560 0 -1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_130
timestamp 1607194124
transform 1 0 5792 0 -1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap7_3
timestamp 1607194124
transform 1 0 6656 0 1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap7_3
timestamp 1607194124
transform 1 0 6560 0 1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_125
timestamp 1607194124
transform 1 0 5792 0 1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_131
timestamp 1607194124
transform 1 0 7040 0 -1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_124
timestamp 1607194124
transform 1 0 7040 0 1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_132
timestamp 1607194124
transform 1 0 8288 0 -1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap8_4
timestamp 1607194124
transform 1 0 7904 0 -1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap8_4
timestamp 1607194124
transform 1 0 7808 0 -1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_123
timestamp 1607194124
transform 1 0 8288 0 1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap7_4
timestamp 1607194124
transform 1 0 7904 0 1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap7_4
timestamp 1607194124
transform 1 0 7808 0 1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap8_5
timestamp 1607194124
transform 1 0 9152 0 -1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap8_5
timestamp 1607194124
transform 1 0 9056 0 -1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap7_5
timestamp 1607194124
transform 1 0 9152 0 1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap7_5
timestamp 1607194124
transform 1 0 9056 0 1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap8_6
timestamp 1607194124
transform 1 0 10400 0 -1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap8_6
timestamp 1607194124
transform 1 0 10304 0 -1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_133
timestamp 1607194124
transform 1 0 9536 0 -1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap7_6
timestamp 1607194124
transform 1 0 10400 0 1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap7_6
timestamp 1607194124
transform 1 0 10304 0 1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_122
timestamp 1607194124
transform 1 0 9536 0 1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_134
timestamp 1607194124
transform 1 0 10784 0 -1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_121
timestamp 1607194124
transform 1 0 10784 0 1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_135
timestamp 1607194124
transform 1 0 12032 0 -1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap8_7
timestamp 1607194124
transform 1 0 11648 0 -1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap8_7
timestamp 1607194124
transform 1 0 11552 0 -1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_120
timestamp 1607194124
transform 1 0 12032 0 1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap7_7
timestamp 1607194124
transform 1 0 11648 0 1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap7_7
timestamp 1607194124
transform 1 0 11552 0 1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap8_8
timestamp 1607194124
transform 1 0 12896 0 -1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap8_8
timestamp 1607194124
transform 1 0 12800 0 -1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap7_8
timestamp 1607194124
transform 1 0 12896 0 1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap7_8
timestamp 1607194124
transform 1 0 12800 0 1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap8_9
timestamp 1607194124
transform 1 0 14144 0 -1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap8_9
timestamp 1607194124
transform 1 0 14048 0 -1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_136
timestamp 1607194124
transform 1 0 13280 0 -1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap7_9
timestamp 1607194124
transform 1 0 14144 0 1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap7_9
timestamp 1607194124
transform 1 0 14048 0 1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_119
timestamp 1607194124
transform 1 0 13280 0 1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_137
timestamp 1607194124
transform 1 0 14528 0 -1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_118
timestamp 1607194124
transform 1 0 14528 0 1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_138
timestamp 1607194124
transform 1 0 15776 0 -1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap8_10
timestamp 1607194124
transform 1 0 15392 0 -1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap8_10
timestamp 1607194124
transform 1 0 15296 0 -1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_117
timestamp 1607194124
transform 1 0 15776 0 1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap7_10
timestamp 1607194124
transform 1 0 15392 0 1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap7_10
timestamp 1607194124
transform 1 0 15296 0 1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap8_11
timestamp 1607194124
transform 1 0 16640 0 -1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap8_11
timestamp 1607194124
transform 1 0 16544 0 -1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap7_11
timestamp 1607194124
transform 1 0 16640 0 1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap7_11
timestamp 1607194124
transform 1 0 16544 0 1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap8_12
timestamp 1607194124
transform 1 0 17888 0 -1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap8_12
timestamp 1607194124
transform 1 0 17792 0 -1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_139
timestamp 1607194124
transform 1 0 17024 0 -1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap7_12
timestamp 1607194124
transform 1 0 17888 0 1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap7_12
timestamp 1607194124
transform 1 0 17792 0 1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_116
timestamp 1607194124
transform 1 0 17024 0 1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_140
timestamp 1607194124
transform 1 0 18272 0 -1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_115
timestamp 1607194124
transform 1 0 18272 0 1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_141
timestamp 1607194124
transform 1 0 19520 0 -1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap8_13
timestamp 1607194124
transform 1 0 19136 0 -1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap8_13
timestamp 1607194124
transform 1 0 19040 0 -1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_114
timestamp 1607194124
transform 1 0 19520 0 1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap7_13
timestamp 1607194124
transform 1 0 19136 0 1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap7_13
timestamp 1607194124
transform 1 0 19040 0 1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_142
timestamp 1607194124
transform 1 0 20768 0 -1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap8_14
timestamp 1607194124
transform 1 0 20384 0 -1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap8_14
timestamp 1607194124
transform 1 0 20288 0 -1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_113
timestamp 1607194124
transform 1 0 20768 0 1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap7_14
timestamp 1607194124
transform 1 0 20384 0 1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap7_14
timestamp 1607194124
transform 1 0 20288 0 1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap8_15
timestamp 1607194124
transform 1 0 21632 0 -1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap8_15
timestamp 1607194124
transform 1 0 21536 0 -1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap7_15
timestamp 1607194124
transform 1 0 21632 0 1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap7_15
timestamp 1607194124
transform 1 0 21536 0 1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_143
timestamp 1607194124
transform 1 0 22016 0 -1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_112
timestamp 1607194124
transform 1 0 22016 0 1 5722
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap8_16
timestamp 1607194124
transform 1 0 22880 0 -1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap8_16
timestamp 1607194124
transform 1 0 22784 0 -1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap7_16
timestamp 1607194124
transform 1 0 22880 0 1 5722
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap7_16
timestamp 1607194124
transform 1 0 22784 0 1 5722
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap9_0
timestamp 1607194124
transform 1 0 2816 0 1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_19
timestamp 1607194124
transform 1 0 2048 0 1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_18
timestamp 1607194124
transform 1 0 1952 0 1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_159
timestamp 1607194124
transform 1 0 3296 0 1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap9_0
timestamp 1607194124
transform 1 0 2912 0 1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_158
timestamp 1607194124
transform 1 0 4544 0 1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap9_1
timestamp 1607194124
transform 1 0 4160 0 1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap9_1
timestamp 1607194124
transform 1 0 4064 0 1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap9_2
timestamp 1607194124
transform 1 0 5408 0 1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap9_2
timestamp 1607194124
transform 1 0 5312 0 1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap9_3
timestamp 1607194124
transform 1 0 6656 0 1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap9_3
timestamp 1607194124
transform 1 0 6560 0 1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_157
timestamp 1607194124
transform 1 0 5792 0 1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_156
timestamp 1607194124
transform 1 0 7040 0 1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_155
timestamp 1607194124
transform 1 0 8288 0 1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap9_4
timestamp 1607194124
transform 1 0 7904 0 1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap9_4
timestamp 1607194124
transform 1 0 7808 0 1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap9_5
timestamp 1607194124
transform 1 0 9152 0 1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap9_5
timestamp 1607194124
transform 1 0 9056 0 1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap9_6
timestamp 1607194124
transform 1 0 10400 0 1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap9_6
timestamp 1607194124
transform 1 0 10304 0 1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_154
timestamp 1607194124
transform 1 0 9536 0 1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_153
timestamp 1607194124
transform 1 0 10784 0 1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_152
timestamp 1607194124
transform 1 0 12032 0 1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap9_7
timestamp 1607194124
transform 1 0 11648 0 1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap9_7
timestamp 1607194124
transform 1 0 11552 0 1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap9_8
timestamp 1607194124
transform 1 0 12896 0 1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap9_8
timestamp 1607194124
transform 1 0 12800 0 1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap9_9
timestamp 1607194124
transform 1 0 14144 0 1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap9_9
timestamp 1607194124
transform 1 0 14048 0 1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_151
timestamp 1607194124
transform 1 0 13280 0 1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_150
timestamp 1607194124
transform 1 0 14528 0 1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_149
timestamp 1607194124
transform 1 0 15776 0 1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap9_10
timestamp 1607194124
transform 1 0 15392 0 1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap9_10
timestamp 1607194124
transform 1 0 15296 0 1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap9_11
timestamp 1607194124
transform 1 0 16640 0 1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap9_11
timestamp 1607194124
transform 1 0 16544 0 1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap9_12
timestamp 1607194124
transform 1 0 17888 0 1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap9_12
timestamp 1607194124
transform 1 0 17792 0 1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_148
timestamp 1607194124
transform 1 0 17024 0 1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_147
timestamp 1607194124
transform 1 0 18272 0 1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_146
timestamp 1607194124
transform 1 0 19520 0 1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap9_13
timestamp 1607194124
transform 1 0 19136 0 1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap9_13
timestamp 1607194124
transform 1 0 19040 0 1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_145
timestamp 1607194124
transform 1 0 20768 0 1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap9_14
timestamp 1607194124
transform 1 0 20384 0 1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap9_14
timestamp 1607194124
transform 1 0 20288 0 1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap9_15
timestamp 1607194124
transform 1 0 21632 0 1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap9_15
timestamp 1607194124
transform 1 0 21536 0 1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_144
timestamp 1607194124
transform 1 0 22016 0 1 7054
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap9_16
timestamp 1607194124
transform 1 0 22880 0 1 7054
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap9_16
timestamp 1607194124
transform 1 0 22784 0 1 7054
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap10_0
timestamp 1607194124
transform 1 0 2816 0 -1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_21
timestamp 1607194124
transform 1 0 2048 0 -1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_20
timestamp 1607194124
transform 1 0 1952 0 -1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_160
timestamp 1607194124
transform 1 0 3296 0 -1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap10_0
timestamp 1607194124
transform 1 0 2912 0 -1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_161
timestamp 1607194124
transform 1 0 4544 0 -1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap10_1
timestamp 1607194124
transform 1 0 4160 0 -1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap10_1
timestamp 1607194124
transform 1 0 4064 0 -1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap10_2
timestamp 1607194124
transform 1 0 5408 0 -1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap10_2
timestamp 1607194124
transform 1 0 5312 0 -1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap10_3
timestamp 1607194124
transform 1 0 6656 0 -1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap10_3
timestamp 1607194124
transform 1 0 6560 0 -1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_162
timestamp 1607194124
transform 1 0 5792 0 -1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_163
timestamp 1607194124
transform 1 0 7040 0 -1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_164
timestamp 1607194124
transform 1 0 8288 0 -1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap10_4
timestamp 1607194124
transform 1 0 7904 0 -1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap10_4
timestamp 1607194124
transform 1 0 7808 0 -1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap10_5
timestamp 1607194124
transform 1 0 9152 0 -1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap10_5
timestamp 1607194124
transform 1 0 9056 0 -1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap10_6
timestamp 1607194124
transform 1 0 10400 0 -1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap10_6
timestamp 1607194124
transform 1 0 10304 0 -1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_165
timestamp 1607194124
transform 1 0 9536 0 -1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_166
timestamp 1607194124
transform 1 0 10784 0 -1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_167
timestamp 1607194124
transform 1 0 12032 0 -1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap10_7
timestamp 1607194124
transform 1 0 11648 0 -1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap10_7
timestamp 1607194124
transform 1 0 11552 0 -1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap10_8
timestamp 1607194124
transform 1 0 12896 0 -1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap10_8
timestamp 1607194124
transform 1 0 12800 0 -1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap10_9
timestamp 1607194124
transform 1 0 14144 0 -1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap10_9
timestamp 1607194124
transform 1 0 14048 0 -1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_168
timestamp 1607194124
transform 1 0 13280 0 -1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_169
timestamp 1607194124
transform 1 0 14528 0 -1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_170
timestamp 1607194124
transform 1 0 15776 0 -1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap10_10
timestamp 1607194124
transform 1 0 15392 0 -1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap10_10
timestamp 1607194124
transform 1 0 15296 0 -1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap10_11
timestamp 1607194124
transform 1 0 16640 0 -1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap10_11
timestamp 1607194124
transform 1 0 16544 0 -1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap10_12
timestamp 1607194124
transform 1 0 17888 0 -1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap10_12
timestamp 1607194124
transform 1 0 17792 0 -1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_171
timestamp 1607194124
transform 1 0 17024 0 -1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_172
timestamp 1607194124
transform 1 0 18272 0 -1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_173
timestamp 1607194124
transform 1 0 19520 0 -1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap10_13
timestamp 1607194124
transform 1 0 19136 0 -1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap10_13
timestamp 1607194124
transform 1 0 19040 0 -1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_174
timestamp 1607194124
transform 1 0 20768 0 -1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap10_14
timestamp 1607194124
transform 1 0 20384 0 -1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap10_14
timestamp 1607194124
transform 1 0 20288 0 -1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap10_15
timestamp 1607194124
transform 1 0 21632 0 -1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap10_15
timestamp 1607194124
transform 1 0 21536 0 -1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_175
timestamp 1607194124
transform 1 0 22016 0 -1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap10_16
timestamp 1607194124
transform 1 0 22880 0 -1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap10_16
timestamp 1607194124
transform 1 0 22784 0 -1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap11_0
timestamp 1607194124
transform 1 0 2816 0 1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_23
timestamp 1607194124
transform 1 0 2048 0 1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_22
timestamp 1607194124
transform 1 0 1952 0 1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_191
timestamp 1607194124
transform 1 0 3296 0 1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap11_0
timestamp 1607194124
transform 1 0 2912 0 1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_190
timestamp 1607194124
transform 1 0 4544 0 1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap11_1
timestamp 1607194124
transform 1 0 4160 0 1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap11_1
timestamp 1607194124
transform 1 0 4064 0 1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap11_2
timestamp 1607194124
transform 1 0 5408 0 1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap11_2
timestamp 1607194124
transform 1 0 5312 0 1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap11_3
timestamp 1607194124
transform 1 0 6656 0 1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap11_3
timestamp 1607194124
transform 1 0 6560 0 1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_189
timestamp 1607194124
transform 1 0 5792 0 1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_188
timestamp 1607194124
transform 1 0 7040 0 1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_187
timestamp 1607194124
transform 1 0 8288 0 1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap11_4
timestamp 1607194124
transform 1 0 7904 0 1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap11_4
timestamp 1607194124
transform 1 0 7808 0 1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap11_5
timestamp 1607194124
transform 1 0 9152 0 1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap11_5
timestamp 1607194124
transform 1 0 9056 0 1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap11_6
timestamp 1607194124
transform 1 0 10400 0 1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap11_6
timestamp 1607194124
transform 1 0 10304 0 1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_186
timestamp 1607194124
transform 1 0 9536 0 1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_185
timestamp 1607194124
transform 1 0 10784 0 1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_184
timestamp 1607194124
transform 1 0 12032 0 1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap11_7
timestamp 1607194124
transform 1 0 11648 0 1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap11_7
timestamp 1607194124
transform 1 0 11552 0 1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap11_8
timestamp 1607194124
transform 1 0 12896 0 1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap11_8
timestamp 1607194124
transform 1 0 12800 0 1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap11_9
timestamp 1607194124
transform 1 0 14144 0 1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap11_9
timestamp 1607194124
transform 1 0 14048 0 1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_183
timestamp 1607194124
transform 1 0 13280 0 1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_182
timestamp 1607194124
transform 1 0 14528 0 1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_181
timestamp 1607194124
transform 1 0 15776 0 1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap11_10
timestamp 1607194124
transform 1 0 15392 0 1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap11_10
timestamp 1607194124
transform 1 0 15296 0 1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap11_11
timestamp 1607194124
transform 1 0 16640 0 1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap11_11
timestamp 1607194124
transform 1 0 16544 0 1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap11_12
timestamp 1607194124
transform 1 0 17888 0 1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap11_12
timestamp 1607194124
transform 1 0 17792 0 1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_180
timestamp 1607194124
transform 1 0 17024 0 1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_179
timestamp 1607194124
transform 1 0 18272 0 1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_178
timestamp 1607194124
transform 1 0 19520 0 1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap11_13
timestamp 1607194124
transform 1 0 19136 0 1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap11_13
timestamp 1607194124
transform 1 0 19040 0 1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_177
timestamp 1607194124
transform 1 0 20768 0 1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap11_14
timestamp 1607194124
transform 1 0 20384 0 1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap11_14
timestamp 1607194124
transform 1 0 20288 0 1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap11_15
timestamp 1607194124
transform 1 0 21632 0 1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap11_15
timestamp 1607194124
transform 1 0 21536 0 1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_176
timestamp 1607194124
transform 1 0 22016 0 1 8386
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap11_16
timestamp 1607194124
transform 1 0 22880 0 1 8386
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap11_16
timestamp 1607194124
transform 1 0 22784 0 1 8386
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap12_0
timestamp 1607194124
transform 1 0 2816 0 -1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_25
timestamp 1607194124
transform 1 0 2048 0 -1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_24
timestamp 1607194124
transform 1 0 1952 0 -1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_192
timestamp 1607194124
transform 1 0 3296 0 -1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap12_0
timestamp 1607194124
transform 1 0 2912 0 -1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_193
timestamp 1607194124
transform 1 0 4544 0 -1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap12_1
timestamp 1607194124
transform 1 0 4160 0 -1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap12_1
timestamp 1607194124
transform 1 0 4064 0 -1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap12_2
timestamp 1607194124
transform 1 0 5408 0 -1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap12_2
timestamp 1607194124
transform 1 0 5312 0 -1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap12_3
timestamp 1607194124
transform 1 0 6656 0 -1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap12_3
timestamp 1607194124
transform 1 0 6560 0 -1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_194
timestamp 1607194124
transform 1 0 5792 0 -1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_195
timestamp 1607194124
transform 1 0 7040 0 -1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_196
timestamp 1607194124
transform 1 0 8288 0 -1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap12_4
timestamp 1607194124
transform 1 0 7904 0 -1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap12_4
timestamp 1607194124
transform 1 0 7808 0 -1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap12_5
timestamp 1607194124
transform 1 0 9152 0 -1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap12_5
timestamp 1607194124
transform 1 0 9056 0 -1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap12_6
timestamp 1607194124
transform 1 0 10400 0 -1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap12_6
timestamp 1607194124
transform 1 0 10304 0 -1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_197
timestamp 1607194124
transform 1 0 9536 0 -1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_198
timestamp 1607194124
transform 1 0 10784 0 -1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_199
timestamp 1607194124
transform 1 0 12032 0 -1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap12_7
timestamp 1607194124
transform 1 0 11648 0 -1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap12_7
timestamp 1607194124
transform 1 0 11552 0 -1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap12_8
timestamp 1607194124
transform 1 0 12896 0 -1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap12_8
timestamp 1607194124
transform 1 0 12800 0 -1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap12_9
timestamp 1607194124
transform 1 0 14144 0 -1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap12_9
timestamp 1607194124
transform 1 0 14048 0 -1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_200
timestamp 1607194124
transform 1 0 13280 0 -1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_201
timestamp 1607194124
transform 1 0 14528 0 -1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_202
timestamp 1607194124
transform 1 0 15776 0 -1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap12_10
timestamp 1607194124
transform 1 0 15392 0 -1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap12_10
timestamp 1607194124
transform 1 0 15296 0 -1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap12_11
timestamp 1607194124
transform 1 0 16640 0 -1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap12_11
timestamp 1607194124
transform 1 0 16544 0 -1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap12_12
timestamp 1607194124
transform 1 0 17888 0 -1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap12_12
timestamp 1607194124
transform 1 0 17792 0 -1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_203
timestamp 1607194124
transform 1 0 17024 0 -1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_204
timestamp 1607194124
transform 1 0 18272 0 -1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_205
timestamp 1607194124
transform 1 0 19520 0 -1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap12_13
timestamp 1607194124
transform 1 0 19136 0 -1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap12_13
timestamp 1607194124
transform 1 0 19040 0 -1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_206
timestamp 1607194124
transform 1 0 20768 0 -1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap12_14
timestamp 1607194124
transform 1 0 20384 0 -1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap12_14
timestamp 1607194124
transform 1 0 20288 0 -1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap12_15
timestamp 1607194124
transform 1 0 21632 0 -1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap12_15
timestamp 1607194124
transform 1 0 21536 0 -1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_207
timestamp 1607194124
transform 1 0 22016 0 -1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap12_16
timestamp 1607194124
transform 1 0 22880 0 -1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap12_16
timestamp 1607194124
transform 1 0 22784 0 -1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap13_0
timestamp 1607194124
transform 1 0 2816 0 1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_27
timestamp 1607194124
transform 1 0 2048 0 1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_26
timestamp 1607194124
transform 1 0 1952 0 1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_223
timestamp 1607194124
transform 1 0 3296 0 1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap13_0
timestamp 1607194124
transform 1 0 2912 0 1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_222
timestamp 1607194124
transform 1 0 4544 0 1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap13_1
timestamp 1607194124
transform 1 0 4160 0 1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap13_1
timestamp 1607194124
transform 1 0 4064 0 1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap13_2
timestamp 1607194124
transform 1 0 5408 0 1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap13_2
timestamp 1607194124
transform 1 0 5312 0 1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap13_3
timestamp 1607194124
transform 1 0 6656 0 1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap13_3
timestamp 1607194124
transform 1 0 6560 0 1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_221
timestamp 1607194124
transform 1 0 5792 0 1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_220
timestamp 1607194124
transform 1 0 7040 0 1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_219
timestamp 1607194124
transform 1 0 8288 0 1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap13_4
timestamp 1607194124
transform 1 0 7904 0 1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap13_4
timestamp 1607194124
transform 1 0 7808 0 1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap13_5
timestamp 1607194124
transform 1 0 9152 0 1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap13_5
timestamp 1607194124
transform 1 0 9056 0 1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap13_6
timestamp 1607194124
transform 1 0 10400 0 1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap13_6
timestamp 1607194124
transform 1 0 10304 0 1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_218
timestamp 1607194124
transform 1 0 9536 0 1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_217
timestamp 1607194124
transform 1 0 10784 0 1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_216
timestamp 1607194124
transform 1 0 12032 0 1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap13_7
timestamp 1607194124
transform 1 0 11648 0 1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap13_7
timestamp 1607194124
transform 1 0 11552 0 1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap13_8
timestamp 1607194124
transform 1 0 12896 0 1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap13_8
timestamp 1607194124
transform 1 0 12800 0 1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap13_9
timestamp 1607194124
transform 1 0 14144 0 1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap13_9
timestamp 1607194124
transform 1 0 14048 0 1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_215
timestamp 1607194124
transform 1 0 13280 0 1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_214
timestamp 1607194124
transform 1 0 14528 0 1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_213
timestamp 1607194124
transform 1 0 15776 0 1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap13_10
timestamp 1607194124
transform 1 0 15392 0 1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap13_10
timestamp 1607194124
transform 1 0 15296 0 1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap13_11
timestamp 1607194124
transform 1 0 16640 0 1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap13_11
timestamp 1607194124
transform 1 0 16544 0 1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap13_12
timestamp 1607194124
transform 1 0 17888 0 1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap13_12
timestamp 1607194124
transform 1 0 17792 0 1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_212
timestamp 1607194124
transform 1 0 17024 0 1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_211
timestamp 1607194124
transform 1 0 18272 0 1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_210
timestamp 1607194124
transform 1 0 19520 0 1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap13_13
timestamp 1607194124
transform 1 0 19136 0 1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap13_13
timestamp 1607194124
transform 1 0 19040 0 1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_209
timestamp 1607194124
transform 1 0 20768 0 1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap13_14
timestamp 1607194124
transform 1 0 20384 0 1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap13_14
timestamp 1607194124
transform 1 0 20288 0 1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap13_15
timestamp 1607194124
transform 1 0 21632 0 1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap13_15
timestamp 1607194124
transform 1 0 21536 0 1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_208
timestamp 1607194124
transform 1 0 22016 0 1 9718
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap13_16
timestamp 1607194124
transform 1 0 22880 0 1 9718
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap13_16
timestamp 1607194124
transform 1 0 22784 0 1 9718
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap14_0
timestamp 1607194124
transform 1 0 2816 0 -1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_29
timestamp 1607194124
transform 1 0 2048 0 -1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_28
timestamp 1607194124
transform 1 0 1952 0 -1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_224
timestamp 1607194124
transform 1 0 3296 0 -1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap14_0
timestamp 1607194124
transform 1 0 2912 0 -1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_225
timestamp 1607194124
transform 1 0 4544 0 -1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap14_1
timestamp 1607194124
transform 1 0 4160 0 -1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap14_1
timestamp 1607194124
transform 1 0 4064 0 -1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap14_2
timestamp 1607194124
transform 1 0 5408 0 -1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap14_2
timestamp 1607194124
transform 1 0 5312 0 -1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap14_3
timestamp 1607194124
transform 1 0 6656 0 -1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap14_3
timestamp 1607194124
transform 1 0 6560 0 -1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_226
timestamp 1607194124
transform 1 0 5792 0 -1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_227
timestamp 1607194124
transform 1 0 7040 0 -1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_228
timestamp 1607194124
transform 1 0 8288 0 -1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap14_4
timestamp 1607194124
transform 1 0 7904 0 -1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap14_4
timestamp 1607194124
transform 1 0 7808 0 -1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap14_5
timestamp 1607194124
transform 1 0 9152 0 -1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap14_5
timestamp 1607194124
transform 1 0 9056 0 -1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap14_6
timestamp 1607194124
transform 1 0 10400 0 -1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap14_6
timestamp 1607194124
transform 1 0 10304 0 -1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_229
timestamp 1607194124
transform 1 0 9536 0 -1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_230
timestamp 1607194124
transform 1 0 10784 0 -1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_231
timestamp 1607194124
transform 1 0 12032 0 -1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap14_7
timestamp 1607194124
transform 1 0 11648 0 -1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap14_7
timestamp 1607194124
transform 1 0 11552 0 -1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap14_8
timestamp 1607194124
transform 1 0 12896 0 -1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap14_8
timestamp 1607194124
transform 1 0 12800 0 -1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap14_9
timestamp 1607194124
transform 1 0 14144 0 -1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap14_9
timestamp 1607194124
transform 1 0 14048 0 -1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_232
timestamp 1607194124
transform 1 0 13280 0 -1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_233
timestamp 1607194124
transform 1 0 14528 0 -1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_234
timestamp 1607194124
transform 1 0 15776 0 -1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap14_10
timestamp 1607194124
transform 1 0 15392 0 -1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap14_10
timestamp 1607194124
transform 1 0 15296 0 -1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap14_11
timestamp 1607194124
transform 1 0 16640 0 -1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap14_11
timestamp 1607194124
transform 1 0 16544 0 -1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap14_12
timestamp 1607194124
transform 1 0 17888 0 -1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap14_12
timestamp 1607194124
transform 1 0 17792 0 -1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_235
timestamp 1607194124
transform 1 0 17024 0 -1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_236
timestamp 1607194124
transform 1 0 18272 0 -1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_237
timestamp 1607194124
transform 1 0 19520 0 -1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap14_13
timestamp 1607194124
transform 1 0 19136 0 -1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap14_13
timestamp 1607194124
transform 1 0 19040 0 -1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_238
timestamp 1607194124
transform 1 0 20768 0 -1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap14_14
timestamp 1607194124
transform 1 0 20384 0 -1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap14_14
timestamp 1607194124
transform 1 0 20288 0 -1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap14_15
timestamp 1607194124
transform 1 0 21632 0 -1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap14_15
timestamp 1607194124
transform 1 0 21536 0 -1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_239
timestamp 1607194124
transform 1 0 22016 0 -1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap14_16
timestamp 1607194124
transform 1 0 22880 0 -1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap14_16
timestamp 1607194124
transform 1 0 22784 0 -1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap16_0
timestamp 1607194124
transform 1 0 2816 0 -1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_31
timestamp 1607194124
transform 1 0 2048 0 -1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_30
timestamp 1607194124
transform 1 0 1952 0 -1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap15_0
timestamp 1607194124
transform 1 0 2816 0 1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__mux2_1  mux_8 $PDKPATH/libs.ref/sky130_fd_sc_ms/mag
timestamp 1607194124
transform 1 0 1952 0 1 11050
box -38 -49 902 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_0
timestamp 1607194124
transform 1 0 3296 0 -1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap16_0
timestamp 1607194124
transform 1 0 2912 0 -1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_255
timestamp 1607194124
transform 1 0 3296 0 1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap15_0
timestamp 1607194124
transform 1 0 2912 0 1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_1
timestamp 1607194124
transform 1 0 4544 0 -1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap16_1
timestamp 1607194124
transform 1 0 4160 0 -1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap16_1
timestamp 1607194124
transform 1 0 4064 0 -1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_254
timestamp 1607194124
transform 1 0 4544 0 1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap15_1
timestamp 1607194124
transform 1 0 4160 0 1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap15_1
timestamp 1607194124
transform 1 0 4064 0 1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap16_2
timestamp 1607194124
transform 1 0 5408 0 -1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap16_2
timestamp 1607194124
transform 1 0 5312 0 -1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap15_2
timestamp 1607194124
transform 1 0 5408 0 1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap15_2
timestamp 1607194124
transform 1 0 5312 0 1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap16_3
timestamp 1607194124
transform 1 0 6656 0 -1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap16_3
timestamp 1607194124
transform 1 0 6560 0 -1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_2
timestamp 1607194124
transform 1 0 5792 0 -1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap15_3
timestamp 1607194124
transform 1 0 6656 0 1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap15_3
timestamp 1607194124
transform 1 0 6560 0 1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_253
timestamp 1607194124
transform 1 0 5792 0 1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_3
timestamp 1607194124
transform 1 0 7040 0 -1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_252
timestamp 1607194124
transform 1 0 7040 0 1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_4
timestamp 1607194124
transform 1 0 8288 0 -1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap16_4
timestamp 1607194124
transform 1 0 7904 0 -1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap16_4
timestamp 1607194124
transform 1 0 7808 0 -1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_251
timestamp 1607194124
transform 1 0 8288 0 1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap15_4
timestamp 1607194124
transform 1 0 7904 0 1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap15_4
timestamp 1607194124
transform 1 0 7808 0 1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap16_5
timestamp 1607194124
transform 1 0 9152 0 -1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap16_5
timestamp 1607194124
transform 1 0 9056 0 -1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap15_5
timestamp 1607194124
transform 1 0 9152 0 1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap15_5
timestamp 1607194124
transform 1 0 9056 0 1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap16_6
timestamp 1607194124
transform 1 0 10400 0 -1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap16_6
timestamp 1607194124
transform 1 0 10304 0 -1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_5
timestamp 1607194124
transform 1 0 9536 0 -1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap15_6
timestamp 1607194124
transform 1 0 10400 0 1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap15_6
timestamp 1607194124
transform 1 0 10304 0 1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_250
timestamp 1607194124
transform 1 0 9536 0 1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_6
timestamp 1607194124
transform 1 0 10784 0 -1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_249
timestamp 1607194124
transform 1 0 10784 0 1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_7
timestamp 1607194124
transform 1 0 12032 0 -1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap16_7
timestamp 1607194124
transform 1 0 11648 0 -1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap16_7
timestamp 1607194124
transform 1 0 11552 0 -1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_248
timestamp 1607194124
transform 1 0 12032 0 1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap15_7
timestamp 1607194124
transform 1 0 11648 0 1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap15_7
timestamp 1607194124
transform 1 0 11552 0 1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap16_8
timestamp 1607194124
transform 1 0 12896 0 -1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap16_8
timestamp 1607194124
transform 1 0 12800 0 -1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap15_8
timestamp 1607194124
transform 1 0 12896 0 1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap15_8
timestamp 1607194124
transform 1 0 12800 0 1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap16_9
timestamp 1607194124
transform 1 0 14144 0 -1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap16_9
timestamp 1607194124
transform 1 0 14048 0 -1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_8
timestamp 1607194124
transform 1 0 13280 0 -1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap15_9
timestamp 1607194124
transform 1 0 14144 0 1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap15_9
timestamp 1607194124
transform 1 0 14048 0 1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_247
timestamp 1607194124
transform 1 0 13280 0 1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_9
timestamp 1607194124
transform 1 0 14528 0 -1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_246
timestamp 1607194124
transform 1 0 14528 0 1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_10
timestamp 1607194124
transform 1 0 15776 0 -1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap16_10
timestamp 1607194124
transform 1 0 15392 0 -1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap16_10
timestamp 1607194124
transform 1 0 15296 0 -1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_245
timestamp 1607194124
transform 1 0 15776 0 1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap15_10
timestamp 1607194124
transform 1 0 15392 0 1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap15_10
timestamp 1607194124
transform 1 0 15296 0 1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap16_11
timestamp 1607194124
transform 1 0 16640 0 -1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap16_11
timestamp 1607194124
transform 1 0 16544 0 -1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap15_11
timestamp 1607194124
transform 1 0 16640 0 1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap15_11
timestamp 1607194124
transform 1 0 16544 0 1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap16_12
timestamp 1607194124
transform 1 0 17888 0 -1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap16_12
timestamp 1607194124
transform 1 0 17792 0 -1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_11
timestamp 1607194124
transform 1 0 17024 0 -1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap15_12
timestamp 1607194124
transform 1 0 17888 0 1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap15_12
timestamp 1607194124
transform 1 0 17792 0 1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_244
timestamp 1607194124
transform 1 0 17024 0 1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_12
timestamp 1607194124
transform 1 0 18272 0 -1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_243
timestamp 1607194124
transform 1 0 18272 0 1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_13
timestamp 1607194124
transform 1 0 19520 0 -1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap16_13
timestamp 1607194124
transform 1 0 19136 0 -1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap16_13
timestamp 1607194124
transform 1 0 19040 0 -1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_242
timestamp 1607194124
transform 1 0 19520 0 1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap15_13
timestamp 1607194124
transform 1 0 19136 0 1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap15_13
timestamp 1607194124
transform 1 0 19040 0 1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_14
timestamp 1607194124
transform 1 0 20768 0 -1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap16_14
timestamp 1607194124
transform 1 0 20384 0 -1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap16_14
timestamp 1607194124
transform 1 0 20288 0 -1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_241
timestamp 1607194124
transform 1 0 20768 0 1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap15_14
timestamp 1607194124
transform 1 0 20384 0 1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap15_14
timestamp 1607194124
transform 1 0 20288 0 1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap16_15
timestamp 1607194124
transform 1 0 21632 0 -1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap16_15
timestamp 1607194124
transform 1 0 21536 0 -1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap15_15
timestamp 1607194124
transform 1 0 21632 0 1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap15_15
timestamp 1607194124
transform 1 0 21536 0 1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_15
timestamp 1607194124
transform 1 0 22016 0 -1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_8_240
timestamp 1607194124
transform 1 0 22016 0 1 11050
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap16_16
timestamp 1607194124
transform 1 0 22880 0 -1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap16_16
timestamp 1607194124
transform 1 0 22784 0 -1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap15_16
timestamp 1607194124
transform 1 0 22880 0 1 11050
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap15_16
timestamp 1607194124
transform 1 0 22784 0 1 11050
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap17_0
timestamp 1607194124
transform 1 0 2816 0 1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_33
timestamp 1607194124
transform 1 0 2048 0 1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_32
timestamp 1607194124
transform 1 0 1952 0 1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_31
timestamp 1607194124
transform 1 0 3296 0 1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap17_0
timestamp 1607194124
transform 1 0 2912 0 1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_30
timestamp 1607194124
transform 1 0 4544 0 1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap17_1
timestamp 1607194124
transform 1 0 4160 0 1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap17_1
timestamp 1607194124
transform 1 0 4064 0 1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap17_2
timestamp 1607194124
transform 1 0 5408 0 1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap17_2
timestamp 1607194124
transform 1 0 5312 0 1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap17_3
timestamp 1607194124
transform 1 0 6656 0 1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap17_3
timestamp 1607194124
transform 1 0 6560 0 1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_29
timestamp 1607194124
transform 1 0 5792 0 1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_28
timestamp 1607194124
transform 1 0 7040 0 1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_27
timestamp 1607194124
transform 1 0 8288 0 1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap17_4
timestamp 1607194124
transform 1 0 7904 0 1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap17_4
timestamp 1607194124
transform 1 0 7808 0 1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap17_5
timestamp 1607194124
transform 1 0 9152 0 1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap17_5
timestamp 1607194124
transform 1 0 9056 0 1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap17_6
timestamp 1607194124
transform 1 0 10400 0 1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap17_6
timestamp 1607194124
transform 1 0 10304 0 1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_26
timestamp 1607194124
transform 1 0 9536 0 1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_25
timestamp 1607194124
transform 1 0 10784 0 1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_24
timestamp 1607194124
transform 1 0 12032 0 1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap17_7
timestamp 1607194124
transform 1 0 11648 0 1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap17_7
timestamp 1607194124
transform 1 0 11552 0 1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap17_8
timestamp 1607194124
transform 1 0 12896 0 1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap17_8
timestamp 1607194124
transform 1 0 12800 0 1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap17_9
timestamp 1607194124
transform 1 0 14144 0 1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap17_9
timestamp 1607194124
transform 1 0 14048 0 1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_23
timestamp 1607194124
transform 1 0 13280 0 1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_22
timestamp 1607194124
transform 1 0 14528 0 1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_21
timestamp 1607194124
transform 1 0 15776 0 1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap17_10
timestamp 1607194124
transform 1 0 15392 0 1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap17_10
timestamp 1607194124
transform 1 0 15296 0 1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap17_11
timestamp 1607194124
transform 1 0 16640 0 1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap17_11
timestamp 1607194124
transform 1 0 16544 0 1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap17_12
timestamp 1607194124
transform 1 0 17888 0 1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap17_12
timestamp 1607194124
transform 1 0 17792 0 1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_20
timestamp 1607194124
transform 1 0 17024 0 1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_19
timestamp 1607194124
transform 1 0 18272 0 1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_18
timestamp 1607194124
transform 1 0 19520 0 1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap17_13
timestamp 1607194124
transform 1 0 19136 0 1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap17_13
timestamp 1607194124
transform 1 0 19040 0 1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_17
timestamp 1607194124
transform 1 0 20768 0 1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap17_14
timestamp 1607194124
transform 1 0 20384 0 1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap17_14
timestamp 1607194124
transform 1 0 20288 0 1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap17_15
timestamp 1607194124
transform 1 0 21632 0 1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap17_15
timestamp 1607194124
transform 1 0 21536 0 1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_16
timestamp 1607194124
transform 1 0 22016 0 1 12382
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap17_16
timestamp 1607194124
transform 1 0 22880 0 1 12382
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap17_16
timestamp 1607194124
transform 1 0 22784 0 1 12382
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap18_0
timestamp 1607194124
transform 1 0 2816 0 -1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_35
timestamp 1607194124
transform 1 0 2048 0 -1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_34
timestamp 1607194124
transform 1 0 1952 0 -1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_32
timestamp 1607194124
transform 1 0 3296 0 -1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap18_0
timestamp 1607194124
transform 1 0 2912 0 -1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_33
timestamp 1607194124
transform 1 0 4544 0 -1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap18_1
timestamp 1607194124
transform 1 0 4160 0 -1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap18_1
timestamp 1607194124
transform 1 0 4064 0 -1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap18_2
timestamp 1607194124
transform 1 0 5408 0 -1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap18_2
timestamp 1607194124
transform 1 0 5312 0 -1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap18_3
timestamp 1607194124
transform 1 0 6656 0 -1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap18_3
timestamp 1607194124
transform 1 0 6560 0 -1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_34
timestamp 1607194124
transform 1 0 5792 0 -1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_35
timestamp 1607194124
transform 1 0 7040 0 -1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_36
timestamp 1607194124
transform 1 0 8288 0 -1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap18_4
timestamp 1607194124
transform 1 0 7904 0 -1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap18_4
timestamp 1607194124
transform 1 0 7808 0 -1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap18_5
timestamp 1607194124
transform 1 0 9152 0 -1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap18_5
timestamp 1607194124
transform 1 0 9056 0 -1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap18_6
timestamp 1607194124
transform 1 0 10400 0 -1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap18_6
timestamp 1607194124
transform 1 0 10304 0 -1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_37
timestamp 1607194124
transform 1 0 9536 0 -1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_38
timestamp 1607194124
transform 1 0 10784 0 -1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_39
timestamp 1607194124
transform 1 0 12032 0 -1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap18_7
timestamp 1607194124
transform 1 0 11648 0 -1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap18_7
timestamp 1607194124
transform 1 0 11552 0 -1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap18_8
timestamp 1607194124
transform 1 0 12896 0 -1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap18_8
timestamp 1607194124
transform 1 0 12800 0 -1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap18_9
timestamp 1607194124
transform 1 0 14144 0 -1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap18_9
timestamp 1607194124
transform 1 0 14048 0 -1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_40
timestamp 1607194124
transform 1 0 13280 0 -1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_41
timestamp 1607194124
transform 1 0 14528 0 -1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_42
timestamp 1607194124
transform 1 0 15776 0 -1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap18_10
timestamp 1607194124
transform 1 0 15392 0 -1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap18_10
timestamp 1607194124
transform 1 0 15296 0 -1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap18_11
timestamp 1607194124
transform 1 0 16640 0 -1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap18_11
timestamp 1607194124
transform 1 0 16544 0 -1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap18_12
timestamp 1607194124
transform 1 0 17888 0 -1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap18_12
timestamp 1607194124
transform 1 0 17792 0 -1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_43
timestamp 1607194124
transform 1 0 17024 0 -1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_44
timestamp 1607194124
transform 1 0 18272 0 -1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_45
timestamp 1607194124
transform 1 0 19520 0 -1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap18_13
timestamp 1607194124
transform 1 0 19136 0 -1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap18_13
timestamp 1607194124
transform 1 0 19040 0 -1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_46
timestamp 1607194124
transform 1 0 20768 0 -1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap18_14
timestamp 1607194124
transform 1 0 20384 0 -1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap18_14
timestamp 1607194124
transform 1 0 20288 0 -1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap18_15
timestamp 1607194124
transform 1 0 21632 0 -1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap18_15
timestamp 1607194124
transform 1 0 21536 0 -1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_47
timestamp 1607194124
transform 1 0 22016 0 -1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap18_16
timestamp 1607194124
transform 1 0 22880 0 -1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap18_16
timestamp 1607194124
transform 1 0 22784 0 -1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap19_0
timestamp 1607194124
transform 1 0 2816 0 1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_37
timestamp 1607194124
transform 1 0 2048 0 1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_36
timestamp 1607194124
transform 1 0 1952 0 1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_63
timestamp 1607194124
transform 1 0 3296 0 1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap19_0
timestamp 1607194124
transform 1 0 2912 0 1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_62
timestamp 1607194124
transform 1 0 4544 0 1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap19_1
timestamp 1607194124
transform 1 0 4160 0 1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap19_1
timestamp 1607194124
transform 1 0 4064 0 1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap19_2
timestamp 1607194124
transform 1 0 5408 0 1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap19_2
timestamp 1607194124
transform 1 0 5312 0 1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap19_3
timestamp 1607194124
transform 1 0 6656 0 1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap19_3
timestamp 1607194124
transform 1 0 6560 0 1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_61
timestamp 1607194124
transform 1 0 5792 0 1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_60
timestamp 1607194124
transform 1 0 7040 0 1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_59
timestamp 1607194124
transform 1 0 8288 0 1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap19_4
timestamp 1607194124
transform 1 0 7904 0 1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap19_4
timestamp 1607194124
transform 1 0 7808 0 1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap19_5
timestamp 1607194124
transform 1 0 9152 0 1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap19_5
timestamp 1607194124
transform 1 0 9056 0 1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap19_6
timestamp 1607194124
transform 1 0 10400 0 1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap19_6
timestamp 1607194124
transform 1 0 10304 0 1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_58
timestamp 1607194124
transform 1 0 9536 0 1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_57
timestamp 1607194124
transform 1 0 10784 0 1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_56
timestamp 1607194124
transform 1 0 12032 0 1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap19_7
timestamp 1607194124
transform 1 0 11648 0 1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap19_7
timestamp 1607194124
transform 1 0 11552 0 1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap19_8
timestamp 1607194124
transform 1 0 12896 0 1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap19_8
timestamp 1607194124
transform 1 0 12800 0 1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap19_9
timestamp 1607194124
transform 1 0 14144 0 1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap19_9
timestamp 1607194124
transform 1 0 14048 0 1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_55
timestamp 1607194124
transform 1 0 13280 0 1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_54
timestamp 1607194124
transform 1 0 14528 0 1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_53
timestamp 1607194124
transform 1 0 15776 0 1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap19_10
timestamp 1607194124
transform 1 0 15392 0 1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap19_10
timestamp 1607194124
transform 1 0 15296 0 1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap19_11
timestamp 1607194124
transform 1 0 16640 0 1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap19_11
timestamp 1607194124
transform 1 0 16544 0 1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap19_12
timestamp 1607194124
transform 1 0 17888 0 1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap19_12
timestamp 1607194124
transform 1 0 17792 0 1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_52
timestamp 1607194124
transform 1 0 17024 0 1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_51
timestamp 1607194124
transform 1 0 18272 0 1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_50
timestamp 1607194124
transform 1 0 19520 0 1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap19_13
timestamp 1607194124
transform 1 0 19136 0 1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap19_13
timestamp 1607194124
transform 1 0 19040 0 1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_49
timestamp 1607194124
transform 1 0 20768 0 1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap19_14
timestamp 1607194124
transform 1 0 20384 0 1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap19_14
timestamp 1607194124
transform 1 0 20288 0 1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap19_15
timestamp 1607194124
transform 1 0 21632 0 1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap19_15
timestamp 1607194124
transform 1 0 21536 0 1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_48
timestamp 1607194124
transform 1 0 22016 0 1 13714
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap19_16
timestamp 1607194124
transform 1 0 22880 0 1 13714
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap19_16
timestamp 1607194124
transform 1 0 22784 0 1 13714
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap20_0
timestamp 1607194124
transform 1 0 2816 0 -1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_39
timestamp 1607194124
transform 1 0 2048 0 -1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_38
timestamp 1607194124
transform 1 0 1952 0 -1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_64
timestamp 1607194124
transform 1 0 3296 0 -1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap20_0
timestamp 1607194124
transform 1 0 2912 0 -1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_65
timestamp 1607194124
transform 1 0 4544 0 -1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap20_1
timestamp 1607194124
transform 1 0 4160 0 -1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap20_1
timestamp 1607194124
transform 1 0 4064 0 -1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap20_2
timestamp 1607194124
transform 1 0 5408 0 -1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap20_2
timestamp 1607194124
transform 1 0 5312 0 -1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap20_3
timestamp 1607194124
transform 1 0 6656 0 -1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap20_3
timestamp 1607194124
transform 1 0 6560 0 -1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_66
timestamp 1607194124
transform 1 0 5792 0 -1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_67
timestamp 1607194124
transform 1 0 7040 0 -1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_68
timestamp 1607194124
transform 1 0 8288 0 -1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap20_4
timestamp 1607194124
transform 1 0 7904 0 -1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap20_4
timestamp 1607194124
transform 1 0 7808 0 -1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap20_5
timestamp 1607194124
transform 1 0 9152 0 -1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap20_5
timestamp 1607194124
transform 1 0 9056 0 -1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap20_6
timestamp 1607194124
transform 1 0 10400 0 -1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap20_6
timestamp 1607194124
transform 1 0 10304 0 -1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_69
timestamp 1607194124
transform 1 0 9536 0 -1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_70
timestamp 1607194124
transform 1 0 10784 0 -1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_71
timestamp 1607194124
transform 1 0 12032 0 -1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap20_7
timestamp 1607194124
transform 1 0 11648 0 -1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap20_7
timestamp 1607194124
transform 1 0 11552 0 -1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap20_8
timestamp 1607194124
transform 1 0 12896 0 -1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap20_8
timestamp 1607194124
transform 1 0 12800 0 -1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap20_9
timestamp 1607194124
transform 1 0 14144 0 -1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap20_9
timestamp 1607194124
transform 1 0 14048 0 -1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_72
timestamp 1607194124
transform 1 0 13280 0 -1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_73
timestamp 1607194124
transform 1 0 14528 0 -1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_74
timestamp 1607194124
transform 1 0 15776 0 -1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap20_10
timestamp 1607194124
transform 1 0 15392 0 -1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap20_10
timestamp 1607194124
transform 1 0 15296 0 -1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap20_11
timestamp 1607194124
transform 1 0 16640 0 -1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap20_11
timestamp 1607194124
transform 1 0 16544 0 -1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap20_12
timestamp 1607194124
transform 1 0 17888 0 -1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap20_12
timestamp 1607194124
transform 1 0 17792 0 -1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_75
timestamp 1607194124
transform 1 0 17024 0 -1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_76
timestamp 1607194124
transform 1 0 18272 0 -1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_77
timestamp 1607194124
transform 1 0 19520 0 -1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap20_13
timestamp 1607194124
transform 1 0 19136 0 -1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap20_13
timestamp 1607194124
transform 1 0 19040 0 -1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_78
timestamp 1607194124
transform 1 0 20768 0 -1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap20_14
timestamp 1607194124
transform 1 0 20384 0 -1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap20_14
timestamp 1607194124
transform 1 0 20288 0 -1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap20_15
timestamp 1607194124
transform 1 0 21632 0 -1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap20_15
timestamp 1607194124
transform 1 0 21536 0 -1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_79
timestamp 1607194124
transform 1 0 22016 0 -1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap20_16
timestamp 1607194124
transform 1 0 22880 0 -1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap20_16
timestamp 1607194124
transform 1 0 22784 0 -1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap21_0
timestamp 1607194124
transform 1 0 2816 0 1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_41
timestamp 1607194124
transform 1 0 2048 0 1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_40
timestamp 1607194124
transform 1 0 1952 0 1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_95
timestamp 1607194124
transform 1 0 3296 0 1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap21_0
timestamp 1607194124
transform 1 0 2912 0 1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_94
timestamp 1607194124
transform 1 0 4544 0 1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap21_1
timestamp 1607194124
transform 1 0 4160 0 1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap21_1
timestamp 1607194124
transform 1 0 4064 0 1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap21_2
timestamp 1607194124
transform 1 0 5408 0 1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap21_2
timestamp 1607194124
transform 1 0 5312 0 1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap21_3
timestamp 1607194124
transform 1 0 6656 0 1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap21_3
timestamp 1607194124
transform 1 0 6560 0 1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_93
timestamp 1607194124
transform 1 0 5792 0 1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_92
timestamp 1607194124
transform 1 0 7040 0 1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_91
timestamp 1607194124
transform 1 0 8288 0 1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap21_4
timestamp 1607194124
transform 1 0 7904 0 1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap21_4
timestamp 1607194124
transform 1 0 7808 0 1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap21_5
timestamp 1607194124
transform 1 0 9152 0 1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap21_5
timestamp 1607194124
transform 1 0 9056 0 1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap21_6
timestamp 1607194124
transform 1 0 10400 0 1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap21_6
timestamp 1607194124
transform 1 0 10304 0 1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_90
timestamp 1607194124
transform 1 0 9536 0 1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_89
timestamp 1607194124
transform 1 0 10784 0 1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_88
timestamp 1607194124
transform 1 0 12032 0 1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap21_7
timestamp 1607194124
transform 1 0 11648 0 1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap21_7
timestamp 1607194124
transform 1 0 11552 0 1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap21_8
timestamp 1607194124
transform 1 0 12896 0 1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap21_8
timestamp 1607194124
transform 1 0 12800 0 1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap21_9
timestamp 1607194124
transform 1 0 14144 0 1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap21_9
timestamp 1607194124
transform 1 0 14048 0 1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_87
timestamp 1607194124
transform 1 0 13280 0 1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_86
timestamp 1607194124
transform 1 0 14528 0 1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_85
timestamp 1607194124
transform 1 0 15776 0 1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap21_10
timestamp 1607194124
transform 1 0 15392 0 1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap21_10
timestamp 1607194124
transform 1 0 15296 0 1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap21_11
timestamp 1607194124
transform 1 0 16640 0 1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap21_11
timestamp 1607194124
transform 1 0 16544 0 1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap21_12
timestamp 1607194124
transform 1 0 17888 0 1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap21_12
timestamp 1607194124
transform 1 0 17792 0 1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_84
timestamp 1607194124
transform 1 0 17024 0 1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_83
timestamp 1607194124
transform 1 0 18272 0 1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_82
timestamp 1607194124
transform 1 0 19520 0 1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap21_13
timestamp 1607194124
transform 1 0 19136 0 1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap21_13
timestamp 1607194124
transform 1 0 19040 0 1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_81
timestamp 1607194124
transform 1 0 20768 0 1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap21_14
timestamp 1607194124
transform 1 0 20384 0 1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap21_14
timestamp 1607194124
transform 1 0 20288 0 1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap21_15
timestamp 1607194124
transform 1 0 21632 0 1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap21_15
timestamp 1607194124
transform 1 0 21536 0 1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_80
timestamp 1607194124
transform 1 0 22016 0 1 15046
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap21_16
timestamp 1607194124
transform 1 0 22880 0 1 15046
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap21_16
timestamp 1607194124
transform 1 0 22784 0 1 15046
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap22_0
timestamp 1607194124
transform 1 0 2816 0 -1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_43
timestamp 1607194124
transform 1 0 2048 0 -1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_42
timestamp 1607194124
transform 1 0 1952 0 -1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_96
timestamp 1607194124
transform 1 0 3296 0 -1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap22_0
timestamp 1607194124
transform 1 0 2912 0 -1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_97
timestamp 1607194124
transform 1 0 4544 0 -1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap22_1
timestamp 1607194124
transform 1 0 4160 0 -1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap22_1
timestamp 1607194124
transform 1 0 4064 0 -1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap22_2
timestamp 1607194124
transform 1 0 5408 0 -1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap22_2
timestamp 1607194124
transform 1 0 5312 0 -1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap22_3
timestamp 1607194124
transform 1 0 6656 0 -1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap22_3
timestamp 1607194124
transform 1 0 6560 0 -1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_98
timestamp 1607194124
transform 1 0 5792 0 -1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_99
timestamp 1607194124
transform 1 0 7040 0 -1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_100
timestamp 1607194124
transform 1 0 8288 0 -1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap22_4
timestamp 1607194124
transform 1 0 7904 0 -1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap22_4
timestamp 1607194124
transform 1 0 7808 0 -1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap22_5
timestamp 1607194124
transform 1 0 9152 0 -1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap22_5
timestamp 1607194124
transform 1 0 9056 0 -1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap22_6
timestamp 1607194124
transform 1 0 10400 0 -1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap22_6
timestamp 1607194124
transform 1 0 10304 0 -1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_101
timestamp 1607194124
transform 1 0 9536 0 -1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_102
timestamp 1607194124
transform 1 0 10784 0 -1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_103
timestamp 1607194124
transform 1 0 12032 0 -1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap22_7
timestamp 1607194124
transform 1 0 11648 0 -1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap22_7
timestamp 1607194124
transform 1 0 11552 0 -1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap22_8
timestamp 1607194124
transform 1 0 12896 0 -1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap22_8
timestamp 1607194124
transform 1 0 12800 0 -1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap22_9
timestamp 1607194124
transform 1 0 14144 0 -1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap22_9
timestamp 1607194124
transform 1 0 14048 0 -1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_104
timestamp 1607194124
transform 1 0 13280 0 -1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_105
timestamp 1607194124
transform 1 0 14528 0 -1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_106
timestamp 1607194124
transform 1 0 15776 0 -1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap22_10
timestamp 1607194124
transform 1 0 15392 0 -1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap22_10
timestamp 1607194124
transform 1 0 15296 0 -1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap22_11
timestamp 1607194124
transform 1 0 16640 0 -1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap22_11
timestamp 1607194124
transform 1 0 16544 0 -1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap22_12
timestamp 1607194124
transform 1 0 17888 0 -1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap22_12
timestamp 1607194124
transform 1 0 17792 0 -1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_107
timestamp 1607194124
transform 1 0 17024 0 -1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_108
timestamp 1607194124
transform 1 0 18272 0 -1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_109
timestamp 1607194124
transform 1 0 19520 0 -1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap22_13
timestamp 1607194124
transform 1 0 19136 0 -1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap22_13
timestamp 1607194124
transform 1 0 19040 0 -1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_110
timestamp 1607194124
transform 1 0 20768 0 -1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap22_14
timestamp 1607194124
transform 1 0 20384 0 -1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap22_14
timestamp 1607194124
transform 1 0 20288 0 -1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap22_15
timestamp 1607194124
transform 1 0 21632 0 -1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap22_15
timestamp 1607194124
transform 1 0 21536 0 -1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_111
timestamp 1607194124
transform 1 0 22016 0 -1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap22_16
timestamp 1607194124
transform 1 0 22880 0 -1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap22_16
timestamp 1607194124
transform 1 0 22784 0 -1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap24_0
timestamp 1607194124
transform 1 0 2816 0 -1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_45
timestamp 1607194124
transform 1 0 2048 0 -1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_44
timestamp 1607194124
transform 1 0 1952 0 -1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap23_0
timestamp 1607194124
transform 1 0 2816 0 1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__mux2_1  mux_7
timestamp 1607194124
transform 1 0 1952 0 1 16378
box -38 -49 902 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_0
timestamp 1607194124
transform 1 0 3296 0 -1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap24_0
timestamp 1607194124
transform 1 0 2912 0 -1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_127
timestamp 1607194124
transform 1 0 3296 0 1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap23_0
timestamp 1607194124
transform 1 0 2912 0 1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_1
timestamp 1607194124
transform 1 0 4544 0 -1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap24_1
timestamp 1607194124
transform 1 0 4160 0 -1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap24_1
timestamp 1607194124
transform 1 0 4064 0 -1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_126
timestamp 1607194124
transform 1 0 4544 0 1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap23_1
timestamp 1607194124
transform 1 0 4160 0 1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap23_1
timestamp 1607194124
transform 1 0 4064 0 1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap24_2
timestamp 1607194124
transform 1 0 5408 0 -1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap24_2
timestamp 1607194124
transform 1 0 5312 0 -1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap23_2
timestamp 1607194124
transform 1 0 5408 0 1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap23_2
timestamp 1607194124
transform 1 0 5312 0 1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap24_3
timestamp 1607194124
transform 1 0 6656 0 -1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap24_3
timestamp 1607194124
transform 1 0 6560 0 -1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_2
timestamp 1607194124
transform 1 0 5792 0 -1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap23_3
timestamp 1607194124
transform 1 0 6656 0 1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap23_3
timestamp 1607194124
transform 1 0 6560 0 1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_125
timestamp 1607194124
transform 1 0 5792 0 1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_3
timestamp 1607194124
transform 1 0 7040 0 -1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_124
timestamp 1607194124
transform 1 0 7040 0 1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_4
timestamp 1607194124
transform 1 0 8288 0 -1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap24_4
timestamp 1607194124
transform 1 0 7904 0 -1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap24_4
timestamp 1607194124
transform 1 0 7808 0 -1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_123
timestamp 1607194124
transform 1 0 8288 0 1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap23_4
timestamp 1607194124
transform 1 0 7904 0 1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap23_4
timestamp 1607194124
transform 1 0 7808 0 1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap24_5
timestamp 1607194124
transform 1 0 9152 0 -1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap24_5
timestamp 1607194124
transform 1 0 9056 0 -1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap23_5
timestamp 1607194124
transform 1 0 9152 0 1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap23_5
timestamp 1607194124
transform 1 0 9056 0 1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap24_6
timestamp 1607194124
transform 1 0 10400 0 -1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap24_6
timestamp 1607194124
transform 1 0 10304 0 -1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_5
timestamp 1607194124
transform 1 0 9536 0 -1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap23_6
timestamp 1607194124
transform 1 0 10400 0 1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap23_6
timestamp 1607194124
transform 1 0 10304 0 1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_122
timestamp 1607194124
transform 1 0 9536 0 1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_6
timestamp 1607194124
transform 1 0 10784 0 -1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_121
timestamp 1607194124
transform 1 0 10784 0 1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_7
timestamp 1607194124
transform 1 0 12032 0 -1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap24_7
timestamp 1607194124
transform 1 0 11648 0 -1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap24_7
timestamp 1607194124
transform 1 0 11552 0 -1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_120
timestamp 1607194124
transform 1 0 12032 0 1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap23_7
timestamp 1607194124
transform 1 0 11648 0 1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap23_7
timestamp 1607194124
transform 1 0 11552 0 1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap24_8
timestamp 1607194124
transform 1 0 12896 0 -1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap24_8
timestamp 1607194124
transform 1 0 12800 0 -1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap23_8
timestamp 1607194124
transform 1 0 12896 0 1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap23_8
timestamp 1607194124
transform 1 0 12800 0 1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap24_9
timestamp 1607194124
transform 1 0 14144 0 -1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap24_9
timestamp 1607194124
transform 1 0 14048 0 -1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_8
timestamp 1607194124
transform 1 0 13280 0 -1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap23_9
timestamp 1607194124
transform 1 0 14144 0 1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap23_9
timestamp 1607194124
transform 1 0 14048 0 1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_119
timestamp 1607194124
transform 1 0 13280 0 1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_9
timestamp 1607194124
transform 1 0 14528 0 -1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_118
timestamp 1607194124
transform 1 0 14528 0 1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_10
timestamp 1607194124
transform 1 0 15776 0 -1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap24_10
timestamp 1607194124
transform 1 0 15392 0 -1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap24_10
timestamp 1607194124
transform 1 0 15296 0 -1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_117
timestamp 1607194124
transform 1 0 15776 0 1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap23_10
timestamp 1607194124
transform 1 0 15392 0 1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap23_10
timestamp 1607194124
transform 1 0 15296 0 1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap24_11
timestamp 1607194124
transform 1 0 16640 0 -1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap24_11
timestamp 1607194124
transform 1 0 16544 0 -1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap23_11
timestamp 1607194124
transform 1 0 16640 0 1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap23_11
timestamp 1607194124
transform 1 0 16544 0 1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap24_12
timestamp 1607194124
transform 1 0 17888 0 -1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap24_12
timestamp 1607194124
transform 1 0 17792 0 -1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_11
timestamp 1607194124
transform 1 0 17024 0 -1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap23_12
timestamp 1607194124
transform 1 0 17888 0 1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap23_12
timestamp 1607194124
transform 1 0 17792 0 1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_116
timestamp 1607194124
transform 1 0 17024 0 1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_12
timestamp 1607194124
transform 1 0 18272 0 -1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_115
timestamp 1607194124
transform 1 0 18272 0 1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_13
timestamp 1607194124
transform 1 0 19520 0 -1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap24_13
timestamp 1607194124
transform 1 0 19136 0 -1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap24_13
timestamp 1607194124
transform 1 0 19040 0 -1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_114
timestamp 1607194124
transform 1 0 19520 0 1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap23_13
timestamp 1607194124
transform 1 0 19136 0 1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap23_13
timestamp 1607194124
transform 1 0 19040 0 1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_14
timestamp 1607194124
transform 1 0 20768 0 -1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap24_14
timestamp 1607194124
transform 1 0 20384 0 -1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap24_14
timestamp 1607194124
transform 1 0 20288 0 -1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_113
timestamp 1607194124
transform 1 0 20768 0 1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap23_14
timestamp 1607194124
transform 1 0 20384 0 1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap23_14
timestamp 1607194124
transform 1 0 20288 0 1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap24_15
timestamp 1607194124
transform 1 0 21632 0 -1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap24_15
timestamp 1607194124
transform 1 0 21536 0 -1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap23_15
timestamp 1607194124
transform 1 0 21632 0 1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap23_15
timestamp 1607194124
transform 1 0 21536 0 1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_15
timestamp 1607194124
transform 1 0 22016 0 -1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_7_112
timestamp 1607194124
transform 1 0 22016 0 1 16378
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap24_16
timestamp 1607194124
transform 1 0 22880 0 -1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap24_16
timestamp 1607194124
transform 1 0 22784 0 -1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap23_16
timestamp 1607194124
transform 1 0 22880 0 1 16378
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap23_16
timestamp 1607194124
transform 1 0 22784 0 1 16378
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap25_0
timestamp 1607194124
transform 1 0 2816 0 1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_47
timestamp 1607194124
transform 1 0 2048 0 1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_46
timestamp 1607194124
transform 1 0 1952 0 1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_31
timestamp 1607194124
transform 1 0 3296 0 1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap25_0
timestamp 1607194124
transform 1 0 2912 0 1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_30
timestamp 1607194124
transform 1 0 4544 0 1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap25_1
timestamp 1607194124
transform 1 0 4160 0 1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap25_1
timestamp 1607194124
transform 1 0 4064 0 1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap25_2
timestamp 1607194124
transform 1 0 5408 0 1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap25_2
timestamp 1607194124
transform 1 0 5312 0 1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap25_3
timestamp 1607194124
transform 1 0 6656 0 1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap25_3
timestamp 1607194124
transform 1 0 6560 0 1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_29
timestamp 1607194124
transform 1 0 5792 0 1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_28
timestamp 1607194124
transform 1 0 7040 0 1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_27
timestamp 1607194124
transform 1 0 8288 0 1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap25_4
timestamp 1607194124
transform 1 0 7904 0 1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap25_4
timestamp 1607194124
transform 1 0 7808 0 1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap25_5
timestamp 1607194124
transform 1 0 9152 0 1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap25_5
timestamp 1607194124
transform 1 0 9056 0 1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap25_6
timestamp 1607194124
transform 1 0 10400 0 1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap25_6
timestamp 1607194124
transform 1 0 10304 0 1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_26
timestamp 1607194124
transform 1 0 9536 0 1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_25
timestamp 1607194124
transform 1 0 10784 0 1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_24
timestamp 1607194124
transform 1 0 12032 0 1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap25_7
timestamp 1607194124
transform 1 0 11648 0 1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap25_7
timestamp 1607194124
transform 1 0 11552 0 1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap25_8
timestamp 1607194124
transform 1 0 12896 0 1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap25_8
timestamp 1607194124
transform 1 0 12800 0 1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap25_9
timestamp 1607194124
transform 1 0 14144 0 1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap25_9
timestamp 1607194124
transform 1 0 14048 0 1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_23
timestamp 1607194124
transform 1 0 13280 0 1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_22
timestamp 1607194124
transform 1 0 14528 0 1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_21
timestamp 1607194124
transform 1 0 15776 0 1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap25_10
timestamp 1607194124
transform 1 0 15392 0 1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap25_10
timestamp 1607194124
transform 1 0 15296 0 1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap25_11
timestamp 1607194124
transform 1 0 16640 0 1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap25_11
timestamp 1607194124
transform 1 0 16544 0 1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap25_12
timestamp 1607194124
transform 1 0 17888 0 1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap25_12
timestamp 1607194124
transform 1 0 17792 0 1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_20
timestamp 1607194124
transform 1 0 17024 0 1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_19
timestamp 1607194124
transform 1 0 18272 0 1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_18
timestamp 1607194124
transform 1 0 19520 0 1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap25_13
timestamp 1607194124
transform 1 0 19136 0 1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap25_13
timestamp 1607194124
transform 1 0 19040 0 1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_17
timestamp 1607194124
transform 1 0 20768 0 1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap25_14
timestamp 1607194124
transform 1 0 20384 0 1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap25_14
timestamp 1607194124
transform 1 0 20288 0 1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap25_15
timestamp 1607194124
transform 1 0 21632 0 1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap25_15
timestamp 1607194124
transform 1 0 21536 0 1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_16
timestamp 1607194124
transform 1 0 22016 0 1 17710
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap25_16
timestamp 1607194124
transform 1 0 22880 0 1 17710
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap25_16
timestamp 1607194124
transform 1 0 22784 0 1 17710
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap26_0
timestamp 1607194124
transform 1 0 2816 0 -1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_49
timestamp 1607194124
transform 1 0 2048 0 -1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_48
timestamp 1607194124
transform 1 0 1952 0 -1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_32
timestamp 1607194124
transform 1 0 3296 0 -1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap26_0
timestamp 1607194124
transform 1 0 2912 0 -1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_33
timestamp 1607194124
transform 1 0 4544 0 -1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap26_1
timestamp 1607194124
transform 1 0 4160 0 -1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap26_1
timestamp 1607194124
transform 1 0 4064 0 -1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap26_2
timestamp 1607194124
transform 1 0 5408 0 -1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap26_2
timestamp 1607194124
transform 1 0 5312 0 -1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap26_3
timestamp 1607194124
transform 1 0 6656 0 -1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap26_3
timestamp 1607194124
transform 1 0 6560 0 -1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_34
timestamp 1607194124
transform 1 0 5792 0 -1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_35
timestamp 1607194124
transform 1 0 7040 0 -1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_36
timestamp 1607194124
transform 1 0 8288 0 -1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap26_4
timestamp 1607194124
transform 1 0 7904 0 -1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap26_4
timestamp 1607194124
transform 1 0 7808 0 -1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap26_5
timestamp 1607194124
transform 1 0 9152 0 -1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap26_5
timestamp 1607194124
transform 1 0 9056 0 -1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap26_6
timestamp 1607194124
transform 1 0 10400 0 -1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap26_6
timestamp 1607194124
transform 1 0 10304 0 -1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_37
timestamp 1607194124
transform 1 0 9536 0 -1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_38
timestamp 1607194124
transform 1 0 10784 0 -1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_39
timestamp 1607194124
transform 1 0 12032 0 -1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap26_7
timestamp 1607194124
transform 1 0 11648 0 -1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap26_7
timestamp 1607194124
transform 1 0 11552 0 -1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap26_8
timestamp 1607194124
transform 1 0 12896 0 -1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap26_8
timestamp 1607194124
transform 1 0 12800 0 -1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap26_9
timestamp 1607194124
transform 1 0 14144 0 -1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap26_9
timestamp 1607194124
transform 1 0 14048 0 -1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_40
timestamp 1607194124
transform 1 0 13280 0 -1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_41
timestamp 1607194124
transform 1 0 14528 0 -1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_42
timestamp 1607194124
transform 1 0 15776 0 -1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap26_10
timestamp 1607194124
transform 1 0 15392 0 -1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap26_10
timestamp 1607194124
transform 1 0 15296 0 -1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap26_11
timestamp 1607194124
transform 1 0 16640 0 -1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap26_11
timestamp 1607194124
transform 1 0 16544 0 -1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap26_12
timestamp 1607194124
transform 1 0 17888 0 -1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap26_12
timestamp 1607194124
transform 1 0 17792 0 -1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_43
timestamp 1607194124
transform 1 0 17024 0 -1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_44
timestamp 1607194124
transform 1 0 18272 0 -1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_45
timestamp 1607194124
transform 1 0 19520 0 -1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap26_13
timestamp 1607194124
transform 1 0 19136 0 -1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap26_13
timestamp 1607194124
transform 1 0 19040 0 -1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_46
timestamp 1607194124
transform 1 0 20768 0 -1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap26_14
timestamp 1607194124
transform 1 0 20384 0 -1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap26_14
timestamp 1607194124
transform 1 0 20288 0 -1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap26_15
timestamp 1607194124
transform 1 0 21632 0 -1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap26_15
timestamp 1607194124
transform 1 0 21536 0 -1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_47
timestamp 1607194124
transform 1 0 22016 0 -1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap26_16
timestamp 1607194124
transform 1 0 22880 0 -1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap26_16
timestamp 1607194124
transform 1 0 22784 0 -1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap27_0
timestamp 1607194124
transform 1 0 2816 0 1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__mux2_1  mux_6
timestamp 1607194124
transform 1 0 1952 0 1 19042
box -38 -49 902 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_63
timestamp 1607194124
transform 1 0 3296 0 1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap27_0
timestamp 1607194124
transform 1 0 2912 0 1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_62
timestamp 1607194124
transform 1 0 4544 0 1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap27_1
timestamp 1607194124
transform 1 0 4160 0 1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap27_1
timestamp 1607194124
transform 1 0 4064 0 1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap27_2
timestamp 1607194124
transform 1 0 5408 0 1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap27_2
timestamp 1607194124
transform 1 0 5312 0 1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap27_3
timestamp 1607194124
transform 1 0 6656 0 1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap27_3
timestamp 1607194124
transform 1 0 6560 0 1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_61
timestamp 1607194124
transform 1 0 5792 0 1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_60
timestamp 1607194124
transform 1 0 7040 0 1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_59
timestamp 1607194124
transform 1 0 8288 0 1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap27_4
timestamp 1607194124
transform 1 0 7904 0 1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap27_4
timestamp 1607194124
transform 1 0 7808 0 1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap27_5
timestamp 1607194124
transform 1 0 9152 0 1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap27_5
timestamp 1607194124
transform 1 0 9056 0 1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap27_6
timestamp 1607194124
transform 1 0 10400 0 1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap27_6
timestamp 1607194124
transform 1 0 10304 0 1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_58
timestamp 1607194124
transform 1 0 9536 0 1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_57
timestamp 1607194124
transform 1 0 10784 0 1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_56
timestamp 1607194124
transform 1 0 12032 0 1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap27_7
timestamp 1607194124
transform 1 0 11648 0 1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap27_7
timestamp 1607194124
transform 1 0 11552 0 1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap27_8
timestamp 1607194124
transform 1 0 12896 0 1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap27_8
timestamp 1607194124
transform 1 0 12800 0 1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap27_9
timestamp 1607194124
transform 1 0 14144 0 1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap27_9
timestamp 1607194124
transform 1 0 14048 0 1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_55
timestamp 1607194124
transform 1 0 13280 0 1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_54
timestamp 1607194124
transform 1 0 14528 0 1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_53
timestamp 1607194124
transform 1 0 15776 0 1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap27_10
timestamp 1607194124
transform 1 0 15392 0 1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap27_10
timestamp 1607194124
transform 1 0 15296 0 1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap27_11
timestamp 1607194124
transform 1 0 16640 0 1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap27_11
timestamp 1607194124
transform 1 0 16544 0 1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap27_12
timestamp 1607194124
transform 1 0 17888 0 1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap27_12
timestamp 1607194124
transform 1 0 17792 0 1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_52
timestamp 1607194124
transform 1 0 17024 0 1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_51
timestamp 1607194124
transform 1 0 18272 0 1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_50
timestamp 1607194124
transform 1 0 19520 0 1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap27_13
timestamp 1607194124
transform 1 0 19136 0 1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap27_13
timestamp 1607194124
transform 1 0 19040 0 1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_49
timestamp 1607194124
transform 1 0 20768 0 1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap27_14
timestamp 1607194124
transform 1 0 20384 0 1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap27_14
timestamp 1607194124
transform 1 0 20288 0 1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap27_15
timestamp 1607194124
transform 1 0 21632 0 1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap27_15
timestamp 1607194124
transform 1 0 21536 0 1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_6_48
timestamp 1607194124
transform 1 0 22016 0 1 19042
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap27_16
timestamp 1607194124
transform 1 0 22880 0 1 19042
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap27_16
timestamp 1607194124
transform 1 0 22784 0 1 19042
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap28_0
timestamp 1607194124
transform 1 0 2816 0 -1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_51
timestamp 1607194124
transform 1 0 2048 0 -1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_50
timestamp 1607194124
transform 1 0 1952 0 -1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_0
timestamp 1607194124
transform 1 0 3296 0 -1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap28_0
timestamp 1607194124
transform 1 0 2912 0 -1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_1
timestamp 1607194124
transform 1 0 4544 0 -1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap28_1
timestamp 1607194124
transform 1 0 4160 0 -1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap28_1
timestamp 1607194124
transform 1 0 4064 0 -1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap28_2
timestamp 1607194124
transform 1 0 5408 0 -1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap28_2
timestamp 1607194124
transform 1 0 5312 0 -1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap28_3
timestamp 1607194124
transform 1 0 6656 0 -1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap28_3
timestamp 1607194124
transform 1 0 6560 0 -1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_2
timestamp 1607194124
transform 1 0 5792 0 -1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_3
timestamp 1607194124
transform 1 0 7040 0 -1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_4
timestamp 1607194124
transform 1 0 8288 0 -1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap28_4
timestamp 1607194124
transform 1 0 7904 0 -1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap28_4
timestamp 1607194124
transform 1 0 7808 0 -1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap28_5
timestamp 1607194124
transform 1 0 9152 0 -1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap28_5
timestamp 1607194124
transform 1 0 9056 0 -1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap28_6
timestamp 1607194124
transform 1 0 10400 0 -1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap28_6
timestamp 1607194124
transform 1 0 10304 0 -1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_5
timestamp 1607194124
transform 1 0 9536 0 -1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_6
timestamp 1607194124
transform 1 0 10784 0 -1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_7
timestamp 1607194124
transform 1 0 12032 0 -1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap28_7
timestamp 1607194124
transform 1 0 11648 0 -1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap28_7
timestamp 1607194124
transform 1 0 11552 0 -1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap28_8
timestamp 1607194124
transform 1 0 12896 0 -1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap28_8
timestamp 1607194124
transform 1 0 12800 0 -1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap28_9
timestamp 1607194124
transform 1 0 14144 0 -1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap28_9
timestamp 1607194124
transform 1 0 14048 0 -1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_8
timestamp 1607194124
transform 1 0 13280 0 -1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_9
timestamp 1607194124
transform 1 0 14528 0 -1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_10
timestamp 1607194124
transform 1 0 15776 0 -1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap28_10
timestamp 1607194124
transform 1 0 15392 0 -1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap28_10
timestamp 1607194124
transform 1 0 15296 0 -1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap28_11
timestamp 1607194124
transform 1 0 16640 0 -1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap28_11
timestamp 1607194124
transform 1 0 16544 0 -1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap28_12
timestamp 1607194124
transform 1 0 17888 0 -1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap28_12
timestamp 1607194124
transform 1 0 17792 0 -1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_11
timestamp 1607194124
transform 1 0 17024 0 -1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_12
timestamp 1607194124
transform 1 0 18272 0 -1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_13
timestamp 1607194124
transform 1 0 19520 0 -1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap28_13
timestamp 1607194124
transform 1 0 19136 0 -1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap28_13
timestamp 1607194124
transform 1 0 19040 0 -1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_14
timestamp 1607194124
transform 1 0 20768 0 -1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap28_14
timestamp 1607194124
transform 1 0 20384 0 -1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap28_14
timestamp 1607194124
transform 1 0 20288 0 -1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap28_15
timestamp 1607194124
transform 1 0 21632 0 -1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap28_15
timestamp 1607194124
transform 1 0 21536 0 -1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_15
timestamp 1607194124
transform 1 0 22016 0 -1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap28_16
timestamp 1607194124
transform 1 0 22880 0 -1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap28_16
timestamp 1607194124
transform 1 0 22784 0 -1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap29_0
timestamp 1607194124
transform 1 0 2816 0 1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__mux2_1  mux_5
timestamp 1607194124
transform 1 0 1952 0 1 20374
box -38 -49 902 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_31
timestamp 1607194124
transform 1 0 3296 0 1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap29_0
timestamp 1607194124
transform 1 0 2912 0 1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_30
timestamp 1607194124
transform 1 0 4544 0 1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap29_1
timestamp 1607194124
transform 1 0 4160 0 1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap29_1
timestamp 1607194124
transform 1 0 4064 0 1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap29_2
timestamp 1607194124
transform 1 0 5408 0 1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap29_2
timestamp 1607194124
transform 1 0 5312 0 1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap29_3
timestamp 1607194124
transform 1 0 6656 0 1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap29_3
timestamp 1607194124
transform 1 0 6560 0 1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_29
timestamp 1607194124
transform 1 0 5792 0 1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_28
timestamp 1607194124
transform 1 0 7040 0 1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_27
timestamp 1607194124
transform 1 0 8288 0 1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap29_4
timestamp 1607194124
transform 1 0 7904 0 1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap29_4
timestamp 1607194124
transform 1 0 7808 0 1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap29_5
timestamp 1607194124
transform 1 0 9152 0 1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap29_5
timestamp 1607194124
transform 1 0 9056 0 1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap29_6
timestamp 1607194124
transform 1 0 10400 0 1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap29_6
timestamp 1607194124
transform 1 0 10304 0 1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_26
timestamp 1607194124
transform 1 0 9536 0 1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_25
timestamp 1607194124
transform 1 0 10784 0 1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_24
timestamp 1607194124
transform 1 0 12032 0 1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap29_7
timestamp 1607194124
transform 1 0 11648 0 1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap29_7
timestamp 1607194124
transform 1 0 11552 0 1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap29_8
timestamp 1607194124
transform 1 0 12896 0 1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap29_8
timestamp 1607194124
transform 1 0 12800 0 1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap29_9
timestamp 1607194124
transform 1 0 14144 0 1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap29_9
timestamp 1607194124
transform 1 0 14048 0 1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_23
timestamp 1607194124
transform 1 0 13280 0 1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_22
timestamp 1607194124
transform 1 0 14528 0 1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_21
timestamp 1607194124
transform 1 0 15776 0 1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap29_10
timestamp 1607194124
transform 1 0 15392 0 1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap29_10
timestamp 1607194124
transform 1 0 15296 0 1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap29_11
timestamp 1607194124
transform 1 0 16640 0 1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap29_11
timestamp 1607194124
transform 1 0 16544 0 1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap29_12
timestamp 1607194124
transform 1 0 17888 0 1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap29_12
timestamp 1607194124
transform 1 0 17792 0 1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_20
timestamp 1607194124
transform 1 0 17024 0 1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_19
timestamp 1607194124
transform 1 0 18272 0 1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_18
timestamp 1607194124
transform 1 0 19520 0 1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap29_13
timestamp 1607194124
transform 1 0 19136 0 1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap29_13
timestamp 1607194124
transform 1 0 19040 0 1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_17
timestamp 1607194124
transform 1 0 20768 0 1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap29_14
timestamp 1607194124
transform 1 0 20384 0 1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap29_14
timestamp 1607194124
transform 1 0 20288 0 1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap29_15
timestamp 1607194124
transform 1 0 21632 0 1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap29_15
timestamp 1607194124
transform 1 0 21536 0 1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_5_16
timestamp 1607194124
transform 1 0 22016 0 1 20374
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap29_16
timestamp 1607194124
transform 1 0 22880 0 1 20374
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap29_16
timestamp 1607194124
transform 1 0 22784 0 1 20374
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap31_0
timestamp 1607194124
transform 1 0 2816 0 1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__mux2_1  mux_4
timestamp 1607194124
transform 1 0 1952 0 1 21706
box -38 -49 902 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap30_0
timestamp 1607194124
transform 1 0 2816 0 -1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_53
timestamp 1607194124
transform 1 0 2048 0 -1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_52
timestamp 1607194124
transform 1 0 1952 0 -1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_4_15
timestamp 1607194124
transform 1 0 3296 0 1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap31_0
timestamp 1607194124
transform 1 0 2912 0 1 21706
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_4_0
timestamp 1607194124
transform 1 0 3296 0 -1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap30_0
timestamp 1607194124
transform 1 0 2912 0 -1 21706
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_4_14
timestamp 1607194124
transform 1 0 4544 0 1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap31_1
timestamp 1607194124
transform 1 0 4160 0 1 21706
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap31_1
timestamp 1607194124
transform 1 0 4064 0 1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_4_1
timestamp 1607194124
transform 1 0 4544 0 -1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap30_1
timestamp 1607194124
transform 1 0 4160 0 -1 21706
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap30_1
timestamp 1607194124
transform 1 0 4064 0 -1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap31_2
timestamp 1607194124
transform 1 0 5408 0 1 21706
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap31_2
timestamp 1607194124
transform 1 0 5312 0 1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap30_2
timestamp 1607194124
transform 1 0 5408 0 -1 21706
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap30_2
timestamp 1607194124
transform 1 0 5312 0 -1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap31_3
timestamp 1607194124
transform 1 0 6656 0 1 21706
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap31_3
timestamp 1607194124
transform 1 0 6560 0 1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_4_13
timestamp 1607194124
transform 1 0 5792 0 1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap30_3
timestamp 1607194124
transform 1 0 6656 0 -1 21706
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap30_3
timestamp 1607194124
transform 1 0 6560 0 -1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_4_2
timestamp 1607194124
transform 1 0 5792 0 -1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_4_12
timestamp 1607194124
transform 1 0 7040 0 1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_4_3
timestamp 1607194124
transform 1 0 7040 0 -1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_4_11
timestamp 1607194124
transform 1 0 8288 0 1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap31_4
timestamp 1607194124
transform 1 0 7904 0 1 21706
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap31_4
timestamp 1607194124
transform 1 0 7808 0 1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_4_4
timestamp 1607194124
transform 1 0 8288 0 -1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap30_4
timestamp 1607194124
transform 1 0 7904 0 -1 21706
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap30_4
timestamp 1607194124
transform 1 0 7808 0 -1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap31_5
timestamp 1607194124
transform 1 0 9152 0 1 21706
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap31_5
timestamp 1607194124
transform 1 0 9056 0 1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap30_5
timestamp 1607194124
transform 1 0 9152 0 -1 21706
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap30_5
timestamp 1607194124
transform 1 0 9056 0 -1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap31_6
timestamp 1607194124
transform 1 0 10400 0 1 21706
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap31_6
timestamp 1607194124
transform 1 0 10304 0 1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_4_10
timestamp 1607194124
transform 1 0 9536 0 1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap30_6
timestamp 1607194124
transform 1 0 10400 0 -1 21706
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap30_6
timestamp 1607194124
transform 1 0 10304 0 -1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_4_5
timestamp 1607194124
transform 1 0 9536 0 -1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_4_9
timestamp 1607194124
transform 1 0 10784 0 1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_4_6
timestamp 1607194124
transform 1 0 10784 0 -1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_4_8
timestamp 1607194124
transform 1 0 12032 0 1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap31_7
timestamp 1607194124
transform 1 0 11648 0 1 21706
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap31_7
timestamp 1607194124
transform 1 0 11552 0 1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_4_7
timestamp 1607194124
transform 1 0 12032 0 -1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap30_7
timestamp 1607194124
transform 1 0 11648 0 -1 21706
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap30_7
timestamp 1607194124
transform 1 0 11552 0 -1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap31_8
timestamp 1607194124
transform 1 0 12896 0 1 21706
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap31_8
timestamp 1607194124
transform 1 0 12800 0 1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap30_8
timestamp 1607194124
transform 1 0 12896 0 -1 21706
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap30_8
timestamp 1607194124
transform 1 0 12800 0 -1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_86
timestamp 1607194124
transform 1 0 14144 0 1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_85
timestamp 1607194124
transform 1 0 13376 0 1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_84
timestamp 1607194124
transform 1 0 13280 0 1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_62
timestamp 1607194124
transform 1 0 14144 0 -1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_61
timestamp 1607194124
transform 1 0 13376 0 -1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_60
timestamp 1607194124
transform 1 0 13280 0 -1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_89
timestamp 1607194124
transform 1 0 15104 0 1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_88
timestamp 1607194124
transform 1 0 15008 0 1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_87
timestamp 1607194124
transform 1 0 14240 0 1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__fill_8  FILL_65
timestamp 1607194124
transform 1 0 15104 0 -1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_64
timestamp 1607194124
transform 1 0 15008 0 -1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_63
timestamp 1607194124
transform 1 0 14240 0 -1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__fill_8  FILL_91
timestamp 1607194124
transform 1 0 15968 0 1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_90
timestamp 1607194124
transform 1 0 15872 0 1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_67
timestamp 1607194124
transform 1 0 15968 0 -1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_66
timestamp 1607194124
transform 1 0 15872 0 -1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_93
timestamp 1607194124
transform 1 0 16832 0 1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_92
timestamp 1607194124
transform 1 0 16736 0 1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_69
timestamp 1607194124
transform 1 0 16832 0 -1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_68
timestamp 1607194124
transform 1 0 16736 0 -1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_95
timestamp 1607194124
transform 1 0 17696 0 1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_94
timestamp 1607194124
transform 1 0 17600 0 1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_71
timestamp 1607194124
transform 1 0 17696 0 -1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_70
timestamp 1607194124
transform 1 0 17600 0 -1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_97
timestamp 1607194124
transform 1 0 18560 0 1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_96
timestamp 1607194124
transform 1 0 18464 0 1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_73
timestamp 1607194124
transform 1 0 18560 0 -1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_72
timestamp 1607194124
transform 1 0 18464 0 -1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_99
timestamp 1607194124
transform 1 0 19424 0 1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_98
timestamp 1607194124
transform 1 0 19328 0 1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_75
timestamp 1607194124
transform 1 0 19424 0 -1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_74
timestamp 1607194124
transform 1 0 19328 0 -1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_101
timestamp 1607194124
transform 1 0 20288 0 1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_100
timestamp 1607194124
transform 1 0 20192 0 1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_77
timestamp 1607194124
transform 1 0 20288 0 -1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_76
timestamp 1607194124
transform 1 0 20192 0 -1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_103
timestamp 1607194124
transform 1 0 21152 0 1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_102
timestamp 1607194124
transform 1 0 21056 0 1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_79
timestamp 1607194124
transform 1 0 21152 0 -1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_78
timestamp 1607194124
transform 1 0 21056 0 -1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_105
timestamp 1607194124
transform 1 0 22016 0 1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_104
timestamp 1607194124
transform 1 0 21920 0 1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_81
timestamp 1607194124
transform 1 0 22016 0 -1 21706
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_80
timestamp 1607194124
transform 1 0 21920 0 -1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_1  FILL_107 $PDKPATH/libs.ref/sky130_fd_sc_ms/mag
timestamp 1607194124
transform 1 0 23168 0 1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_4  FILL_106 $PDKPATH/libs.ref/sky130_fd_sc_ms/mag
timestamp 1607194124
transform 1 0 22784 0 1 21706
box -38 -49 422 715
use sky130_fd_sc_ms__fill_1  FILL_83
timestamp 1607194124
transform 1 0 23168 0 -1 21706
box -38 -49 134 715
use sky130_fd_sc_ms__fill_4  FILL_82
timestamp 1607194124
transform 1 0 22784 0 -1 21706
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap32_0
timestamp 1607194124
transform 1 0 2816 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_55
timestamp 1607194124
transform 1 0 2048 0 -1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_54
timestamp 1607194124
transform 1 0 1952 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_3_0
timestamp 1607194124
transform 1 0 3296 0 -1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap32_0
timestamp 1607194124
transform 1 0 2912 0 -1 23038
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_3_1
timestamp 1607194124
transform 1 0 4544 0 -1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap32_1
timestamp 1607194124
transform 1 0 4160 0 -1 23038
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap32_1
timestamp 1607194124
transform 1 0 4064 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap32_2
timestamp 1607194124
transform 1 0 5408 0 -1 23038
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap32_2
timestamp 1607194124
transform 1 0 5312 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap32_3
timestamp 1607194124
transform 1 0 6656 0 -1 23038
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap32_3
timestamp 1607194124
transform 1 0 6560 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_3_2
timestamp 1607194124
transform 1 0 5792 0 -1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_3_3
timestamp 1607194124
transform 1 0 7040 0 -1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__fill_8  FILL_109
timestamp 1607194124
transform 1 0 8384 0 -1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_108
timestamp 1607194124
transform 1 0 8288 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap32_4
timestamp 1607194124
transform 1 0 7904 0 -1 23038
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap32_4
timestamp 1607194124
transform 1 0 7808 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_111
timestamp 1607194124
transform 1 0 9248 0 -1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_110
timestamp 1607194124
transform 1 0 9152 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_113
timestamp 1607194124
transform 1 0 10112 0 -1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_112
timestamp 1607194124
transform 1 0 10016 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_115
timestamp 1607194124
transform 1 0 10976 0 -1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_114
timestamp 1607194124
transform 1 0 10880 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_117
timestamp 1607194124
transform 1 0 11840 0 -1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_116
timestamp 1607194124
transform 1 0 11744 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_119
timestamp 1607194124
transform 1 0 12704 0 -1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_118
timestamp 1607194124
transform 1 0 12608 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_121
timestamp 1607194124
transform 1 0 13568 0 -1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_120
timestamp 1607194124
transform 1 0 13472 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_123
timestamp 1607194124
transform 1 0 14432 0 -1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_122
timestamp 1607194124
transform 1 0 14336 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_126
timestamp 1607194124
transform 1 0 16064 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_125
timestamp 1607194124
transform 1 0 15296 0 -1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_124
timestamp 1607194124
transform 1 0 15200 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_128
timestamp 1607194124
transform 1 0 16928 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_127
timestamp 1607194124
transform 1 0 16160 0 -1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__fill_8  FILL_131
timestamp 1607194124
transform 1 0 17888 0 -1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_130
timestamp 1607194124
transform 1 0 17792 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_129
timestamp 1607194124
transform 1 0 17024 0 -1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__fill_8  FILL_133
timestamp 1607194124
transform 1 0 18752 0 -1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_132
timestamp 1607194124
transform 1 0 18656 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_135
timestamp 1607194124
transform 1 0 19616 0 -1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_134
timestamp 1607194124
transform 1 0 19520 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_137
timestamp 1607194124
transform 1 0 20480 0 -1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_136
timestamp 1607194124
transform 1 0 20384 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_139
timestamp 1607194124
transform 1 0 21344 0 -1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_138
timestamp 1607194124
transform 1 0 21248 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_141
timestamp 1607194124
transform 1 0 22208 0 -1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_140
timestamp 1607194124
transform 1 0 22112 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_1  FILL_143
timestamp 1607194124
transform 1 0 23168 0 -1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_2  FILL_142 $PDKPATH/libs.ref/sky130_fd_sc_ms/mag
timestamp 1607194124
transform 1 0 22976 0 -1 23038
box -38 -49 230 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap33_0
timestamp 1607194124
transform 1 0 2816 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__mux2_1  mux_3
timestamp 1607194124
transform 1 0 1952 0 1 23038
box -38 -49 902 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_3_7
timestamp 1607194124
transform 1 0 3296 0 1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap33_0
timestamp 1607194124
transform 1 0 2912 0 1 23038
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_3_6
timestamp 1607194124
transform 1 0 4544 0 1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap33_1
timestamp 1607194124
transform 1 0 4160 0 1 23038
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap33_1
timestamp 1607194124
transform 1 0 4064 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap33_2
timestamp 1607194124
transform 1 0 5408 0 1 23038
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap33_2
timestamp 1607194124
transform 1 0 5312 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap33_3
timestamp 1607194124
transform 1 0 6656 0 1 23038
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap33_3
timestamp 1607194124
transform 1 0 6560 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_3_5
timestamp 1607194124
transform 1 0 5792 0 1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_3_4
timestamp 1607194124
transform 1 0 7040 0 1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__fill_8  FILL_145
timestamp 1607194124
transform 1 0 8384 0 1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_144
timestamp 1607194124
transform 1 0 8288 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap33_4
timestamp 1607194124
transform 1 0 7904 0 1 23038
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap33_4
timestamp 1607194124
transform 1 0 7808 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_147
timestamp 1607194124
transform 1 0 9248 0 1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_146
timestamp 1607194124
transform 1 0 9152 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_149
timestamp 1607194124
transform 1 0 10112 0 1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_148
timestamp 1607194124
transform 1 0 10016 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_151
timestamp 1607194124
transform 1 0 10976 0 1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_150
timestamp 1607194124
transform 1 0 10880 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_153
timestamp 1607194124
transform 1 0 11840 0 1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_152
timestamp 1607194124
transform 1 0 11744 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_155
timestamp 1607194124
transform 1 0 12704 0 1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_154
timestamp 1607194124
transform 1 0 12608 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_157
timestamp 1607194124
transform 1 0 13568 0 1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_156
timestamp 1607194124
transform 1 0 13472 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_159
timestamp 1607194124
transform 1 0 14432 0 1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_158
timestamp 1607194124
transform 1 0 14336 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_162
timestamp 1607194124
transform 1 0 16064 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_161
timestamp 1607194124
transform 1 0 15296 0 1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_160
timestamp 1607194124
transform 1 0 15200 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_164
timestamp 1607194124
transform 1 0 16928 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_163
timestamp 1607194124
transform 1 0 16160 0 1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__fill_8  FILL_167
timestamp 1607194124
transform 1 0 17888 0 1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_166
timestamp 1607194124
transform 1 0 17792 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_165
timestamp 1607194124
transform 1 0 17024 0 1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__fill_8  FILL_169
timestamp 1607194124
transform 1 0 18752 0 1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_168
timestamp 1607194124
transform 1 0 18656 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_171
timestamp 1607194124
transform 1 0 19616 0 1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_170
timestamp 1607194124
transform 1 0 19520 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_173
timestamp 1607194124
transform 1 0 20480 0 1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_172
timestamp 1607194124
transform 1 0 20384 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_175
timestamp 1607194124
transform 1 0 21344 0 1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_174
timestamp 1607194124
transform 1 0 21248 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_177
timestamp 1607194124
transform 1 0 22208 0 1 23038
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_176
timestamp 1607194124
transform 1 0 22112 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_1  FILL_179
timestamp 1607194124
transform 1 0 23168 0 1 23038
box -38 -49 134 715
use sky130_fd_sc_ms__fill_2  FILL_178
timestamp 1607194124
transform 1 0 22976 0 1 23038
box -38 -49 230 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap34_0
timestamp 1607194124
transform 1 0 2816 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_57
timestamp 1607194124
transform 1 0 2048 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_56
timestamp 1607194124
transform 1 0 1952 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_2_0
timestamp 1607194124
transform 1 0 3296 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap34_0
timestamp 1607194124
transform 1 0 2912 0 -1 24370
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_2_1
timestamp 1607194124
transform 1 0 4544 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap34_1
timestamp 1607194124
transform 1 0 4160 0 -1 24370
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap34_1
timestamp 1607194124
transform 1 0 4064 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap34_2
timestamp 1607194124
transform 1 0 5408 0 -1 24370
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap34_2
timestamp 1607194124
transform 1 0 5312 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_182
timestamp 1607194124
transform 1 0 6656 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_181
timestamp 1607194124
transform 1 0 5888 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_180
timestamp 1607194124
transform 1 0 5792 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_184
timestamp 1607194124
transform 1 0 7520 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_183
timestamp 1607194124
transform 1 0 6752 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__fill_8  FILL_187
timestamp 1607194124
transform 1 0 8480 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_186
timestamp 1607194124
transform 1 0 8384 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_185
timestamp 1607194124
transform 1 0 7616 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__fill_8  FILL_189
timestamp 1607194124
transform 1 0 9344 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_188
timestamp 1607194124
transform 1 0 9248 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_191
timestamp 1607194124
transform 1 0 10208 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_190
timestamp 1607194124
transform 1 0 10112 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_193
timestamp 1607194124
transform 1 0 11072 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_192
timestamp 1607194124
transform 1 0 10976 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_195
timestamp 1607194124
transform 1 0 11936 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_194
timestamp 1607194124
transform 1 0 11840 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_197
timestamp 1607194124
transform 1 0 12800 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_196
timestamp 1607194124
transform 1 0 12704 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_199
timestamp 1607194124
transform 1 0 13664 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_198
timestamp 1607194124
transform 1 0 13568 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_201
timestamp 1607194124
transform 1 0 14528 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_200
timestamp 1607194124
transform 1 0 14432 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_203
timestamp 1607194124
transform 1 0 15392 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_202
timestamp 1607194124
transform 1 0 15296 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_205
timestamp 1607194124
transform 1 0 16256 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_204
timestamp 1607194124
transform 1 0 16160 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_208
timestamp 1607194124
transform 1 0 17888 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_207
timestamp 1607194124
transform 1 0 17120 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_206
timestamp 1607194124
transform 1 0 17024 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_211
timestamp 1607194124
transform 1 0 18848 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_210
timestamp 1607194124
transform 1 0 18752 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_209
timestamp 1607194124
transform 1 0 17984 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__fill_8  FILL_213
timestamp 1607194124
transform 1 0 19712 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_212
timestamp 1607194124
transform 1 0 19616 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_215
timestamp 1607194124
transform 1 0 20576 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_214
timestamp 1607194124
transform 1 0 20480 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_217
timestamp 1607194124
transform 1 0 21440 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_216
timestamp 1607194124
transform 1 0 21344 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_219
timestamp 1607194124
transform 1 0 22304 0 -1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_218
timestamp 1607194124
transform 1 0 22208 0 -1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_2  FILL_220
timestamp 1607194124
transform 1 0 23072 0 -1 24370
box -38 -49 230 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap35_0
timestamp 1607194124
transform 1 0 2816 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__mux2_1  mux_2
timestamp 1607194124
transform 1 0 1952 0 1 24370
box -38 -49 902 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_2_3
timestamp 1607194124
transform 1 0 3296 0 1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap35_0
timestamp 1607194124
transform 1 0 2912 0 1 24370
box -38 -49 422 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_2_2
timestamp 1607194124
transform 1 0 4544 0 1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap35_1
timestamp 1607194124
transform 1 0 4160 0 1 24370
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap35_1
timestamp 1607194124
transform 1 0 4064 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap35_2
timestamp 1607194124
transform 1 0 5408 0 1 24370
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap35_2
timestamp 1607194124
transform 1 0 5312 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_223
timestamp 1607194124
transform 1 0 6656 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_222
timestamp 1607194124
transform 1 0 5888 0 1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_221
timestamp 1607194124
transform 1 0 5792 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_225
timestamp 1607194124
transform 1 0 7520 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_224
timestamp 1607194124
transform 1 0 6752 0 1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__fill_8  FILL_228
timestamp 1607194124
transform 1 0 8480 0 1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_227
timestamp 1607194124
transform 1 0 8384 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_226
timestamp 1607194124
transform 1 0 7616 0 1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__fill_8  FILL_230
timestamp 1607194124
transform 1 0 9344 0 1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_229
timestamp 1607194124
transform 1 0 9248 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_232
timestamp 1607194124
transform 1 0 10208 0 1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_231
timestamp 1607194124
transform 1 0 10112 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_234
timestamp 1607194124
transform 1 0 11072 0 1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_233
timestamp 1607194124
transform 1 0 10976 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_236
timestamp 1607194124
transform 1 0 11936 0 1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_235
timestamp 1607194124
transform 1 0 11840 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_238
timestamp 1607194124
transform 1 0 12800 0 1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_237
timestamp 1607194124
transform 1 0 12704 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_240
timestamp 1607194124
transform 1 0 13664 0 1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_239
timestamp 1607194124
transform 1 0 13568 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_242
timestamp 1607194124
transform 1 0 14528 0 1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_241
timestamp 1607194124
transform 1 0 14432 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_244
timestamp 1607194124
transform 1 0 15392 0 1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_243
timestamp 1607194124
transform 1 0 15296 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_246
timestamp 1607194124
transform 1 0 16256 0 1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_245
timestamp 1607194124
transform 1 0 16160 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_249
timestamp 1607194124
transform 1 0 17888 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_248
timestamp 1607194124
transform 1 0 17120 0 1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_247
timestamp 1607194124
transform 1 0 17024 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_252
timestamp 1607194124
transform 1 0 18848 0 1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_251
timestamp 1607194124
transform 1 0 18752 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_250
timestamp 1607194124
transform 1 0 17984 0 1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__fill_8  FILL_254
timestamp 1607194124
transform 1 0 19712 0 1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_253
timestamp 1607194124
transform 1 0 19616 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_256
timestamp 1607194124
transform 1 0 20576 0 1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_255
timestamp 1607194124
transform 1 0 20480 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_258
timestamp 1607194124
transform 1 0 21440 0 1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_257
timestamp 1607194124
transform 1 0 21344 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_260
timestamp 1607194124
transform 1 0 22304 0 1 24370
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_259
timestamp 1607194124
transform 1 0 22208 0 1 24370
box -38 -49 134 715
use sky130_fd_sc_ms__fill_2  FILL_261
timestamp 1607194124
transform 1 0 23072 0 1 24370
box -38 -49 230 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap36_0
timestamp 1607194124
transform 1 0 2816 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_59
timestamp 1607194124
transform 1 0 2048 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_58
timestamp 1607194124
transform 1 0 1952 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_1_0
timestamp 1607194124
transform 1 0 3296 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap36_0
timestamp 1607194124
transform 1 0 2912 0 -1 25702
box -38 -49 422 715
use sky130_fd_sc_ms__fill_8  FILL_263
timestamp 1607194124
transform 1 0 4640 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_262
timestamp 1607194124
transform 1 0 4544 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap36_1
timestamp 1607194124
transform 1 0 4160 0 -1 25702
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap36_1
timestamp 1607194124
transform 1 0 4064 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_265
timestamp 1607194124
transform 1 0 5504 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_264
timestamp 1607194124
transform 1 0 5408 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_267
timestamp 1607194124
transform 1 0 6368 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_266
timestamp 1607194124
transform 1 0 6272 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_269
timestamp 1607194124
transform 1 0 7232 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_268
timestamp 1607194124
transform 1 0 7136 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_271
timestamp 1607194124
transform 1 0 8096 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_270
timestamp 1607194124
transform 1 0 8000 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_273
timestamp 1607194124
transform 1 0 8960 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_272
timestamp 1607194124
transform 1 0 8864 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_275
timestamp 1607194124
transform 1 0 9824 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_274
timestamp 1607194124
transform 1 0 9728 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_277
timestamp 1607194124
transform 1 0 10688 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_276
timestamp 1607194124
transform 1 0 10592 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_279
timestamp 1607194124
transform 1 0 11552 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_278
timestamp 1607194124
transform 1 0 11456 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_282
timestamp 1607194124
transform 1 0 13184 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_281
timestamp 1607194124
transform 1 0 12416 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_280
timestamp 1607194124
transform 1 0 12320 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_285
timestamp 1607194124
transform 1 0 14144 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_284
timestamp 1607194124
transform 1 0 14048 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_283
timestamp 1607194124
transform 1 0 13280 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__fill_8  FILL_287
timestamp 1607194124
transform 1 0 15008 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_286
timestamp 1607194124
transform 1 0 14912 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_289
timestamp 1607194124
transform 1 0 15872 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_288
timestamp 1607194124
transform 1 0 15776 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_291
timestamp 1607194124
transform 1 0 16736 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_290
timestamp 1607194124
transform 1 0 16640 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_293
timestamp 1607194124
transform 1 0 17600 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_292
timestamp 1607194124
transform 1 0 17504 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_295
timestamp 1607194124
transform 1 0 18464 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_294
timestamp 1607194124
transform 1 0 18368 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_297
timestamp 1607194124
transform 1 0 19328 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_296
timestamp 1607194124
transform 1 0 19232 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_299
timestamp 1607194124
transform 1 0 20192 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_298
timestamp 1607194124
transform 1 0 20096 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_301
timestamp 1607194124
transform 1 0 21056 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_300
timestamp 1607194124
transform 1 0 20960 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_303
timestamp 1607194124
transform 1 0 21920 0 -1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_302
timestamp 1607194124
transform 1 0 21824 0 -1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_2  FILL_305
timestamp 1607194124
transform 1 0 23072 0 -1 25702
box -38 -49 230 715
use sky130_fd_sc_ms__fill_4  FILL_304
timestamp 1607194124
transform 1 0 22688 0 -1 25702
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap37_0
timestamp 1607194124
transform 1 0 2816 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__mux2_1  mux_1
timestamp 1607194124
transform 1 0 1952 0 1 25702
box -38 -49 902 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_1_1
timestamp 1607194124
transform 1 0 3296 0 1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap37_0
timestamp 1607194124
transform 1 0 2912 0 1 25702
box -38 -49 422 715
use sky130_fd_sc_ms__fill_8  FILL_307
timestamp 1607194124
transform 1 0 4640 0 1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_306
timestamp 1607194124
transform 1 0 4544 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap37_1
timestamp 1607194124
transform 1 0 4160 0 1 25702
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap37_1
timestamp 1607194124
transform 1 0 4064 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_309
timestamp 1607194124
transform 1 0 5504 0 1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_308
timestamp 1607194124
transform 1 0 5408 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_311
timestamp 1607194124
transform 1 0 6368 0 1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_310
timestamp 1607194124
transform 1 0 6272 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_313
timestamp 1607194124
transform 1 0 7232 0 1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_312
timestamp 1607194124
transform 1 0 7136 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_315
timestamp 1607194124
transform 1 0 8096 0 1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_314
timestamp 1607194124
transform 1 0 8000 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_317
timestamp 1607194124
transform 1 0 8960 0 1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_316
timestamp 1607194124
transform 1 0 8864 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_319
timestamp 1607194124
transform 1 0 9824 0 1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_318
timestamp 1607194124
transform 1 0 9728 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_321
timestamp 1607194124
transform 1 0 10688 0 1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_320
timestamp 1607194124
transform 1 0 10592 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_323
timestamp 1607194124
transform 1 0 11552 0 1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_322
timestamp 1607194124
transform 1 0 11456 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_326
timestamp 1607194124
transform 1 0 13184 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_325
timestamp 1607194124
transform 1 0 12416 0 1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_324
timestamp 1607194124
transform 1 0 12320 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_329
timestamp 1607194124
transform 1 0 14144 0 1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_328
timestamp 1607194124
transform 1 0 14048 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_327
timestamp 1607194124
transform 1 0 13280 0 1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__fill_8  FILL_331
timestamp 1607194124
transform 1 0 15008 0 1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_330
timestamp 1607194124
transform 1 0 14912 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_333
timestamp 1607194124
transform 1 0 15872 0 1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_332
timestamp 1607194124
transform 1 0 15776 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_335
timestamp 1607194124
transform 1 0 16736 0 1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_334
timestamp 1607194124
transform 1 0 16640 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_337
timestamp 1607194124
transform 1 0 17600 0 1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_336
timestamp 1607194124
transform 1 0 17504 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_339
timestamp 1607194124
transform 1 0 18464 0 1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_338
timestamp 1607194124
transform 1 0 18368 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_341
timestamp 1607194124
transform 1 0 19328 0 1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_340
timestamp 1607194124
transform 1 0 19232 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_343
timestamp 1607194124
transform 1 0 20192 0 1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_342
timestamp 1607194124
transform 1 0 20096 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_345
timestamp 1607194124
transform 1 0 21056 0 1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_344
timestamp 1607194124
transform 1 0 20960 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_347
timestamp 1607194124
transform 1 0 21920 0 1 25702
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_346
timestamp 1607194124
transform 1 0 21824 0 1 25702
box -38 -49 134 715
use sky130_fd_sc_ms__fill_2  FILL_349
timestamp 1607194124
transform 1 0 23072 0 1 25702
box -38 -49 230 715
use sky130_fd_sc_ms__fill_4  FILL_348
timestamp 1607194124
transform 1 0 22688 0 1 25702
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap38_0
timestamp 1607194124
transform 1 0 2816 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__mux2_1  mux_0
timestamp 1607194124
transform 1 0 1952 0 -1 27034
box -38 -49 902 715
use sky130_fd_sc_ms__dlygate4sd1_1  delay_0_0
timestamp 1607194124
transform 1 0 3296 0 -1 27034
box -38 -49 806 715
use sky130_fd_sc_ms__decap_4  decap38_0
timestamp 1607194124
transform 1 0 2912 0 -1 27034
box -38 -49 422 715
use sky130_fd_sc_ms__fill_8  FILL_351
timestamp 1607194124
transform 1 0 4640 0 -1 27034
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_350
timestamp 1607194124
transform 1 0 4544 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__decap_4  decap38_1
timestamp 1607194124
transform 1 0 4160 0 -1 27034
box -38 -49 422 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  tap38_1
timestamp 1607194124
transform 1 0 4064 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_353
timestamp 1607194124
transform 1 0 5504 0 -1 27034
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_352
timestamp 1607194124
transform 1 0 5408 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_355
timestamp 1607194124
transform 1 0 6368 0 -1 27034
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_354
timestamp 1607194124
transform 1 0 6272 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_357
timestamp 1607194124
transform 1 0 7232 0 -1 27034
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_356
timestamp 1607194124
transform 1 0 7136 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_359
timestamp 1607194124
transform 1 0 8096 0 -1 27034
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_358
timestamp 1607194124
transform 1 0 8000 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_361
timestamp 1607194124
transform 1 0 8960 0 -1 27034
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_360
timestamp 1607194124
transform 1 0 8864 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_363
timestamp 1607194124
transform 1 0 9824 0 -1 27034
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_362
timestamp 1607194124
transform 1 0 9728 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_365
timestamp 1607194124
transform 1 0 10688 0 -1 27034
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_364
timestamp 1607194124
transform 1 0 10592 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_367
timestamp 1607194124
transform 1 0 11552 0 -1 27034
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_366
timestamp 1607194124
transform 1 0 11456 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_370
timestamp 1607194124
transform 1 0 13184 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_369
timestamp 1607194124
transform 1 0 12416 0 -1 27034
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_368
timestamp 1607194124
transform 1 0 12320 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_373
timestamp 1607194124
transform 1 0 14144 0 -1 27034
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_372
timestamp 1607194124
transform 1 0 14048 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_371
timestamp 1607194124
transform 1 0 13280 0 -1 27034
box -38 -49 806 715
use sky130_fd_sc_ms__fill_8  FILL_375
timestamp 1607194124
transform 1 0 15008 0 -1 27034
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_374
timestamp 1607194124
transform 1 0 14912 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_377
timestamp 1607194124
transform 1 0 15872 0 -1 27034
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_376
timestamp 1607194124
transform 1 0 15776 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_379
timestamp 1607194124
transform 1 0 16736 0 -1 27034
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_378
timestamp 1607194124
transform 1 0 16640 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_381
timestamp 1607194124
transform 1 0 17600 0 -1 27034
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_380
timestamp 1607194124
transform 1 0 17504 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_383
timestamp 1607194124
transform 1 0 18464 0 -1 27034
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_382
timestamp 1607194124
transform 1 0 18368 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_385
timestamp 1607194124
transform 1 0 19328 0 -1 27034
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_384
timestamp 1607194124
transform 1 0 19232 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_387
timestamp 1607194124
transform 1 0 20192 0 -1 27034
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_386
timestamp 1607194124
transform 1 0 20096 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_389
timestamp 1607194124
transform 1 0 21056 0 -1 27034
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_388
timestamp 1607194124
transform 1 0 20960 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__fill_8  FILL_391
timestamp 1607194124
transform 1 0 21920 0 -1 27034
box -38 -49 806 715
use sky130_fd_sc_ms__tapvpwrvgnd_1  FILL_390
timestamp 1607194124
transform 1 0 21824 0 -1 27034
box -38 -49 134 715
use sky130_fd_sc_ms__fill_2  FILL_393
timestamp 1607194124
transform 1 0 23072 0 -1 27034
box -38 -49 230 715
use sky130_fd_sc_ms__fill_4  FILL_392
timestamp 1607194124
transform 1 0 22688 0 -1 27034
box -38 -49 422 715
<< labels >>
rlabel metal3 s 800 960 920 1216 6 inp_i
port 0 nsew default input
rlabel metal3 s 800 26936 920 27192 6 out_o
port 1 nsew default tristate
rlabel metal3 s 800 10888 920 11144 6 en_i[8]
port 2 nsew default input
rlabel metal3 s 800 16192 920 16448 6 en_i[7]
port 3 nsew default input
rlabel metal3 s 800 18912 920 19168 6 en_i[6]
port 4 nsew default input
rlabel metal3 s 800 20272 920 20528 6 en_i[5]
port 5 nsew default input
rlabel metal3 s 800 21632 920 21888 6 en_i[4]
port 6 nsew default input
rlabel metal3 s 800 22856 920 23112 6 en_i[3]
port 7 nsew default input
rlabel metal3 s 800 24216 920 24472 6 en_i[2]
port 8 nsew default input
rlabel metal3 s 800 25576 920 25832 6 en_i[1]
port 9 nsew default input
rlabel metal3 s 800 26256 920 26512 6 en_i[0]
port 10 nsew default input
rlabel metal5 s 1952 2692 23264 3012 6 VPWR
port 11 nsew default input
rlabel metal5 s 1952 20692 23264 21012 6 VGND
port 12 nsew default input
<< properties >>
string FIXED_BBOX 0 1 24102 28167
<< end >>
